magic
tech sky130A
magscale 1 2
timestamp 1758168748
<< metal1 >>
rect 333731 591775 338393 591829
rect 333731 591539 338103 591775
rect 338097 591485 338103 591539
rect 338393 591485 338399 591775
rect 257406 590510 257726 590516
rect 287844 590510 288164 590516
rect 257726 590190 287844 590510
rect 257406 590184 257726 590190
rect 287844 590184 288164 590190
rect 307105 590319 307275 590325
rect 307275 590149 307822 590319
rect 307105 590143 307275 590149
rect 338103 588877 338393 591485
rect 338097 588587 338103 588877
rect 338393 588587 338399 588877
rect 338103 588035 338393 588587
rect 338103 587739 338393 587745
rect 255190 510813 258688 510819
rect 148121 506934 255190 510813
rect 257054 507309 258688 507315
rect 148121 443358 151619 506934
rect 255190 506928 257054 506934
rect 306098 473946 310898 473952
rect 288563 472816 288569 473346
rect 289099 472816 291278 473346
rect 290878 469712 291518 472036
rect 296870 471945 306098 473946
rect 296158 471575 297401 471945
rect 297771 471575 306098 471945
rect 290872 469072 290878 469712
rect 291518 469072 291524 469712
rect 296870 469146 306098 471575
rect 306098 469140 310898 469146
rect 149102 437806 149422 443358
rect 149096 437486 149102 437806
rect 149422 437486 149428 437806
rect 149102 435938 149422 437486
rect 8362 261315 8493 261350
rect 8362 261245 8387 261315
rect 8457 261245 10882 261315
rect 8362 261225 8493 261245
rect 495812 140997 496688 141003
rect 488766 140867 489382 140873
rect 489382 140251 493474 140867
rect 494090 140251 495812 140867
rect 488766 140245 489382 140251
rect 496688 140121 501754 140997
rect 502630 140121 502636 140997
rect 495812 140115 496688 140121
rect 461961 139194 462131 139200
rect 462131 139024 462371 139194
rect 461961 139018 462131 139024
<< via1 >>
rect 338103 591485 338393 591775
rect 257406 590190 257726 590510
rect 287844 590190 288164 590510
rect 307105 590149 307275 590319
rect 338103 588587 338393 588877
rect 338103 587745 338393 588035
rect 255190 507315 258688 510813
rect 255190 506934 257054 507315
rect 288569 472816 289099 473346
rect 297401 471575 297771 471945
rect 290878 469072 291518 469712
rect 306098 469146 310898 473946
rect 149102 437486 149422 437806
rect 8387 261245 8457 261315
rect 488766 140251 489382 140867
rect 493474 140251 494090 140867
rect 495812 140121 496688 140997
rect 501754 140121 502630 140997
rect 461961 139024 462131 139194
<< metal2 >>
rect 306258 599752 344106 600184
rect 274222 595025 276722 595030
rect 274218 592535 274227 595025
rect 276717 593088 276726 595025
rect 306439 593349 306509 599752
rect 289209 593279 306509 593349
rect 307105 594295 308461 594465
rect 308631 594295 308640 594465
rect 275898 592535 276506 592538
rect 276717 592535 279366 593088
rect 274222 592520 279366 592535
rect 288821 592520 289156 592524
rect 274222 592515 289161 592520
rect 274222 592180 288821 592515
rect 289156 592180 289161 592515
rect 298334 592459 298404 593279
rect 274222 592175 289161 592180
rect 274222 590588 279366 592175
rect 288821 592171 289156 592175
rect 288674 591491 289634 591502
rect 291314 591491 291424 592202
rect 288674 591381 291424 591491
rect 257406 590510 257726 590519
rect 287849 590510 288159 590514
rect 257400 590190 257406 590510
rect 257726 590190 257732 590510
rect 287838 590190 287844 590510
rect 288164 590190 288170 590510
rect 257406 590181 257726 590190
rect 287849 590186 288159 590190
rect 288674 588421 289634 591381
rect 307105 590319 307275 594295
rect 338103 591775 338393 591784
rect 338103 591331 338393 591485
rect 338103 590554 338393 591041
rect 270797 587584 270806 588421
rect 271643 587584 289634 588421
rect 291314 587871 291404 590312
rect 307099 590149 307105 590319
rect 307275 590149 307281 590319
rect 338099 590274 338108 590554
rect 338388 590274 338397 590554
rect 338103 588877 338393 590274
rect 338103 588035 338393 588587
rect 288674 587574 289634 587584
rect 289849 587781 291404 587871
rect 234629 587111 234719 587120
rect 289849 587111 289939 587781
rect 338097 587745 338103 588035
rect 338393 587745 338399 588035
rect 234719 587021 289939 587111
rect 234629 587012 234719 587021
rect 236793 586799 236883 586808
rect 291983 586799 292073 587312
rect 236883 586709 292073 586799
rect 338103 586744 338393 587745
rect 236793 586700 236883 586709
rect 338099 586655 338108 586744
rect 338388 586655 338397 586744
rect 338099 586464 338103 586655
rect 338393 586464 338397 586655
rect 338103 586356 338393 586365
rect 240447 584312 240537 584321
rect 240537 584222 292101 584312
rect 240447 584213 240537 584222
rect 306322 583870 308492 584118
rect 265881 578736 265890 579201
rect 266355 579114 286811 579201
rect 266355 578822 286432 579114
rect 286724 578822 286811 579114
rect 266355 578736 286811 578822
rect 243956 571852 244176 571861
rect 291821 571852 292031 571856
rect 244176 571847 292036 571852
rect 244176 571637 291821 571847
rect 292031 571637 292036 571847
rect 244176 571632 292036 571637
rect 243956 571623 244176 571632
rect 291821 571628 292031 571632
rect 291888 570930 292326 571124
rect 247634 570925 292326 570930
rect 247634 570715 291977 570925
rect 292187 570715 292326 570925
rect 247634 570710 292326 570715
rect 249200 570363 249420 570710
rect 291888 570506 292326 570710
rect 249200 570274 249279 570363
rect 249381 570274 249420 570363
rect 249200 570045 249420 570054
rect 292245 568142 292455 568146
rect 229961 567922 229970 568142
rect 230190 568137 292460 568142
rect 230190 567927 292245 568137
rect 292455 567927 292460 568137
rect 230190 567922 292460 567927
rect 292245 567918 292455 567922
rect 255190 532282 258688 532287
rect 255186 528794 255195 532282
rect 258683 528794 258692 532282
rect 255190 528682 258688 528794
rect 257054 526818 258688 528682
rect 255190 510813 258688 526818
rect 255184 506934 255190 510813
rect 258688 507315 258694 510813
rect 257054 506934 257060 507315
rect 293564 478336 293674 583267
rect 306322 581858 306570 583870
rect 303290 581610 306570 581858
rect 308191 579849 308912 580019
rect 308191 575685 308361 579849
rect 332634 575685 332643 575847
rect 308191 575515 332643 575685
rect 332634 575353 332643 575515
rect 333137 575353 333146 575847
rect 343674 486512 344106 599752
rect 347632 585517 347792 585521
rect 461812 585517 461821 585645
rect 347627 585512 461821 585517
rect 347627 585352 347632 585512
rect 347792 585352 461821 585512
rect 347627 585347 461821 585352
rect 347632 585343 347792 585347
rect 461812 585219 461821 585347
rect 462247 585219 462256 585645
rect 371804 575847 372288 575851
rect 371799 575842 444605 575847
rect 371799 575358 371804 575842
rect 372288 575358 444605 575842
rect 371799 575353 444605 575358
rect 445099 575353 445333 575847
rect 371804 575349 372288 575353
rect 343674 485880 344106 486080
rect 415673 478336 416703 478340
rect 152395 477296 152404 478336
rect 153444 478331 416708 478336
rect 153444 477925 415673 478331
rect 153444 477735 291713 477925
rect 291903 477735 415673 477925
rect 153444 477301 415673 477735
rect 416703 477301 416708 478331
rect 153444 477296 416708 477301
rect 415673 477292 416703 477296
rect 343674 475891 344106 475896
rect 343670 475469 343679 475891
rect 344101 475469 344110 475891
rect 343674 475103 344106 475469
rect 153674 475079 422144 475103
rect 431840 475079 432768 475083
rect 153674 475074 432773 475079
rect 153674 474979 431840 475074
rect 153674 474789 292223 474979
rect 292413 474789 431840 474979
rect 153674 474666 431840 474789
rect 153737 472745 154377 474666
rect 343674 474096 344106 474666
rect 417287 474146 431840 474666
rect 432768 474146 432773 475074
rect 417287 474141 432773 474146
rect 431840 474137 432768 474141
rect 309343 473946 314133 473950
rect 288569 473346 289099 473352
rect 288560 472816 288569 473346
rect 289099 472816 289108 473346
rect 288569 472810 289099 472816
rect 153733 472115 153742 472745
rect 154372 472115 154381 472745
rect 153737 472110 154377 472115
rect 290878 469712 291518 469718
rect 290869 469072 290878 469712
rect 291518 469072 291527 469712
rect 290878 469066 291518 469072
rect 294388 464776 294498 472185
rect 296388 471302 296498 472203
rect 297401 471945 297771 471951
rect 297392 471575 297401 471945
rect 297771 471575 297780 471945
rect 297401 471569 297771 471575
rect 296388 471185 301718 471302
rect 296392 468802 301718 471185
rect 306092 469146 306098 473946
rect 310898 473941 314138 473946
rect 314133 469151 314138 473941
rect 310898 469146 314138 469151
rect 309343 469142 314133 469146
rect 299218 467044 301718 468802
rect 466781 467044 469271 467048
rect 299218 467039 469276 467044
rect 294170 459648 296431 464776
rect 299218 464549 466781 467039
rect 469271 464549 469276 467039
rect 299218 464544 469276 464549
rect 466781 464540 469271 464544
rect 453211 459648 455701 459652
rect 294050 459643 455706 459648
rect 294050 457153 453211 459643
rect 455701 457153 455706 459643
rect 294050 457148 455706 457153
rect 453211 457144 455701 457148
rect 151524 442682 151761 442691
rect 150755 442559 151009 442568
rect 150755 441805 151009 442305
rect 150827 441143 150937 441805
rect 151524 440952 151761 442445
rect 140131 439680 140241 439689
rect 140241 439570 141469 439680
rect 140131 439561 140241 439570
rect 149102 437806 149422 437812
rect 149102 437229 149422 437486
rect 149098 436919 149107 437229
rect 149417 436919 149426 437229
rect 149102 436914 149422 436919
rect 149102 436485 149422 436496
rect 149098 436175 149107 436485
rect 149417 436175 149426 436485
rect 149102 436164 149422 436175
rect 5660 336789 5772 336794
rect 5656 336687 5665 336789
rect 5767 336687 5776 336789
rect 5660 327595 5772 336687
rect 5660 327474 5772 327483
rect 8362 261315 8493 261350
rect 8362 261245 8387 261315
rect 8457 261245 8493 261315
rect 8362 261225 8493 261245
rect 9016 191337 9126 191346
rect 9126 191227 10882 191337
rect 9016 191218 9126 191227
rect 501754 140997 502630 141003
rect 493474 140867 494090 140873
rect 495806 140867 495812 140997
rect 488760 140251 488766 140867
rect 489382 140251 493474 140867
rect 494090 140251 495812 140867
rect 493474 140245 494090 140251
rect 495806 140121 495812 140251
rect 496688 140121 501754 140997
rect 502630 140121 503862 140997
rect 501754 140115 502630 140121
rect 461961 139833 462131 139842
rect 461961 139194 462131 139663
rect 461955 139024 461961 139194
rect 462131 139024 462137 139194
rect 126336 133775 127424 133780
rect 126332 132697 126341 133775
rect 127419 132697 127428 133775
rect 456062 133482 463212 133662
rect 462900 132745 463148 133482
rect 126336 129154 127424 132697
rect 144651 129154 145729 129158
rect 127424 129149 146798 129154
rect 127424 128071 144651 129149
rect 145729 128071 146798 129149
rect 460671 128894 460841 128903
rect 460841 128724 463461 128894
rect 460671 128715 460841 128724
rect 127424 128066 146798 128071
rect 126336 127220 127424 128066
rect 144651 128062 145729 128066
rect 19138 125184 19258 125193
rect 19138 118686 19258 125064
rect 21326 124954 21446 124963
rect 21326 120178 21446 124834
rect 27250 124898 27370 124907
rect 130318 124898 130428 124902
rect 27370 124893 130433 124898
rect 27370 124783 130318 124893
rect 130428 124783 130433 124893
rect 27370 124778 130433 124783
rect 27250 124769 27370 124778
rect 130318 124774 130428 124778
rect 24558 123672 24678 123681
rect 24678 123552 124366 123672
rect 24558 123543 24678 123552
rect 124246 120770 124366 123552
rect 134262 120770 134372 120774
rect 124246 120765 134377 120770
rect 124246 120655 134262 120765
rect 134372 120655 134377 120765
rect 124246 120650 134377 120655
rect 134262 120646 134372 120650
rect 138342 120178 138452 120182
rect 21326 120173 138457 120178
rect 21326 120063 138342 120173
rect 138452 120063 138457 120173
rect 21326 120058 138457 120063
rect 138342 120054 138452 120058
rect 142286 118686 142396 118690
rect 19138 118681 142401 118686
rect 19138 118571 142286 118681
rect 142396 118571 142401 118681
rect 19138 118566 142401 118571
rect 142286 118562 142396 118566
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 274227 592538 276717 595025
rect 308461 594295 308631 594465
rect 274227 592535 275898 592538
rect 276506 592535 276717 592538
rect 288821 592180 289156 592515
rect 257406 590190 257726 590510
rect 287849 590195 288159 590505
rect 338103 591485 338393 591775
rect 338103 591041 338393 591331
rect 270806 587584 271643 588421
rect 338108 590274 338388 590554
rect 234629 587021 234719 587111
rect 236793 586709 236883 586799
rect 338108 586655 338388 586744
rect 338103 586365 338393 586655
rect 240447 584222 240537 584312
rect 265890 578736 266355 579201
rect 286432 578822 286724 579114
rect 243956 571632 244176 571852
rect 291821 571637 292031 571847
rect 291977 570715 292187 570925
rect 249279 570274 249381 570363
rect 249200 570054 249420 570274
rect 229970 567922 230190 568142
rect 292245 567927 292455 568137
rect 255195 528794 258683 532282
rect 255190 526818 257054 528682
rect 332643 575353 333137 575847
rect 347632 585352 347792 585512
rect 461821 585219 462247 585645
rect 371804 575358 372288 575842
rect 444605 575353 445099 575847
rect 343674 486080 344106 486512
rect 152404 477296 153444 478336
rect 291713 477735 291903 477925
rect 415673 477301 416703 478331
rect 343679 475469 344101 475891
rect 292223 474789 292413 474979
rect 431840 474146 432768 475074
rect 288569 472816 289099 473346
rect 153742 472115 154372 472745
rect 290878 469072 291518 469712
rect 297401 471575 297771 471945
rect 309343 469151 310898 473941
rect 310898 469151 314133 473941
rect 466781 464549 469271 467039
rect 453211 457153 455701 459643
rect 150755 442305 151009 442559
rect 151524 442445 151761 442682
rect 140131 439570 140241 439680
rect 149107 436919 149417 437229
rect 149107 436175 149417 436485
rect 5665 336687 5767 336789
rect 5660 327483 5772 327595
rect 8387 261245 8457 261315
rect 9016 191227 9126 191337
rect 501754 140121 502630 140997
rect 461961 139663 462131 139833
rect 126341 132697 127419 133775
rect 126336 128066 127424 129154
rect 144651 128071 145729 129149
rect 460671 128724 460841 128894
rect 19138 125064 19258 125184
rect 21326 124834 21446 124954
rect 27250 124778 27370 124898
rect 130318 124783 130428 124893
rect 24558 123552 24678 123672
rect 134262 120655 134372 120765
rect 138342 120063 138452 120173
rect 142286 118571 142396 118681
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703390 418394 704800
rect 413394 703190 427730 703390
rect 413394 702300 418394 703190
rect 18694 696582 21194 702300
rect 18694 694082 66444 696582
rect 18694 693414 21194 694082
rect -800 682742 1700 685242
rect 63944 684066 66444 694082
rect 68940 690186 71440 702300
rect 122330 696788 124830 702300
rect 122330 696678 126146 696788
rect 122330 696013 124830 696678
rect 126036 696013 126146 696678
rect 122330 693513 173102 696013
rect 126036 690672 126146 693513
rect 68940 687686 168136 690186
rect -800 680242 61598 682742
rect 63944 681566 158432 684066
rect 59098 676618 61598 680242
rect 59098 674118 150778 676618
rect 6330 658270 8830 672796
rect 6330 655770 12018 658270
rect -800 643842 5110 648642
rect 148278 645006 150778 674118
rect 155932 650340 158432 681566
rect 165636 662826 168136 687686
rect 170602 669306 173102 693513
rect 177230 680264 179730 702300
rect 228438 698529 229478 698530
rect 228433 697491 228439 698529
rect 229477 697491 229483 698529
rect 331191 698285 332129 698286
rect 228438 686814 229478 697491
rect 331186 697349 331192 698285
rect 332128 697349 332134 698285
rect 228438 685774 316158 686814
rect 177230 677764 284582 680264
rect 170602 666806 276722 669306
rect 165636 660326 272166 662826
rect 155932 647840 265150 650340
rect 148278 642506 258688 645006
rect -800 633842 5110 638642
rect 256188 590510 258688 642506
rect 256188 590190 257406 590510
rect 257726 590190 258688 590510
rect 234624 587111 234724 587116
rect 234624 587021 234629 587111
rect 234719 587021 234724 587111
rect 234624 587016 234724 587021
rect 229965 568142 230195 568147
rect 229965 567922 229970 568142
rect 230190 567922 230195 568142
rect 229965 567917 230195 567922
rect -800 561902 1660 564242
rect -800 559442 1754 561902
rect -800 551902 1660 554242
rect -800 549442 1754 551902
rect 80622 533334 80734 533362
rect 229970 533334 230190 567917
rect 75398 533114 230190 533334
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 891 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect 1366 464931 1478 465323
rect 80622 464931 80734 533114
rect 234629 528757 234719 587016
rect 236788 586799 236888 586804
rect 236788 586709 236793 586799
rect 236883 586709 236888 586799
rect 236788 586704 236888 586709
rect 84431 528667 234719 528757
rect 1366 464874 80766 464931
rect -800 464819 80766 464874
rect -800 464762 1478 464819
rect -800 463580 480 463692
rect -800 462398 702 462510
rect 817 462376 1034 462476
rect 1134 462376 1140 462476
rect -800 425086 803 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 27458 421652
rect -800 420358 591 420470
rect 604 419288 690 419310
rect -800 419276 690 419288
rect -800 419176 717 419276
rect 817 419176 1034 419276
rect 1134 419176 1140 419276
rect -800 381864 979 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect 5660 379054 5772 419818
rect 1356 378430 1468 378793
rect -800 378318 1468 378430
rect 1356 377248 1468 378318
rect 24558 377248 24678 377756
rect -800 377136 824 377248
rect 1285 377136 24682 377248
rect 604 376076 690 376110
rect 604 376066 717 376076
rect -800 375976 717 376066
rect 817 375976 1034 376076
rect 1134 375976 1140 376076
rect -800 375954 690 375976
rect -800 338642 480 338754
rect -800 337460 480 337572
rect 5660 336789 5772 376032
rect 5660 336687 5665 336789
rect 5767 336687 5772 336789
rect 5660 336682 5772 336687
rect -800 336278 480 336390
rect 21326 335208 21446 335228
rect -800 335096 21476 335208
rect -800 333914 480 334026
rect -800 332810 654 332844
rect -800 332776 690 332810
rect -800 332732 717 332776
rect 542 332676 717 332732
rect 817 332676 1034 332776
rect 1134 332676 1140 332776
rect 542 332632 690 332676
rect 578 332608 690 332632
rect 5655 327595 5777 327600
rect 5655 327483 5660 327595
rect 5772 327483 5777 327595
rect 5655 327478 5777 327483
rect -800 295420 680 295532
rect -800 294238 480 294350
rect 5660 293381 5772 327478
rect 5660 293263 5772 293269
rect -800 293056 480 293168
rect 3192 291986 3304 292104
rect -800 291874 3840 291986
rect 3694 290804 3806 291874
rect -800 290692 1908 290804
rect 3672 290692 9839 290804
rect -800 289610 654 289622
rect -800 289576 690 289610
rect -800 289510 717 289576
rect 604 289498 717 289510
rect 660 289476 717 289498
rect 817 289476 1034 289576
rect 1134 289476 1140 289576
rect 9727 289082 9839 290692
rect 19138 289082 19258 291172
rect 9482 288962 19286 289082
rect 9727 288921 9839 288962
rect 8362 261320 8493 261350
rect 8362 261250 8382 261320
rect 8462 261250 8493 261320
rect 8362 261245 8387 261250
rect 8457 261245 8493 261250
rect 8362 261225 8493 261245
rect 19138 253335 19258 288962
rect 21326 253341 21446 335096
rect 24558 260523 24678 377136
rect 24553 260405 24559 260523
rect 24677 260405 24683 260523
rect 24558 260404 24678 260405
rect 27250 258973 27370 421540
rect 27245 258855 27251 258973
rect 27369 258855 27375 258973
rect 27250 258854 27370 258855
rect 19133 253217 19139 253335
rect 19257 253217 19263 253335
rect 21321 253223 21327 253341
rect 21445 253223 21451 253341
rect 21326 253222 21446 253223
rect 19138 253216 19258 253217
rect 5661 253173 5771 253178
rect 5660 253172 10882 253173
rect 5660 253062 5661 253172
rect 5771 253062 10882 253172
rect 5660 253061 10882 253062
rect 5661 253056 5771 253061
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect 84431 248964 84521 528667
rect 236793 525413 236883 586704
rect 240442 584312 240542 584317
rect 240442 584222 240447 584312
rect 240537 584222 240542 584312
rect 240442 584217 240542 584222
rect 90569 525323 236883 525413
rect -800 248852 84746 248964
rect 84431 248166 84521 248852
rect -800 247670 480 247782
rect 19138 247348 19258 247668
rect 604 246600 690 246610
rect -800 246576 690 246600
rect -800 246488 717 246576
rect 588 246476 717 246488
rect 817 246476 1034 246576
rect 1134 246476 1140 246576
rect 588 246407 690 246476
rect 7127 243720 7217 243726
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 7127 200580 7217 243630
rect 7127 200490 10882 200580
rect 10674 191537 10784 191543
rect 10784 191427 10882 191537
rect 10674 191421 10784 191427
rect 9011 191342 9131 191348
rect 9011 191227 9016 191232
rect 9126 191227 9131 191232
rect 9011 191222 9131 191227
rect 2175 177688 3090 177800
rect -800 172888 3090 177688
rect 2175 167688 3090 172888
rect -800 162888 3090 167688
rect 19138 125189 19258 247228
rect 21326 247552 21446 247558
rect 19133 125184 19263 125189
rect 19133 125064 19138 125184
rect 19258 125064 19263 125184
rect 19133 125059 19263 125064
rect 21326 124959 21446 247432
rect 24558 245562 24678 245568
rect 21321 124954 21451 124959
rect -800 124776 480 124888
rect 21321 124834 21326 124954
rect 21446 124834 21451 124954
rect 21321 124829 21451 124834
rect -800 123594 480 123706
rect 24558 123677 24678 245442
rect 27250 244826 27370 244832
rect 27250 124903 27370 244706
rect 27245 124898 27375 124903
rect 27245 124778 27250 124898
rect 27370 124778 27375 124898
rect 27245 124773 27375 124778
rect 24553 123672 24683 123677
rect 24553 123552 24558 123672
rect 24678 123552 24683 123672
rect 24553 123547 24683 123552
rect -800 122412 480 122524
rect 90569 121342 90659 525323
rect 240447 524479 240537 584217
rect 256188 578600 258688 590190
rect 243951 571852 244181 571857
rect 243951 571632 243956 571852
rect 244176 571632 244181 571852
rect 243951 571627 244181 571632
rect -800 121230 90659 121342
rect -800 120048 480 120160
rect 604 118984 690 119010
rect 445 118978 690 118984
rect -800 118976 690 118978
rect -800 118876 717 118976
rect 817 118876 1034 118976
rect 1134 118876 1140 118976
rect -800 118866 480 118876
rect 90569 113839 90659 121230
rect 96745 524389 240537 524479
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect 96745 78120 96835 524389
rect 243956 520756 244176 571627
rect 249200 570363 249420 570892
rect 249200 570279 249279 570363
rect 249195 570274 249279 570279
rect 249381 570279 249420 570363
rect 249381 570274 249425 570279
rect 249195 570054 249200 570274
rect 249420 570054 249425 570274
rect 249195 570049 249425 570054
rect 249200 569732 249420 570049
rect 102724 520536 244176 520756
rect -800 78008 96840 78120
rect -800 76826 480 76938
rect 604 75776 690 75810
rect 604 75756 717 75776
rect -800 75676 717 75756
rect 817 75676 1034 75776
rect 1134 75676 1140 75776
rect -800 75644 662 75676
rect 96745 71505 96835 78008
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect 102724 34898 102944 520536
rect 249274 518820 249386 569732
rect 255190 532282 258688 578600
rect 255190 528794 255195 532282
rect 258683 528794 258688 532282
rect 255190 528789 258688 528794
rect 262650 579201 265150 647840
rect 269666 588421 272166 660326
rect 269406 587584 270806 588421
rect 271643 587584 272166 588421
rect 269666 587380 272166 587584
rect 265885 579201 266360 579206
rect 262650 578736 265890 579201
rect 266355 578736 266360 579201
rect 255190 528687 257054 528789
rect 255185 528682 257059 528687
rect 255185 526818 255190 528682
rect 257054 526818 257059 528682
rect 255185 526813 257059 526818
rect -800 34786 102944 34898
rect 102724 34178 102944 34786
rect 110138 518708 249386 518820
rect -800 33604 480 33716
rect 604 32534 690 32577
rect -800 32422 690 32534
rect 604 32376 690 32422
rect 604 32298 717 32376
rect 660 32276 717 32298
rect 817 32276 1034 32376
rect 1134 32276 1140 32376
rect -800 16910 480 17022
rect 110138 16048 110250 518708
rect 262650 500548 265150 578736
rect 265885 578731 266360 578736
rect 137358 498048 265150 500548
rect 137784 441645 139433 498048
rect 269658 496755 272166 587380
rect 125868 439996 139433 441645
rect 139873 496322 272166 496755
rect 274222 595025 276722 666806
rect 274222 592535 274227 595025
rect 275898 592535 276506 592538
rect 276717 592535 276722 595025
rect 139873 496129 272158 496322
rect 125868 133775 127897 439996
rect 139873 439680 140499 496129
rect 269658 496118 272158 496129
rect 274222 494642 276722 592535
rect 282082 581021 284582 677764
rect 315118 608532 316158 685774
rect 331191 627679 332129 697349
rect 415894 693150 418394 702300
rect 427530 693150 427730 703190
rect 465394 702300 470394 704800
rect 415894 690650 456486 693150
rect 427530 688862 427730 690650
rect 331191 626741 432773 627679
rect 315118 607492 416708 608532
rect 308456 594465 308636 594470
rect 308456 594295 308461 594465
rect 308631 594295 347797 594465
rect 308456 594290 308636 594295
rect 288816 592515 289161 592520
rect 288816 592402 288821 592515
rect 288522 592292 288821 592402
rect 288816 592180 288821 592292
rect 289156 592402 289161 592515
rect 289696 592402 289804 592407
rect 289156 592401 289805 592402
rect 289156 592293 289696 592401
rect 289804 592293 289805 592401
rect 289156 592292 289805 592293
rect 289156 592180 289161 592292
rect 289696 592287 289804 592292
rect 288816 592175 289161 592180
rect 338103 592197 338393 592203
rect 338103 591780 338393 591907
rect 338098 591775 338398 591780
rect 338098 591485 338103 591775
rect 338393 591485 338398 591775
rect 338098 591480 338398 591485
rect 338103 591336 338393 591480
rect 338098 591331 338398 591336
rect 338098 591041 338103 591331
rect 338393 591041 338398 591331
rect 338098 591036 338398 591041
rect 338103 590554 338393 591036
rect 287845 590510 288163 590515
rect 287844 590509 288164 590510
rect 287844 590191 287845 590509
rect 288163 590191 288164 590509
rect 287844 590190 288164 590191
rect 338103 590274 338108 590554
rect 338388 590274 338393 590554
rect 287845 590185 288163 590190
rect 338103 586744 338393 590274
rect 338103 586660 338108 586744
rect 338098 586655 338108 586660
rect 338388 586660 338393 586744
rect 338388 586655 338398 586660
rect 338098 586365 338103 586655
rect 338393 586365 338398 586655
rect 338098 586360 338398 586365
rect 347627 585512 347797 594295
rect 347627 585352 347632 585512
rect 347792 585352 347797 585512
rect 347627 585347 347797 585352
rect 293114 581021 293204 584901
rect 282082 580719 293310 581021
rect 282082 576984 284582 580719
rect 293114 579712 293204 580719
rect 289792 579119 290092 579124
rect 286427 579118 290093 579119
rect 286427 579114 289792 579118
rect 286427 578822 286432 579114
rect 286724 578822 289792 579114
rect 286427 578818 289792 578822
rect 290092 578818 290093 579118
rect 286427 578817 290093 578818
rect 289792 578812 290092 578817
rect 308982 578275 309667 578281
rect 308982 577584 309667 577590
rect 282082 574484 291184 576984
rect 332638 575847 333142 575852
rect 332638 575353 332643 575847
rect 333137 575842 372293 575847
rect 333137 575358 371804 575842
rect 372288 575358 372293 575842
rect 333137 575353 372293 575358
rect 332638 575348 333142 575353
rect 141510 493746 276986 494642
rect 141510 441759 142406 493746
rect 274222 493676 276722 493746
rect 288684 490736 291184 574484
rect 291817 571852 292035 571857
rect 291816 571851 292036 571852
rect 291816 571633 291817 571851
rect 292035 571633 292036 571851
rect 291816 571632 292036 571633
rect 291817 571627 292035 571632
rect 291888 570929 292326 571124
rect 291888 570711 291973 570929
rect 292191 570711 292326 570929
rect 291888 570506 292326 570711
rect 292241 568142 292459 568147
rect 292240 568141 292460 568142
rect 292240 567923 292241 568141
rect 292459 567923 292460 568141
rect 292240 567922 292460 567923
rect 292241 567917 292459 567922
rect 148059 489641 291184 490736
rect 141510 441500 141829 441759
rect 142088 441500 142406 441759
rect 141510 440950 142406 441500
rect 148349 441443 148864 489641
rect 150248 478336 151288 484306
rect 152399 478336 153449 478341
rect 149648 477296 152404 478336
rect 153444 477296 153449 478336
rect 150248 442824 151288 477296
rect 152399 477291 153449 477296
rect 288684 473608 291184 489641
rect 343669 486512 344111 486517
rect 343669 486080 343674 486512
rect 344106 486080 344111 486512
rect 343669 486075 344111 486080
rect 291708 477925 291908 477930
rect 291708 477735 291713 477925
rect 291903 477735 291908 477925
rect 153737 472745 154377 473120
rect 288558 472811 288564 473351
rect 289094 473346 289104 473351
rect 289099 472816 289104 473346
rect 289718 473208 290319 473608
rect 289094 472811 289104 472816
rect 153737 472115 153742 472745
rect 154372 472115 154377 472745
rect 150755 442564 151009 442824
rect 151519 442682 151766 442687
rect 153737 442682 154377 472115
rect 289973 471179 290063 473208
rect 291708 472920 291908 477735
rect 343674 475891 344106 486075
rect 415668 478331 416708 607492
rect 415668 477301 415673 478331
rect 416703 477301 416708 478331
rect 415668 477296 416708 477301
rect 343674 475469 343679 475891
rect 344101 475469 344106 475891
rect 343674 475464 344106 475469
rect 431835 475074 432773 626741
rect 444600 575847 445104 575852
rect 453206 575847 455706 690650
rect 461816 585645 462252 585650
rect 466776 585645 469276 702300
rect 510594 698160 515394 704800
rect 520594 698160 525394 704800
rect 566594 702300 571594 704800
rect 566594 690142 571476 702300
rect 554148 689282 571476 690142
rect 547286 669777 548114 669782
rect 561083 669777 561913 689282
rect 566594 674025 571476 689282
rect 574600 682984 582176 683000
rect 574600 682800 584800 682984
rect 574440 682402 584800 682800
rect 574440 678818 575238 682402
rect 582000 678818 584800 682402
rect 574440 678370 584800 678818
rect 582300 677984 584800 678370
rect 547285 669776 561913 669777
rect 547285 668948 547286 669776
rect 548114 668948 561913 669776
rect 566588 669143 566594 674025
rect 571476 669143 571482 674025
rect 547285 668947 561913 668948
rect 547286 668942 548114 668947
rect 534554 639784 536034 644584
rect 540834 639784 584800 644584
rect 534554 629784 536768 634584
rect 541568 629784 584800 634584
rect 577935 625014 578045 629784
rect 577930 624906 577936 625014
rect 578044 624906 578050 625014
rect 577935 624905 578045 624906
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 461816 585219 461821 585645
rect 462247 585219 469276 585645
rect 461816 585214 462252 585219
rect 444600 575353 444605 575847
rect 445099 575353 455706 575847
rect 444600 575348 445104 575353
rect 292218 474979 292418 474984
rect 292218 474789 292223 474979
rect 292413 474789 292418 474979
rect 292218 472964 292418 474789
rect 431835 474146 431840 475074
rect 432768 474146 432773 475074
rect 431835 474141 432773 474146
rect 314131 473946 318929 473951
rect 309338 473945 318930 473946
rect 309338 473941 314131 473945
rect 291188 471179 291278 472125
rect 297396 471945 297406 471950
rect 297396 471575 297401 471945
rect 297396 471570 297406 471575
rect 297776 471570 297782 471950
rect 289973 471089 291278 471179
rect 290873 469712 290883 469717
rect 290873 469072 290878 469712
rect 290873 469067 290883 469072
rect 291523 469067 291529 469717
rect 309338 469151 309343 473941
rect 309338 469147 314131 469151
rect 318929 469147 318930 473945
rect 309338 469146 318930 469147
rect 314131 469141 318929 469146
rect 453206 462143 455706 575353
rect 466776 467039 469276 585219
rect 583520 584744 584800 584856
rect 581085 583562 584800 583674
rect 582340 555352 584800 555362
rect 581085 554285 584800 555352
rect 578987 550570 584800 554285
rect 582340 550562 584800 550570
rect 581085 544277 584800 545362
rect 578987 540562 584800 544277
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 534554 494140 584800 494252
rect 466776 464549 466781 467039
rect 469271 464549 469276 467039
rect 453206 459643 461052 462143
rect 453206 457153 453211 459643
rect 455701 457153 455706 459643
rect 453206 457148 455706 457153
rect 150750 442559 151014 442564
rect 150750 442305 150755 442559
rect 151009 442305 151014 442559
rect 151519 442445 151524 442682
rect 151761 442445 154377 442682
rect 151519 442440 151766 442445
rect 150750 442300 151014 442305
rect 153737 442243 154377 442445
rect 148349 441353 150467 441443
rect 148349 441141 148864 441353
rect 139873 439570 140131 439680
rect 140241 439570 140499 439680
rect 139873 439312 140499 439570
rect 149102 437233 149422 437234
rect 149097 436915 149103 437233
rect 149421 436915 149427 437233
rect 149102 436914 149422 436915
rect 149102 436489 149422 436490
rect 149097 436171 149103 436489
rect 149421 436171 149427 436489
rect 149102 436170 149422 436171
rect 125868 132697 126341 133775
rect 127419 132697 127897 133775
rect 125868 129154 127897 132697
rect 125868 128636 126336 129154
rect 126331 128066 126336 128636
rect 127424 128636 127897 129154
rect 127424 128066 127429 128636
rect 126331 128061 127429 128066
rect 130313 124893 130433 131530
rect 130313 124783 130318 124893
rect 130428 124783 130433 124893
rect 130313 124778 130433 124783
rect 134257 120765 134377 131548
rect 134257 120655 134262 120765
rect 134372 120655 134377 120765
rect 134257 120650 134377 120655
rect 138337 120173 138457 131448
rect 138337 120063 138342 120173
rect 138452 120063 138457 120173
rect 138337 120058 138457 120063
rect 142281 118681 142401 131424
rect 144647 129154 145733 129159
rect 144646 129153 145734 129154
rect 144646 128067 144647 129153
rect 145733 128067 145734 129153
rect 460671 128899 460841 459643
rect 466776 459040 469276 464549
rect 461524 456540 469276 459040
rect 461823 139833 462269 456540
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 534554 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 582476 364801 582546 364886
rect 582482 364786 582546 364801
rect 582646 364786 582787 364886
rect 582918 364784 584800 364896
rect 583520 363602 584800 363714
rect 534554 362420 584800 362532
rect 503116 141266 504528 141271
rect 499369 139852 499375 141266
rect 500789 141265 504529 141266
rect 500789 140997 503116 141265
rect 500789 140121 501754 140997
rect 502630 140121 503116 140997
rect 500789 139853 503116 140121
rect 504528 140997 504529 141265
rect 504528 140121 505628 140997
rect 506504 140121 506510 140997
rect 504528 139853 504529 140121
rect 500789 139852 504529 139853
rect 503116 139847 504528 139852
rect 461823 139663 461961 139833
rect 462131 139663 462269 139833
rect 461823 139525 462269 139663
rect 460666 128894 460846 128899
rect 456132 128660 458042 128780
rect 460666 128724 460671 128894
rect 460841 128724 460846 128894
rect 460666 128719 460846 128724
rect 144646 128066 145734 128067
rect 144647 128061 145733 128066
rect 457922 126066 458042 128660
rect 463525 126465 463531 127150
rect 464216 126465 464222 127150
rect 534554 126066 534666 362420
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583093 358874 584800 358986
rect 542712 344507 542832 344508
rect 542640 344387 570754 344507
rect 457922 125946 534814 126066
rect 542712 124836 542832 344387
rect 570634 317310 570754 344387
rect 583138 319656 584800 319674
rect 582918 319646 584800 319656
rect 582476 319561 582546 319646
rect 582482 319546 582546 319561
rect 582646 319546 582787 319646
rect 582887 319562 584800 319646
rect 582887 319546 583364 319562
rect 582918 319544 583364 319546
rect 583520 318380 584800 318492
rect 570463 317198 584800 317310
rect 570634 316193 570754 317198
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 581256 313652 584800 313764
rect 456202 124716 542832 124836
rect 544022 276244 580683 276364
rect 544022 120756 544142 276244
rect 580563 272888 580683 276244
rect 582918 275252 583364 275256
rect 582918 275246 584800 275252
rect 582476 275161 582546 275246
rect 582482 275146 582546 275161
rect 582646 275146 582787 275246
rect 582887 275146 584800 275246
rect 582918 275144 584800 275146
rect 583156 275140 584800 275144
rect 583520 273958 584800 274070
rect 580563 272776 584800 272888
rect 580563 272105 580683 272776
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 582310 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 578645 198242 579069 198298
rect 552812 196966 579468 198242
rect 552812 196230 554140 196966
rect 550944 191768 554140 196230
rect 578296 196230 579468 196966
rect 578296 191768 584800 196230
rect 550944 191430 584800 191768
rect 552812 190928 579468 191430
rect 553276 187154 558076 190928
rect 551320 186340 579660 187154
rect 551320 186230 553050 186340
rect 550944 181430 553050 186230
rect 551320 181150 553050 181430
rect 576862 186230 579660 186340
rect 576862 181430 584800 186230
rect 576862 181150 579660 181430
rect 551320 180540 579660 181150
rect 553276 164626 558076 180540
rect 552718 164209 558786 164626
rect 552718 159411 553277 164209
rect 558075 159411 558786 164209
rect 552718 158880 558786 159411
rect 582340 149347 584800 151630
rect 576060 146887 584800 149347
rect 582340 146830 584800 146887
rect 582340 139290 584800 141630
rect 576060 136830 584800 139290
rect 456280 120636 544278 120756
rect 544022 120620 544142 120636
rect 461464 119798 571679 119918
rect 142281 118571 142286 118681
rect 142396 118571 142401 118681
rect 142281 118566 142401 118571
rect 461620 116812 461740 119798
rect 456242 116692 461740 116812
rect 571559 92866 571679 119798
rect 582918 95246 583364 95256
rect 582476 95161 582546 95246
rect 582482 95146 582546 95161
rect 582646 95146 582787 95246
rect 582887 95230 583364 95246
rect 582887 95146 584800 95230
rect 582918 95144 584800 95146
rect 583184 95118 584800 95144
rect 583520 93936 584800 94048
rect 570398 92754 584800 92866
rect 571559 89505 571679 92754
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 583520 16910 584800 17022
rect 10662 15936 110250 16048
rect -800 15728 480 15840
rect -800 14546 480 14658
rect 10662 13476 10774 15936
rect 583520 15728 584800 15840
rect 583520 14546 584800 14658
rect -800 13364 10882 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11010 674 11112
rect -800 11000 690 11010
rect 583520 11000 584800 11112
rect 562 10976 690 11000
rect 562 10876 717 10976
rect 817 10876 1034 10976
rect 1134 10876 1140 10976
rect 562 10868 674 10876
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 1849 8748
rect 583520 8636 584800 8748
rect -800 7454 584 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 354 4020
rect 466 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 717 419176 817 419276
rect 717 375976 817 376076
rect 717 332676 817 332776
rect 717 289476 817 289576
rect 717 246476 817 246576
rect 717 118876 817 118976
rect 717 75676 817 75776
rect 717 32276 817 32376
rect 582787 319546 582887 319646
rect 582787 275146 582887 275246
rect 582787 95146 582887 95246
rect 717 10876 817 10976
<< via3 >>
rect 228439 697491 229477 698529
rect 331192 697349 332128 698285
rect 1034 462376 1134 462476
rect 1034 419176 1134 419276
rect 1034 375976 1134 376076
rect 1034 332676 1134 332776
rect 5660 293269 5772 293381
rect 1034 289476 1134 289576
rect 8382 261315 8462 261320
rect 8382 261250 8387 261315
rect 8387 261250 8457 261315
rect 8457 261250 8462 261315
rect 24559 260405 24677 260523
rect 27251 258855 27369 258973
rect 19139 253217 19257 253335
rect 21327 253223 21445 253341
rect 5661 253062 5771 253172
rect 19138 247228 19258 247348
rect 1034 246476 1134 246576
rect 7127 243630 7217 243720
rect 10674 191427 10784 191537
rect 9011 191337 9131 191342
rect 9011 191232 9016 191337
rect 9016 191232 9126 191337
rect 9126 191232 9131 191337
rect 21326 247432 21446 247552
rect 24558 245442 24678 245562
rect 27250 244706 27370 244826
rect 1034 118876 1134 118976
rect 1034 75676 1134 75776
rect 1034 32276 1134 32376
rect 289696 592293 289804 592401
rect 338103 591907 338393 592197
rect 287845 590505 288163 590509
rect 287845 590195 287849 590505
rect 287849 590195 288159 590505
rect 288159 590195 288163 590505
rect 287845 590191 288163 590195
rect 289792 578818 290092 579118
rect 308982 577590 309667 578275
rect 291817 571847 292035 571851
rect 291817 571637 291821 571847
rect 291821 571637 292031 571847
rect 292031 571637 292035 571847
rect 291817 571633 292035 571637
rect 291973 570925 292191 570929
rect 291973 570715 291977 570925
rect 291977 570715 292187 570925
rect 292187 570715 292191 570925
rect 291973 570711 292191 570715
rect 292241 568137 292459 568141
rect 292241 567927 292245 568137
rect 292245 567927 292455 568137
rect 292455 567927 292459 568137
rect 292241 567923 292459 567927
rect 141829 441500 142088 441759
rect 288564 473346 289094 473351
rect 288564 472816 288569 473346
rect 288569 472816 289094 473346
rect 288564 472811 289094 472816
rect 575238 678818 582000 682402
rect 547286 668948 548114 669776
rect 566594 669143 571476 674025
rect 536034 639784 540834 644584
rect 536768 629784 541568 634584
rect 577936 624906 578044 625014
rect 314131 473941 318929 473945
rect 297406 471945 297776 471950
rect 297406 471575 297771 471945
rect 297771 471575 297776 471945
rect 297406 471570 297776 471575
rect 290883 469712 291523 469717
rect 290883 469072 291518 469712
rect 291518 469072 291523 469712
rect 290883 469067 291523 469072
rect 314131 469151 314133 473941
rect 314133 469151 318929 473941
rect 314131 469147 318929 469151
rect 149103 437229 149421 437233
rect 149103 436919 149107 437229
rect 149107 436919 149417 437229
rect 149417 436919 149421 437229
rect 149103 436915 149421 436919
rect 149103 436485 149421 436489
rect 149103 436175 149107 436485
rect 149107 436175 149417 436485
rect 149417 436175 149421 436485
rect 149103 436171 149421 436175
rect 144647 129149 145733 129153
rect 144647 128071 144651 129149
rect 144651 128071 145729 129149
rect 145729 128071 145733 129149
rect 144647 128067 145733 128071
rect 582546 364786 582646 364886
rect 499375 139852 500789 141266
rect 503116 139853 504528 141265
rect 505628 140121 506504 140997
rect 463531 126465 464216 127150
rect 582546 319546 582646 319646
rect 582546 275146 582646 275246
rect 554140 191768 578296 196966
rect 553050 181150 576862 186340
rect 553277 159411 558075 164209
rect 582546 95146 582646 95246
rect 1034 10876 1134 10976
rect 354 3908 466 4020
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329590 701834 334030 701858
rect 229190 699708 231180 699960
rect 229190 698530 229597 699708
rect 228350 698529 229597 698530
rect 228350 697491 228439 698529
rect 229477 697552 229597 698529
rect 229477 697491 231180 697552
rect 228350 697490 231180 697491
rect 229190 697460 231180 697490
rect 329590 697442 329614 701834
rect 334006 697442 334030 701834
rect 329590 697349 331192 697442
rect 332128 697349 334030 697442
rect 329590 694172 334030 697349
rect 574553 682650 577887 682687
rect 574553 682402 582200 682650
rect 574553 678818 575238 682402
rect 582000 678818 582200 682402
rect 574553 678570 582200 678818
rect 566593 674025 571477 674026
rect 1033 462476 1135 462477
rect 2440 462476 2540 462606
rect 1033 462376 1034 462476
rect 1134 462376 2540 462476
rect 1033 462375 1135 462376
rect 2440 422228 2540 462376
rect 8387 422228 8457 672796
rect 9016 422228 9126 672796
rect 10674 422228 10784 672796
rect 478811 669776 566594 674025
rect 478811 668948 547286 669776
rect 548114 669143 566594 669776
rect 571476 669143 571477 674025
rect 548114 668948 548311 669143
rect 566593 669142 571477 669143
rect 478811 668947 548311 668948
rect 478811 597477 483889 668947
rect 574553 665164 577887 678570
rect 303894 592806 304214 596286
rect 339885 593924 483889 597477
rect 335215 593094 483889 593924
rect 303894 592534 303918 592806
rect 304190 592534 304214 592806
rect 303894 592510 304214 592534
rect 289695 592401 292013 592402
rect 289695 592293 289696 592401
rect 289804 592293 292013 592401
rect 339885 592399 483889 593094
rect 490227 661830 577887 665164
rect 289695 592292 292013 592293
rect 338102 592197 338394 592198
rect 338102 591907 338103 592197
rect 338393 591907 338394 592197
rect 338102 591906 338394 591907
rect 287844 591878 292634 591902
rect 287844 591606 292338 591878
rect 292610 591606 292634 591878
rect 287844 591582 292634 591606
rect 287844 590509 288164 591582
rect 287844 590191 287845 590509
rect 288163 590191 288164 590509
rect 287844 590190 288164 590191
rect 338103 586460 338393 591906
rect 293834 579119 293944 582037
rect 289791 579118 294040 579119
rect 289791 578818 289792 579118
rect 290092 578818 294040 579118
rect 289791 578817 294040 578818
rect 294534 571852 294754 581972
rect 291816 571851 294754 571852
rect 291816 571633 291817 571851
rect 292035 571633 294754 571851
rect 291816 571632 294754 571633
rect 291888 570930 292326 571124
rect 297534 570930 297754 582004
rect 291888 570929 297754 570930
rect 291888 570711 291973 570929
rect 292191 570711 297754 570929
rect 291888 570710 297754 570711
rect 291888 570506 292326 570710
rect 300534 568142 300754 582016
rect 308981 578275 309668 578276
rect 308981 577590 308982 578275
rect 309667 577590 309668 578275
rect 308981 577589 309668 577590
rect 292240 568141 300754 568142
rect 292240 567923 292241 568141
rect 292459 567923 300754 568141
rect 292240 567922 300754 567923
rect 308982 557285 309667 577589
rect 314130 473945 339500 473946
rect 289093 473351 289095 473352
rect 289094 472811 289095 473351
rect 289093 472810 289095 472811
rect 297405 471950 297407 471951
rect 297405 471570 297406 471950
rect 297405 471569 297407 471570
rect 290882 469717 290884 469718
rect 290882 469067 290883 469717
rect 314130 469147 314131 473945
rect 318929 473922 339500 473945
rect 318929 469170 334724 473922
rect 339476 469170 339500 473922
rect 318929 469147 339500 469170
rect 314130 469146 339500 469147
rect 290882 469066 290884 469067
rect 141828 441759 142089 441760
rect 141828 441500 141829 441759
rect 142088 441500 142089 441759
rect 141828 439981 142089 441500
rect 149102 437233 149422 437234
rect 149102 436915 149103 437233
rect 149421 436915 149422 437233
rect 149102 436914 149422 436915
rect 149102 436489 149422 436490
rect 149102 436171 149103 436489
rect 149421 436171 149422 436489
rect 149102 436170 149422 436171
rect 1033 419276 1135 419277
rect 2440 419276 2540 419818
rect 1033 419176 1034 419276
rect 1134 419176 2540 419276
rect 1033 419175 1135 419176
rect 1033 376076 1135 376077
rect 2440 376076 2540 419176
rect 8387 379054 8457 419818
rect 9016 379054 9126 419818
rect 10674 379054 10784 419818
rect 1033 375976 1034 376076
rect 1134 375976 2540 376076
rect 1033 375975 1135 375976
rect 1033 332776 1135 332777
rect 2440 332776 2540 375976
rect 1033 332676 1034 332776
rect 1134 332676 2540 332776
rect 1033 332675 1135 332676
rect 1033 289576 1135 289577
rect 2440 289576 2540 332676
rect 5659 293381 5773 293382
rect 5659 293269 5660 293381
rect 5772 293269 5773 293381
rect 5659 293268 5773 293269
rect 1033 289476 1034 289576
rect 1134 289476 2540 289576
rect 1033 289475 1135 289476
rect 1033 246576 1135 246577
rect 2440 246576 2540 289476
rect 5660 253172 5772 293268
rect 8387 261321 8457 376032
rect 8381 261320 8463 261321
rect 8381 261250 8382 261320
rect 8462 261250 8463 261320
rect 8381 261249 8463 261250
rect 5660 253062 5661 253172
rect 5771 253062 5772 253172
rect 5660 253061 5772 253062
rect 1033 246476 1034 246576
rect 1134 246476 2540 246576
rect 1033 246475 1135 246476
rect 2440 178862 2540 246476
rect 9016 191343 9126 376032
rect 10674 191538 10784 376032
rect 24558 260523 24678 260524
rect 24558 260405 24559 260523
rect 24677 260405 24678 260523
rect 19138 253335 19258 254086
rect 19138 253217 19139 253335
rect 19257 253217 19258 253335
rect 19138 247349 19258 253217
rect 21326 253341 21446 253342
rect 21326 253223 21327 253341
rect 21445 253223 21446 253341
rect 21326 247553 21446 253223
rect 21325 247552 21447 247553
rect 21325 247432 21326 247552
rect 21446 247432 21447 247552
rect 21325 247431 21447 247432
rect 19137 247348 19259 247349
rect 19137 247228 19138 247348
rect 19258 247228 19259 247348
rect 19137 247227 19259 247228
rect 24558 245563 24678 260405
rect 27250 258973 27370 258974
rect 27250 258855 27251 258973
rect 27369 258855 27370 258973
rect 24557 245562 24679 245563
rect 24557 245442 24558 245562
rect 24678 245442 24679 245562
rect 24557 245441 24679 245442
rect 27250 244827 27370 258855
rect 27249 244826 27371 244827
rect 27249 244706 27250 244826
rect 27370 244706 27371 244826
rect 27249 244705 27371 244706
rect 10673 191537 10785 191538
rect 10673 191427 10674 191537
rect 10784 191427 10785 191537
rect 10673 191426 10785 191427
rect 9010 191342 9132 191343
rect 9010 191232 9011 191342
rect 9131 191232 9132 191342
rect 9010 191231 9132 191232
rect 4379 181780 4624 184240
rect 2440 178762 4664 178862
rect 1919 164695 3090 178276
rect 2175 163346 3090 164695
rect 4564 160876 4664 178762
rect 2622 160776 4664 160876
rect 1033 118976 1135 118977
rect 2622 118976 2722 160776
rect 490227 145105 493561 661830
rect 540833 644584 540835 644585
rect 540834 639784 540835 644584
rect 540833 639783 540835 639784
rect 541567 634584 541569 634585
rect 541568 629784 541569 634584
rect 541567 629783 541569 629784
rect 577935 625014 578045 625015
rect 577935 624906 577936 625014
rect 578044 624906 578045 625014
rect 508868 559006 533522 559030
rect 508868 557261 528746 559006
rect 508868 556624 509895 557261
rect 510532 556624 528746 557261
rect 508868 554254 528746 556624
rect 533498 554254 533522 559006
rect 508868 554230 533522 554254
rect 577935 539255 578045 624906
rect 577935 539145 582651 539255
rect 511640 473922 537996 473946
rect 511640 469170 533220 473922
rect 537972 469170 537996 473922
rect 511640 469146 537996 469170
rect 507116 457972 534522 457996
rect 507116 453220 507140 457972
rect 511892 453220 534522 457972
rect 507116 453196 534522 453220
rect 582541 364996 582651 539145
rect 582436 364886 582756 364996
rect 582436 364786 582546 364886
rect 582646 364786 582756 364886
rect 582436 364676 582756 364786
rect 582541 319756 582651 364676
rect 582436 319646 582756 319756
rect 582436 319546 582546 319646
rect 582646 319546 582756 319646
rect 582436 319436 582756 319546
rect 582541 275356 582651 319436
rect 582436 275246 582756 275356
rect 582436 275146 582546 275246
rect 582646 275146 582756 275246
rect 582436 275036 582756 275146
rect 580888 242005 581188 245316
rect 582541 242005 582651 275036
rect 580888 241895 582651 242005
rect 552812 196966 579468 198242
rect 552812 191768 554140 196966
rect 578296 191768 579468 196966
rect 552812 190928 579468 191768
rect 551320 186340 579660 187154
rect 551320 181150 553050 186340
rect 576862 181150 579660 186340
rect 551320 180540 579660 181150
rect 552718 164209 558786 164626
rect 552718 159411 553277 164209
rect 558075 159411 558786 164209
rect 552718 158880 558786 159411
rect 580888 159120 581188 241895
rect 582541 241680 582651 241895
rect 580888 158290 581422 159120
rect 462379 141771 493561 145105
rect 499374 141266 500790 141267
rect 494841 141242 499375 141266
rect 494841 139876 495525 141242
rect 496891 139876 499375 141242
rect 494841 139852 499375 139876
rect 500789 141265 507515 141266
rect 500789 139853 503116 141265
rect 504528 140997 507515 141265
rect 504528 140121 505628 140997
rect 506504 140121 507515 140997
rect 504528 139853 507515 140121
rect 500789 139852 507515 139853
rect 499374 139851 500790 139852
rect 459182 134644 459867 134700
rect 453395 134620 461504 134644
rect 453395 134348 453419 134620
rect 453691 134348 461504 134620
rect 453395 134324 461504 134348
rect 144646 129153 145734 129154
rect 144646 128067 144647 129153
rect 145733 128067 145734 129153
rect 144646 128066 145734 128067
rect 459182 127150 459867 134324
rect 581122 132708 581422 158290
rect 582515 132708 582625 134578
rect 581122 132408 582720 132708
rect 463530 127150 464217 127151
rect 459182 126465 463531 127150
rect 464216 126465 557323 127150
rect 463530 126464 464217 126465
rect 1033 118876 1034 118976
rect 1134 118876 2722 118976
rect 1033 118875 1135 118876
rect 1033 75776 1135 75777
rect 2622 75776 2722 118876
rect 1033 75676 1034 75776
rect 1134 75676 2722 75776
rect 1033 75675 1135 75676
rect 1033 32376 1135 32377
rect 2622 32376 2722 75676
rect 1033 32276 1034 32376
rect 1134 32276 2722 32376
rect 1033 32275 1135 32276
rect 1033 10976 1135 10977
rect 2622 10976 2722 32276
rect 1033 10876 1034 10976
rect 1134 10876 2722 10976
rect 1033 10875 1135 10876
rect 2622 7266 2722 10876
rect 582420 95356 582720 132408
rect 582420 95246 582756 95356
rect 582420 95146 582546 95246
rect 582646 95146 582756 95246
rect 582420 95036 582756 95146
rect 2324 6966 2866 7266
rect 353 4020 467 4021
rect 353 3908 354 4020
rect 466 3908 467 4020
rect 353 3907 467 3908
rect 2324 3730 2624 6966
rect 582420 3730 582720 95036
rect 2324 3430 582720 3730
<< via4 >>
rect 229597 697552 231180 699708
rect 329614 698285 334006 701834
rect 329614 697442 331192 698285
rect 331192 697442 332128 698285
rect 332128 697442 334006 698285
rect 303894 596286 304214 596606
rect 303918 592534 304190 592806
rect 292338 591606 292610 591878
rect 338088 586140 338408 586460
rect 308982 556600 309667 557285
rect 288563 473351 289093 473352
rect 288563 472811 288564 473351
rect 288564 472811 289093 473351
rect 288563 472810 289093 472811
rect 297407 471950 297777 471951
rect 297407 471570 297776 471950
rect 297776 471570 297777 471950
rect 297407 471569 297777 471570
rect 290884 469717 291524 469718
rect 290884 469067 291523 469717
rect 291523 469067 291524 469717
rect 334724 469170 339476 473922
rect 290884 469066 291524 469067
rect 149126 436938 149398 437210
rect 149126 436194 149398 436466
rect 7012 243720 7332 243835
rect 7012 243630 7127 243720
rect 7127 243630 7217 243720
rect 7217 243630 7332 243720
rect 7012 243515 7332 243630
rect 536033 644584 540833 644585
rect 536033 639784 536034 644584
rect 536034 639784 540833 644584
rect 536033 639783 540833 639784
rect 536767 634584 541567 634585
rect 536767 629784 536768 634584
rect 536768 629784 541567 634584
rect 536767 629783 541567 629784
rect 504068 554230 508868 559030
rect 509895 556624 510532 557261
rect 528746 554254 533498 559006
rect 506840 469146 511640 473946
rect 533220 469170 537972 473922
rect 507140 453220 511892 457972
rect 534522 453196 539322 457996
rect 554140 191768 578296 196966
rect 553050 181150 576862 186340
rect 553300 159434 558052 164186
rect 495525 139876 496891 141242
rect 507515 139852 510119 141266
rect 453419 134348 453691 134620
rect 557323 126465 558008 127150
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 229160 699708 231660 702300
rect 229160 697552 229597 699708
rect 231180 697552 231660 699708
rect 229160 697490 231660 697552
rect 329590 701834 334230 702300
rect 329590 697442 329614 701834
rect 334006 700360 334230 701834
rect 334006 697442 334030 700360
rect 329590 697418 334030 697442
rect 7012 422228 7332 672796
rect 518241 644584 520957 646724
rect 536009 644585 540857 644609
rect 536009 644584 536033 644585
rect 518241 639784 536033 644584
rect 518241 634584 520957 639784
rect 536009 639783 536033 639784
rect 540833 639783 540857 644585
rect 536009 639759 540857 639783
rect 536743 634585 541591 634609
rect 536743 634584 536767 634585
rect 518241 629784 536767 634584
rect 303870 596606 304238 596630
rect 303870 596286 303894 596606
rect 304214 596286 340720 596606
rect 303870 596262 304238 596286
rect 304812 594242 307352 594562
rect 303894 592806 304214 592830
rect 303894 592534 303918 592806
rect 304190 592534 304214 592806
rect 303894 592510 304214 592534
rect 292314 591878 292634 591902
rect 292314 591606 292338 591878
rect 292610 591606 292634 591878
rect 292314 591582 292634 591606
rect 337754 588588 340470 596286
rect 518241 588588 520957 629784
rect 536743 629783 536767 629784
rect 541567 629783 541591 634585
rect 536743 629759 541591 629783
rect 337754 586460 520957 588588
rect 337754 586140 338088 586460
rect 338408 586140 520957 586460
rect 337754 585872 520957 586140
rect 290594 559030 290914 582110
rect 304924 559030 305244 580778
rect 504044 559030 508892 559054
rect 283960 557285 504068 559030
rect 283960 556600 308982 557285
rect 309667 556600 504068 557285
rect 283960 554230 504068 556600
rect 508868 557285 508892 559030
rect 508868 557261 510556 557285
rect 508868 556624 509895 557261
rect 510532 556624 510556 557261
rect 508868 556600 510556 556624
rect 508868 554230 508892 556600
rect 504044 554206 508892 554230
rect 518241 489282 520957 585872
rect 528722 559006 552198 559030
rect 528722 554254 528746 559006
rect 533498 554254 558076 559006
rect 528722 554230 558076 554254
rect 284208 486566 520957 489282
rect 284208 473346 286924 486566
rect 506816 473946 511664 473970
rect 296978 473922 506840 473946
rect 288539 473352 289117 473376
rect 288539 473346 288563 473352
rect 284208 472816 288563 473346
rect 284208 471752 286924 472816
rect 288539 472810 288563 472816
rect 289093 472810 289117 473352
rect 288539 472786 289117 472810
rect 296978 471951 334724 473922
rect 296978 471569 297407 471951
rect 297777 471569 334724 471951
rect 290860 469718 291548 469742
rect 290860 469066 290884 469718
rect 291524 469712 291548 469718
rect 296978 469712 334724 471569
rect 291524 469170 334724 469712
rect 339476 469170 506840 473922
rect 291524 469146 506840 469170
rect 511640 469146 511664 473946
rect 291524 469072 302376 469146
rect 506816 469122 511664 469146
rect 291524 469066 291548 469072
rect 290860 469042 291548 469066
rect 96586 457972 511916 457996
rect 96586 453220 507140 457972
rect 511892 453220 511916 457972
rect 96586 453196 511916 453220
rect 7012 379054 7332 419818
rect 7012 243859 7332 376032
rect 6988 243835 7356 243859
rect 6988 243515 7012 243835
rect 7332 243515 7356 243835
rect 6988 243491 7356 243515
rect 96586 92376 101386 453196
rect 518241 446868 520957 486566
rect 553276 473946 558076 554230
rect 533196 473922 558076 473946
rect 533196 469170 533220 473922
rect 537972 469170 558076 473922
rect 533196 469146 558076 469170
rect 534498 457996 539346 458020
rect 553276 457996 558076 469146
rect 534498 453196 534522 457996
rect 539322 453196 558076 457996
rect 534498 453172 539346 453196
rect 118982 444152 520957 446868
rect 118982 109188 121698 444152
rect 518241 437454 520957 444152
rect 149102 437210 149422 437234
rect 149102 436938 149126 437210
rect 149398 436938 149422 437210
rect 454905 437134 520957 437454
rect 149102 436466 149422 436938
rect 149102 436194 149126 436466
rect 149398 436194 149422 436466
rect 149102 434728 149422 436194
rect 149102 434408 149964 434728
rect 518241 427454 520957 437134
rect 454905 427134 520957 427454
rect 518241 417454 520957 427134
rect 454905 417134 520957 417454
rect 518241 407454 520957 417134
rect 454905 407134 520957 407454
rect 518241 397454 520957 407134
rect 454905 397134 520957 397454
rect 518241 387454 520957 397134
rect 454905 387134 520957 387454
rect 518241 377454 520957 387134
rect 454905 377134 520957 377454
rect 518241 367454 520957 377134
rect 454905 367134 520957 367454
rect 518241 357454 520957 367134
rect 454905 357134 520957 357454
rect 518241 347454 520957 357134
rect 454905 347134 520957 347454
rect 518241 337454 520957 347134
rect 454905 337134 520957 337454
rect 518241 327454 520957 337134
rect 454905 327134 520957 327454
rect 518241 317454 520957 327134
rect 454905 317134 520957 317454
rect 518241 307454 520957 317134
rect 454905 307134 520957 307454
rect 518241 297454 520957 307134
rect 454905 297134 520957 297454
rect 518241 287454 520957 297134
rect 454905 287134 520957 287454
rect 518241 277454 520957 287134
rect 454905 277134 520957 277454
rect 518241 267454 520957 277134
rect 454905 267134 520957 267454
rect 518241 257454 520957 267134
rect 454905 257134 520957 257454
rect 518241 247454 520957 257134
rect 454905 247134 520957 247454
rect 518241 237454 520957 247134
rect 454905 237134 520957 237454
rect 518241 227454 520957 237134
rect 454905 227134 520957 227454
rect 518241 217454 520957 227134
rect 454905 217134 520957 217454
rect 518241 207454 520957 217134
rect 454905 207134 520957 207454
rect 518241 197454 520957 207134
rect 553276 198242 558076 453196
rect 454905 197134 520957 197454
rect 518241 187454 520957 197134
rect 552812 196966 579468 198242
rect 552812 191768 554140 196966
rect 578296 191768 579468 196966
rect 552812 190928 579468 191768
rect 454905 187134 520957 187454
rect 553276 187154 558076 190928
rect 518241 177454 520957 187134
rect 551320 186340 579660 187154
rect 551320 181150 553050 186340
rect 576862 181150 579660 186340
rect 551320 180540 579660 181150
rect 454905 177134 520957 177454
rect 518241 167454 520957 177134
rect 553276 167476 558076 180540
rect 454905 167134 520957 167454
rect 518241 157454 520957 167134
rect 550944 164186 571790 167476
rect 550944 162676 553300 164186
rect 454905 157134 520957 157454
rect 518241 147454 520957 157134
rect 454905 147134 520957 147454
rect 518241 141320 520957 147134
rect 494530 141266 520957 141320
rect 494530 141242 507515 141266
rect 494530 139876 495525 141242
rect 496891 139876 507515 141242
rect 494530 139852 507515 139876
rect 510119 139852 520957 141266
rect 494530 139799 520957 139852
rect 453395 134620 453715 134644
rect 453395 134348 453419 134620
rect 453691 134348 453715 134620
rect 453395 134324 453715 134348
rect 518241 109188 520957 139799
rect 553276 159434 553300 162676
rect 558052 162676 571790 164186
rect 558052 159434 558076 162676
rect 553276 127150 558076 159434
rect 553276 126465 557323 127150
rect 558008 126465 558076 127150
rect 118982 106472 525544 109188
rect 553276 92376 558076 126465
rect 96586 87576 558076 92376
use array_SR  array_SR_0
timestamp 1758153220
transform 1 0 149469 0 1 114190
box -21072 586 308046 327366
use bias  bias_1
timestamp 1758153220
transform 1 0 289348 0 1 473566
box 790 -2236 7180 -220
use opamp_wrapper  opamp_wrapper_0
timestamp 1758069660
transform 1 0 464481 0 1 129134
box -2280 -2669 27441 13665
use opamp_wrapper  opamp_wrapper_1
timestamp 1758069660
transform 1 0 309932 0 1 580259
box -2280 -2669 27441 13665
use pixel_array  pixel_array_0
timestamp 1758143320
transform 1 0 294314 0 1 588742
box -3720 -8600 11230 5820
use sky130_fd_pr__res_generic_m3_3NNQKJ  sky130_fd_pr__res_generic_m3_3NNQKJ_0
timestamp 1758069660
transform 0 1 582837 -1 0 364836
box -50 -107 50 107
use sky130_fd_pr__res_generic_m3_3NNQKJ  sky130_fd_pr__res_generic_m3_3NNQKJ_1
timestamp 1758069660
transform 0 1 767 -1 0 462426
box -50 -107 50 107
<< labels >>
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
