magic
tech sky130A
timestamp 1758224069
<< metal5 >>
rect 19600 27800 20800 28000
rect 21400 27800 22600 28000
rect 41800 27800 42700 28000
rect 19600 27200 20900 27800
rect 21400 27200 22700 27800
rect 41800 27500 42800 27800
rect 19700 27000 20800 27200
rect 21400 27000 22600 27200
rect 41800 27000 43000 27500
rect 43800 27200 45200 28000
rect 43900 27000 45200 27200
rect 46900 27000 47500 28800
rect 19900 24600 20300 27000
rect 21800 24600 22300 27000
rect 42200 26400 43100 27000
rect 24400 25900 25200 26200
rect 29300 25900 29600 26200
rect 33000 25900 33400 26200
rect 42200 25900 43200 26400
rect 23900 25700 25400 25900
rect 27400 25700 28300 25900
rect 28900 25700 30000 25900
rect 31100 25700 32000 25900
rect 32600 25700 33700 25900
rect 23600 25400 25700 25700
rect 23600 25100 25800 25400
rect 27200 25100 28300 25700
rect 28800 25400 30100 25700
rect 28600 25100 30200 25400
rect 31000 25100 32000 25700
rect 32500 25400 33800 25700
rect 32300 25100 34000 25400
rect 23600 24900 24400 25100
rect 25100 24900 25800 25100
rect 27400 24900 28300 25100
rect 28460 24900 29340 25100
rect 29500 24900 30200 25100
rect 31100 24900 32000 25100
rect 32200 24900 33100 25100
rect 33260 24900 34000 25100
rect 34600 25100 35800 25900
rect 36600 25100 37800 25900
rect 34600 24900 35600 25100
rect 36700 24900 37800 25100
rect 42200 25700 43300 25900
rect 42200 24940 42640 25700
rect 42800 25100 43400 25700
rect 23600 24600 23900 24900
rect 25300 24600 25900 24900
rect 19900 23600 22300 24600
rect 24500 23600 25200 23800
rect 25400 23600 25900 24600
rect 19900 20700 20300 23600
rect 21800 20700 22300 23600
rect 23900 23300 25900 23600
rect 23600 23100 25900 23300
rect 23500 22800 25900 23100
rect 23400 22500 24400 22800
rect 25200 22500 25900 22800
rect 23400 22300 24100 22500
rect 23300 22000 23900 22300
rect 23300 21200 23800 22000
rect 25400 21500 25900 22500
rect 25200 21200 25900 21500
rect 23300 21000 23900 21200
rect 25100 21000 25900 21200
rect 23400 20700 24000 21000
rect 24800 20700 25900 21000
rect 28000 24600 29200 24900
rect 29800 24600 30100 24900
rect 31700 24600 32900 24900
rect 33500 24600 33800 24900
rect 34800 24600 35400 24900
rect 28000 24400 28900 24600
rect 31700 24400 32600 24600
rect 34900 24400 35400 24600
rect 37000 24600 37600 24900
rect 37000 24400 37400 24600
rect 28000 24100 28800 24400
rect 31700 24100 32500 24400
rect 34900 24100 35500 24400
rect 28000 23800 28700 24100
rect 31700 23800 32400 24100
rect 35000 23800 35500 24100
rect 36800 24100 37400 24400
rect 36800 23800 37300 24100
rect 28000 23600 28600 23800
rect 31700 23600 32300 23800
rect 35000 23600 35600 23800
rect 28000 20700 28300 23600
rect 31700 20700 32000 23600
rect 35200 23300 35600 23600
rect 36700 23600 37300 23800
rect 36700 23300 37200 23600
rect 35200 23100 35800 23300
rect 35300 22800 35800 23100
rect 36600 23100 37200 23300
rect 36600 22800 37100 23100
rect 35300 22500 35900 22800
rect 35400 22300 35900 22500
rect 36500 22500 37100 22800
rect 36500 22300 37000 22500
rect 35400 22000 36000 22300
rect 35500 21800 36000 22000
rect 36400 22000 37000 22300
rect 36400 21800 36800 22000
rect 35500 21500 36100 21800
rect 35600 21200 36100 21500
rect 36260 21500 36800 21800
rect 36260 21200 36700 21500
rect 35600 21000 36700 21200
rect 19400 20400 20800 20700
rect 21400 20400 22700 20700
rect 23400 20400 26400 20700
rect 19400 19900 20900 20400
rect 21400 19900 22800 20400
rect 23500 20200 26400 20400
rect 23600 19900 25300 20200
rect 25460 19900 26400 20200
rect 27100 19900 29600 20700
rect 30800 19900 33400 20700
rect 35800 20400 36600 21000
rect 42200 20700 42700 24940
rect 43000 24900 43600 25100
rect 43100 24600 43600 24900
rect 43100 24400 43700 24600
rect 43200 23800 43800 24400
rect 43300 23600 43900 23800
rect 43400 23300 43900 23600
rect 43400 23100 44000 23300
rect 43600 22500 44200 23100
rect 43700 22300 44240 22500
rect 43800 22000 44240 22300
rect 44400 22000 44900 27000
rect 46200 24900 47500 25900
rect 43800 21800 44900 22000
rect 43900 21200 44900 21800
rect 44000 20700 44900 21200
rect 47000 20700 47500 24900
rect 35900 20200 36600 20400
rect 23800 19700 25000 19900
rect 35900 19700 36500 20200
rect 41900 19900 43300 20700
rect 44200 20400 44900 20700
rect 44300 19900 44900 20400
rect 46000 19900 48700 20700
rect 35800 19100 36400 19700
rect 35600 18600 36200 19100
rect 35600 18400 36100 18600
rect 35500 18100 36100 18400
rect 34600 17800 36500 18100
rect 34600 17600 36600 17800
rect 34600 17300 36500 17600
rect 10100 13900 12100 14200
rect 10000 13700 12500 13900
rect 10000 13400 12700 13700
rect 10100 13100 12800 13400
rect 26300 13100 26900 15000
rect 45100 14700 45600 15000
rect 52700 14700 53200 15000
rect 56400 14700 56900 15000
rect 44600 14400 46000 14700
rect 48100 14400 50200 14700
rect 52300 14400 53500 14700
rect 56000 14400 57200 14700
rect 42700 14200 42920 14220
rect 44500 14200 46200 14400
rect 37300 13900 38600 14200
rect 37100 13700 38840 13900
rect 39000 13700 39400 14200
rect 41000 13900 42400 14200
rect 42700 14060 43100 14200
rect 42760 13900 43100 14060
rect 44400 13900 46300 14200
rect 48100 13900 50300 14400
rect 52200 14200 53600 14400
rect 55900 14200 57500 14400
rect 52100 13900 53800 14200
rect 55800 13900 57600 14200
rect 40800 13700 42600 13900
rect 42760 13700 43200 13900
rect 44300 13700 45100 13900
rect 45600 13700 46400 13900
rect 37000 13400 39400 13700
rect 40700 13400 43200 13700
rect 36800 13100 37800 13400
rect 38200 13100 39400 13400
rect 40600 13100 41500 13400
rect 41900 13100 43200 13400
rect 44200 13400 44900 13700
rect 45800 13400 46400 13700
rect 48100 13700 50200 13900
rect 52000 13700 52700 13900
rect 53000 13700 53900 13900
rect 55800 13700 56500 13900
rect 56900 13700 57700 13900
rect 44200 13100 44800 13400
rect 46000 13100 46600 13400
rect 10600 10300 10900 13100
rect 12100 12900 12800 13100
rect 36700 12900 37400 13100
rect 38500 12900 39400 13100
rect 12200 12600 13000 12900
rect 12500 12400 13000 12600
rect 36600 12600 37300 12900
rect 38600 12600 39400 12900
rect 40400 12900 41300 13100
rect 42200 12900 43200 13100
rect 40400 12600 41000 12900
rect 42500 12600 43200 12900
rect 36600 12400 37200 12600
rect 38800 12400 39400 12600
rect 40300 12400 40900 12600
rect 12500 12100 13100 12400
rect 15000 12100 15800 12400
rect 18800 12100 19600 12400
rect 22700 12100 23500 12400
rect 30200 12100 31000 12400
rect 12600 11600 13100 12100
rect 14600 11800 16200 12100
rect 18500 11800 19900 12100
rect 20060 11800 20400 12100
rect 14400 11600 16300 11800
rect 18200 11600 20400 11800
rect 12500 11300 13100 11600
rect 14300 11300 16600 11600
rect 18100 11300 20400 11600
rect 21100 11600 22100 12100
rect 22300 11800 23800 12100
rect 22260 11600 24000 11800
rect 21100 11300 24100 11600
rect 25600 11300 26900 12100
rect 12500 11100 13000 11300
rect 12400 10800 13000 11100
rect 14200 11100 15100 11300
rect 15700 11100 16700 11300
rect 14200 10800 14900 11100
rect 16000 10800 16700 11100
rect 18000 11100 18800 11300
rect 19600 11100 20400 11300
rect 21200 11100 22800 11300
rect 23400 11100 24200 11300
rect 25700 11100 26900 11300
rect 28900 11800 29600 12100
rect 29900 11800 31200 12100
rect 36500 11800 37100 12400
rect 38900 11800 39400 12400
rect 28900 11300 31400 11800
rect 36400 11600 37000 11800
rect 39000 11600 39400 11800
rect 40200 11800 40800 12400
rect 42600 12100 43200 12600
rect 44000 12900 44600 13100
rect 44000 12400 44500 12900
rect 44200 12100 44400 12400
rect 28900 11100 30200 11300
rect 30800 11100 31600 11300
rect 18000 10800 18600 11100
rect 19800 10800 20400 11100
rect 12100 10500 13000 10800
rect 11500 10300 12800 10500
rect 14000 10300 14600 10800
rect 16200 10300 16800 10800
rect 18000 10300 18500 10800
rect 19900 10300 20400 10800
rect 10600 10000 12700 10300
rect 13900 10000 14500 10300
rect 16300 10000 16900 10300
rect 18000 10000 18600 10300
rect 20000 10000 20400 10300
rect 21600 10800 22600 11100
rect 23600 10800 24400 11100
rect 21600 10500 22400 10800
rect 23800 10500 24400 10800
rect 21600 10300 22300 10500
rect 23900 10300 24500 10500
rect 21600 10000 22200 10300
rect 10600 9800 12500 10000
rect 13900 9800 14400 10000
rect 16400 9800 16900 10000
rect 10600 9500 12400 9800
rect 10600 6900 10900 9500
rect 11600 9200 12500 9500
rect 11900 9000 12600 9200
rect 12000 8700 12700 9000
rect 13900 8700 16900 9800
rect 18100 9800 19000 10000
rect 18100 9500 19800 9800
rect 18200 9200 20000 9500
rect 18500 9000 20300 9200
rect 19100 8700 20400 9000
rect 12100 8400 12800 8700
rect 12200 8200 12800 8400
rect 13900 8200 14400 8700
rect 19700 8400 20500 8700
rect 19900 8200 20500 8400
rect 12400 7900 13000 8200
rect 13900 7900 14500 8200
rect 17900 7900 18200 8200
rect 12500 7400 13100 7900
rect 14000 7400 14600 7900
rect 16600 7400 16800 7700
rect 17900 7400 18400 7900
rect 20000 7400 20500 8200
rect 12600 6900 13200 7400
rect 14200 7100 14900 7400
rect 16400 7100 16900 7400
rect 14200 6900 15000 7100
rect 16100 6900 16900 7100
rect 10100 6600 11500 6900
rect 12700 6600 13600 6900
rect 14300 6600 16900 6900
rect 17900 7100 18500 7400
rect 19900 7100 20500 7400
rect 17900 6900 18600 7100
rect 19800 6900 20500 7100
rect 21600 8400 22100 10000
rect 24000 9500 24500 10300
rect 24100 9200 24500 9500
rect 24100 9000 24600 9200
rect 21600 8200 22200 8400
rect 24000 8200 24500 9000
rect 21600 7700 22300 8200
rect 23900 7900 24500 8200
rect 23800 7700 24400 7900
rect 21600 7400 22600 7700
rect 23600 7400 24400 7700
rect 21600 7100 22700 7400
rect 23400 7100 24200 7400
rect 21600 6900 24100 7100
rect 26500 6900 26900 11100
rect 29300 10800 30100 11100
rect 31000 10800 31600 11100
rect 29300 10500 30000 10800
rect 31100 10500 31700 10800
rect 29300 10300 29900 10500
rect 29300 6900 29800 10300
rect 31200 6900 31700 10500
rect 32800 9500 35600 10500
rect 36400 8700 36800 11600
rect 39100 11300 39260 11600
rect 40200 11300 40700 11800
rect 42700 11600 43200 12100
rect 46100 11600 46600 13100
rect 42800 11300 43100 11600
rect 46000 11300 46600 11600
rect 48100 11600 48600 13700
rect 51800 13400 52600 13700
rect 53300 13400 53900 13700
rect 55700 13400 56300 13700
rect 57100 13400 57700 13700
rect 51800 13100 52400 13400
rect 53400 13100 54000 13400
rect 55700 13100 56200 13400
rect 57200 13100 57800 13400
rect 51700 12600 52300 13100
rect 53500 12900 54000 13100
rect 55600 12900 56200 13100
rect 57400 12900 57800 13100
rect 51700 12100 52200 12600
rect 53500 12400 54100 12900
rect 51600 11800 52200 12100
rect 48800 11600 49700 11800
rect 48100 11300 49900 11600
rect 40100 8700 40600 11300
rect 45800 11100 46400 11300
rect 45700 10800 46400 11100
rect 48100 11100 50000 11300
rect 48100 10800 50200 11100
rect 45600 10500 46300 10800
rect 48100 10500 48800 10800
rect 49600 10500 50300 10800
rect 45500 10300 46200 10500
rect 48100 10300 48600 10500
rect 49700 10300 50400 10500
rect 45400 10000 46100 10300
rect 49800 10000 50400 10300
rect 45200 9800 46000 10000
rect 49900 9800 50400 10000
rect 45100 9500 45800 9800
rect 50000 9500 50400 9800
rect 45000 9200 45700 9500
rect 44900 9000 45600 9200
rect 44800 8700 45500 9000
rect 36400 8400 37000 8700
rect 36500 8200 37000 8400
rect 40200 8200 40700 8700
rect 44600 8400 45400 8700
rect 44500 8200 45200 8400
rect 50000 8200 50500 9500
rect 51600 8700 52100 11800
rect 53600 11600 54100 12400
rect 53800 9500 54100 11600
rect 55600 11100 56000 12900
rect 57400 12600 58000 12900
rect 57500 11800 58000 12600
rect 57500 11600 58100 11800
rect 57400 11100 58100 11600
rect 55600 10800 56200 11100
rect 57200 10800 58100 11100
rect 55700 10500 56300 10800
rect 57100 10500 58100 10800
rect 55700 10300 56400 10500
rect 57000 10300 58100 10500
rect 55800 10000 58100 10300
rect 55800 9800 57500 10000
rect 56000 9500 57400 9800
rect 57660 9640 58100 10000
rect 36500 7900 37100 8200
rect 39100 7900 39500 8200
rect 40200 7900 40800 8200
rect 43000 7900 43200 8200
rect 44400 7900 45100 8200
rect 36500 7700 37200 7900
rect 39000 7700 39500 7900
rect 36600 7400 37200 7700
rect 38900 7400 39500 7700
rect 40300 7700 40900 7900
rect 42700 7700 43200 7900
rect 44300 7700 45000 7900
rect 49900 7700 50400 8200
rect 51700 7900 52200 8700
rect 53600 8200 54100 9500
rect 56200 9200 57100 9500
rect 57600 9200 58100 9640
rect 57500 9000 58100 9200
rect 57500 8400 58000 9000
rect 57400 8200 58000 8400
rect 51700 7700 52300 7900
rect 53500 7700 54100 8200
rect 57200 7900 57800 8200
rect 57100 7700 57800 7900
rect 40300 7400 41000 7700
rect 42600 7400 43200 7700
rect 44200 7400 44900 7700
rect 47800 7400 48200 7700
rect 49800 7400 50400 7700
rect 51800 7400 52300 7700
rect 36700 7100 37400 7400
rect 38800 7100 39500 7400
rect 40400 7100 41200 7400
rect 42500 7100 43200 7400
rect 44000 7100 44800 7400
rect 46200 7100 46600 7400
rect 47800 7100 48500 7400
rect 49700 7100 50300 7400
rect 51800 7100 52400 7400
rect 53400 7100 54000 7700
rect 57000 7400 57700 7700
rect 56900 7100 57600 7400
rect 36800 6900 37600 7100
rect 38500 6900 39400 7100
rect 40600 6900 41400 7100
rect 42400 6900 43100 7100
rect 43900 6900 44600 7100
rect 46200 6900 46700 7100
rect 47800 6900 48600 7100
rect 49400 6900 50300 7100
rect 52000 6900 52600 7100
rect 53300 6900 53900 7100
rect 56600 6900 57600 7100
rect 17900 6600 19200 6900
rect 19360 6600 20400 6900
rect 10000 6400 11600 6600
rect 10100 6100 11600 6400
rect 12800 6100 13700 6600
rect 14400 6400 16800 6600
rect 17900 6400 20300 6600
rect 21600 6440 22040 6900
rect 22200 6600 24000 6900
rect 14600 6100 16600 6400
rect 17900 6100 20200 6400
rect 14900 5800 16200 6100
rect 18600 5800 19900 6100
rect 21600 4300 22100 6440
rect 22300 6400 23900 6600
rect 22600 6100 23500 6400
rect 25300 6100 28100 6900
rect 28800 6100 30100 6900
rect 30800 6100 32000 6900
rect 37000 6600 38000 6900
rect 38200 6600 39200 6900
rect 40700 6600 41800 6900
rect 41960 6600 43000 6900
rect 37100 6400 39100 6600
rect 40800 6400 42800 6600
rect 37200 6100 38900 6400
rect 40900 6100 42700 6400
rect 43900 6100 46700 6900
rect 47900 6600 50200 6900
rect 52000 6600 53800 6900
rect 48000 6400 50000 6600
rect 52100 6400 53800 6600
rect 55600 6600 57400 6900
rect 55600 6400 57200 6600
rect 48200 6100 49900 6400
rect 52200 6100 53500 6400
rect 55600 6100 57000 6400
rect 37400 5800 38600 6100
rect 41200 5800 42500 6100
rect 48500 5800 49700 6100
rect 52400 5800 53400 6100
rect 55700 5800 56800 6100
rect 21100 3500 22800 4300
<< properties >>
string GDS_END 2458154
string GDS_FILE /home/hni/TopmetalSe-Respin/mag/text.gds
string GDS_START 102
<< end >>
