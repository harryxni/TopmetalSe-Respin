* NGSPICE file created from pixel_array_fill.ext - technology: sky130A

.subckt pixel_fill gring VDD GND VREF ROW_SEL NB1 VBIAS NB2 AMP_IN SF_IB PIX_OUT CSA_VREF
X0 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5 pd=7.5 as=24.809025 ps=56.34 w=2 l=1.44
X1 a_4120_n520# VBIAS a_4120_n750# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.995 ps=8.8 w=1 l=0.8
X2 a_5720_n730# a_4600_n810# GND VDD sky130_fd_pr__pfet_01v8_lvt ad=0.25 pd=1.5 as=0.35 ps=2.7 w=1 l=1
X3 a_4330_n30# a_3852_n32# a_3852_n32# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.23 pd=1.65 as=0.3927 ps=2.8 w=1 l=2
X4 VDD SF_IB a_5720_n730# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.25 ps=1.5 w=1 l=1
X5 a_5460_10# a_4330_n30# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X6 a_3852_n32# VBIAS a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.76 ps=8.8 w=1 l=0.8
X7 VDD a_4120_n520# a_4600_n810# GND sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=1
X8 a_4120_n750# AMP_IN a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=1.995 pd=8.8 as=1.4 ps=7.4 w=7 l=0.15
X9 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.119375 pd=7.15 as=0 ps=0 w=2 l=3.35
X10 a_4120_n520# a_3852_n32# a_5460_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X11 AMP_IN a_4600_n810# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 GND NB1 a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0.42 pd=3.1 as=0.42 ps=3.1 w=1.2 l=1
X13 a_5750_n920# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=0.6 pd=2.95 as=5.4 ps=9.4 w=2 l=1
X14 a_4050_n2590# VREF a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=1.4 pd=7.4 as=1.76 ps=8.8 w=7 l=0.15
X15 a_4600_n810# NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1.15
X16 VDD a_4330_n30# a_4330_n30# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.23 ps=1.65 w=1 l=2
X17 VDD a_5720_n730# a_5750_n920# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.6 ps=2.95 w=1 l=0.15
X18 AMP_IN CSA_VREF a_4600_n810# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.294 pd=2.24 as=0.273 ps=2.14 w=0.42 l=8
X19 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=10.715 pd=15.9 as=0 ps=0 w=2.6 l=0.35
.ends

.subckt pixel_array_fill VBIAS VREF NB2 VDD SF_IB CSA_VREF NB1 ROW_SEL0 GND ROW_SEL1
+ ROW_SEL2 PIX0_IN GRING PIX1_IN PIX2_IN PIX3_IN PIX4_IN PIX5_IN PIX6_IN PIX_OUT0
+ PIX7_IN PIX_OUT1 PIX8_IN PIX_OUT2 ARRAY_OUT COL_SEL0 COL_SEl1 COL_SEL2
Xpixel_fill_1 GRING VDD GND VREF ROW_SEL0 NB1 VBIAS NB2 PIX1_IN SF_IB PIX_OUT1 CSA_VREF
+ pixel_fill
Xpixel_fill_0 GRING VDD GND VREF ROW_SEL0 NB1 VBIAS NB2 PIX0_IN SF_IB PIX_OUT0 CSA_VREF
+ pixel_fill
Xpixel_fill_2 GRING VDD GND VREF ROW_SEL0 NB1 VBIAS NB2 PIX2_IN SF_IB PIX_OUT2 CSA_VREF
+ pixel_fill
Xpixel_fill_3 GRING VDD GND VREF ROW_SEL1 NB1 VBIAS NB2 PIX3_IN SF_IB PIX_OUT0 CSA_VREF
+ pixel_fill
Xpixel_fill_4 GRING VDD GND VREF ROW_SEL1 NB1 VBIAS NB2 PIX4_IN SF_IB PIX_OUT1 CSA_VREF
+ pixel_fill
Xpixel_fill_5 GRING VDD GND VREF ROW_SEL1 NB1 VBIAS NB2 PIX5_IN SF_IB PIX_OUT2 CSA_VREF
+ pixel_fill
Xpixel_fill_6 GRING VDD GND VREF ROW_SEL2 NB1 VBIAS NB2 PIX6_IN SF_IB PIX_OUT0 CSA_VREF
+ pixel_fill
Xpixel_fill_7 GRING VDD GND VREF ROW_SEL2 NB1 VBIAS NB2 PIX7_IN SF_IB PIX_OUT1 CSA_VREF
+ pixel_fill
Xpixel_fill_8 GRING VDD GND VREF ROW_SEL2 NB1 VBIAS NB2 PIX8_IN SF_IB PIX_OUT2 CSA_VREF
+ pixel_fill
X0 PIX_OUT2 COL_SEL2 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X1 PIX_OUT1 COL_SEl1 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X2 PIX_OUT0 COL_SEL0 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
.ends

