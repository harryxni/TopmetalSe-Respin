magic
tech sky130A
magscale 1 2
timestamp 1758069660
<< metal3 >>
rect -50 50 50 107
rect -50 -107 50 -50
<< rmetal3 >>
rect -50 -50 50 50
<< properties >>
string gencell sky130_fd_pr__res_generic_m3
string library sky130
string parameters w 0.500 l 0.500 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 47.0m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
