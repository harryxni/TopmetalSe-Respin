magic
tech sky130A
timestamp 1758310990
<< metal5 >>
rect 19800 18900 20000 19000
rect 19400 18800 20000 18900
rect 19100 18700 20000 18800
rect 18700 18600 19800 18700
rect 18500 18500 19600 18600
rect 18100 18400 19300 18500
rect 17700 18300 18900 18400
rect 17200 18200 18500 18300
rect 0 18100 400 18200
rect 16800 18100 18100 18200
rect 0 18060 600 18100
rect 0 18000 760 18060
rect 16500 18000 17900 18100
rect 200 17900 1100 18000
rect 16000 17900 17400 18000
rect 600 17800 1600 17900
rect 15500 17800 17000 17900
rect 900 17700 2100 17800
rect 12200 17700 12360 17800
rect 14900 17700 16500 17800
rect 1400 17600 2800 17700
rect 11900 17600 12700 17700
rect 14300 17600 16000 17700
rect 1700 17500 3200 17600
rect 11800 17500 12700 17600
rect 13900 17500 15700 17600
rect 2200 17400 4000 17500
rect 11600 17400 12800 17500
rect 13200 17400 15200 17500
rect 2800 17300 5100 17400
rect 8800 17300 9600 17400
rect 11500 17300 14600 17400
rect 3600 17200 6600 17300
rect 8600 17200 9800 17300
rect 10900 17200 13800 17300
rect 4400 17100 13100 17200
rect 5000 17000 12800 17100
rect 6300 16900 12600 17000
rect 8400 16800 10100 16900
rect 8600 16700 10100 16800
rect 11300 16800 12200 16900
rect 11300 16700 12100 16800
rect 9200 16500 10200 16700
rect 9300 15900 10200 16500
rect 9200 15500 10200 15900
rect 9100 15200 10200 15500
rect 9000 15000 10200 15200
rect 8900 14500 10200 15000
rect 8800 13700 10200 14500
rect 11200 16100 12100 16700
rect 11200 15700 12200 16100
rect 11200 15300 12300 15700
rect 11200 14900 12400 15300
rect 11200 14700 12500 14900
rect 11200 14300 12600 14700
rect 11300 13900 12600 14300
rect 8800 12800 10100 13700
rect 11300 12900 12700 13900
rect 5600 12300 6600 12400
rect 5200 12200 6900 12300
rect 8800 12200 10200 12800
rect 11300 12700 12600 12900
rect 11200 12600 12600 12700
rect 11100 12500 12600 12600
rect 10800 12400 12600 12500
rect 10700 12300 12600 12400
rect 10600 12200 12600 12300
rect 4900 12100 7100 12200
rect 4800 12000 7100 12100
rect 4600 11900 7300 12000
rect 4500 11800 7400 11900
rect 8800 11884 10239 12200
rect 10539 11884 12600 12200
rect 8800 11800 12600 11884
rect 4400 11700 5400 11800
rect 6600 11700 7500 11800
rect 8900 11700 12600 11800
rect 4300 11600 5200 11700
rect 6800 11600 7600 11700
rect 4300 11500 5100 11600
rect 6900 11500 7700 11600
rect 8900 11500 12500 11700
rect 4200 11400 4900 11500
rect 7000 11400 7800 11500
rect 8900 11400 12600 11500
rect 4100 11300 4800 11400
rect 7100 11300 7800 11400
rect 9000 11300 12600 11400
rect 4100 11200 4700 11300
rect 7200 11200 7900 11300
rect 9000 11200 12700 11300
rect 4100 11100 4600 11200
rect 4000 11000 4600 11100
rect 7300 11000 8000 11200
rect 9100 11000 12800 11200
rect 4000 10900 4400 11000
rect 3900 10800 4400 10900
rect 7400 10800 8100 11000
rect 9200 10900 12900 11000
rect 9300 10800 12900 10900
rect 3900 10500 4300 10800
rect 7400 10700 8200 10800
rect 3900 10400 4200 10500
rect 7500 10400 8200 10700
rect 9300 10600 12800 10800
rect 9300 10552 12700 10600
rect 9300 10400 11896 10552
rect 12256 10500 12700 10552
rect 12256 10400 12600 10500
rect 4000 10300 4200 10400
rect 7600 9700 8200 10400
rect 9200 10204 11896 10400
rect 9200 9900 12100 10204
rect 7500 9500 8200 9700
rect 9100 9800 12100 9900
rect 7500 9400 8100 9500
rect 9100 9400 12200 9800
rect 7400 9100 8100 9400
rect 9000 9100 12200 9400
rect 7400 9000 8000 9100
rect 7300 8900 8000 9000
rect 7300 8500 7900 8900
rect 8900 8800 12200 9100
rect 8900 8600 12100 8800
rect 7300 8000 7800 8500
rect 8900 8400 12000 8600
rect 8900 8200 11900 8400
rect 8900 8100 11800 8200
rect 7300 7800 7900 8000
rect 8900 7900 11700 8100
rect 8900 7800 11600 7900
rect 7400 7700 7900 7800
rect 8800 7700 11500 7800
rect 7400 7600 8000 7700
rect 7400 7500 8100 7600
rect 7500 7400 8100 7500
rect 7600 7300 8300 7400
rect 8800 7300 11400 7700
rect 7600 7200 8400 7300
rect 8700 7200 11500 7300
rect 7700 7100 11700 7200
rect 7800 7000 11700 7100
rect 7900 6900 11900 7000
rect 8100 6800 12100 6900
rect 8200 6758 12300 6800
rect 8405 6700 12300 6758
rect 8405 6600 12500 6700
rect 8405 6524 12600 6600
rect 8300 6500 12600 6524
rect 8300 6400 12800 6500
rect 8200 6300 13000 6400
rect 8200 6200 13200 6300
rect 8100 6100 13300 6200
rect 8100 6000 13400 6100
rect 8100 5900 13500 6000
rect 8000 5800 9800 5900
rect 10000 5800 13600 5900
rect 7900 5700 9700 5800
rect 10300 5700 13700 5800
rect 7800 5600 9600 5700
rect 10900 5600 13700 5700
rect 7700 5500 9600 5600
rect 11200 5500 13800 5600
rect 6000 5400 9500 5500
rect 11800 5400 13800 5500
rect 5600 5300 9400 5400
rect 12200 5300 13800 5400
rect 5400 5200 9400 5300
rect 12500 5200 13800 5300
rect 5300 5000 9300 5200
rect 5300 4900 9200 5000
rect 5300 4800 9100 4900
rect 12600 4800 13900 5200
rect 5300 4700 9000 4800
rect 5300 4600 8900 4700
rect 5300 4500 8800 4600
rect 5300 4400 8600 4500
rect 5300 4300 8200 4400
rect 5300 4100 6300 4300
rect 6900 4200 7300 4300
rect 12700 4200 13900 4800
rect 5400 3900 6300 4100
rect 5400 3700 6400 3900
rect 5500 3600 6600 3700
rect 5600 3500 6600 3600
rect 12800 3600 13900 4200
rect 14900 3869 15600 3900
rect 14900 3800 15700 3869
rect 14400 3700 15700 3800
rect 14100 3600 15600 3700
rect 12800 3500 15600 3600
rect 5600 3400 6700 3500
rect 12900 3400 15500 3500
rect 5700 3300 6900 3400
rect 12900 3300 15300 3400
rect 5900 3200 7000 3300
rect 12900 3200 15100 3300
rect 6300 3100 7100 3200
rect 12900 3100 14800 3200
rect 6400 3000 7200 3100
rect 12900 3000 14600 3100
rect 6600 2960 7200 3000
rect 6600 2900 7300 2960
rect 13000 2900 14300 3000
rect 6900 2800 7300 2900
rect 13100 2800 13900 2900
rect 13200 2700 13600 2800
<< properties >>
<< end >>
