** sch_path: /home/hni/TopmetalSe-Respin/xschem/array_SR.sch
.subckt array_SR ARRAY_OUT SF_IB gring VBIAS VDD VREF GND NB2 NB1 CSA_VREF ROW_ENA COL_ENA ROW_RST COL_RST ROW_DIN COL_DIN ROW_CLK
+ COL_CLK
*.PININFO ARRAY_OUT:O COL_ENA:I COL_RST:I COL_DIN:I COL_CLK:I ROW_ENA:I ROW_RST:I ROW_DIN:I ROW_CLK:I VBIAS:I VREF:I NB1:I gring:I
*+ CSA_VREF:I NB2:I SF_IB:I VDD:I GND:I
x1 VDD GND SF_IB gring VBIAS ARRAY_OUT ROW_SEL[0] ROW_SEL[1] ROW_SEL[2] ROW_SEL[3] ROW_SEL[4] ROW_SEL[5] ROW_SEL[6] ROW_SEL[7]
+ ROW_SEL[8] ROW_SEL[9] ROW_SEL[10] ROW_SEL[11] ROW_SEL[12] ROW_SEL[13] ROW_SEL[14] ROW_SEL[15] ROW_SEL[16] ROW_SEL[17] ROW_SEL[18]
+ ROW_SEL[19] ROW_SEL[20] ROW_SEL[21] ROW_SEL[22] ROW_SEL[23] ROW_SEL[24] ROW_SEL[25] ROW_SEL[26] ROW_SEL[27] ROW_SEL[28] ROW_SEL[29]
+ ROW_SEL[30] ROW_SEL[31] ROW_SEL[32] ROW_SEL[33] ROW_SEL[34] ROW_SEL[35] ROW_SEL[36] ROW_SEL[37] ROW_SEL[38] ROW_SEL[39] ROW_SEL[40]
+ ROW_SEL[41] ROW_SEL[42] ROW_SEL[43] ROW_SEL[44] ROW_SEL[45] ROW_SEL[46] ROW_SEL[47] ROW_SEL[48] ROW_SEL[49] ROW_SEL[50] ROW_SEL[51]
+ ROW_SEL[52] ROW_SEL[53] ROW_SEL[54] ROW_SEL[55] ROW_SEL[56] ROW_SEL[57] ROW_SEL[58] ROW_SEL[59] ROW_SEL[60] ROW_SEL[61] ROW_SEL[62]
+ ROW_SEL[63] ROW_SEL[64] ROW_SEL[65] ROW_SEL[66] ROW_SEL[67] ROW_SEL[68] ROW_SEL[69] ROW_SEL[70] ROW_SEL[71] ROW_SEL[72] ROW_SEL[73]
+ ROW_SEL[74] ROW_SEL[75] ROW_SEL[76] ROW_SEL[77] ROW_SEL[78] ROW_SEL[79] ROW_SEL[80] ROW_SEL[81] ROW_SEL[82] ROW_SEL[83] ROW_SEL[84]
+ ROW_SEL[85] ROW_SEL[86] ROW_SEL[87] ROW_SEL[88] ROW_SEL[89] ROW_SEL[90] ROW_SEL[91] ROW_SEL[92] ROW_SEL[93] ROW_SEL[94] ROW_SEL[95]
+ ROW_SEL[96] ROW_SEL[97] ROW_SEL[98] ROW_SEL[99] VREF NB2 NB1 CSA_VREF COL_SEL[0] COL_SEL[1] COL_SEL[2] COL_SEL[3] COL_SEL[4] COL_SEL[5]
+ COL_SEL[6] COL_SEL[7] COL_SEL[8] COL_SEL[9] COL_SEL[10] COL_SEL[11] COL_SEL[12] COL_SEL[13] COL_SEL[14] COL_SEL[15] COL_SEL[16] COL_SEL[17]
+ COL_SEL[18] COL_SEL[19] COL_SEL[20] COL_SEL[21] COL_SEL[22] COL_SEL[23] COL_SEL[24] COL_SEL[25] COL_SEL[26] COL_SEL[27] COL_SEL[28]
+ COL_SEL[29] COL_SEL[30] COL_SEL[31] COL_SEL[32] COL_SEL[33] COL_SEL[34] COL_SEL[35] COL_SEL[36] COL_SEL[37] COL_SEL[38] COL_SEL[39]
+ COL_SEL[40] COL_SEL[41] COL_SEL[42] COL_SEL[43] COL_SEL[44] COL_SEL[45] COL_SEL[46] COL_SEL[47] COL_SEL[48] COL_SEL[49] COL_SEL[50]
+ COL_SEL[51] COL_SEL[52] COL_SEL[53] COL_SEL[54] COL_SEL[55] COL_SEL[56] COL_SEL[57] COL_SEL[58] COL_SEL[59] COL_SEL[60] COL_SEL[61]
+ COL_SEL[62] COL_SEL[63] COL_SEL[64] COL_SEL[65] COL_SEL[66] COL_SEL[67] COL_SEL[68] COL_SEL[69] COL_SEL[70] COL_SEL[71] COL_SEL[72]
+ COL_SEL[73] COL_SEL[74] COL_SEL[75] COL_SEL[76] COL_SEL[77] COL_SEL[78] COL_SEL[79] COL_SEL[80] COL_SEL[81] COL_SEL[82] COL_SEL[83]
+ COL_SEL[84] COL_SEL[85] COL_SEL[86] COL_SEL[87] COL_SEL[88] COL_SEL[89] COL_SEL[90] COL_SEL[91] COL_SEL[92] COL_SEL[93] COL_SEL[94]
+ COL_SEL[95] COL_SEL[96] COL_SEL[97] COL_SEL[98] COL_SEL[99] array100
x3 GND VDD ROW_CLK ROW_DIN net1 ROW_ENA ROW_RST ROW_SEL[99] ROW_SEL[98] ROW_SEL[97] ROW_SEL[96] ROW_SEL[95] ROW_SEL[94]
+ ROW_SEL[93] ROW_SEL[92] ROW_SEL[91] ROW_SEL[90] ROW_SEL[89] ROW_SEL[88] ROW_SEL[87] ROW_SEL[86] ROW_SEL[85] ROW_SEL[84] ROW_SEL[83]
+ ROW_SEL[82] ROW_SEL[81] ROW_SEL[80] ROW_SEL[79] ROW_SEL[78] ROW_SEL[77] ROW_SEL[76] ROW_SEL[75] ROW_SEL[74] ROW_SEL[73] ROW_SEL[72]
+ ROW_SEL[71] ROW_SEL[70] ROW_SEL[69] ROW_SEL[68] ROW_SEL[67] ROW_SEL[66] ROW_SEL[65] ROW_SEL[64] ROW_SEL[63] ROW_SEL[62] ROW_SEL[61]
+ ROW_SEL[60] ROW_SEL[59] ROW_SEL[58] ROW_SEL[57] ROW_SEL[56] ROW_SEL[55] ROW_SEL[54] ROW_SEL[53] ROW_SEL[52] ROW_SEL[51] ROW_SEL[50]
+ ROW_SEL[49] ROW_SEL[48] ROW_SEL[47] ROW_SEL[46] ROW_SEL[45] ROW_SEL[44] ROW_SEL[43] ROW_SEL[42] ROW_SEL[41] ROW_SEL[40] ROW_SEL[39]
+ ROW_SEL[38] ROW_SEL[37] ROW_SEL[36] ROW_SEL[35] ROW_SEL[34] ROW_SEL[33] ROW_SEL[32] ROW_SEL[31] ROW_SEL[30] ROW_SEL[29] ROW_SEL[28]
+ ROW_SEL[27] ROW_SEL[26] ROW_SEL[25] ROW_SEL[24] ROW_SEL[23] ROW_SEL[22] ROW_SEL[21] ROW_SEL[20] ROW_SEL[19] ROW_SEL[18] ROW_SEL[17]
+ ROW_SEL[16] ROW_SEL[15] ROW_SEL[14] ROW_SEL[13] ROW_SEL[12] ROW_SEL[11] ROW_SEL[10] ROW_SEL[9] ROW_SEL[8] ROW_SEL[7] ROW_SEL[6] ROW_SEL[5]
+ ROW_SEL[4] ROW_SEL[3] ROW_SEL[2] ROW_SEL[1] ROW_SEL[0] shift_register
x2 GND VDD COL_CLK COL_DIN net2 COL_ENA COL_RST COL_SEL[99] COL_SEL[98] COL_SEL[97] COL_SEL[96] COL_SEL[95] COL_SEL[94]
+ COL_SEL[93] COL_SEL[92] COL_SEL[91] COL_SEL[90] COL_SEL[89] COL_SEL[88] COL_SEL[87] COL_SEL[86] COL_SEL[85] COL_SEL[84] COL_SEL[83]
+ COL_SEL[82] COL_SEL[81] COL_SEL[80] COL_SEL[79] COL_SEL[78] COL_SEL[77] COL_SEL[76] COL_SEL[75] COL_SEL[74] COL_SEL[73] COL_SEL[72]
+ COL_SEL[71] COL_SEL[70] COL_SEL[69] COL_SEL[68] COL_SEL[67] COL_SEL[66] COL_SEL[65] COL_SEL[64] COL_SEL[63] COL_SEL[62] COL_SEL[61]
+ COL_SEL[60] COL_SEL[59] COL_SEL[58] COL_SEL[57] COL_SEL[56] COL_SEL[55] COL_SEL[54] COL_SEL[53] COL_SEL[52] COL_SEL[51] COL_SEL[50]
+ COL_SEL[49] COL_SEL[48] COL_SEL[47] COL_SEL[46] COL_SEL[45] COL_SEL[44] COL_SEL[43] COL_SEL[42] COL_SEL[41] COL_SEL[40] COL_SEL[39]
+ COL_SEL[38] COL_SEL[37] COL_SEL[36] COL_SEL[35] COL_SEL[34] COL_SEL[33] COL_SEL[32] COL_SEL[31] COL_SEL[30] COL_SEL[29] COL_SEL[28]
+ COL_SEL[27] COL_SEL[26] COL_SEL[25] COL_SEL[24] COL_SEL[23] COL_SEL[22] COL_SEL[21] COL_SEL[20] COL_SEL[19] COL_SEL[18] COL_SEL[17]
+ COL_SEL[16] COL_SEL[15] COL_SEL[14] COL_SEL[13] COL_SEL[12] COL_SEL[11] COL_SEL[10] COL_SEL[9] COL_SEL[8] COL_SEL[7] COL_SEL[6] COL_SEL[5]
+ COL_SEL[4] COL_SEL[3] COL_SEL[2] COL_SEL[1] COL_SEL[0] shift_registerC
.ends

* expanding   symbol:  array100.sym # of pins=12
** sym_path: /home/hni/TopmetalSe-Respin/xschem/array100.sym
** sch_path: /home/hni/TopmetalSe-Respin/xschem/array100.sch
.subckt array100 VDD GND SF_IB gring VBIAS ARRAY_OUT ROW_SEL[0] ROW_SEL[1] ROW_SEL[2] ROW_SEL[3] ROW_SEL[4] ROW_SEL[5] ROW_SEL[6]
+ ROW_SEL[7] ROW_SEL[8] ROW_SEL[9] ROW_SEL[10] ROW_SEL[11] ROW_SEL[12] ROW_SEL[13] ROW_SEL[14] ROW_SEL[15] ROW_SEL[16] ROW_SEL[17] ROW_SEL[18]
+ ROW_SEL[19] ROW_SEL[20] ROW_SEL[21] ROW_SEL[22] ROW_SEL[23] ROW_SEL[24] ROW_SEL[25] ROW_SEL[26] ROW_SEL[27] ROW_SEL[28] ROW_SEL[29]
+ ROW_SEL[30] ROW_SEL[31] ROW_SEL[32] ROW_SEL[33] ROW_SEL[34] ROW_SEL[35] ROW_SEL[36] ROW_SEL[37] ROW_SEL[38] ROW_SEL[39] ROW_SEL[40]
+ ROW_SEL[41] ROW_SEL[42] ROW_SEL[43] ROW_SEL[44] ROW_SEL[45] ROW_SEL[46] ROW_SEL[47] ROW_SEL[48] ROW_SEL[49] ROW_SEL[50] ROW_SEL[51]
+ ROW_SEL[52] ROW_SEL[53] ROW_SEL[54] ROW_SEL[55] ROW_SEL[56] ROW_SEL[57] ROW_SEL[58] ROW_SEL[59] ROW_SEL[60] ROW_SEL[61] ROW_SEL[62]
+ ROW_SEL[63] ROW_SEL[64] ROW_SEL[65] ROW_SEL[66] ROW_SEL[67] ROW_SEL[68] ROW_SEL[69] ROW_SEL[70] ROW_SEL[71] ROW_SEL[72] ROW_SEL[73]
+ ROW_SEL[74] ROW_SEL[75] ROW_SEL[76] ROW_SEL[77] ROW_SEL[78] ROW_SEL[79] ROW_SEL[80] ROW_SEL[81] ROW_SEL[82] ROW_SEL[83] ROW_SEL[84]
+ ROW_SEL[85] ROW_SEL[86] ROW_SEL[87] ROW_SEL[88] ROW_SEL[89] ROW_SEL[90] ROW_SEL[91] ROW_SEL[92] ROW_SEL[93] ROW_SEL[94] ROW_SEL[95]
+ ROW_SEL[96] ROW_SEL[97] ROW_SEL[98] ROW_SEL[99] VREF NB2 NB1 CSA_VREF COL_SEL[0] COL_SEL[1] COL_SEL[2] COL_SEL[3] COL_SEL[4] COL_SEL[5]
+ COL_SEL[6] COL_SEL[7] COL_SEL[8] COL_SEL[9] COL_SEL[10] COL_SEL[11] COL_SEL[12] COL_SEL[13] COL_SEL[14] COL_SEL[15] COL_SEL[16] COL_SEL[17]
+ COL_SEL[18] COL_SEL[19] COL_SEL[20] COL_SEL[21] COL_SEL[22] COL_SEL[23] COL_SEL[24] COL_SEL[25] COL_SEL[26] COL_SEL[27] COL_SEL[28]
+ COL_SEL[29] COL_SEL[30] COL_SEL[31] COL_SEL[32] COL_SEL[33] COL_SEL[34] COL_SEL[35] COL_SEL[36] COL_SEL[37] COL_SEL[38] COL_SEL[39]
+ COL_SEL[40] COL_SEL[41] COL_SEL[42] COL_SEL[43] COL_SEL[44] COL_SEL[45] COL_SEL[46] COL_SEL[47] COL_SEL[48] COL_SEL[49] COL_SEL[50]
+ COL_SEL[51] COL_SEL[52] COL_SEL[53] COL_SEL[54] COL_SEL[55] COL_SEL[56] COL_SEL[57] COL_SEL[58] COL_SEL[59] COL_SEL[60] COL_SEL[61]
+ COL_SEL[62] COL_SEL[63] COL_SEL[64] COL_SEL[65] COL_SEL[66] COL_SEL[67] COL_SEL[68] COL_SEL[69] COL_SEL[70] COL_SEL[71] COL_SEL[72]
+ COL_SEL[73] COL_SEL[74] COL_SEL[75] COL_SEL[76] COL_SEL[77] COL_SEL[78] COL_SEL[79] COL_SEL[80] COL_SEL[81] COL_SEL[82] COL_SEL[83]
+ COL_SEL[84] COL_SEL[85] COL_SEL[86] COL_SEL[87] COL_SEL[88] COL_SEL[89] COL_SEL[90] COL_SEL[91] COL_SEL[92] COL_SEL[93] COL_SEL[94]
+ COL_SEL[95] COL_SEL[96] COL_SEL[97] COL_SEL[98] COL_SEL[99]
*.PININFO VDD:I GND:I SF_IB:I gring:I VBIAS:I ARRAY_OUT:O ROW_SEL[0:99]:I VREF:I NB2:I NB1:I CSA_VREF:I COL_SEL[0:99]:I
xPix0 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[0] VREF PIX_IN[0] NB2 NB1 CSA_VREF pixel
xPix1 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[0] VREF PIX_IN[1] NB2 NB1 CSA_VREF pixel
xPix2 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[0] VREF PIX_IN[2] NB2 NB1 CSA_VREF pixel
xPix3 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[0] VREF PIX_IN[3] NB2 NB1 CSA_VREF pixel
xPix4 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[0] VREF PIX_IN[4] NB2 NB1 CSA_VREF pixel
xPix5 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[0] VREF PIX_IN[5] NB2 NB1 CSA_VREF pixel
xPix6 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[0] VREF PIX_IN[6] NB2 NB1 CSA_VREF pixel
xPix7 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[0] VREF PIX_IN[7] NB2 NB1 CSA_VREF pixel
xPix8 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[0] VREF PIX_IN[8] NB2 NB1 CSA_VREF pixel
xPix9 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[0] VREF PIX_IN[9] NB2 NB1 CSA_VREF pixel
xPix10 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[0] VREF PIX_IN[10] NB2 NB1 CSA_VREF pixel
xPix11 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[0] VREF PIX_IN[11] NB2 NB1 CSA_VREF pixel
xPix12 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[0] VREF PIX_IN[12] NB2 NB1 CSA_VREF pixel
xPix13 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[0] VREF PIX_IN[13] NB2 NB1 CSA_VREF pixel
xPix14 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[0] VREF PIX_IN[14] NB2 NB1 CSA_VREF pixel
xPix15 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[0] VREF PIX_IN[15] NB2 NB1 CSA_VREF pixel
xPix16 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[0] VREF PIX_IN[16] NB2 NB1 CSA_VREF pixel
xPix17 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[0] VREF PIX_IN[17] NB2 NB1 CSA_VREF pixel
xPix18 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[0] VREF PIX_IN[18] NB2 NB1 CSA_VREF pixel
xPix19 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[0] VREF PIX_IN[19] NB2 NB1 CSA_VREF pixel
xPix20 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[0] VREF PIX_IN[20] NB2 NB1 CSA_VREF pixel
xPix21 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[0] VREF PIX_IN[21] NB2 NB1 CSA_VREF pixel
xPix22 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[0] VREF PIX_IN[22] NB2 NB1 CSA_VREF pixel
xPix23 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[0] VREF PIX_IN[23] NB2 NB1 CSA_VREF pixel
xPix24 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[0] VREF PIX_IN[24] NB2 NB1 CSA_VREF pixel
xPix25 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[0] VREF PIX_IN[25] NB2 NB1 CSA_VREF pixel
xPix26 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[0] VREF PIX_IN[26] NB2 NB1 CSA_VREF pixel
xPix27 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[0] VREF PIX_IN[27] NB2 NB1 CSA_VREF pixel
xPix28 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[0] VREF PIX_IN[28] NB2 NB1 CSA_VREF pixel
xPix29 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[0] VREF PIX_IN[29] NB2 NB1 CSA_VREF pixel
xPix30 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[0] VREF PIX_IN[30] NB2 NB1 CSA_VREF pixel
xPix31 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[0] VREF PIX_IN[31] NB2 NB1 CSA_VREF pixel
xPix32 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[0] VREF PIX_IN[32] NB2 NB1 CSA_VREF pixel
xPix33 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[0] VREF PIX_IN[33] NB2 NB1 CSA_VREF pixel
xPix34 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[0] VREF PIX_IN[34] NB2 NB1 CSA_VREF pixel
xPix35 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[0] VREF PIX_IN[35] NB2 NB1 CSA_VREF pixel
xPix36 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[0] VREF PIX_IN[36] NB2 NB1 CSA_VREF pixel
xPix37 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[0] VREF PIX_IN[37] NB2 NB1 CSA_VREF pixel
xPix38 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[0] VREF PIX_IN[38] NB2 NB1 CSA_VREF pixel
xPix39 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[0] VREF PIX_IN[39] NB2 NB1 CSA_VREF pixel
xPix40 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[0] VREF PIX_IN[40] NB2 NB1 CSA_VREF pixel
xPix41 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[0] VREF PIX_IN[41] NB2 NB1 CSA_VREF pixel
xPix42 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[0] VREF PIX_IN[42] NB2 NB1 CSA_VREF pixel
xPix43 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[0] VREF PIX_IN[43] NB2 NB1 CSA_VREF pixel
xPix44 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[0] VREF PIX_IN[44] NB2 NB1 CSA_VREF pixel
xPix45 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[0] VREF PIX_IN[45] NB2 NB1 CSA_VREF pixel
xPix46 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[0] VREF PIX_IN[46] NB2 NB1 CSA_VREF pixel
xPix47 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[0] VREF PIX_IN[47] NB2 NB1 CSA_VREF pixel
xPix48 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[0] VREF PIX_IN[48] NB2 NB1 CSA_VREF pixel
xPix49 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[0] VREF PIX_IN[49] NB2 NB1 CSA_VREF pixel
xPix50 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[0] VREF PIX_IN[50] NB2 NB1 CSA_VREF pixel
xPix51 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[0] VREF PIX_IN[51] NB2 NB1 CSA_VREF pixel
xPix52 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[0] VREF PIX_IN[52] NB2 NB1 CSA_VREF pixel
xPix53 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[0] VREF PIX_IN[53] NB2 NB1 CSA_VREF pixel
xPix54 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[0] VREF PIX_IN[54] NB2 NB1 CSA_VREF pixel
xPix55 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[0] VREF PIX_IN[55] NB2 NB1 CSA_VREF pixel
xPix56 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[0] VREF PIX_IN[56] NB2 NB1 CSA_VREF pixel
xPix57 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[0] VREF PIX_IN[57] NB2 NB1 CSA_VREF pixel
xPix58 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[0] VREF PIX_IN[58] NB2 NB1 CSA_VREF pixel
xPix59 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[0] VREF PIX_IN[59] NB2 NB1 CSA_VREF pixel
xPix60 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[0] VREF PIX_IN[60] NB2 NB1 CSA_VREF pixel
xPix61 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[0] VREF PIX_IN[61] NB2 NB1 CSA_VREF pixel
xPix62 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[0] VREF PIX_IN[62] NB2 NB1 CSA_VREF pixel
xPix63 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[0] VREF PIX_IN[63] NB2 NB1 CSA_VREF pixel
xPix64 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[0] VREF PIX_IN[64] NB2 NB1 CSA_VREF pixel
xPix65 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[0] VREF PIX_IN[65] NB2 NB1 CSA_VREF pixel
xPix66 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[0] VREF PIX_IN[66] NB2 NB1 CSA_VREF pixel
xPix67 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[0] VREF PIX_IN[67] NB2 NB1 CSA_VREF pixel
xPix68 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[0] VREF PIX_IN[68] NB2 NB1 CSA_VREF pixel
xPix69 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[0] VREF PIX_IN[69] NB2 NB1 CSA_VREF pixel
xPix70 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[0] VREF PIX_IN[70] NB2 NB1 CSA_VREF pixel
xPix71 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[0] VREF PIX_IN[71] NB2 NB1 CSA_VREF pixel
xPix72 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[0] VREF PIX_IN[72] NB2 NB1 CSA_VREF pixel
xPix73 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[0] VREF PIX_IN[73] NB2 NB1 CSA_VREF pixel
xPix74 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[0] VREF PIX_IN[74] NB2 NB1 CSA_VREF pixel
xPix75 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[0] VREF PIX_IN[75] NB2 NB1 CSA_VREF pixel
xPix76 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[0] VREF PIX_IN[76] NB2 NB1 CSA_VREF pixel
xPix77 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[0] VREF PIX_IN[77] NB2 NB1 CSA_VREF pixel
xPix78 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[0] VREF PIX_IN[78] NB2 NB1 CSA_VREF pixel
xPix79 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[0] VREF PIX_IN[79] NB2 NB1 CSA_VREF pixel
xPix80 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[0] VREF PIX_IN[80] NB2 NB1 CSA_VREF pixel
xPix81 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[0] VREF PIX_IN[81] NB2 NB1 CSA_VREF pixel
xPix82 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[0] VREF PIX_IN[82] NB2 NB1 CSA_VREF pixel
xPix83 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[0] VREF PIX_IN[83] NB2 NB1 CSA_VREF pixel
xPix84 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[0] VREF PIX_IN[84] NB2 NB1 CSA_VREF pixel
xPix85 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[0] VREF PIX_IN[85] NB2 NB1 CSA_VREF pixel
xPix86 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[0] VREF PIX_IN[86] NB2 NB1 CSA_VREF pixel
xPix87 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[0] VREF PIX_IN[87] NB2 NB1 CSA_VREF pixel
xPix88 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[0] VREF PIX_IN[88] NB2 NB1 CSA_VREF pixel
xPix89 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[0] VREF PIX_IN[89] NB2 NB1 CSA_VREF pixel
xPix90 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[0] VREF PIX_IN[90] NB2 NB1 CSA_VREF pixel
xPix91 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[0] VREF PIX_IN[91] NB2 NB1 CSA_VREF pixel
xPix92 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[0] VREF PIX_IN[92] NB2 NB1 CSA_VREF pixel
xPix93 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[0] VREF PIX_IN[93] NB2 NB1 CSA_VREF pixel
xPix94 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[0] VREF PIX_IN[94] NB2 NB1 CSA_VREF pixel
xPix95 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[0] VREF PIX_IN[95] NB2 NB1 CSA_VREF pixel
xPix96 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[0] VREF PIX_IN[96] NB2 NB1 CSA_VREF pixel
xPix97 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[0] VREF PIX_IN[97] NB2 NB1 CSA_VREF pixel
xPix98 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[0] VREF PIX_IN[98] NB2 NB1 CSA_VREF pixel
xPix99 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[0] VREF PIX_IN[99] NB2 NB1 CSA_VREF pixel
xPix100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[1] VREF PIX_IN[100] NB2 NB1 CSA_VREF pixel
xPix101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[1] VREF PIX_IN[101] NB2 NB1 CSA_VREF pixel
xPix102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[1] VREF PIX_IN[102] NB2 NB1 CSA_VREF pixel
xPix103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[1] VREF PIX_IN[103] NB2 NB1 CSA_VREF pixel
xPix104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[1] VREF PIX_IN[104] NB2 NB1 CSA_VREF pixel
xPix105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[1] VREF PIX_IN[105] NB2 NB1 CSA_VREF pixel
xPix106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[1] VREF PIX_IN[106] NB2 NB1 CSA_VREF pixel
xPix107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[1] VREF PIX_IN[107] NB2 NB1 CSA_VREF pixel
xPix108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[1] VREF PIX_IN[108] NB2 NB1 CSA_VREF pixel
xPix109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[1] VREF PIX_IN[109] NB2 NB1 CSA_VREF pixel
xPix110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[1] VREF PIX_IN[110] NB2 NB1 CSA_VREF pixel
xPix111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[1] VREF PIX_IN[111] NB2 NB1 CSA_VREF pixel
xPix112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[1] VREF PIX_IN[112] NB2 NB1 CSA_VREF pixel
xPix113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[1] VREF PIX_IN[113] NB2 NB1 CSA_VREF pixel
xPix114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[1] VREF PIX_IN[114] NB2 NB1 CSA_VREF pixel
xPix115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[1] VREF PIX_IN[115] NB2 NB1 CSA_VREF pixel
xPix116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[1] VREF PIX_IN[116] NB2 NB1 CSA_VREF pixel
xPix117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[1] VREF PIX_IN[117] NB2 NB1 CSA_VREF pixel
xPix118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[1] VREF PIX_IN[118] NB2 NB1 CSA_VREF pixel
xPix119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[1] VREF PIX_IN[119] NB2 NB1 CSA_VREF pixel
xPix120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[1] VREF PIX_IN[120] NB2 NB1 CSA_VREF pixel
xPix121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[1] VREF PIX_IN[121] NB2 NB1 CSA_VREF pixel
xPix122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[1] VREF PIX_IN[122] NB2 NB1 CSA_VREF pixel
xPix123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[1] VREF PIX_IN[123] NB2 NB1 CSA_VREF pixel
xPix124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[1] VREF PIX_IN[124] NB2 NB1 CSA_VREF pixel
xPix125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[1] VREF PIX_IN[125] NB2 NB1 CSA_VREF pixel
xPix126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[1] VREF PIX_IN[126] NB2 NB1 CSA_VREF pixel
xPix127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[1] VREF PIX_IN[127] NB2 NB1 CSA_VREF pixel
xPix128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[1] VREF PIX_IN[128] NB2 NB1 CSA_VREF pixel
xPix129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[1] VREF PIX_IN[129] NB2 NB1 CSA_VREF pixel
xPix130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[1] VREF PIX_IN[130] NB2 NB1 CSA_VREF pixel
xPix131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[1] VREF PIX_IN[131] NB2 NB1 CSA_VREF pixel
xPix132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[1] VREF PIX_IN[132] NB2 NB1 CSA_VREF pixel
xPix133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[1] VREF PIX_IN[133] NB2 NB1 CSA_VREF pixel
xPix134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[1] VREF PIX_IN[134] NB2 NB1 CSA_VREF pixel
xPix135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[1] VREF PIX_IN[135] NB2 NB1 CSA_VREF pixel
xPix136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[1] VREF PIX_IN[136] NB2 NB1 CSA_VREF pixel
xPix137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[1] VREF PIX_IN[137] NB2 NB1 CSA_VREF pixel
xPix138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[1] VREF PIX_IN[138] NB2 NB1 CSA_VREF pixel
xPix139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[1] VREF PIX_IN[139] NB2 NB1 CSA_VREF pixel
xPix140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[1] VREF PIX_IN[140] NB2 NB1 CSA_VREF pixel
xPix141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[1] VREF PIX_IN[141] NB2 NB1 CSA_VREF pixel
xPix142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[1] VREF PIX_IN[142] NB2 NB1 CSA_VREF pixel
xPix143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[1] VREF PIX_IN[143] NB2 NB1 CSA_VREF pixel
xPix144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[1] VREF PIX_IN[144] NB2 NB1 CSA_VREF pixel
xPix145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[1] VREF PIX_IN[145] NB2 NB1 CSA_VREF pixel
xPix146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[1] VREF PIX_IN[146] NB2 NB1 CSA_VREF pixel
xPix147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[1] VREF PIX_IN[147] NB2 NB1 CSA_VREF pixel
xPix148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[1] VREF PIX_IN[148] NB2 NB1 CSA_VREF pixel
xPix149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[1] VREF PIX_IN[149] NB2 NB1 CSA_VREF pixel
xPix150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[1] VREF PIX_IN[150] NB2 NB1 CSA_VREF pixel
xPix151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[1] VREF PIX_IN[151] NB2 NB1 CSA_VREF pixel
xPix152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[1] VREF PIX_IN[152] NB2 NB1 CSA_VREF pixel
xPix153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[1] VREF PIX_IN[153] NB2 NB1 CSA_VREF pixel
xPix154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[1] VREF PIX_IN[154] NB2 NB1 CSA_VREF pixel
xPix155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[1] VREF PIX_IN[155] NB2 NB1 CSA_VREF pixel
xPix156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[1] VREF PIX_IN[156] NB2 NB1 CSA_VREF pixel
xPix157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[1] VREF PIX_IN[157] NB2 NB1 CSA_VREF pixel
xPix158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[1] VREF PIX_IN[158] NB2 NB1 CSA_VREF pixel
xPix159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[1] VREF PIX_IN[159] NB2 NB1 CSA_VREF pixel
xPix160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[1] VREF PIX_IN[160] NB2 NB1 CSA_VREF pixel
xPix161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[1] VREF PIX_IN[161] NB2 NB1 CSA_VREF pixel
xPix162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[1] VREF PIX_IN[162] NB2 NB1 CSA_VREF pixel
xPix163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[1] VREF PIX_IN[163] NB2 NB1 CSA_VREF pixel
xPix164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[1] VREF PIX_IN[164] NB2 NB1 CSA_VREF pixel
xPix165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[1] VREF PIX_IN[165] NB2 NB1 CSA_VREF pixel
xPix166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[1] VREF PIX_IN[166] NB2 NB1 CSA_VREF pixel
xPix167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[1] VREF PIX_IN[167] NB2 NB1 CSA_VREF pixel
xPix168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[1] VREF PIX_IN[168] NB2 NB1 CSA_VREF pixel
xPix169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[1] VREF PIX_IN[169] NB2 NB1 CSA_VREF pixel
xPix170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[1] VREF PIX_IN[170] NB2 NB1 CSA_VREF pixel
xPix171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[1] VREF PIX_IN[171] NB2 NB1 CSA_VREF pixel
xPix172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[1] VREF PIX_IN[172] NB2 NB1 CSA_VREF pixel
xPix173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[1] VREF PIX_IN[173] NB2 NB1 CSA_VREF pixel
xPix174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[1] VREF PIX_IN[174] NB2 NB1 CSA_VREF pixel
xPix175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[1] VREF PIX_IN[175] NB2 NB1 CSA_VREF pixel
xPix176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[1] VREF PIX_IN[176] NB2 NB1 CSA_VREF pixel
xPix177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[1] VREF PIX_IN[177] NB2 NB1 CSA_VREF pixel
xPix178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[1] VREF PIX_IN[178] NB2 NB1 CSA_VREF pixel
xPix179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[1] VREF PIX_IN[179] NB2 NB1 CSA_VREF pixel
xPix180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[1] VREF PIX_IN[180] NB2 NB1 CSA_VREF pixel
xPix181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[1] VREF PIX_IN[181] NB2 NB1 CSA_VREF pixel
xPix182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[1] VREF PIX_IN[182] NB2 NB1 CSA_VREF pixel
xPix183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[1] VREF PIX_IN[183] NB2 NB1 CSA_VREF pixel
xPix184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[1] VREF PIX_IN[184] NB2 NB1 CSA_VREF pixel
xPix185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[1] VREF PIX_IN[185] NB2 NB1 CSA_VREF pixel
xPix186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[1] VREF PIX_IN[186] NB2 NB1 CSA_VREF pixel
xPix187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[1] VREF PIX_IN[187] NB2 NB1 CSA_VREF pixel
xPix188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[1] VREF PIX_IN[188] NB2 NB1 CSA_VREF pixel
xPix189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[1] VREF PIX_IN[189] NB2 NB1 CSA_VREF pixel
xPix190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[1] VREF PIX_IN[190] NB2 NB1 CSA_VREF pixel
xPix191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[1] VREF PIX_IN[191] NB2 NB1 CSA_VREF pixel
xPix192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[1] VREF PIX_IN[192] NB2 NB1 CSA_VREF pixel
xPix193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[1] VREF PIX_IN[193] NB2 NB1 CSA_VREF pixel
xPix194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[1] VREF PIX_IN[194] NB2 NB1 CSA_VREF pixel
xPix195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[1] VREF PIX_IN[195] NB2 NB1 CSA_VREF pixel
xPix196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[1] VREF PIX_IN[196] NB2 NB1 CSA_VREF pixel
xPix197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[1] VREF PIX_IN[197] NB2 NB1 CSA_VREF pixel
xPix198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[1] VREF PIX_IN[198] NB2 NB1 CSA_VREF pixel
xPix199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[1] VREF PIX_IN[199] NB2 NB1 CSA_VREF pixel
xPix200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[2] VREF PIX_IN[200] NB2 NB1 CSA_VREF pixel
xPix201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[2] VREF PIX_IN[201] NB2 NB1 CSA_VREF pixel
xPix202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[2] VREF PIX_IN[202] NB2 NB1 CSA_VREF pixel
xPix203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[2] VREF PIX_IN[203] NB2 NB1 CSA_VREF pixel
xPix204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[2] VREF PIX_IN[204] NB2 NB1 CSA_VREF pixel
xPix205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[2] VREF PIX_IN[205] NB2 NB1 CSA_VREF pixel
xPix206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[2] VREF PIX_IN[206] NB2 NB1 CSA_VREF pixel
xPix207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[2] VREF PIX_IN[207] NB2 NB1 CSA_VREF pixel
xPix208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[2] VREF PIX_IN[208] NB2 NB1 CSA_VREF pixel
xPix209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[2] VREF PIX_IN[209] NB2 NB1 CSA_VREF pixel
xPix210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[2] VREF PIX_IN[210] NB2 NB1 CSA_VREF pixel
xPix211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[2] VREF PIX_IN[211] NB2 NB1 CSA_VREF pixel
xPix212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[2] VREF PIX_IN[212] NB2 NB1 CSA_VREF pixel
xPix213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[2] VREF PIX_IN[213] NB2 NB1 CSA_VREF pixel
xPix214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[2] VREF PIX_IN[214] NB2 NB1 CSA_VREF pixel
xPix215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[2] VREF PIX_IN[215] NB2 NB1 CSA_VREF pixel
xPix216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[2] VREF PIX_IN[216] NB2 NB1 CSA_VREF pixel
xPix217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[2] VREF PIX_IN[217] NB2 NB1 CSA_VREF pixel
xPix218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[2] VREF PIX_IN[218] NB2 NB1 CSA_VREF pixel
xPix219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[2] VREF PIX_IN[219] NB2 NB1 CSA_VREF pixel
xPix220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[2] VREF PIX_IN[220] NB2 NB1 CSA_VREF pixel
xPix221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[2] VREF PIX_IN[221] NB2 NB1 CSA_VREF pixel
xPix222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[2] VREF PIX_IN[222] NB2 NB1 CSA_VREF pixel
xPix223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[2] VREF PIX_IN[223] NB2 NB1 CSA_VREF pixel
xPix224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[2] VREF PIX_IN[224] NB2 NB1 CSA_VREF pixel
xPix225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[2] VREF PIX_IN[225] NB2 NB1 CSA_VREF pixel
xPix226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[2] VREF PIX_IN[226] NB2 NB1 CSA_VREF pixel
xPix227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[2] VREF PIX_IN[227] NB2 NB1 CSA_VREF pixel
xPix228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[2] VREF PIX_IN[228] NB2 NB1 CSA_VREF pixel
xPix229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[2] VREF PIX_IN[229] NB2 NB1 CSA_VREF pixel
xPix230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[2] VREF PIX_IN[230] NB2 NB1 CSA_VREF pixel
xPix231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[2] VREF PIX_IN[231] NB2 NB1 CSA_VREF pixel
xPix232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[2] VREF PIX_IN[232] NB2 NB1 CSA_VREF pixel
xPix233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[2] VREF PIX_IN[233] NB2 NB1 CSA_VREF pixel
xPix234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[2] VREF PIX_IN[234] NB2 NB1 CSA_VREF pixel
xPix235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[2] VREF PIX_IN[235] NB2 NB1 CSA_VREF pixel
xPix236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[2] VREF PIX_IN[236] NB2 NB1 CSA_VREF pixel
xPix237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[2] VREF PIX_IN[237] NB2 NB1 CSA_VREF pixel
xPix238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[2] VREF PIX_IN[238] NB2 NB1 CSA_VREF pixel
xPix239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[2] VREF PIX_IN[239] NB2 NB1 CSA_VREF pixel
xPix240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[2] VREF PIX_IN[240] NB2 NB1 CSA_VREF pixel
xPix241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[2] VREF PIX_IN[241] NB2 NB1 CSA_VREF pixel
xPix242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[2] VREF PIX_IN[242] NB2 NB1 CSA_VREF pixel
xPix243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[2] VREF PIX_IN[243] NB2 NB1 CSA_VREF pixel
xPix244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[2] VREF PIX_IN[244] NB2 NB1 CSA_VREF pixel
xPix245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[2] VREF PIX_IN[245] NB2 NB1 CSA_VREF pixel
xPix246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[2] VREF PIX_IN[246] NB2 NB1 CSA_VREF pixel
xPix247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[2] VREF PIX_IN[247] NB2 NB1 CSA_VREF pixel
xPix248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[2] VREF PIX_IN[248] NB2 NB1 CSA_VREF pixel
xPix249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[2] VREF PIX_IN[249] NB2 NB1 CSA_VREF pixel
xPix250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[2] VREF PIX_IN[250] NB2 NB1 CSA_VREF pixel
xPix251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[2] VREF PIX_IN[251] NB2 NB1 CSA_VREF pixel
xPix252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[2] VREF PIX_IN[252] NB2 NB1 CSA_VREF pixel
xPix253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[2] VREF PIX_IN[253] NB2 NB1 CSA_VREF pixel
xPix254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[2] VREF PIX_IN[254] NB2 NB1 CSA_VREF pixel
xPix255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[2] VREF PIX_IN[255] NB2 NB1 CSA_VREF pixel
xPix256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[2] VREF PIX_IN[256] NB2 NB1 CSA_VREF pixel
xPix257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[2] VREF PIX_IN[257] NB2 NB1 CSA_VREF pixel
xPix258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[2] VREF PIX_IN[258] NB2 NB1 CSA_VREF pixel
xPix259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[2] VREF PIX_IN[259] NB2 NB1 CSA_VREF pixel
xPix260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[2] VREF PIX_IN[260] NB2 NB1 CSA_VREF pixel
xPix261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[2] VREF PIX_IN[261] NB2 NB1 CSA_VREF pixel
xPix262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[2] VREF PIX_IN[262] NB2 NB1 CSA_VREF pixel
xPix263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[2] VREF PIX_IN[263] NB2 NB1 CSA_VREF pixel
xPix264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[2] VREF PIX_IN[264] NB2 NB1 CSA_VREF pixel
xPix265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[2] VREF PIX_IN[265] NB2 NB1 CSA_VREF pixel
xPix266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[2] VREF PIX_IN[266] NB2 NB1 CSA_VREF pixel
xPix267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[2] VREF PIX_IN[267] NB2 NB1 CSA_VREF pixel
xPix268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[2] VREF PIX_IN[268] NB2 NB1 CSA_VREF pixel
xPix269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[2] VREF PIX_IN[269] NB2 NB1 CSA_VREF pixel
xPix270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[2] VREF PIX_IN[270] NB2 NB1 CSA_VREF pixel
xPix271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[2] VREF PIX_IN[271] NB2 NB1 CSA_VREF pixel
xPix272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[2] VREF PIX_IN[272] NB2 NB1 CSA_VREF pixel
xPix273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[2] VREF PIX_IN[273] NB2 NB1 CSA_VREF pixel
xPix274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[2] VREF PIX_IN[274] NB2 NB1 CSA_VREF pixel
xPix275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[2] VREF PIX_IN[275] NB2 NB1 CSA_VREF pixel
xPix276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[2] VREF PIX_IN[276] NB2 NB1 CSA_VREF pixel
xPix277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[2] VREF PIX_IN[277] NB2 NB1 CSA_VREF pixel
xPix278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[2] VREF PIX_IN[278] NB2 NB1 CSA_VREF pixel
xPix279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[2] VREF PIX_IN[279] NB2 NB1 CSA_VREF pixel
xPix280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[2] VREF PIX_IN[280] NB2 NB1 CSA_VREF pixel
xPix281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[2] VREF PIX_IN[281] NB2 NB1 CSA_VREF pixel
xPix282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[2] VREF PIX_IN[282] NB2 NB1 CSA_VREF pixel
xPix283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[2] VREF PIX_IN[283] NB2 NB1 CSA_VREF pixel
xPix284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[2] VREF PIX_IN[284] NB2 NB1 CSA_VREF pixel
xPix285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[2] VREF PIX_IN[285] NB2 NB1 CSA_VREF pixel
xPix286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[2] VREF PIX_IN[286] NB2 NB1 CSA_VREF pixel
xPix287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[2] VREF PIX_IN[287] NB2 NB1 CSA_VREF pixel
xPix288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[2] VREF PIX_IN[288] NB2 NB1 CSA_VREF pixel
xPix289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[2] VREF PIX_IN[289] NB2 NB1 CSA_VREF pixel
xPix290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[2] VREF PIX_IN[290] NB2 NB1 CSA_VREF pixel
xPix291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[2] VREF PIX_IN[291] NB2 NB1 CSA_VREF pixel
xPix292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[2] VREF PIX_IN[292] NB2 NB1 CSA_VREF pixel
xPix293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[2] VREF PIX_IN[293] NB2 NB1 CSA_VREF pixel
xPix294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[2] VREF PIX_IN[294] NB2 NB1 CSA_VREF pixel
xPix295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[2] VREF PIX_IN[295] NB2 NB1 CSA_VREF pixel
xPix296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[2] VREF PIX_IN[296] NB2 NB1 CSA_VREF pixel
xPix297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[2] VREF PIX_IN[297] NB2 NB1 CSA_VREF pixel
xPix298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[2] VREF PIX_IN[298] NB2 NB1 CSA_VREF pixel
xPix299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[2] VREF PIX_IN[299] NB2 NB1 CSA_VREF pixel
xPix300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[3] VREF PIX_IN[300] NB2 NB1 CSA_VREF pixel
xPix301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[3] VREF PIX_IN[301] NB2 NB1 CSA_VREF pixel
xPix302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[3] VREF PIX_IN[302] NB2 NB1 CSA_VREF pixel
xPix303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[3] VREF PIX_IN[303] NB2 NB1 CSA_VREF pixel
xPix304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[3] VREF PIX_IN[304] NB2 NB1 CSA_VREF pixel
xPix305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[3] VREF PIX_IN[305] NB2 NB1 CSA_VREF pixel
xPix306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[3] VREF PIX_IN[306] NB2 NB1 CSA_VREF pixel
xPix307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[3] VREF PIX_IN[307] NB2 NB1 CSA_VREF pixel
xPix308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[3] VREF PIX_IN[308] NB2 NB1 CSA_VREF pixel
xPix309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[3] VREF PIX_IN[309] NB2 NB1 CSA_VREF pixel
xPix310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[3] VREF PIX_IN[310] NB2 NB1 CSA_VREF pixel
xPix311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[3] VREF PIX_IN[311] NB2 NB1 CSA_VREF pixel
xPix312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[3] VREF PIX_IN[312] NB2 NB1 CSA_VREF pixel
xPix313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[3] VREF PIX_IN[313] NB2 NB1 CSA_VREF pixel
xPix314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[3] VREF PIX_IN[314] NB2 NB1 CSA_VREF pixel
xPix315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[3] VREF PIX_IN[315] NB2 NB1 CSA_VREF pixel
xPix316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[3] VREF PIX_IN[316] NB2 NB1 CSA_VREF pixel
xPix317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[3] VREF PIX_IN[317] NB2 NB1 CSA_VREF pixel
xPix318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[3] VREF PIX_IN[318] NB2 NB1 CSA_VREF pixel
xPix319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[3] VREF PIX_IN[319] NB2 NB1 CSA_VREF pixel
xPix320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[3] VREF PIX_IN[320] NB2 NB1 CSA_VREF pixel
xPix321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[3] VREF PIX_IN[321] NB2 NB1 CSA_VREF pixel
xPix322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[3] VREF PIX_IN[322] NB2 NB1 CSA_VREF pixel
xPix323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[3] VREF PIX_IN[323] NB2 NB1 CSA_VREF pixel
xPix324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[3] VREF PIX_IN[324] NB2 NB1 CSA_VREF pixel
xPix325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[3] VREF PIX_IN[325] NB2 NB1 CSA_VREF pixel
xPix326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[3] VREF PIX_IN[326] NB2 NB1 CSA_VREF pixel
xPix327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[3] VREF PIX_IN[327] NB2 NB1 CSA_VREF pixel
xPix328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[3] VREF PIX_IN[328] NB2 NB1 CSA_VREF pixel
xPix329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[3] VREF PIX_IN[329] NB2 NB1 CSA_VREF pixel
xPix330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[3] VREF PIX_IN[330] NB2 NB1 CSA_VREF pixel
xPix331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[3] VREF PIX_IN[331] NB2 NB1 CSA_VREF pixel
xPix332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[3] VREF PIX_IN[332] NB2 NB1 CSA_VREF pixel
xPix333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[3] VREF PIX_IN[333] NB2 NB1 CSA_VREF pixel
xPix334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[3] VREF PIX_IN[334] NB2 NB1 CSA_VREF pixel
xPix335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[3] VREF PIX_IN[335] NB2 NB1 CSA_VREF pixel
xPix336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[3] VREF PIX_IN[336] NB2 NB1 CSA_VREF pixel
xPix337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[3] VREF PIX_IN[337] NB2 NB1 CSA_VREF pixel
xPix338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[3] VREF PIX_IN[338] NB2 NB1 CSA_VREF pixel
xPix339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[3] VREF PIX_IN[339] NB2 NB1 CSA_VREF pixel
xPix340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[3] VREF PIX_IN[340] NB2 NB1 CSA_VREF pixel
xPix341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[3] VREF PIX_IN[341] NB2 NB1 CSA_VREF pixel
xPix342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[3] VREF PIX_IN[342] NB2 NB1 CSA_VREF pixel
xPix343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[3] VREF PIX_IN[343] NB2 NB1 CSA_VREF pixel
xPix344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[3] VREF PIX_IN[344] NB2 NB1 CSA_VREF pixel
xPix345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[3] VREF PIX_IN[345] NB2 NB1 CSA_VREF pixel
xPix346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[3] VREF PIX_IN[346] NB2 NB1 CSA_VREF pixel
xPix347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[3] VREF PIX_IN[347] NB2 NB1 CSA_VREF pixel
xPix348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[3] VREF PIX_IN[348] NB2 NB1 CSA_VREF pixel
xPix349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[3] VREF PIX_IN[349] NB2 NB1 CSA_VREF pixel
xPix350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[3] VREF PIX_IN[350] NB2 NB1 CSA_VREF pixel
xPix351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[3] VREF PIX_IN[351] NB2 NB1 CSA_VREF pixel
xPix352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[3] VREF PIX_IN[352] NB2 NB1 CSA_VREF pixel
xPix353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[3] VREF PIX_IN[353] NB2 NB1 CSA_VREF pixel
xPix354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[3] VREF PIX_IN[354] NB2 NB1 CSA_VREF pixel
xPix355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[3] VREF PIX_IN[355] NB2 NB1 CSA_VREF pixel
xPix356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[3] VREF PIX_IN[356] NB2 NB1 CSA_VREF pixel
xPix357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[3] VREF PIX_IN[357] NB2 NB1 CSA_VREF pixel
xPix358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[3] VREF PIX_IN[358] NB2 NB1 CSA_VREF pixel
xPix359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[3] VREF PIX_IN[359] NB2 NB1 CSA_VREF pixel
xPix360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[3] VREF PIX_IN[360] NB2 NB1 CSA_VREF pixel
xPix361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[3] VREF PIX_IN[361] NB2 NB1 CSA_VREF pixel
xPix362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[3] VREF PIX_IN[362] NB2 NB1 CSA_VREF pixel
xPix363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[3] VREF PIX_IN[363] NB2 NB1 CSA_VREF pixel
xPix364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[3] VREF PIX_IN[364] NB2 NB1 CSA_VREF pixel
xPix365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[3] VREF PIX_IN[365] NB2 NB1 CSA_VREF pixel
xPix366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[3] VREF PIX_IN[366] NB2 NB1 CSA_VREF pixel
xPix367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[3] VREF PIX_IN[367] NB2 NB1 CSA_VREF pixel
xPix368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[3] VREF PIX_IN[368] NB2 NB1 CSA_VREF pixel
xPix369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[3] VREF PIX_IN[369] NB2 NB1 CSA_VREF pixel
xPix370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[3] VREF PIX_IN[370] NB2 NB1 CSA_VREF pixel
xPix371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[3] VREF PIX_IN[371] NB2 NB1 CSA_VREF pixel
xPix372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[3] VREF PIX_IN[372] NB2 NB1 CSA_VREF pixel
xPix373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[3] VREF PIX_IN[373] NB2 NB1 CSA_VREF pixel
xPix374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[3] VREF PIX_IN[374] NB2 NB1 CSA_VREF pixel
xPix375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[3] VREF PIX_IN[375] NB2 NB1 CSA_VREF pixel
xPix376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[3] VREF PIX_IN[376] NB2 NB1 CSA_VREF pixel
xPix377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[3] VREF PIX_IN[377] NB2 NB1 CSA_VREF pixel
xPix378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[3] VREF PIX_IN[378] NB2 NB1 CSA_VREF pixel
xPix379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[3] VREF PIX_IN[379] NB2 NB1 CSA_VREF pixel
xPix380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[3] VREF PIX_IN[380] NB2 NB1 CSA_VREF pixel
xPix381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[3] VREF PIX_IN[381] NB2 NB1 CSA_VREF pixel
xPix382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[3] VREF PIX_IN[382] NB2 NB1 CSA_VREF pixel
xPix383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[3] VREF PIX_IN[383] NB2 NB1 CSA_VREF pixel
xPix384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[3] VREF PIX_IN[384] NB2 NB1 CSA_VREF pixel
xPix385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[3] VREF PIX_IN[385] NB2 NB1 CSA_VREF pixel
xPix386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[3] VREF PIX_IN[386] NB2 NB1 CSA_VREF pixel
xPix387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[3] VREF PIX_IN[387] NB2 NB1 CSA_VREF pixel
xPix388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[3] VREF PIX_IN[388] NB2 NB1 CSA_VREF pixel
xPix389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[3] VREF PIX_IN[389] NB2 NB1 CSA_VREF pixel
xPix390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[3] VREF PIX_IN[390] NB2 NB1 CSA_VREF pixel
xPix391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[3] VREF PIX_IN[391] NB2 NB1 CSA_VREF pixel
xPix392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[3] VREF PIX_IN[392] NB2 NB1 CSA_VREF pixel
xPix393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[3] VREF PIX_IN[393] NB2 NB1 CSA_VREF pixel
xPix394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[3] VREF PIX_IN[394] NB2 NB1 CSA_VREF pixel
xPix395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[3] VREF PIX_IN[395] NB2 NB1 CSA_VREF pixel
xPix396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[3] VREF PIX_IN[396] NB2 NB1 CSA_VREF pixel
xPix397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[3] VREF PIX_IN[397] NB2 NB1 CSA_VREF pixel
xPix398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[3] VREF PIX_IN[398] NB2 NB1 CSA_VREF pixel
xPix399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[3] VREF PIX_IN[399] NB2 NB1 CSA_VREF pixel
xPix400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[4] VREF PIX_IN[400] NB2 NB1 CSA_VREF pixel
xPix401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[4] VREF PIX_IN[401] NB2 NB1 CSA_VREF pixel
xPix402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[4] VREF PIX_IN[402] NB2 NB1 CSA_VREF pixel
xPix403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[4] VREF PIX_IN[403] NB2 NB1 CSA_VREF pixel
xPix404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[4] VREF PIX_IN[404] NB2 NB1 CSA_VREF pixel
xPix405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[4] VREF PIX_IN[405] NB2 NB1 CSA_VREF pixel
xPix406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[4] VREF PIX_IN[406] NB2 NB1 CSA_VREF pixel
xPix407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[4] VREF PIX_IN[407] NB2 NB1 CSA_VREF pixel
xPix408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[4] VREF PIX_IN[408] NB2 NB1 CSA_VREF pixel
xPix409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[4] VREF PIX_IN[409] NB2 NB1 CSA_VREF pixel
xPix410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[4] VREF PIX_IN[410] NB2 NB1 CSA_VREF pixel
xPix411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[4] VREF PIX_IN[411] NB2 NB1 CSA_VREF pixel
xPix412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[4] VREF PIX_IN[412] NB2 NB1 CSA_VREF pixel
xPix413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[4] VREF PIX_IN[413] NB2 NB1 CSA_VREF pixel
xPix414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[4] VREF PIX_IN[414] NB2 NB1 CSA_VREF pixel
xPix415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[4] VREF PIX_IN[415] NB2 NB1 CSA_VREF pixel
xPix416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[4] VREF PIX_IN[416] NB2 NB1 CSA_VREF pixel
xPix417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[4] VREF PIX_IN[417] NB2 NB1 CSA_VREF pixel
xPix418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[4] VREF PIX_IN[418] NB2 NB1 CSA_VREF pixel
xPix419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[4] VREF PIX_IN[419] NB2 NB1 CSA_VREF pixel
xPix420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[4] VREF PIX_IN[420] NB2 NB1 CSA_VREF pixel
xPix421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[4] VREF PIX_IN[421] NB2 NB1 CSA_VREF pixel
xPix422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[4] VREF PIX_IN[422] NB2 NB1 CSA_VREF pixel
xPix423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[4] VREF PIX_IN[423] NB2 NB1 CSA_VREF pixel
xPix424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[4] VREF PIX_IN[424] NB2 NB1 CSA_VREF pixel
xPix425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[4] VREF PIX_IN[425] NB2 NB1 CSA_VREF pixel
xPix426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[4] VREF PIX_IN[426] NB2 NB1 CSA_VREF pixel
xPix427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[4] VREF PIX_IN[427] NB2 NB1 CSA_VREF pixel
xPix428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[4] VREF PIX_IN[428] NB2 NB1 CSA_VREF pixel
xPix429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[4] VREF PIX_IN[429] NB2 NB1 CSA_VREF pixel
xPix430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[4] VREF PIX_IN[430] NB2 NB1 CSA_VREF pixel
xPix431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[4] VREF PIX_IN[431] NB2 NB1 CSA_VREF pixel
xPix432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[4] VREF PIX_IN[432] NB2 NB1 CSA_VREF pixel
xPix433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[4] VREF PIX_IN[433] NB2 NB1 CSA_VREF pixel
xPix434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[4] VREF PIX_IN[434] NB2 NB1 CSA_VREF pixel
xPix435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[4] VREF PIX_IN[435] NB2 NB1 CSA_VREF pixel
xPix436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[4] VREF PIX_IN[436] NB2 NB1 CSA_VREF pixel
xPix437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[4] VREF PIX_IN[437] NB2 NB1 CSA_VREF pixel
xPix438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[4] VREF PIX_IN[438] NB2 NB1 CSA_VREF pixel
xPix439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[4] VREF PIX_IN[439] NB2 NB1 CSA_VREF pixel
xPix440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[4] VREF PIX_IN[440] NB2 NB1 CSA_VREF pixel
xPix441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[4] VREF PIX_IN[441] NB2 NB1 CSA_VREF pixel
xPix442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[4] VREF PIX_IN[442] NB2 NB1 CSA_VREF pixel
xPix443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[4] VREF PIX_IN[443] NB2 NB1 CSA_VREF pixel
xPix444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[4] VREF PIX_IN[444] NB2 NB1 CSA_VREF pixel
xPix445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[4] VREF PIX_IN[445] NB2 NB1 CSA_VREF pixel
xPix446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[4] VREF PIX_IN[446] NB2 NB1 CSA_VREF pixel
xPix447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[4] VREF PIX_IN[447] NB2 NB1 CSA_VREF pixel
xPix448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[4] VREF PIX_IN[448] NB2 NB1 CSA_VREF pixel
xPix449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[4] VREF PIX_IN[449] NB2 NB1 CSA_VREF pixel
xPix450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[4] VREF PIX_IN[450] NB2 NB1 CSA_VREF pixel
xPix451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[4] VREF PIX_IN[451] NB2 NB1 CSA_VREF pixel
xPix452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[4] VREF PIX_IN[452] NB2 NB1 CSA_VREF pixel
xPix453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[4] VREF PIX_IN[453] NB2 NB1 CSA_VREF pixel
xPix454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[4] VREF PIX_IN[454] NB2 NB1 CSA_VREF pixel
xPix455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[4] VREF PIX_IN[455] NB2 NB1 CSA_VREF pixel
xPix456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[4] VREF PIX_IN[456] NB2 NB1 CSA_VREF pixel
xPix457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[4] VREF PIX_IN[457] NB2 NB1 CSA_VREF pixel
xPix458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[4] VREF PIX_IN[458] NB2 NB1 CSA_VREF pixel
xPix459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[4] VREF PIX_IN[459] NB2 NB1 CSA_VREF pixel
xPix460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[4] VREF PIX_IN[460] NB2 NB1 CSA_VREF pixel
xPix461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[4] VREF PIX_IN[461] NB2 NB1 CSA_VREF pixel
xPix462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[4] VREF PIX_IN[462] NB2 NB1 CSA_VREF pixel
xPix463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[4] VREF PIX_IN[463] NB2 NB1 CSA_VREF pixel
xPix464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[4] VREF PIX_IN[464] NB2 NB1 CSA_VREF pixel
xPix465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[4] VREF PIX_IN[465] NB2 NB1 CSA_VREF pixel
xPix466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[4] VREF PIX_IN[466] NB2 NB1 CSA_VREF pixel
xPix467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[4] VREF PIX_IN[467] NB2 NB1 CSA_VREF pixel
xPix468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[4] VREF PIX_IN[468] NB2 NB1 CSA_VREF pixel
xPix469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[4] VREF PIX_IN[469] NB2 NB1 CSA_VREF pixel
xPix470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[4] VREF PIX_IN[470] NB2 NB1 CSA_VREF pixel
xPix471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[4] VREF PIX_IN[471] NB2 NB1 CSA_VREF pixel
xPix472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[4] VREF PIX_IN[472] NB2 NB1 CSA_VREF pixel
xPix473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[4] VREF PIX_IN[473] NB2 NB1 CSA_VREF pixel
xPix474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[4] VREF PIX_IN[474] NB2 NB1 CSA_VREF pixel
xPix475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[4] VREF PIX_IN[475] NB2 NB1 CSA_VREF pixel
xPix476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[4] VREF PIX_IN[476] NB2 NB1 CSA_VREF pixel
xPix477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[4] VREF PIX_IN[477] NB2 NB1 CSA_VREF pixel
xPix478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[4] VREF PIX_IN[478] NB2 NB1 CSA_VREF pixel
xPix479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[4] VREF PIX_IN[479] NB2 NB1 CSA_VREF pixel
xPix480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[4] VREF PIX_IN[480] NB2 NB1 CSA_VREF pixel
xPix481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[4] VREF PIX_IN[481] NB2 NB1 CSA_VREF pixel
xPix482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[4] VREF PIX_IN[482] NB2 NB1 CSA_VREF pixel
xPix483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[4] VREF PIX_IN[483] NB2 NB1 CSA_VREF pixel
xPix484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[4] VREF PIX_IN[484] NB2 NB1 CSA_VREF pixel
xPix485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[4] VREF PIX_IN[485] NB2 NB1 CSA_VREF pixel
xPix486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[4] VREF PIX_IN[486] NB2 NB1 CSA_VREF pixel
xPix487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[4] VREF PIX_IN[487] NB2 NB1 CSA_VREF pixel
xPix488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[4] VREF PIX_IN[488] NB2 NB1 CSA_VREF pixel
xPix489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[4] VREF PIX_IN[489] NB2 NB1 CSA_VREF pixel
xPix490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[4] VREF PIX_IN[490] NB2 NB1 CSA_VREF pixel
xPix491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[4] VREF PIX_IN[491] NB2 NB1 CSA_VREF pixel
xPix492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[4] VREF PIX_IN[492] NB2 NB1 CSA_VREF pixel
xPix493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[4] VREF PIX_IN[493] NB2 NB1 CSA_VREF pixel
xPix494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[4] VREF PIX_IN[494] NB2 NB1 CSA_VREF pixel
xPix495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[4] VREF PIX_IN[495] NB2 NB1 CSA_VREF pixel
xPix496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[4] VREF PIX_IN[496] NB2 NB1 CSA_VREF pixel
xPix497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[4] VREF PIX_IN[497] NB2 NB1 CSA_VREF pixel
xPix498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[4] VREF PIX_IN[498] NB2 NB1 CSA_VREF pixel
xPix499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[4] VREF PIX_IN[499] NB2 NB1 CSA_VREF pixel
xPix500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[5] VREF PIX_IN[500] NB2 NB1 CSA_VREF pixel
xPix501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[5] VREF PIX_IN[501] NB2 NB1 CSA_VREF pixel
xPix502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[5] VREF PIX_IN[502] NB2 NB1 CSA_VREF pixel
xPix503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[5] VREF PIX_IN[503] NB2 NB1 CSA_VREF pixel
xPix504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[5] VREF PIX_IN[504] NB2 NB1 CSA_VREF pixel
xPix505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[5] VREF PIX_IN[505] NB2 NB1 CSA_VREF pixel
xPix506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[5] VREF PIX_IN[506] NB2 NB1 CSA_VREF pixel
xPix507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[5] VREF PIX_IN[507] NB2 NB1 CSA_VREF pixel
xPix508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[5] VREF PIX_IN[508] NB2 NB1 CSA_VREF pixel
xPix509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[5] VREF PIX_IN[509] NB2 NB1 CSA_VREF pixel
xPix510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[5] VREF PIX_IN[510] NB2 NB1 CSA_VREF pixel
xPix511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[5] VREF PIX_IN[511] NB2 NB1 CSA_VREF pixel
xPix512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[5] VREF PIX_IN[512] NB2 NB1 CSA_VREF pixel
xPix513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[5] VREF PIX_IN[513] NB2 NB1 CSA_VREF pixel
xPix514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[5] VREF PIX_IN[514] NB2 NB1 CSA_VREF pixel
xPix515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[5] VREF PIX_IN[515] NB2 NB1 CSA_VREF pixel
xPix516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[5] VREF PIX_IN[516] NB2 NB1 CSA_VREF pixel
xPix517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[5] VREF PIX_IN[517] NB2 NB1 CSA_VREF pixel
xPix518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[5] VREF PIX_IN[518] NB2 NB1 CSA_VREF pixel
xPix519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[5] VREF PIX_IN[519] NB2 NB1 CSA_VREF pixel
xPix520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[5] VREF PIX_IN[520] NB2 NB1 CSA_VREF pixel
xPix521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[5] VREF PIX_IN[521] NB2 NB1 CSA_VREF pixel
xPix522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[5] VREF PIX_IN[522] NB2 NB1 CSA_VREF pixel
xPix523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[5] VREF PIX_IN[523] NB2 NB1 CSA_VREF pixel
xPix524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[5] VREF PIX_IN[524] NB2 NB1 CSA_VREF pixel
xPix525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[5] VREF PIX_IN[525] NB2 NB1 CSA_VREF pixel
xPix526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[5] VREF PIX_IN[526] NB2 NB1 CSA_VREF pixel
xPix527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[5] VREF PIX_IN[527] NB2 NB1 CSA_VREF pixel
xPix528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[5] VREF PIX_IN[528] NB2 NB1 CSA_VREF pixel
xPix529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[5] VREF PIX_IN[529] NB2 NB1 CSA_VREF pixel
xPix530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[5] VREF PIX_IN[530] NB2 NB1 CSA_VREF pixel
xPix531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[5] VREF PIX_IN[531] NB2 NB1 CSA_VREF pixel
xPix532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[5] VREF PIX_IN[532] NB2 NB1 CSA_VREF pixel
xPix533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[5] VREF PIX_IN[533] NB2 NB1 CSA_VREF pixel
xPix534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[5] VREF PIX_IN[534] NB2 NB1 CSA_VREF pixel
xPix535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[5] VREF PIX_IN[535] NB2 NB1 CSA_VREF pixel
xPix536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[5] VREF PIX_IN[536] NB2 NB1 CSA_VREF pixel
xPix537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[5] VREF PIX_IN[537] NB2 NB1 CSA_VREF pixel
xPix538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[5] VREF PIX_IN[538] NB2 NB1 CSA_VREF pixel
xPix539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[5] VREF PIX_IN[539] NB2 NB1 CSA_VREF pixel
xPix540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[5] VREF PIX_IN[540] NB2 NB1 CSA_VREF pixel
xPix541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[5] VREF PIX_IN[541] NB2 NB1 CSA_VREF pixel
xPix542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[5] VREF PIX_IN[542] NB2 NB1 CSA_VREF pixel
xPix543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[5] VREF PIX_IN[543] NB2 NB1 CSA_VREF pixel
xPix544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[5] VREF PIX_IN[544] NB2 NB1 CSA_VREF pixel
xPix545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[5] VREF PIX_IN[545] NB2 NB1 CSA_VREF pixel
xPix546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[5] VREF PIX_IN[546] NB2 NB1 CSA_VREF pixel
xPix547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[5] VREF PIX_IN[547] NB2 NB1 CSA_VREF pixel
xPix548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[5] VREF PIX_IN[548] NB2 NB1 CSA_VREF pixel
xPix549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[5] VREF PIX_IN[549] NB2 NB1 CSA_VREF pixel
xPix550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[5] VREF PIX_IN[550] NB2 NB1 CSA_VREF pixel
xPix551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[5] VREF PIX_IN[551] NB2 NB1 CSA_VREF pixel
xPix552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[5] VREF PIX_IN[552] NB2 NB1 CSA_VREF pixel
xPix553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[5] VREF PIX_IN[553] NB2 NB1 CSA_VREF pixel
xPix554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[5] VREF PIX_IN[554] NB2 NB1 CSA_VREF pixel
xPix555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[5] VREF PIX_IN[555] NB2 NB1 CSA_VREF pixel
xPix556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[5] VREF PIX_IN[556] NB2 NB1 CSA_VREF pixel
xPix557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[5] VREF PIX_IN[557] NB2 NB1 CSA_VREF pixel
xPix558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[5] VREF PIX_IN[558] NB2 NB1 CSA_VREF pixel
xPix559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[5] VREF PIX_IN[559] NB2 NB1 CSA_VREF pixel
xPix560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[5] VREF PIX_IN[560] NB2 NB1 CSA_VREF pixel
xPix561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[5] VREF PIX_IN[561] NB2 NB1 CSA_VREF pixel
xPix562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[5] VREF PIX_IN[562] NB2 NB1 CSA_VREF pixel
xPix563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[5] VREF PIX_IN[563] NB2 NB1 CSA_VREF pixel
xPix564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[5] VREF PIX_IN[564] NB2 NB1 CSA_VREF pixel
xPix565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[5] VREF PIX_IN[565] NB2 NB1 CSA_VREF pixel
xPix566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[5] VREF PIX_IN[566] NB2 NB1 CSA_VREF pixel
xPix567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[5] VREF PIX_IN[567] NB2 NB1 CSA_VREF pixel
xPix568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[5] VREF PIX_IN[568] NB2 NB1 CSA_VREF pixel
xPix569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[5] VREF PIX_IN[569] NB2 NB1 CSA_VREF pixel
xPix570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[5] VREF PIX_IN[570] NB2 NB1 CSA_VREF pixel
xPix571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[5] VREF PIX_IN[571] NB2 NB1 CSA_VREF pixel
xPix572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[5] VREF PIX_IN[572] NB2 NB1 CSA_VREF pixel
xPix573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[5] VREF PIX_IN[573] NB2 NB1 CSA_VREF pixel
xPix574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[5] VREF PIX_IN[574] NB2 NB1 CSA_VREF pixel
xPix575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[5] VREF PIX_IN[575] NB2 NB1 CSA_VREF pixel
xPix576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[5] VREF PIX_IN[576] NB2 NB1 CSA_VREF pixel
xPix577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[5] VREF PIX_IN[577] NB2 NB1 CSA_VREF pixel
xPix578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[5] VREF PIX_IN[578] NB2 NB1 CSA_VREF pixel
xPix579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[5] VREF PIX_IN[579] NB2 NB1 CSA_VREF pixel
xPix580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[5] VREF PIX_IN[580] NB2 NB1 CSA_VREF pixel
xPix581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[5] VREF PIX_IN[581] NB2 NB1 CSA_VREF pixel
xPix582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[5] VREF PIX_IN[582] NB2 NB1 CSA_VREF pixel
xPix583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[5] VREF PIX_IN[583] NB2 NB1 CSA_VREF pixel
xPix584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[5] VREF PIX_IN[584] NB2 NB1 CSA_VREF pixel
xPix585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[5] VREF PIX_IN[585] NB2 NB1 CSA_VREF pixel
xPix586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[5] VREF PIX_IN[586] NB2 NB1 CSA_VREF pixel
xPix587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[5] VREF PIX_IN[587] NB2 NB1 CSA_VREF pixel
xPix588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[5] VREF PIX_IN[588] NB2 NB1 CSA_VREF pixel
xPix589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[5] VREF PIX_IN[589] NB2 NB1 CSA_VREF pixel
xPix590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[5] VREF PIX_IN[590] NB2 NB1 CSA_VREF pixel
xPix591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[5] VREF PIX_IN[591] NB2 NB1 CSA_VREF pixel
xPix592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[5] VREF PIX_IN[592] NB2 NB1 CSA_VREF pixel
xPix593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[5] VREF PIX_IN[593] NB2 NB1 CSA_VREF pixel
xPix594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[5] VREF PIX_IN[594] NB2 NB1 CSA_VREF pixel
xPix595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[5] VREF PIX_IN[595] NB2 NB1 CSA_VREF pixel
xPix596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[5] VREF PIX_IN[596] NB2 NB1 CSA_VREF pixel
xPix597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[5] VREF PIX_IN[597] NB2 NB1 CSA_VREF pixel
xPix598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[5] VREF PIX_IN[598] NB2 NB1 CSA_VREF pixel
xPix599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[5] VREF PIX_IN[599] NB2 NB1 CSA_VREF pixel
xPix600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[6] VREF PIX_IN[600] NB2 NB1 CSA_VREF pixel
xPix601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[6] VREF PIX_IN[601] NB2 NB1 CSA_VREF pixel
xPix602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[6] VREF PIX_IN[602] NB2 NB1 CSA_VREF pixel
xPix603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[6] VREF PIX_IN[603] NB2 NB1 CSA_VREF pixel
xPix604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[6] VREF PIX_IN[604] NB2 NB1 CSA_VREF pixel
xPix605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[6] VREF PIX_IN[605] NB2 NB1 CSA_VREF pixel
xPix606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[6] VREF PIX_IN[606] NB2 NB1 CSA_VREF pixel
xPix607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[6] VREF PIX_IN[607] NB2 NB1 CSA_VREF pixel
xPix608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[6] VREF PIX_IN[608] NB2 NB1 CSA_VREF pixel
xPix609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[6] VREF PIX_IN[609] NB2 NB1 CSA_VREF pixel
xPix610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[6] VREF PIX_IN[610] NB2 NB1 CSA_VREF pixel
xPix611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[6] VREF PIX_IN[611] NB2 NB1 CSA_VREF pixel
xPix612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[6] VREF PIX_IN[612] NB2 NB1 CSA_VREF pixel
xPix613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[6] VREF PIX_IN[613] NB2 NB1 CSA_VREF pixel
xPix614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[6] VREF PIX_IN[614] NB2 NB1 CSA_VREF pixel
xPix615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[6] VREF PIX_IN[615] NB2 NB1 CSA_VREF pixel
xPix616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[6] VREF PIX_IN[616] NB2 NB1 CSA_VREF pixel
xPix617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[6] VREF PIX_IN[617] NB2 NB1 CSA_VREF pixel
xPix618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[6] VREF PIX_IN[618] NB2 NB1 CSA_VREF pixel
xPix619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[6] VREF PIX_IN[619] NB2 NB1 CSA_VREF pixel
xPix620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[6] VREF PIX_IN[620] NB2 NB1 CSA_VREF pixel
xPix621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[6] VREF PIX_IN[621] NB2 NB1 CSA_VREF pixel
xPix622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[6] VREF PIX_IN[622] NB2 NB1 CSA_VREF pixel
xPix623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[6] VREF PIX_IN[623] NB2 NB1 CSA_VREF pixel
xPix624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[6] VREF PIX_IN[624] NB2 NB1 CSA_VREF pixel
xPix625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[6] VREF PIX_IN[625] NB2 NB1 CSA_VREF pixel
xPix626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[6] VREF PIX_IN[626] NB2 NB1 CSA_VREF pixel
xPix627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[6] VREF PIX_IN[627] NB2 NB1 CSA_VREF pixel
xPix628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[6] VREF PIX_IN[628] NB2 NB1 CSA_VREF pixel
xPix629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[6] VREF PIX_IN[629] NB2 NB1 CSA_VREF pixel
xPix630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[6] VREF PIX_IN[630] NB2 NB1 CSA_VREF pixel
xPix631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[6] VREF PIX_IN[631] NB2 NB1 CSA_VREF pixel
xPix632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[6] VREF PIX_IN[632] NB2 NB1 CSA_VREF pixel
xPix633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[6] VREF PIX_IN[633] NB2 NB1 CSA_VREF pixel
xPix634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[6] VREF PIX_IN[634] NB2 NB1 CSA_VREF pixel
xPix635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[6] VREF PIX_IN[635] NB2 NB1 CSA_VREF pixel
xPix636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[6] VREF PIX_IN[636] NB2 NB1 CSA_VREF pixel
xPix637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[6] VREF PIX_IN[637] NB2 NB1 CSA_VREF pixel
xPix638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[6] VREF PIX_IN[638] NB2 NB1 CSA_VREF pixel
xPix639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[6] VREF PIX_IN[639] NB2 NB1 CSA_VREF pixel
xPix640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[6] VREF PIX_IN[640] NB2 NB1 CSA_VREF pixel
xPix641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[6] VREF PIX_IN[641] NB2 NB1 CSA_VREF pixel
xPix642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[6] VREF PIX_IN[642] NB2 NB1 CSA_VREF pixel
xPix643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[6] VREF PIX_IN[643] NB2 NB1 CSA_VREF pixel
xPix644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[6] VREF PIX_IN[644] NB2 NB1 CSA_VREF pixel
xPix645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[6] VREF PIX_IN[645] NB2 NB1 CSA_VREF pixel
xPix646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[6] VREF PIX_IN[646] NB2 NB1 CSA_VREF pixel
xPix647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[6] VREF PIX_IN[647] NB2 NB1 CSA_VREF pixel
xPix648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[6] VREF PIX_IN[648] NB2 NB1 CSA_VREF pixel
xPix649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[6] VREF PIX_IN[649] NB2 NB1 CSA_VREF pixel
xPix650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[6] VREF PIX_IN[650] NB2 NB1 CSA_VREF pixel
xPix651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[6] VREF PIX_IN[651] NB2 NB1 CSA_VREF pixel
xPix652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[6] VREF PIX_IN[652] NB2 NB1 CSA_VREF pixel
xPix653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[6] VREF PIX_IN[653] NB2 NB1 CSA_VREF pixel
xPix654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[6] VREF PIX_IN[654] NB2 NB1 CSA_VREF pixel
xPix655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[6] VREF PIX_IN[655] NB2 NB1 CSA_VREF pixel
xPix656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[6] VREF PIX_IN[656] NB2 NB1 CSA_VREF pixel
xPix657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[6] VREF PIX_IN[657] NB2 NB1 CSA_VREF pixel
xPix658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[6] VREF PIX_IN[658] NB2 NB1 CSA_VREF pixel
xPix659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[6] VREF PIX_IN[659] NB2 NB1 CSA_VREF pixel
xPix660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[6] VREF PIX_IN[660] NB2 NB1 CSA_VREF pixel
xPix661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[6] VREF PIX_IN[661] NB2 NB1 CSA_VREF pixel
xPix662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[6] VREF PIX_IN[662] NB2 NB1 CSA_VREF pixel
xPix663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[6] VREF PIX_IN[663] NB2 NB1 CSA_VREF pixel
xPix664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[6] VREF PIX_IN[664] NB2 NB1 CSA_VREF pixel
xPix665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[6] VREF PIX_IN[665] NB2 NB1 CSA_VREF pixel
xPix666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[6] VREF PIX_IN[666] NB2 NB1 CSA_VREF pixel
xPix667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[6] VREF PIX_IN[667] NB2 NB1 CSA_VREF pixel
xPix668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[6] VREF PIX_IN[668] NB2 NB1 CSA_VREF pixel
xPix669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[6] VREF PIX_IN[669] NB2 NB1 CSA_VREF pixel
xPix670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[6] VREF PIX_IN[670] NB2 NB1 CSA_VREF pixel
xPix671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[6] VREF PIX_IN[671] NB2 NB1 CSA_VREF pixel
xPix672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[6] VREF PIX_IN[672] NB2 NB1 CSA_VREF pixel
xPix673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[6] VREF PIX_IN[673] NB2 NB1 CSA_VREF pixel
xPix674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[6] VREF PIX_IN[674] NB2 NB1 CSA_VREF pixel
xPix675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[6] VREF PIX_IN[675] NB2 NB1 CSA_VREF pixel
xPix676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[6] VREF PIX_IN[676] NB2 NB1 CSA_VREF pixel
xPix677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[6] VREF PIX_IN[677] NB2 NB1 CSA_VREF pixel
xPix678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[6] VREF PIX_IN[678] NB2 NB1 CSA_VREF pixel
xPix679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[6] VREF PIX_IN[679] NB2 NB1 CSA_VREF pixel
xPix680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[6] VREF PIX_IN[680] NB2 NB1 CSA_VREF pixel
xPix681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[6] VREF PIX_IN[681] NB2 NB1 CSA_VREF pixel
xPix682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[6] VREF PIX_IN[682] NB2 NB1 CSA_VREF pixel
xPix683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[6] VREF PIX_IN[683] NB2 NB1 CSA_VREF pixel
xPix684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[6] VREF PIX_IN[684] NB2 NB1 CSA_VREF pixel
xPix685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[6] VREF PIX_IN[685] NB2 NB1 CSA_VREF pixel
xPix686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[6] VREF PIX_IN[686] NB2 NB1 CSA_VREF pixel
xPix687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[6] VREF PIX_IN[687] NB2 NB1 CSA_VREF pixel
xPix688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[6] VREF PIX_IN[688] NB2 NB1 CSA_VREF pixel
xPix689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[6] VREF PIX_IN[689] NB2 NB1 CSA_VREF pixel
xPix690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[6] VREF PIX_IN[690] NB2 NB1 CSA_VREF pixel
xPix691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[6] VREF PIX_IN[691] NB2 NB1 CSA_VREF pixel
xPix692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[6] VREF PIX_IN[692] NB2 NB1 CSA_VREF pixel
xPix693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[6] VREF PIX_IN[693] NB2 NB1 CSA_VREF pixel
xPix694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[6] VREF PIX_IN[694] NB2 NB1 CSA_VREF pixel
xPix695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[6] VREF PIX_IN[695] NB2 NB1 CSA_VREF pixel
xPix696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[6] VREF PIX_IN[696] NB2 NB1 CSA_VREF pixel
xPix697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[6] VREF PIX_IN[697] NB2 NB1 CSA_VREF pixel
xPix698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[6] VREF PIX_IN[698] NB2 NB1 CSA_VREF pixel
xPix699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[6] VREF PIX_IN[699] NB2 NB1 CSA_VREF pixel
xPix700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[7] VREF PIX_IN[700] NB2 NB1 CSA_VREF pixel
xPix701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[7] VREF PIX_IN[701] NB2 NB1 CSA_VREF pixel
xPix702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[7] VREF PIX_IN[702] NB2 NB1 CSA_VREF pixel
xPix703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[7] VREF PIX_IN[703] NB2 NB1 CSA_VREF pixel
xPix704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[7] VREF PIX_IN[704] NB2 NB1 CSA_VREF pixel
xPix705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[7] VREF PIX_IN[705] NB2 NB1 CSA_VREF pixel
xPix706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[7] VREF PIX_IN[706] NB2 NB1 CSA_VREF pixel
xPix707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[7] VREF PIX_IN[707] NB2 NB1 CSA_VREF pixel
xPix708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[7] VREF PIX_IN[708] NB2 NB1 CSA_VREF pixel
xPix709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[7] VREF PIX_IN[709] NB2 NB1 CSA_VREF pixel
xPix710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[7] VREF PIX_IN[710] NB2 NB1 CSA_VREF pixel
xPix711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[7] VREF PIX_IN[711] NB2 NB1 CSA_VREF pixel
xPix712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[7] VREF PIX_IN[712] NB2 NB1 CSA_VREF pixel
xPix713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[7] VREF PIX_IN[713] NB2 NB1 CSA_VREF pixel
xPix714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[7] VREF PIX_IN[714] NB2 NB1 CSA_VREF pixel
xPix715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[7] VREF PIX_IN[715] NB2 NB1 CSA_VREF pixel
xPix716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[7] VREF PIX_IN[716] NB2 NB1 CSA_VREF pixel
xPix717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[7] VREF PIX_IN[717] NB2 NB1 CSA_VREF pixel
xPix718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[7] VREF PIX_IN[718] NB2 NB1 CSA_VREF pixel
xPix719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[7] VREF PIX_IN[719] NB2 NB1 CSA_VREF pixel
xPix720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[7] VREF PIX_IN[720] NB2 NB1 CSA_VREF pixel
xPix721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[7] VREF PIX_IN[721] NB2 NB1 CSA_VREF pixel
xPix722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[7] VREF PIX_IN[722] NB2 NB1 CSA_VREF pixel
xPix723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[7] VREF PIX_IN[723] NB2 NB1 CSA_VREF pixel
xPix724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[7] VREF PIX_IN[724] NB2 NB1 CSA_VREF pixel
xPix725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[7] VREF PIX_IN[725] NB2 NB1 CSA_VREF pixel
xPix726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[7] VREF PIX_IN[726] NB2 NB1 CSA_VREF pixel
xPix727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[7] VREF PIX_IN[727] NB2 NB1 CSA_VREF pixel
xPix728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[7] VREF PIX_IN[728] NB2 NB1 CSA_VREF pixel
xPix729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[7] VREF PIX_IN[729] NB2 NB1 CSA_VREF pixel
xPix730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[7] VREF PIX_IN[730] NB2 NB1 CSA_VREF pixel
xPix731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[7] VREF PIX_IN[731] NB2 NB1 CSA_VREF pixel
xPix732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[7] VREF PIX_IN[732] NB2 NB1 CSA_VREF pixel
xPix733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[7] VREF PIX_IN[733] NB2 NB1 CSA_VREF pixel
xPix734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[7] VREF PIX_IN[734] NB2 NB1 CSA_VREF pixel
xPix735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[7] VREF PIX_IN[735] NB2 NB1 CSA_VREF pixel
xPix736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[7] VREF PIX_IN[736] NB2 NB1 CSA_VREF pixel
xPix737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[7] VREF PIX_IN[737] NB2 NB1 CSA_VREF pixel
xPix738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[7] VREF PIX_IN[738] NB2 NB1 CSA_VREF pixel
xPix739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[7] VREF PIX_IN[739] NB2 NB1 CSA_VREF pixel
xPix740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[7] VREF PIX_IN[740] NB2 NB1 CSA_VREF pixel
xPix741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[7] VREF PIX_IN[741] NB2 NB1 CSA_VREF pixel
xPix742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[7] VREF PIX_IN[742] NB2 NB1 CSA_VREF pixel
xPix743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[7] VREF PIX_IN[743] NB2 NB1 CSA_VREF pixel
xPix744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[7] VREF PIX_IN[744] NB2 NB1 CSA_VREF pixel
xPix745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[7] VREF PIX_IN[745] NB2 NB1 CSA_VREF pixel
xPix746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[7] VREF PIX_IN[746] NB2 NB1 CSA_VREF pixel
xPix747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[7] VREF PIX_IN[747] NB2 NB1 CSA_VREF pixel
xPix748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[7] VREF PIX_IN[748] NB2 NB1 CSA_VREF pixel
xPix749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[7] VREF PIX_IN[749] NB2 NB1 CSA_VREF pixel
xPix750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[7] VREF PIX_IN[750] NB2 NB1 CSA_VREF pixel
xPix751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[7] VREF PIX_IN[751] NB2 NB1 CSA_VREF pixel
xPix752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[7] VREF PIX_IN[752] NB2 NB1 CSA_VREF pixel
xPix753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[7] VREF PIX_IN[753] NB2 NB1 CSA_VREF pixel
xPix754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[7] VREF PIX_IN[754] NB2 NB1 CSA_VREF pixel
xPix755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[7] VREF PIX_IN[755] NB2 NB1 CSA_VREF pixel
xPix756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[7] VREF PIX_IN[756] NB2 NB1 CSA_VREF pixel
xPix757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[7] VREF PIX_IN[757] NB2 NB1 CSA_VREF pixel
xPix758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[7] VREF PIX_IN[758] NB2 NB1 CSA_VREF pixel
xPix759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[7] VREF PIX_IN[759] NB2 NB1 CSA_VREF pixel
xPix760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[7] VREF PIX_IN[760] NB2 NB1 CSA_VREF pixel
xPix761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[7] VREF PIX_IN[761] NB2 NB1 CSA_VREF pixel
xPix762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[7] VREF PIX_IN[762] NB2 NB1 CSA_VREF pixel
xPix763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[7] VREF PIX_IN[763] NB2 NB1 CSA_VREF pixel
xPix764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[7] VREF PIX_IN[764] NB2 NB1 CSA_VREF pixel
xPix765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[7] VREF PIX_IN[765] NB2 NB1 CSA_VREF pixel
xPix766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[7] VREF PIX_IN[766] NB2 NB1 CSA_VREF pixel
xPix767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[7] VREF PIX_IN[767] NB2 NB1 CSA_VREF pixel
xPix768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[7] VREF PIX_IN[768] NB2 NB1 CSA_VREF pixel
xPix769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[7] VREF PIX_IN[769] NB2 NB1 CSA_VREF pixel
xPix770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[7] VREF PIX_IN[770] NB2 NB1 CSA_VREF pixel
xPix771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[7] VREF PIX_IN[771] NB2 NB1 CSA_VREF pixel
xPix772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[7] VREF PIX_IN[772] NB2 NB1 CSA_VREF pixel
xPix773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[7] VREF PIX_IN[773] NB2 NB1 CSA_VREF pixel
xPix774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[7] VREF PIX_IN[774] NB2 NB1 CSA_VREF pixel
xPix775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[7] VREF PIX_IN[775] NB2 NB1 CSA_VREF pixel
xPix776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[7] VREF PIX_IN[776] NB2 NB1 CSA_VREF pixel
xPix777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[7] VREF PIX_IN[777] NB2 NB1 CSA_VREF pixel
xPix778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[7] VREF PIX_IN[778] NB2 NB1 CSA_VREF pixel
xPix779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[7] VREF PIX_IN[779] NB2 NB1 CSA_VREF pixel
xPix780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[7] VREF PIX_IN[780] NB2 NB1 CSA_VREF pixel
xPix781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[7] VREF PIX_IN[781] NB2 NB1 CSA_VREF pixel
xPix782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[7] VREF PIX_IN[782] NB2 NB1 CSA_VREF pixel
xPix783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[7] VREF PIX_IN[783] NB2 NB1 CSA_VREF pixel
xPix784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[7] VREF PIX_IN[784] NB2 NB1 CSA_VREF pixel
xPix785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[7] VREF PIX_IN[785] NB2 NB1 CSA_VREF pixel
xPix786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[7] VREF PIX_IN[786] NB2 NB1 CSA_VREF pixel
xPix787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[7] VREF PIX_IN[787] NB2 NB1 CSA_VREF pixel
xPix788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[7] VREF PIX_IN[788] NB2 NB1 CSA_VREF pixel
xPix789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[7] VREF PIX_IN[789] NB2 NB1 CSA_VREF pixel
xPix790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[7] VREF PIX_IN[790] NB2 NB1 CSA_VREF pixel
xPix791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[7] VREF PIX_IN[791] NB2 NB1 CSA_VREF pixel
xPix792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[7] VREF PIX_IN[792] NB2 NB1 CSA_VREF pixel
xPix793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[7] VREF PIX_IN[793] NB2 NB1 CSA_VREF pixel
xPix794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[7] VREF PIX_IN[794] NB2 NB1 CSA_VREF pixel
xPix795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[7] VREF PIX_IN[795] NB2 NB1 CSA_VREF pixel
xPix796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[7] VREF PIX_IN[796] NB2 NB1 CSA_VREF pixel
xPix797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[7] VREF PIX_IN[797] NB2 NB1 CSA_VREF pixel
xPix798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[7] VREF PIX_IN[798] NB2 NB1 CSA_VREF pixel
xPix799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[7] VREF PIX_IN[799] NB2 NB1 CSA_VREF pixel
xPix800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[8] VREF PIX_IN[800] NB2 NB1 CSA_VREF pixel
xPix801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[8] VREF PIX_IN[801] NB2 NB1 CSA_VREF pixel
xPix802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[8] VREF PIX_IN[802] NB2 NB1 CSA_VREF pixel
xPix803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[8] VREF PIX_IN[803] NB2 NB1 CSA_VREF pixel
xPix804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[8] VREF PIX_IN[804] NB2 NB1 CSA_VREF pixel
xPix805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[8] VREF PIX_IN[805] NB2 NB1 CSA_VREF pixel
xPix806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[8] VREF PIX_IN[806] NB2 NB1 CSA_VREF pixel
xPix807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[8] VREF PIX_IN[807] NB2 NB1 CSA_VREF pixel
xPix808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[8] VREF PIX_IN[808] NB2 NB1 CSA_VREF pixel
xPix809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[8] VREF PIX_IN[809] NB2 NB1 CSA_VREF pixel
xPix810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[8] VREF PIX_IN[810] NB2 NB1 CSA_VREF pixel
xPix811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[8] VREF PIX_IN[811] NB2 NB1 CSA_VREF pixel
xPix812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[8] VREF PIX_IN[812] NB2 NB1 CSA_VREF pixel
xPix813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[8] VREF PIX_IN[813] NB2 NB1 CSA_VREF pixel
xPix814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[8] VREF PIX_IN[814] NB2 NB1 CSA_VREF pixel
xPix815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[8] VREF PIX_IN[815] NB2 NB1 CSA_VREF pixel
xPix816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[8] VREF PIX_IN[816] NB2 NB1 CSA_VREF pixel
xPix817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[8] VREF PIX_IN[817] NB2 NB1 CSA_VREF pixel
xPix818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[8] VREF PIX_IN[818] NB2 NB1 CSA_VREF pixel
xPix819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[8] VREF PIX_IN[819] NB2 NB1 CSA_VREF pixel
xPix820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[8] VREF PIX_IN[820] NB2 NB1 CSA_VREF pixel
xPix821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[8] VREF PIX_IN[821] NB2 NB1 CSA_VREF pixel
xPix822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[8] VREF PIX_IN[822] NB2 NB1 CSA_VREF pixel
xPix823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[8] VREF PIX_IN[823] NB2 NB1 CSA_VREF pixel
xPix824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[8] VREF PIX_IN[824] NB2 NB1 CSA_VREF pixel
xPix825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[8] VREF PIX_IN[825] NB2 NB1 CSA_VREF pixel
xPix826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[8] VREF PIX_IN[826] NB2 NB1 CSA_VREF pixel
xPix827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[8] VREF PIX_IN[827] NB2 NB1 CSA_VREF pixel
xPix828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[8] VREF PIX_IN[828] NB2 NB1 CSA_VREF pixel
xPix829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[8] VREF PIX_IN[829] NB2 NB1 CSA_VREF pixel
xPix830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[8] VREF PIX_IN[830] NB2 NB1 CSA_VREF pixel
xPix831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[8] VREF PIX_IN[831] NB2 NB1 CSA_VREF pixel
xPix832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[8] VREF PIX_IN[832] NB2 NB1 CSA_VREF pixel
xPix833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[8] VREF PIX_IN[833] NB2 NB1 CSA_VREF pixel
xPix834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[8] VREF PIX_IN[834] NB2 NB1 CSA_VREF pixel
xPix835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[8] VREF PIX_IN[835] NB2 NB1 CSA_VREF pixel
xPix836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[8] VREF PIX_IN[836] NB2 NB1 CSA_VREF pixel
xPix837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[8] VREF PIX_IN[837] NB2 NB1 CSA_VREF pixel
xPix838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[8] VREF PIX_IN[838] NB2 NB1 CSA_VREF pixel
xPix839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[8] VREF PIX_IN[839] NB2 NB1 CSA_VREF pixel
xPix840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[8] VREF PIX_IN[840] NB2 NB1 CSA_VREF pixel
xPix841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[8] VREF PIX_IN[841] NB2 NB1 CSA_VREF pixel
xPix842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[8] VREF PIX_IN[842] NB2 NB1 CSA_VREF pixel
xPix843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[8] VREF PIX_IN[843] NB2 NB1 CSA_VREF pixel
xPix844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[8] VREF PIX_IN[844] NB2 NB1 CSA_VREF pixel
xPix845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[8] VREF PIX_IN[845] NB2 NB1 CSA_VREF pixel
xPix846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[8] VREF PIX_IN[846] NB2 NB1 CSA_VREF pixel
xPix847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[8] VREF PIX_IN[847] NB2 NB1 CSA_VREF pixel
xPix848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[8] VREF PIX_IN[848] NB2 NB1 CSA_VREF pixel
xPix849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[8] VREF PIX_IN[849] NB2 NB1 CSA_VREF pixel
xPix850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[8] VREF PIX_IN[850] NB2 NB1 CSA_VREF pixel
xPix851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[8] VREF PIX_IN[851] NB2 NB1 CSA_VREF pixel
xPix852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[8] VREF PIX_IN[852] NB2 NB1 CSA_VREF pixel
xPix853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[8] VREF PIX_IN[853] NB2 NB1 CSA_VREF pixel
xPix854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[8] VREF PIX_IN[854] NB2 NB1 CSA_VREF pixel
xPix855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[8] VREF PIX_IN[855] NB2 NB1 CSA_VREF pixel
xPix856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[8] VREF PIX_IN[856] NB2 NB1 CSA_VREF pixel
xPix857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[8] VREF PIX_IN[857] NB2 NB1 CSA_VREF pixel
xPix858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[8] VREF PIX_IN[858] NB2 NB1 CSA_VREF pixel
xPix859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[8] VREF PIX_IN[859] NB2 NB1 CSA_VREF pixel
xPix860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[8] VREF PIX_IN[860] NB2 NB1 CSA_VREF pixel
xPix861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[8] VREF PIX_IN[861] NB2 NB1 CSA_VREF pixel
xPix862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[8] VREF PIX_IN[862] NB2 NB1 CSA_VREF pixel
xPix863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[8] VREF PIX_IN[863] NB2 NB1 CSA_VREF pixel
xPix864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[8] VREF PIX_IN[864] NB2 NB1 CSA_VREF pixel
xPix865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[8] VREF PIX_IN[865] NB2 NB1 CSA_VREF pixel
xPix866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[8] VREF PIX_IN[866] NB2 NB1 CSA_VREF pixel
xPix867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[8] VREF PIX_IN[867] NB2 NB1 CSA_VREF pixel
xPix868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[8] VREF PIX_IN[868] NB2 NB1 CSA_VREF pixel
xPix869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[8] VREF PIX_IN[869] NB2 NB1 CSA_VREF pixel
xPix870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[8] VREF PIX_IN[870] NB2 NB1 CSA_VREF pixel
xPix871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[8] VREF PIX_IN[871] NB2 NB1 CSA_VREF pixel
xPix872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[8] VREF PIX_IN[872] NB2 NB1 CSA_VREF pixel
xPix873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[8] VREF PIX_IN[873] NB2 NB1 CSA_VREF pixel
xPix874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[8] VREF PIX_IN[874] NB2 NB1 CSA_VREF pixel
xPix875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[8] VREF PIX_IN[875] NB2 NB1 CSA_VREF pixel
xPix876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[8] VREF PIX_IN[876] NB2 NB1 CSA_VREF pixel
xPix877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[8] VREF PIX_IN[877] NB2 NB1 CSA_VREF pixel
xPix878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[8] VREF PIX_IN[878] NB2 NB1 CSA_VREF pixel
xPix879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[8] VREF PIX_IN[879] NB2 NB1 CSA_VREF pixel
xPix880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[8] VREF PIX_IN[880] NB2 NB1 CSA_VREF pixel
xPix881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[8] VREF PIX_IN[881] NB2 NB1 CSA_VREF pixel
xPix882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[8] VREF PIX_IN[882] NB2 NB1 CSA_VREF pixel
xPix883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[8] VREF PIX_IN[883] NB2 NB1 CSA_VREF pixel
xPix884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[8] VREF PIX_IN[884] NB2 NB1 CSA_VREF pixel
xPix885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[8] VREF PIX_IN[885] NB2 NB1 CSA_VREF pixel
xPix886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[8] VREF PIX_IN[886] NB2 NB1 CSA_VREF pixel
xPix887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[8] VREF PIX_IN[887] NB2 NB1 CSA_VREF pixel
xPix888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[8] VREF PIX_IN[888] NB2 NB1 CSA_VREF pixel
xPix889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[8] VREF PIX_IN[889] NB2 NB1 CSA_VREF pixel
xPix890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[8] VREF PIX_IN[890] NB2 NB1 CSA_VREF pixel
xPix891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[8] VREF PIX_IN[891] NB2 NB1 CSA_VREF pixel
xPix892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[8] VREF PIX_IN[892] NB2 NB1 CSA_VREF pixel
xPix893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[8] VREF PIX_IN[893] NB2 NB1 CSA_VREF pixel
xPix894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[8] VREF PIX_IN[894] NB2 NB1 CSA_VREF pixel
xPix895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[8] VREF PIX_IN[895] NB2 NB1 CSA_VREF pixel
xPix896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[8] VREF PIX_IN[896] NB2 NB1 CSA_VREF pixel
xPix897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[8] VREF PIX_IN[897] NB2 NB1 CSA_VREF pixel
xPix898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[8] VREF PIX_IN[898] NB2 NB1 CSA_VREF pixel
xPix899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[8] VREF PIX_IN[899] NB2 NB1 CSA_VREF pixel
xPix900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[9] VREF PIX_IN[900] NB2 NB1 CSA_VREF pixel
xPix901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[9] VREF PIX_IN[901] NB2 NB1 CSA_VREF pixel
xPix902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[9] VREF PIX_IN[902] NB2 NB1 CSA_VREF pixel
xPix903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[9] VREF PIX_IN[903] NB2 NB1 CSA_VREF pixel
xPix904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[9] VREF PIX_IN[904] NB2 NB1 CSA_VREF pixel
xPix905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[9] VREF PIX_IN[905] NB2 NB1 CSA_VREF pixel
xPix906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[9] VREF PIX_IN[906] NB2 NB1 CSA_VREF pixel
xPix907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[9] VREF PIX_IN[907] NB2 NB1 CSA_VREF pixel
xPix908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[9] VREF PIX_IN[908] NB2 NB1 CSA_VREF pixel
xPix909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[9] VREF PIX_IN[909] NB2 NB1 CSA_VREF pixel
xPix910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[9] VREF PIX_IN[910] NB2 NB1 CSA_VREF pixel
xPix911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[9] VREF PIX_IN[911] NB2 NB1 CSA_VREF pixel
xPix912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[9] VREF PIX_IN[912] NB2 NB1 CSA_VREF pixel
xPix913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[9] VREF PIX_IN[913] NB2 NB1 CSA_VREF pixel
xPix914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[9] VREF PIX_IN[914] NB2 NB1 CSA_VREF pixel
xPix915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[9] VREF PIX_IN[915] NB2 NB1 CSA_VREF pixel
xPix916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[9] VREF PIX_IN[916] NB2 NB1 CSA_VREF pixel
xPix917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[9] VREF PIX_IN[917] NB2 NB1 CSA_VREF pixel
xPix918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[9] VREF PIX_IN[918] NB2 NB1 CSA_VREF pixel
xPix919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[9] VREF PIX_IN[919] NB2 NB1 CSA_VREF pixel
xPix920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[9] VREF PIX_IN[920] NB2 NB1 CSA_VREF pixel
xPix921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[9] VREF PIX_IN[921] NB2 NB1 CSA_VREF pixel
xPix922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[9] VREF PIX_IN[922] NB2 NB1 CSA_VREF pixel
xPix923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[9] VREF PIX_IN[923] NB2 NB1 CSA_VREF pixel
xPix924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[9] VREF PIX_IN[924] NB2 NB1 CSA_VREF pixel
xPix925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[9] VREF PIX_IN[925] NB2 NB1 CSA_VREF pixel
xPix926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[9] VREF PIX_IN[926] NB2 NB1 CSA_VREF pixel
xPix927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[9] VREF PIX_IN[927] NB2 NB1 CSA_VREF pixel
xPix928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[9] VREF PIX_IN[928] NB2 NB1 CSA_VREF pixel
xPix929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[9] VREF PIX_IN[929] NB2 NB1 CSA_VREF pixel
xPix930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[9] VREF PIX_IN[930] NB2 NB1 CSA_VREF pixel
xPix931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[9] VREF PIX_IN[931] NB2 NB1 CSA_VREF pixel
xPix932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[9] VREF PIX_IN[932] NB2 NB1 CSA_VREF pixel
xPix933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[9] VREF PIX_IN[933] NB2 NB1 CSA_VREF pixel
xPix934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[9] VREF PIX_IN[934] NB2 NB1 CSA_VREF pixel
xPix935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[9] VREF PIX_IN[935] NB2 NB1 CSA_VREF pixel
xPix936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[9] VREF PIX_IN[936] NB2 NB1 CSA_VREF pixel
xPix937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[9] VREF PIX_IN[937] NB2 NB1 CSA_VREF pixel
xPix938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[9] VREF PIX_IN[938] NB2 NB1 CSA_VREF pixel
xPix939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[9] VREF PIX_IN[939] NB2 NB1 CSA_VREF pixel
xPix940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[9] VREF PIX_IN[940] NB2 NB1 CSA_VREF pixel
xPix941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[9] VREF PIX_IN[941] NB2 NB1 CSA_VREF pixel
xPix942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[9] VREF PIX_IN[942] NB2 NB1 CSA_VREF pixel
xPix943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[9] VREF PIX_IN[943] NB2 NB1 CSA_VREF pixel
xPix944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[9] VREF PIX_IN[944] NB2 NB1 CSA_VREF pixel
xPix945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[9] VREF PIX_IN[945] NB2 NB1 CSA_VREF pixel
xPix946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[9] VREF PIX_IN[946] NB2 NB1 CSA_VREF pixel
xPix947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[9] VREF PIX_IN[947] NB2 NB1 CSA_VREF pixel
xPix948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[9] VREF PIX_IN[948] NB2 NB1 CSA_VREF pixel
xPix949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[9] VREF PIX_IN[949] NB2 NB1 CSA_VREF pixel
xPix950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[9] VREF PIX_IN[950] NB2 NB1 CSA_VREF pixel
xPix951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[9] VREF PIX_IN[951] NB2 NB1 CSA_VREF pixel
xPix952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[9] VREF PIX_IN[952] NB2 NB1 CSA_VREF pixel
xPix953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[9] VREF PIX_IN[953] NB2 NB1 CSA_VREF pixel
xPix954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[9] VREF PIX_IN[954] NB2 NB1 CSA_VREF pixel
xPix955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[9] VREF PIX_IN[955] NB2 NB1 CSA_VREF pixel
xPix956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[9] VREF PIX_IN[956] NB2 NB1 CSA_VREF pixel
xPix957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[9] VREF PIX_IN[957] NB2 NB1 CSA_VREF pixel
xPix958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[9] VREF PIX_IN[958] NB2 NB1 CSA_VREF pixel
xPix959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[9] VREF PIX_IN[959] NB2 NB1 CSA_VREF pixel
xPix960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[9] VREF PIX_IN[960] NB2 NB1 CSA_VREF pixel
xPix961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[9] VREF PIX_IN[961] NB2 NB1 CSA_VREF pixel
xPix962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[9] VREF PIX_IN[962] NB2 NB1 CSA_VREF pixel
xPix963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[9] VREF PIX_IN[963] NB2 NB1 CSA_VREF pixel
xPix964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[9] VREF PIX_IN[964] NB2 NB1 CSA_VREF pixel
xPix965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[9] VREF PIX_IN[965] NB2 NB1 CSA_VREF pixel
xPix966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[9] VREF PIX_IN[966] NB2 NB1 CSA_VREF pixel
xPix967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[9] VREF PIX_IN[967] NB2 NB1 CSA_VREF pixel
xPix968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[9] VREF PIX_IN[968] NB2 NB1 CSA_VREF pixel
xPix969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[9] VREF PIX_IN[969] NB2 NB1 CSA_VREF pixel
xPix970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[9] VREF PIX_IN[970] NB2 NB1 CSA_VREF pixel
xPix971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[9] VREF PIX_IN[971] NB2 NB1 CSA_VREF pixel
xPix972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[9] VREF PIX_IN[972] NB2 NB1 CSA_VREF pixel
xPix973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[9] VREF PIX_IN[973] NB2 NB1 CSA_VREF pixel
xPix974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[9] VREF PIX_IN[974] NB2 NB1 CSA_VREF pixel
xPix975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[9] VREF PIX_IN[975] NB2 NB1 CSA_VREF pixel
xPix976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[9] VREF PIX_IN[976] NB2 NB1 CSA_VREF pixel
xPix977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[9] VREF PIX_IN[977] NB2 NB1 CSA_VREF pixel
xPix978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[9] VREF PIX_IN[978] NB2 NB1 CSA_VREF pixel
xPix979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[9] VREF PIX_IN[979] NB2 NB1 CSA_VREF pixel
xPix980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[9] VREF PIX_IN[980] NB2 NB1 CSA_VREF pixel
xPix981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[9] VREF PIX_IN[981] NB2 NB1 CSA_VREF pixel
xPix982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[9] VREF PIX_IN[982] NB2 NB1 CSA_VREF pixel
xPix983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[9] VREF PIX_IN[983] NB2 NB1 CSA_VREF pixel
xPix984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[9] VREF PIX_IN[984] NB2 NB1 CSA_VREF pixel
xPix985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[9] VREF PIX_IN[985] NB2 NB1 CSA_VREF pixel
xPix986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[9] VREF PIX_IN[986] NB2 NB1 CSA_VREF pixel
xPix987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[9] VREF PIX_IN[987] NB2 NB1 CSA_VREF pixel
xPix988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[9] VREF PIX_IN[988] NB2 NB1 CSA_VREF pixel
xPix989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[9] VREF PIX_IN[989] NB2 NB1 CSA_VREF pixel
xPix990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[9] VREF PIX_IN[990] NB2 NB1 CSA_VREF pixel
xPix991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[9] VREF PIX_IN[991] NB2 NB1 CSA_VREF pixel
xPix992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[9] VREF PIX_IN[992] NB2 NB1 CSA_VREF pixel
xPix993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[9] VREF PIX_IN[993] NB2 NB1 CSA_VREF pixel
xPix994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[9] VREF PIX_IN[994] NB2 NB1 CSA_VREF pixel
xPix995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[9] VREF PIX_IN[995] NB2 NB1 CSA_VREF pixel
xPix996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[9] VREF PIX_IN[996] NB2 NB1 CSA_VREF pixel
xPix997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[9] VREF PIX_IN[997] NB2 NB1 CSA_VREF pixel
xPix998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[9] VREF PIX_IN[998] NB2 NB1 CSA_VREF pixel
xPix999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[9] VREF PIX_IN[999] NB2 NB1 CSA_VREF pixel
xPix1000 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[10] VREF PIX_IN[1000] NB2 NB1 CSA_VREF pixel
xPix1001 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[10] VREF PIX_IN[1001] NB2 NB1 CSA_VREF pixel
xPix1002 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[10] VREF PIX_IN[1002] NB2 NB1 CSA_VREF pixel
xPix1003 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[10] VREF PIX_IN[1003] NB2 NB1 CSA_VREF pixel
xPix1004 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[10] VREF PIX_IN[1004] NB2 NB1 CSA_VREF pixel
xPix1005 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[10] VREF PIX_IN[1005] NB2 NB1 CSA_VREF pixel
xPix1006 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[10] VREF PIX_IN[1006] NB2 NB1 CSA_VREF pixel
xPix1007 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[10] VREF PIX_IN[1007] NB2 NB1 CSA_VREF pixel
xPix1008 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[10] VREF PIX_IN[1008] NB2 NB1 CSA_VREF pixel
xPix1009 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[10] VREF PIX_IN[1009] NB2 NB1 CSA_VREF pixel
xPix1010 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[10] VREF PIX_IN[1010] NB2 NB1 CSA_VREF pixel
xPix1011 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[10] VREF PIX_IN[1011] NB2 NB1 CSA_VREF pixel
xPix1012 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[10] VREF PIX_IN[1012] NB2 NB1 CSA_VREF pixel
xPix1013 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[10] VREF PIX_IN[1013] NB2 NB1 CSA_VREF pixel
xPix1014 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[10] VREF PIX_IN[1014] NB2 NB1 CSA_VREF pixel
xPix1015 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[10] VREF PIX_IN[1015] NB2 NB1 CSA_VREF pixel
xPix1016 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[10] VREF PIX_IN[1016] NB2 NB1 CSA_VREF pixel
xPix1017 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[10] VREF PIX_IN[1017] NB2 NB1 CSA_VREF pixel
xPix1018 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[10] VREF PIX_IN[1018] NB2 NB1 CSA_VREF pixel
xPix1019 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[10] VREF PIX_IN[1019] NB2 NB1 CSA_VREF pixel
xPix1020 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[10] VREF PIX_IN[1020] NB2 NB1 CSA_VREF pixel
xPix1021 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[10] VREF PIX_IN[1021] NB2 NB1 CSA_VREF pixel
xPix1022 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[10] VREF PIX_IN[1022] NB2 NB1 CSA_VREF pixel
xPix1023 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[10] VREF PIX_IN[1023] NB2 NB1 CSA_VREF pixel
xPix1024 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[10] VREF PIX_IN[1024] NB2 NB1 CSA_VREF pixel
xPix1025 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[10] VREF PIX_IN[1025] NB2 NB1 CSA_VREF pixel
xPix1026 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[10] VREF PIX_IN[1026] NB2 NB1 CSA_VREF pixel
xPix1027 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[10] VREF PIX_IN[1027] NB2 NB1 CSA_VREF pixel
xPix1028 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[10] VREF PIX_IN[1028] NB2 NB1 CSA_VREF pixel
xPix1029 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[10] VREF PIX_IN[1029] NB2 NB1 CSA_VREF pixel
xPix1030 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[10] VREF PIX_IN[1030] NB2 NB1 CSA_VREF pixel
xPix1031 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[10] VREF PIX_IN[1031] NB2 NB1 CSA_VREF pixel
xPix1032 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[10] VREF PIX_IN[1032] NB2 NB1 CSA_VREF pixel
xPix1033 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[10] VREF PIX_IN[1033] NB2 NB1 CSA_VREF pixel
xPix1034 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[10] VREF PIX_IN[1034] NB2 NB1 CSA_VREF pixel
xPix1035 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[10] VREF PIX_IN[1035] NB2 NB1 CSA_VREF pixel
xPix1036 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[10] VREF PIX_IN[1036] NB2 NB1 CSA_VREF pixel
xPix1037 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[10] VREF PIX_IN[1037] NB2 NB1 CSA_VREF pixel
xPix1038 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[10] VREF PIX_IN[1038] NB2 NB1 CSA_VREF pixel
xPix1039 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[10] VREF PIX_IN[1039] NB2 NB1 CSA_VREF pixel
xPix1040 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[10] VREF PIX_IN[1040] NB2 NB1 CSA_VREF pixel
xPix1041 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[10] VREF PIX_IN[1041] NB2 NB1 CSA_VREF pixel
xPix1042 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[10] VREF PIX_IN[1042] NB2 NB1 CSA_VREF pixel
xPix1043 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[10] VREF PIX_IN[1043] NB2 NB1 CSA_VREF pixel
xPix1044 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[10] VREF PIX_IN[1044] NB2 NB1 CSA_VREF pixel
xPix1045 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[10] VREF PIX_IN[1045] NB2 NB1 CSA_VREF pixel
xPix1046 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[10] VREF PIX_IN[1046] NB2 NB1 CSA_VREF pixel
xPix1047 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[10] VREF PIX_IN[1047] NB2 NB1 CSA_VREF pixel
xPix1048 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[10] VREF PIX_IN[1048] NB2 NB1 CSA_VREF pixel
xPix1049 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[10] VREF PIX_IN[1049] NB2 NB1 CSA_VREF pixel
xPix1050 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[10] VREF PIX_IN[1050] NB2 NB1 CSA_VREF pixel
xPix1051 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[10] VREF PIX_IN[1051] NB2 NB1 CSA_VREF pixel
xPix1052 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[10] VREF PIX_IN[1052] NB2 NB1 CSA_VREF pixel
xPix1053 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[10] VREF PIX_IN[1053] NB2 NB1 CSA_VREF pixel
xPix1054 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[10] VREF PIX_IN[1054] NB2 NB1 CSA_VREF pixel
xPix1055 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[10] VREF PIX_IN[1055] NB2 NB1 CSA_VREF pixel
xPix1056 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[10] VREF PIX_IN[1056] NB2 NB1 CSA_VREF pixel
xPix1057 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[10] VREF PIX_IN[1057] NB2 NB1 CSA_VREF pixel
xPix1058 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[10] VREF PIX_IN[1058] NB2 NB1 CSA_VREF pixel
xPix1059 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[10] VREF PIX_IN[1059] NB2 NB1 CSA_VREF pixel
xPix1060 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[10] VREF PIX_IN[1060] NB2 NB1 CSA_VREF pixel
xPix1061 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[10] VREF PIX_IN[1061] NB2 NB1 CSA_VREF pixel
xPix1062 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[10] VREF PIX_IN[1062] NB2 NB1 CSA_VREF pixel
xPix1063 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[10] VREF PIX_IN[1063] NB2 NB1 CSA_VREF pixel
xPix1064 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[10] VREF PIX_IN[1064] NB2 NB1 CSA_VREF pixel
xPix1065 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[10] VREF PIX_IN[1065] NB2 NB1 CSA_VREF pixel
xPix1066 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[10] VREF PIX_IN[1066] NB2 NB1 CSA_VREF pixel
xPix1067 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[10] VREF PIX_IN[1067] NB2 NB1 CSA_VREF pixel
xPix1068 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[10] VREF PIX_IN[1068] NB2 NB1 CSA_VREF pixel
xPix1069 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[10] VREF PIX_IN[1069] NB2 NB1 CSA_VREF pixel
xPix1070 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[10] VREF PIX_IN[1070] NB2 NB1 CSA_VREF pixel
xPix1071 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[10] VREF PIX_IN[1071] NB2 NB1 CSA_VREF pixel
xPix1072 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[10] VREF PIX_IN[1072] NB2 NB1 CSA_VREF pixel
xPix1073 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[10] VREF PIX_IN[1073] NB2 NB1 CSA_VREF pixel
xPix1074 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[10] VREF PIX_IN[1074] NB2 NB1 CSA_VREF pixel
xPix1075 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[10] VREF PIX_IN[1075] NB2 NB1 CSA_VREF pixel
xPix1076 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[10] VREF PIX_IN[1076] NB2 NB1 CSA_VREF pixel
xPix1077 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[10] VREF PIX_IN[1077] NB2 NB1 CSA_VREF pixel
xPix1078 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[10] VREF PIX_IN[1078] NB2 NB1 CSA_VREF pixel
xPix1079 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[10] VREF PIX_IN[1079] NB2 NB1 CSA_VREF pixel
xPix1080 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[10] VREF PIX_IN[1080] NB2 NB1 CSA_VREF pixel
xPix1081 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[10] VREF PIX_IN[1081] NB2 NB1 CSA_VREF pixel
xPix1082 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[10] VREF PIX_IN[1082] NB2 NB1 CSA_VREF pixel
xPix1083 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[10] VREF PIX_IN[1083] NB2 NB1 CSA_VREF pixel
xPix1084 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[10] VREF PIX_IN[1084] NB2 NB1 CSA_VREF pixel
xPix1085 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[10] VREF PIX_IN[1085] NB2 NB1 CSA_VREF pixel
xPix1086 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[10] VREF PIX_IN[1086] NB2 NB1 CSA_VREF pixel
xPix1087 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[10] VREF PIX_IN[1087] NB2 NB1 CSA_VREF pixel
xPix1088 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[10] VREF PIX_IN[1088] NB2 NB1 CSA_VREF pixel
xPix1089 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[10] VREF PIX_IN[1089] NB2 NB1 CSA_VREF pixel
xPix1090 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[10] VREF PIX_IN[1090] NB2 NB1 CSA_VREF pixel
xPix1091 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[10] VREF PIX_IN[1091] NB2 NB1 CSA_VREF pixel
xPix1092 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[10] VREF PIX_IN[1092] NB2 NB1 CSA_VREF pixel
xPix1093 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[10] VREF PIX_IN[1093] NB2 NB1 CSA_VREF pixel
xPix1094 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[10] VREF PIX_IN[1094] NB2 NB1 CSA_VREF pixel
xPix1095 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[10] VREF PIX_IN[1095] NB2 NB1 CSA_VREF pixel
xPix1096 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[10] VREF PIX_IN[1096] NB2 NB1 CSA_VREF pixel
xPix1097 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[10] VREF PIX_IN[1097] NB2 NB1 CSA_VREF pixel
xPix1098 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[10] VREF PIX_IN[1098] NB2 NB1 CSA_VREF pixel
xPix1099 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[10] VREF PIX_IN[1099] NB2 NB1 CSA_VREF pixel
xPix1100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[11] VREF PIX_IN[1100] NB2 NB1 CSA_VREF pixel
xPix1101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[11] VREF PIX_IN[1101] NB2 NB1 CSA_VREF pixel
xPix1102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[11] VREF PIX_IN[1102] NB2 NB1 CSA_VREF pixel
xPix1103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[11] VREF PIX_IN[1103] NB2 NB1 CSA_VREF pixel
xPix1104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[11] VREF PIX_IN[1104] NB2 NB1 CSA_VREF pixel
xPix1105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[11] VREF PIX_IN[1105] NB2 NB1 CSA_VREF pixel
xPix1106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[11] VREF PIX_IN[1106] NB2 NB1 CSA_VREF pixel
xPix1107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[11] VREF PIX_IN[1107] NB2 NB1 CSA_VREF pixel
xPix1108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[11] VREF PIX_IN[1108] NB2 NB1 CSA_VREF pixel
xPix1109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[11] VREF PIX_IN[1109] NB2 NB1 CSA_VREF pixel
xPix1110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[11] VREF PIX_IN[1110] NB2 NB1 CSA_VREF pixel
xPix1111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[11] VREF PIX_IN[1111] NB2 NB1 CSA_VREF pixel
xPix1112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[11] VREF PIX_IN[1112] NB2 NB1 CSA_VREF pixel
xPix1113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[11] VREF PIX_IN[1113] NB2 NB1 CSA_VREF pixel
xPix1114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[11] VREF PIX_IN[1114] NB2 NB1 CSA_VREF pixel
xPix1115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[11] VREF PIX_IN[1115] NB2 NB1 CSA_VREF pixel
xPix1116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[11] VREF PIX_IN[1116] NB2 NB1 CSA_VREF pixel
xPix1117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[11] VREF PIX_IN[1117] NB2 NB1 CSA_VREF pixel
xPix1118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[11] VREF PIX_IN[1118] NB2 NB1 CSA_VREF pixel
xPix1119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[11] VREF PIX_IN[1119] NB2 NB1 CSA_VREF pixel
xPix1120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[11] VREF PIX_IN[1120] NB2 NB1 CSA_VREF pixel
xPix1121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[11] VREF PIX_IN[1121] NB2 NB1 CSA_VREF pixel
xPix1122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[11] VREF PIX_IN[1122] NB2 NB1 CSA_VREF pixel
xPix1123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[11] VREF PIX_IN[1123] NB2 NB1 CSA_VREF pixel
xPix1124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[11] VREF PIX_IN[1124] NB2 NB1 CSA_VREF pixel
xPix1125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[11] VREF PIX_IN[1125] NB2 NB1 CSA_VREF pixel
xPix1126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[11] VREF PIX_IN[1126] NB2 NB1 CSA_VREF pixel
xPix1127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[11] VREF PIX_IN[1127] NB2 NB1 CSA_VREF pixel
xPix1128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[11] VREF PIX_IN[1128] NB2 NB1 CSA_VREF pixel
xPix1129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[11] VREF PIX_IN[1129] NB2 NB1 CSA_VREF pixel
xPix1130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[11] VREF PIX_IN[1130] NB2 NB1 CSA_VREF pixel
xPix1131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[11] VREF PIX_IN[1131] NB2 NB1 CSA_VREF pixel
xPix1132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[11] VREF PIX_IN[1132] NB2 NB1 CSA_VREF pixel
xPix1133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[11] VREF PIX_IN[1133] NB2 NB1 CSA_VREF pixel
xPix1134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[11] VREF PIX_IN[1134] NB2 NB1 CSA_VREF pixel
xPix1135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[11] VREF PIX_IN[1135] NB2 NB1 CSA_VREF pixel
xPix1136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[11] VREF PIX_IN[1136] NB2 NB1 CSA_VREF pixel
xPix1137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[11] VREF PIX_IN[1137] NB2 NB1 CSA_VREF pixel
xPix1138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[11] VREF PIX_IN[1138] NB2 NB1 CSA_VREF pixel
xPix1139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[11] VREF PIX_IN[1139] NB2 NB1 CSA_VREF pixel
xPix1140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[11] VREF PIX_IN[1140] NB2 NB1 CSA_VREF pixel
xPix1141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[11] VREF PIX_IN[1141] NB2 NB1 CSA_VREF pixel
xPix1142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[11] VREF PIX_IN[1142] NB2 NB1 CSA_VREF pixel
xPix1143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[11] VREF PIX_IN[1143] NB2 NB1 CSA_VREF pixel
xPix1144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[11] VREF PIX_IN[1144] NB2 NB1 CSA_VREF pixel
xPix1145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[11] VREF PIX_IN[1145] NB2 NB1 CSA_VREF pixel
xPix1146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[11] VREF PIX_IN[1146] NB2 NB1 CSA_VREF pixel
xPix1147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[11] VREF PIX_IN[1147] NB2 NB1 CSA_VREF pixel
xPix1148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[11] VREF PIX_IN[1148] NB2 NB1 CSA_VREF pixel
xPix1149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[11] VREF PIX_IN[1149] NB2 NB1 CSA_VREF pixel
xPix1150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[11] VREF PIX_IN[1150] NB2 NB1 CSA_VREF pixel
xPix1151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[11] VREF PIX_IN[1151] NB2 NB1 CSA_VREF pixel
xPix1152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[11] VREF PIX_IN[1152] NB2 NB1 CSA_VREF pixel
xPix1153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[11] VREF PIX_IN[1153] NB2 NB1 CSA_VREF pixel
xPix1154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[11] VREF PIX_IN[1154] NB2 NB1 CSA_VREF pixel
xPix1155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[11] VREF PIX_IN[1155] NB2 NB1 CSA_VREF pixel
xPix1156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[11] VREF PIX_IN[1156] NB2 NB1 CSA_VREF pixel
xPix1157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[11] VREF PIX_IN[1157] NB2 NB1 CSA_VREF pixel
xPix1158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[11] VREF PIX_IN[1158] NB2 NB1 CSA_VREF pixel
xPix1159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[11] VREF PIX_IN[1159] NB2 NB1 CSA_VREF pixel
xPix1160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[11] VREF PIX_IN[1160] NB2 NB1 CSA_VREF pixel
xPix1161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[11] VREF PIX_IN[1161] NB2 NB1 CSA_VREF pixel
xPix1162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[11] VREF PIX_IN[1162] NB2 NB1 CSA_VREF pixel
xPix1163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[11] VREF PIX_IN[1163] NB2 NB1 CSA_VREF pixel
xPix1164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[11] VREF PIX_IN[1164] NB2 NB1 CSA_VREF pixel
xPix1165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[11] VREF PIX_IN[1165] NB2 NB1 CSA_VREF pixel
xPix1166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[11] VREF PIX_IN[1166] NB2 NB1 CSA_VREF pixel
xPix1167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[11] VREF PIX_IN[1167] NB2 NB1 CSA_VREF pixel
xPix1168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[11] VREF PIX_IN[1168] NB2 NB1 CSA_VREF pixel
xPix1169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[11] VREF PIX_IN[1169] NB2 NB1 CSA_VREF pixel
xPix1170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[11] VREF PIX_IN[1170] NB2 NB1 CSA_VREF pixel
xPix1171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[11] VREF PIX_IN[1171] NB2 NB1 CSA_VREF pixel
xPix1172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[11] VREF PIX_IN[1172] NB2 NB1 CSA_VREF pixel
xPix1173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[11] VREF PIX_IN[1173] NB2 NB1 CSA_VREF pixel
xPix1174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[11] VREF PIX_IN[1174] NB2 NB1 CSA_VREF pixel
xPix1175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[11] VREF PIX_IN[1175] NB2 NB1 CSA_VREF pixel
xPix1176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[11] VREF PIX_IN[1176] NB2 NB1 CSA_VREF pixel
xPix1177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[11] VREF PIX_IN[1177] NB2 NB1 CSA_VREF pixel
xPix1178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[11] VREF PIX_IN[1178] NB2 NB1 CSA_VREF pixel
xPix1179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[11] VREF PIX_IN[1179] NB2 NB1 CSA_VREF pixel
xPix1180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[11] VREF PIX_IN[1180] NB2 NB1 CSA_VREF pixel
xPix1181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[11] VREF PIX_IN[1181] NB2 NB1 CSA_VREF pixel
xPix1182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[11] VREF PIX_IN[1182] NB2 NB1 CSA_VREF pixel
xPix1183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[11] VREF PIX_IN[1183] NB2 NB1 CSA_VREF pixel
xPix1184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[11] VREF PIX_IN[1184] NB2 NB1 CSA_VREF pixel
xPix1185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[11] VREF PIX_IN[1185] NB2 NB1 CSA_VREF pixel
xPix1186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[11] VREF PIX_IN[1186] NB2 NB1 CSA_VREF pixel
xPix1187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[11] VREF PIX_IN[1187] NB2 NB1 CSA_VREF pixel
xPix1188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[11] VREF PIX_IN[1188] NB2 NB1 CSA_VREF pixel
xPix1189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[11] VREF PIX_IN[1189] NB2 NB1 CSA_VREF pixel
xPix1190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[11] VREF PIX_IN[1190] NB2 NB1 CSA_VREF pixel
xPix1191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[11] VREF PIX_IN[1191] NB2 NB1 CSA_VREF pixel
xPix1192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[11] VREF PIX_IN[1192] NB2 NB1 CSA_VREF pixel
xPix1193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[11] VREF PIX_IN[1193] NB2 NB1 CSA_VREF pixel
xPix1194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[11] VREF PIX_IN[1194] NB2 NB1 CSA_VREF pixel
xPix1195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[11] VREF PIX_IN[1195] NB2 NB1 CSA_VREF pixel
xPix1196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[11] VREF PIX_IN[1196] NB2 NB1 CSA_VREF pixel
xPix1197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[11] VREF PIX_IN[1197] NB2 NB1 CSA_VREF pixel
xPix1198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[11] VREF PIX_IN[1198] NB2 NB1 CSA_VREF pixel
xPix1199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[11] VREF PIX_IN[1199] NB2 NB1 CSA_VREF pixel
xPix1200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[12] VREF PIX_IN[1200] NB2 NB1 CSA_VREF pixel
xPix1201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[12] VREF PIX_IN[1201] NB2 NB1 CSA_VREF pixel
xPix1202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[12] VREF PIX_IN[1202] NB2 NB1 CSA_VREF pixel
xPix1203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[12] VREF PIX_IN[1203] NB2 NB1 CSA_VREF pixel
xPix1204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[12] VREF PIX_IN[1204] NB2 NB1 CSA_VREF pixel
xPix1205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[12] VREF PIX_IN[1205] NB2 NB1 CSA_VREF pixel
xPix1206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[12] VREF PIX_IN[1206] NB2 NB1 CSA_VREF pixel
xPix1207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[12] VREF PIX_IN[1207] NB2 NB1 CSA_VREF pixel
xPix1208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[12] VREF PIX_IN[1208] NB2 NB1 CSA_VREF pixel
xPix1209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[12] VREF PIX_IN[1209] NB2 NB1 CSA_VREF pixel
xPix1210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[12] VREF PIX_IN[1210] NB2 NB1 CSA_VREF pixel
xPix1211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[12] VREF PIX_IN[1211] NB2 NB1 CSA_VREF pixel
xPix1212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[12] VREF PIX_IN[1212] NB2 NB1 CSA_VREF pixel
xPix1213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[12] VREF PIX_IN[1213] NB2 NB1 CSA_VREF pixel
xPix1214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[12] VREF PIX_IN[1214] NB2 NB1 CSA_VREF pixel
xPix1215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[12] VREF PIX_IN[1215] NB2 NB1 CSA_VREF pixel
xPix1216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[12] VREF PIX_IN[1216] NB2 NB1 CSA_VREF pixel
xPix1217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[12] VREF PIX_IN[1217] NB2 NB1 CSA_VREF pixel
xPix1218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[12] VREF PIX_IN[1218] NB2 NB1 CSA_VREF pixel
xPix1219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[12] VREF PIX_IN[1219] NB2 NB1 CSA_VREF pixel
xPix1220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[12] VREF PIX_IN[1220] NB2 NB1 CSA_VREF pixel
xPix1221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[12] VREF PIX_IN[1221] NB2 NB1 CSA_VREF pixel
xPix1222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[12] VREF PIX_IN[1222] NB2 NB1 CSA_VREF pixel
xPix1223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[12] VREF PIX_IN[1223] NB2 NB1 CSA_VREF pixel
xPix1224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[12] VREF PIX_IN[1224] NB2 NB1 CSA_VREF pixel
xPix1225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[12] VREF PIX_IN[1225] NB2 NB1 CSA_VREF pixel
xPix1226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[12] VREF PIX_IN[1226] NB2 NB1 CSA_VREF pixel
xPix1227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[12] VREF PIX_IN[1227] NB2 NB1 CSA_VREF pixel
xPix1228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[12] VREF PIX_IN[1228] NB2 NB1 CSA_VREF pixel
xPix1229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[12] VREF PIX_IN[1229] NB2 NB1 CSA_VREF pixel
xPix1230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[12] VREF PIX_IN[1230] NB2 NB1 CSA_VREF pixel
xPix1231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[12] VREF PIX_IN[1231] NB2 NB1 CSA_VREF pixel
xPix1232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[12] VREF PIX_IN[1232] NB2 NB1 CSA_VREF pixel
xPix1233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[12] VREF PIX_IN[1233] NB2 NB1 CSA_VREF pixel
xPix1234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[12] VREF PIX_IN[1234] NB2 NB1 CSA_VREF pixel
xPix1235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[12] VREF PIX_IN[1235] NB2 NB1 CSA_VREF pixel
xPix1236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[12] VREF PIX_IN[1236] NB2 NB1 CSA_VREF pixel
xPix1237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[12] VREF PIX_IN[1237] NB2 NB1 CSA_VREF pixel
xPix1238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[12] VREF PIX_IN[1238] NB2 NB1 CSA_VREF pixel
xPix1239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[12] VREF PIX_IN[1239] NB2 NB1 CSA_VREF pixel
xPix1240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[12] VREF PIX_IN[1240] NB2 NB1 CSA_VREF pixel
xPix1241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[12] VREF PIX_IN[1241] NB2 NB1 CSA_VREF pixel
xPix1242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[12] VREF PIX_IN[1242] NB2 NB1 CSA_VREF pixel
xPix1243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[12] VREF PIX_IN[1243] NB2 NB1 CSA_VREF pixel
xPix1244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[12] VREF PIX_IN[1244] NB2 NB1 CSA_VREF pixel
xPix1245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[12] VREF PIX_IN[1245] NB2 NB1 CSA_VREF pixel
xPix1246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[12] VREF PIX_IN[1246] NB2 NB1 CSA_VREF pixel
xPix1247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[12] VREF PIX_IN[1247] NB2 NB1 CSA_VREF pixel
xPix1248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[12] VREF PIX_IN[1248] NB2 NB1 CSA_VREF pixel
xPix1249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[12] VREF PIX_IN[1249] NB2 NB1 CSA_VREF pixel
xPix1250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[12] VREF PIX_IN[1250] NB2 NB1 CSA_VREF pixel
xPix1251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[12] VREF PIX_IN[1251] NB2 NB1 CSA_VREF pixel
xPix1252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[12] VREF PIX_IN[1252] NB2 NB1 CSA_VREF pixel
xPix1253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[12] VREF PIX_IN[1253] NB2 NB1 CSA_VREF pixel
xPix1254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[12] VREF PIX_IN[1254] NB2 NB1 CSA_VREF pixel
xPix1255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[12] VREF PIX_IN[1255] NB2 NB1 CSA_VREF pixel
xPix1256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[12] VREF PIX_IN[1256] NB2 NB1 CSA_VREF pixel
xPix1257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[12] VREF PIX_IN[1257] NB2 NB1 CSA_VREF pixel
xPix1258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[12] VREF PIX_IN[1258] NB2 NB1 CSA_VREF pixel
xPix1259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[12] VREF PIX_IN[1259] NB2 NB1 CSA_VREF pixel
xPix1260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[12] VREF PIX_IN[1260] NB2 NB1 CSA_VREF pixel
xPix1261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[12] VREF PIX_IN[1261] NB2 NB1 CSA_VREF pixel
xPix1262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[12] VREF PIX_IN[1262] NB2 NB1 CSA_VREF pixel
xPix1263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[12] VREF PIX_IN[1263] NB2 NB1 CSA_VREF pixel
xPix1264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[12] VREF PIX_IN[1264] NB2 NB1 CSA_VREF pixel
xPix1265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[12] VREF PIX_IN[1265] NB2 NB1 CSA_VREF pixel
xPix1266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[12] VREF PIX_IN[1266] NB2 NB1 CSA_VREF pixel
xPix1267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[12] VREF PIX_IN[1267] NB2 NB1 CSA_VREF pixel
xPix1268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[12] VREF PIX_IN[1268] NB2 NB1 CSA_VREF pixel
xPix1269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[12] VREF PIX_IN[1269] NB2 NB1 CSA_VREF pixel
xPix1270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[12] VREF PIX_IN[1270] NB2 NB1 CSA_VREF pixel
xPix1271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[12] VREF PIX_IN[1271] NB2 NB1 CSA_VREF pixel
xPix1272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[12] VREF PIX_IN[1272] NB2 NB1 CSA_VREF pixel
xPix1273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[12] VREF PIX_IN[1273] NB2 NB1 CSA_VREF pixel
xPix1274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[12] VREF PIX_IN[1274] NB2 NB1 CSA_VREF pixel
xPix1275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[12] VREF PIX_IN[1275] NB2 NB1 CSA_VREF pixel
xPix1276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[12] VREF PIX_IN[1276] NB2 NB1 CSA_VREF pixel
xPix1277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[12] VREF PIX_IN[1277] NB2 NB1 CSA_VREF pixel
xPix1278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[12] VREF PIX_IN[1278] NB2 NB1 CSA_VREF pixel
xPix1279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[12] VREF PIX_IN[1279] NB2 NB1 CSA_VREF pixel
xPix1280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[12] VREF PIX_IN[1280] NB2 NB1 CSA_VREF pixel
xPix1281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[12] VREF PIX_IN[1281] NB2 NB1 CSA_VREF pixel
xPix1282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[12] VREF PIX_IN[1282] NB2 NB1 CSA_VREF pixel
xPix1283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[12] VREF PIX_IN[1283] NB2 NB1 CSA_VREF pixel
xPix1284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[12] VREF PIX_IN[1284] NB2 NB1 CSA_VREF pixel
xPix1285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[12] VREF PIX_IN[1285] NB2 NB1 CSA_VREF pixel
xPix1286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[12] VREF PIX_IN[1286] NB2 NB1 CSA_VREF pixel
xPix1287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[12] VREF PIX_IN[1287] NB2 NB1 CSA_VREF pixel
xPix1288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[12] VREF PIX_IN[1288] NB2 NB1 CSA_VREF pixel
xPix1289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[12] VREF PIX_IN[1289] NB2 NB1 CSA_VREF pixel
xPix1290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[12] VREF PIX_IN[1290] NB2 NB1 CSA_VREF pixel
xPix1291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[12] VREF PIX_IN[1291] NB2 NB1 CSA_VREF pixel
xPix1292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[12] VREF PIX_IN[1292] NB2 NB1 CSA_VREF pixel
xPix1293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[12] VREF PIX_IN[1293] NB2 NB1 CSA_VREF pixel
xPix1294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[12] VREF PIX_IN[1294] NB2 NB1 CSA_VREF pixel
xPix1295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[12] VREF PIX_IN[1295] NB2 NB1 CSA_VREF pixel
xPix1296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[12] VREF PIX_IN[1296] NB2 NB1 CSA_VREF pixel
xPix1297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[12] VREF PIX_IN[1297] NB2 NB1 CSA_VREF pixel
xPix1298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[12] VREF PIX_IN[1298] NB2 NB1 CSA_VREF pixel
xPix1299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[12] VREF PIX_IN[1299] NB2 NB1 CSA_VREF pixel
xPix1300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[13] VREF PIX_IN[1300] NB2 NB1 CSA_VREF pixel
xPix1301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[13] VREF PIX_IN[1301] NB2 NB1 CSA_VREF pixel
xPix1302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[13] VREF PIX_IN[1302] NB2 NB1 CSA_VREF pixel
xPix1303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[13] VREF PIX_IN[1303] NB2 NB1 CSA_VREF pixel
xPix1304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[13] VREF PIX_IN[1304] NB2 NB1 CSA_VREF pixel
xPix1305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[13] VREF PIX_IN[1305] NB2 NB1 CSA_VREF pixel
xPix1306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[13] VREF PIX_IN[1306] NB2 NB1 CSA_VREF pixel
xPix1307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[13] VREF PIX_IN[1307] NB2 NB1 CSA_VREF pixel
xPix1308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[13] VREF PIX_IN[1308] NB2 NB1 CSA_VREF pixel
xPix1309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[13] VREF PIX_IN[1309] NB2 NB1 CSA_VREF pixel
xPix1310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[13] VREF PIX_IN[1310] NB2 NB1 CSA_VREF pixel
xPix1311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[13] VREF PIX_IN[1311] NB2 NB1 CSA_VREF pixel
xPix1312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[13] VREF PIX_IN[1312] NB2 NB1 CSA_VREF pixel
xPix1313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[13] VREF PIX_IN[1313] NB2 NB1 CSA_VREF pixel
xPix1314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[13] VREF PIX_IN[1314] NB2 NB1 CSA_VREF pixel
xPix1315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[13] VREF PIX_IN[1315] NB2 NB1 CSA_VREF pixel
xPix1316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[13] VREF PIX_IN[1316] NB2 NB1 CSA_VREF pixel
xPix1317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[13] VREF PIX_IN[1317] NB2 NB1 CSA_VREF pixel
xPix1318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[13] VREF PIX_IN[1318] NB2 NB1 CSA_VREF pixel
xPix1319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[13] VREF PIX_IN[1319] NB2 NB1 CSA_VREF pixel
xPix1320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[13] VREF PIX_IN[1320] NB2 NB1 CSA_VREF pixel
xPix1321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[13] VREF PIX_IN[1321] NB2 NB1 CSA_VREF pixel
xPix1322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[13] VREF PIX_IN[1322] NB2 NB1 CSA_VREF pixel
xPix1323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[13] VREF PIX_IN[1323] NB2 NB1 CSA_VREF pixel
xPix1324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[13] VREF PIX_IN[1324] NB2 NB1 CSA_VREF pixel
xPix1325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[13] VREF PIX_IN[1325] NB2 NB1 CSA_VREF pixel
xPix1326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[13] VREF PIX_IN[1326] NB2 NB1 CSA_VREF pixel
xPix1327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[13] VREF PIX_IN[1327] NB2 NB1 CSA_VREF pixel
xPix1328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[13] VREF PIX_IN[1328] NB2 NB1 CSA_VREF pixel
xPix1329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[13] VREF PIX_IN[1329] NB2 NB1 CSA_VREF pixel
xPix1330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[13] VREF PIX_IN[1330] NB2 NB1 CSA_VREF pixel
xPix1331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[13] VREF PIX_IN[1331] NB2 NB1 CSA_VREF pixel
xPix1332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[13] VREF PIX_IN[1332] NB2 NB1 CSA_VREF pixel
xPix1333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[13] VREF PIX_IN[1333] NB2 NB1 CSA_VREF pixel
xPix1334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[13] VREF PIX_IN[1334] NB2 NB1 CSA_VREF pixel
xPix1335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[13] VREF PIX_IN[1335] NB2 NB1 CSA_VREF pixel
xPix1336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[13] VREF PIX_IN[1336] NB2 NB1 CSA_VREF pixel
xPix1337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[13] VREF PIX_IN[1337] NB2 NB1 CSA_VREF pixel
xPix1338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[13] VREF PIX_IN[1338] NB2 NB1 CSA_VREF pixel
xPix1339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[13] VREF PIX_IN[1339] NB2 NB1 CSA_VREF pixel
xPix1340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[13] VREF PIX_IN[1340] NB2 NB1 CSA_VREF pixel
xPix1341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[13] VREF PIX_IN[1341] NB2 NB1 CSA_VREF pixel
xPix1342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[13] VREF PIX_IN[1342] NB2 NB1 CSA_VREF pixel
xPix1343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[13] VREF PIX_IN[1343] NB2 NB1 CSA_VREF pixel
xPix1344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[13] VREF PIX_IN[1344] NB2 NB1 CSA_VREF pixel
xPix1345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[13] VREF PIX_IN[1345] NB2 NB1 CSA_VREF pixel
xPix1346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[13] VREF PIX_IN[1346] NB2 NB1 CSA_VREF pixel
xPix1347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[13] VREF PIX_IN[1347] NB2 NB1 CSA_VREF pixel
xPix1348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[13] VREF PIX_IN[1348] NB2 NB1 CSA_VREF pixel
xPix1349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[13] VREF PIX_IN[1349] NB2 NB1 CSA_VREF pixel
xPix1350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[13] VREF PIX_IN[1350] NB2 NB1 CSA_VREF pixel
xPix1351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[13] VREF PIX_IN[1351] NB2 NB1 CSA_VREF pixel
xPix1352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[13] VREF PIX_IN[1352] NB2 NB1 CSA_VREF pixel
xPix1353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[13] VREF PIX_IN[1353] NB2 NB1 CSA_VREF pixel
xPix1354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[13] VREF PIX_IN[1354] NB2 NB1 CSA_VREF pixel
xPix1355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[13] VREF PIX_IN[1355] NB2 NB1 CSA_VREF pixel
xPix1356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[13] VREF PIX_IN[1356] NB2 NB1 CSA_VREF pixel
xPix1357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[13] VREF PIX_IN[1357] NB2 NB1 CSA_VREF pixel
xPix1358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[13] VREF PIX_IN[1358] NB2 NB1 CSA_VREF pixel
xPix1359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[13] VREF PIX_IN[1359] NB2 NB1 CSA_VREF pixel
xPix1360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[13] VREF PIX_IN[1360] NB2 NB1 CSA_VREF pixel
xPix1361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[13] VREF PIX_IN[1361] NB2 NB1 CSA_VREF pixel
xPix1362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[13] VREF PIX_IN[1362] NB2 NB1 CSA_VREF pixel
xPix1363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[13] VREF PIX_IN[1363] NB2 NB1 CSA_VREF pixel
xPix1364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[13] VREF PIX_IN[1364] NB2 NB1 CSA_VREF pixel
xPix1365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[13] VREF PIX_IN[1365] NB2 NB1 CSA_VREF pixel
xPix1366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[13] VREF PIX_IN[1366] NB2 NB1 CSA_VREF pixel
xPix1367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[13] VREF PIX_IN[1367] NB2 NB1 CSA_VREF pixel
xPix1368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[13] VREF PIX_IN[1368] NB2 NB1 CSA_VREF pixel
xPix1369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[13] VREF PIX_IN[1369] NB2 NB1 CSA_VREF pixel
xPix1370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[13] VREF PIX_IN[1370] NB2 NB1 CSA_VREF pixel
xPix1371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[13] VREF PIX_IN[1371] NB2 NB1 CSA_VREF pixel
xPix1372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[13] VREF PIX_IN[1372] NB2 NB1 CSA_VREF pixel
xPix1373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[13] VREF PIX_IN[1373] NB2 NB1 CSA_VREF pixel
xPix1374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[13] VREF PIX_IN[1374] NB2 NB1 CSA_VREF pixel
xPix1375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[13] VREF PIX_IN[1375] NB2 NB1 CSA_VREF pixel
xPix1376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[13] VREF PIX_IN[1376] NB2 NB1 CSA_VREF pixel
xPix1377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[13] VREF PIX_IN[1377] NB2 NB1 CSA_VREF pixel
xPix1378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[13] VREF PIX_IN[1378] NB2 NB1 CSA_VREF pixel
xPix1379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[13] VREF PIX_IN[1379] NB2 NB1 CSA_VREF pixel
xPix1380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[13] VREF PIX_IN[1380] NB2 NB1 CSA_VREF pixel
xPix1381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[13] VREF PIX_IN[1381] NB2 NB1 CSA_VREF pixel
xPix1382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[13] VREF PIX_IN[1382] NB2 NB1 CSA_VREF pixel
xPix1383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[13] VREF PIX_IN[1383] NB2 NB1 CSA_VREF pixel
xPix1384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[13] VREF PIX_IN[1384] NB2 NB1 CSA_VREF pixel
xPix1385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[13] VREF PIX_IN[1385] NB2 NB1 CSA_VREF pixel
xPix1386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[13] VREF PIX_IN[1386] NB2 NB1 CSA_VREF pixel
xPix1387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[13] VREF PIX_IN[1387] NB2 NB1 CSA_VREF pixel
xPix1388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[13] VREF PIX_IN[1388] NB2 NB1 CSA_VREF pixel
xPix1389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[13] VREF PIX_IN[1389] NB2 NB1 CSA_VREF pixel
xPix1390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[13] VREF PIX_IN[1390] NB2 NB1 CSA_VREF pixel
xPix1391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[13] VREF PIX_IN[1391] NB2 NB1 CSA_VREF pixel
xPix1392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[13] VREF PIX_IN[1392] NB2 NB1 CSA_VREF pixel
xPix1393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[13] VREF PIX_IN[1393] NB2 NB1 CSA_VREF pixel
xPix1394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[13] VREF PIX_IN[1394] NB2 NB1 CSA_VREF pixel
xPix1395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[13] VREF PIX_IN[1395] NB2 NB1 CSA_VREF pixel
xPix1396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[13] VREF PIX_IN[1396] NB2 NB1 CSA_VREF pixel
xPix1397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[13] VREF PIX_IN[1397] NB2 NB1 CSA_VREF pixel
xPix1398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[13] VREF PIX_IN[1398] NB2 NB1 CSA_VREF pixel
xPix1399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[13] VREF PIX_IN[1399] NB2 NB1 CSA_VREF pixel
xPix1400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[14] VREF PIX_IN[1400] NB2 NB1 CSA_VREF pixel
xPix1401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[14] VREF PIX_IN[1401] NB2 NB1 CSA_VREF pixel
xPix1402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[14] VREF PIX_IN[1402] NB2 NB1 CSA_VREF pixel
xPix1403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[14] VREF PIX_IN[1403] NB2 NB1 CSA_VREF pixel
xPix1404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[14] VREF PIX_IN[1404] NB2 NB1 CSA_VREF pixel
xPix1405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[14] VREF PIX_IN[1405] NB2 NB1 CSA_VREF pixel
xPix1406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[14] VREF PIX_IN[1406] NB2 NB1 CSA_VREF pixel
xPix1407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[14] VREF PIX_IN[1407] NB2 NB1 CSA_VREF pixel
xPix1408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[14] VREF PIX_IN[1408] NB2 NB1 CSA_VREF pixel
xPix1409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[14] VREF PIX_IN[1409] NB2 NB1 CSA_VREF pixel
xPix1410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[14] VREF PIX_IN[1410] NB2 NB1 CSA_VREF pixel
xPix1411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[14] VREF PIX_IN[1411] NB2 NB1 CSA_VREF pixel
xPix1412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[14] VREF PIX_IN[1412] NB2 NB1 CSA_VREF pixel
xPix1413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[14] VREF PIX_IN[1413] NB2 NB1 CSA_VREF pixel
xPix1414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[14] VREF PIX_IN[1414] NB2 NB1 CSA_VREF pixel
xPix1415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[14] VREF PIX_IN[1415] NB2 NB1 CSA_VREF pixel
xPix1416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[14] VREF PIX_IN[1416] NB2 NB1 CSA_VREF pixel
xPix1417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[14] VREF PIX_IN[1417] NB2 NB1 CSA_VREF pixel
xPix1418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[14] VREF PIX_IN[1418] NB2 NB1 CSA_VREF pixel
xPix1419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[14] VREF PIX_IN[1419] NB2 NB1 CSA_VREF pixel
xPix1420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[14] VREF PIX_IN[1420] NB2 NB1 CSA_VREF pixel
xPix1421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[14] VREF PIX_IN[1421] NB2 NB1 CSA_VREF pixel
xPix1422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[14] VREF PIX_IN[1422] NB2 NB1 CSA_VREF pixel
xPix1423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[14] VREF PIX_IN[1423] NB2 NB1 CSA_VREF pixel
xPix1424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[14] VREF PIX_IN[1424] NB2 NB1 CSA_VREF pixel
xPix1425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[14] VREF PIX_IN[1425] NB2 NB1 CSA_VREF pixel
xPix1426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[14] VREF PIX_IN[1426] NB2 NB1 CSA_VREF pixel
xPix1427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[14] VREF PIX_IN[1427] NB2 NB1 CSA_VREF pixel
xPix1428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[14] VREF PIX_IN[1428] NB2 NB1 CSA_VREF pixel
xPix1429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[14] VREF PIX_IN[1429] NB2 NB1 CSA_VREF pixel
xPix1430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[14] VREF PIX_IN[1430] NB2 NB1 CSA_VREF pixel
xPix1431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[14] VREF PIX_IN[1431] NB2 NB1 CSA_VREF pixel
xPix1432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[14] VREF PIX_IN[1432] NB2 NB1 CSA_VREF pixel
xPix1433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[14] VREF PIX_IN[1433] NB2 NB1 CSA_VREF pixel
xPix1434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[14] VREF PIX_IN[1434] NB2 NB1 CSA_VREF pixel
xPix1435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[14] VREF PIX_IN[1435] NB2 NB1 CSA_VREF pixel
xPix1436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[14] VREF PIX_IN[1436] NB2 NB1 CSA_VREF pixel
xPix1437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[14] VREF PIX_IN[1437] NB2 NB1 CSA_VREF pixel
xPix1438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[14] VREF PIX_IN[1438] NB2 NB1 CSA_VREF pixel
xPix1439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[14] VREF PIX_IN[1439] NB2 NB1 CSA_VREF pixel
xPix1440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[14] VREF PIX_IN[1440] NB2 NB1 CSA_VREF pixel
xPix1441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[14] VREF PIX_IN[1441] NB2 NB1 CSA_VREF pixel
xPix1442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[14] VREF PIX_IN[1442] NB2 NB1 CSA_VREF pixel
xPix1443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[14] VREF PIX_IN[1443] NB2 NB1 CSA_VREF pixel
xPix1444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[14] VREF PIX_IN[1444] NB2 NB1 CSA_VREF pixel
xPix1445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[14] VREF PIX_IN[1445] NB2 NB1 CSA_VREF pixel
xPix1446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[14] VREF PIX_IN[1446] NB2 NB1 CSA_VREF pixel
xPix1447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[14] VREF PIX_IN[1447] NB2 NB1 CSA_VREF pixel
xPix1448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[14] VREF PIX_IN[1448] NB2 NB1 CSA_VREF pixel
xPix1449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[14] VREF PIX_IN[1449] NB2 NB1 CSA_VREF pixel
xPix1450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[14] VREF PIX_IN[1450] NB2 NB1 CSA_VREF pixel
xPix1451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[14] VREF PIX_IN[1451] NB2 NB1 CSA_VREF pixel
xPix1452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[14] VREF PIX_IN[1452] NB2 NB1 CSA_VREF pixel
xPix1453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[14] VREF PIX_IN[1453] NB2 NB1 CSA_VREF pixel
xPix1454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[14] VREF PIX_IN[1454] NB2 NB1 CSA_VREF pixel
xPix1455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[14] VREF PIX_IN[1455] NB2 NB1 CSA_VREF pixel
xPix1456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[14] VREF PIX_IN[1456] NB2 NB1 CSA_VREF pixel
xPix1457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[14] VREF PIX_IN[1457] NB2 NB1 CSA_VREF pixel
xPix1458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[14] VREF PIX_IN[1458] NB2 NB1 CSA_VREF pixel
xPix1459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[14] VREF PIX_IN[1459] NB2 NB1 CSA_VREF pixel
xPix1460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[14] VREF PIX_IN[1460] NB2 NB1 CSA_VREF pixel
xPix1461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[14] VREF PIX_IN[1461] NB2 NB1 CSA_VREF pixel
xPix1462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[14] VREF PIX_IN[1462] NB2 NB1 CSA_VREF pixel
xPix1463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[14] VREF PIX_IN[1463] NB2 NB1 CSA_VREF pixel
xPix1464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[14] VREF PIX_IN[1464] NB2 NB1 CSA_VREF pixel
xPix1465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[14] VREF PIX_IN[1465] NB2 NB1 CSA_VREF pixel
xPix1466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[14] VREF PIX_IN[1466] NB2 NB1 CSA_VREF pixel
xPix1467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[14] VREF PIX_IN[1467] NB2 NB1 CSA_VREF pixel
xPix1468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[14] VREF PIX_IN[1468] NB2 NB1 CSA_VREF pixel
xPix1469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[14] VREF PIX_IN[1469] NB2 NB1 CSA_VREF pixel
xPix1470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[14] VREF PIX_IN[1470] NB2 NB1 CSA_VREF pixel
xPix1471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[14] VREF PIX_IN[1471] NB2 NB1 CSA_VREF pixel
xPix1472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[14] VREF PIX_IN[1472] NB2 NB1 CSA_VREF pixel
xPix1473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[14] VREF PIX_IN[1473] NB2 NB1 CSA_VREF pixel
xPix1474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[14] VREF PIX_IN[1474] NB2 NB1 CSA_VREF pixel
xPix1475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[14] VREF PIX_IN[1475] NB2 NB1 CSA_VREF pixel
xPix1476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[14] VREF PIX_IN[1476] NB2 NB1 CSA_VREF pixel
xPix1477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[14] VREF PIX_IN[1477] NB2 NB1 CSA_VREF pixel
xPix1478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[14] VREF PIX_IN[1478] NB2 NB1 CSA_VREF pixel
xPix1479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[14] VREF PIX_IN[1479] NB2 NB1 CSA_VREF pixel
xPix1480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[14] VREF PIX_IN[1480] NB2 NB1 CSA_VREF pixel
xPix1481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[14] VREF PIX_IN[1481] NB2 NB1 CSA_VREF pixel
xPix1482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[14] VREF PIX_IN[1482] NB2 NB1 CSA_VREF pixel
xPix1483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[14] VREF PIX_IN[1483] NB2 NB1 CSA_VREF pixel
xPix1484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[14] VREF PIX_IN[1484] NB2 NB1 CSA_VREF pixel
xPix1485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[14] VREF PIX_IN[1485] NB2 NB1 CSA_VREF pixel
xPix1486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[14] VREF PIX_IN[1486] NB2 NB1 CSA_VREF pixel
xPix1487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[14] VREF PIX_IN[1487] NB2 NB1 CSA_VREF pixel
xPix1488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[14] VREF PIX_IN[1488] NB2 NB1 CSA_VREF pixel
xPix1489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[14] VREF PIX_IN[1489] NB2 NB1 CSA_VREF pixel
xPix1490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[14] VREF PIX_IN[1490] NB2 NB1 CSA_VREF pixel
xPix1491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[14] VREF PIX_IN[1491] NB2 NB1 CSA_VREF pixel
xPix1492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[14] VREF PIX_IN[1492] NB2 NB1 CSA_VREF pixel
xPix1493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[14] VREF PIX_IN[1493] NB2 NB1 CSA_VREF pixel
xPix1494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[14] VREF PIX_IN[1494] NB2 NB1 CSA_VREF pixel
xPix1495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[14] VREF PIX_IN[1495] NB2 NB1 CSA_VREF pixel
xPix1496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[14] VREF PIX_IN[1496] NB2 NB1 CSA_VREF pixel
xPix1497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[14] VREF PIX_IN[1497] NB2 NB1 CSA_VREF pixel
xPix1498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[14] VREF PIX_IN[1498] NB2 NB1 CSA_VREF pixel
xPix1499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[14] VREF PIX_IN[1499] NB2 NB1 CSA_VREF pixel
xPix1500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[15] VREF PIX_IN[1500] NB2 NB1 CSA_VREF pixel
xPix1501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[15] VREF PIX_IN[1501] NB2 NB1 CSA_VREF pixel
xPix1502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[15] VREF PIX_IN[1502] NB2 NB1 CSA_VREF pixel
xPix1503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[15] VREF PIX_IN[1503] NB2 NB1 CSA_VREF pixel
xPix1504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[15] VREF PIX_IN[1504] NB2 NB1 CSA_VREF pixel
xPix1505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[15] VREF PIX_IN[1505] NB2 NB1 CSA_VREF pixel
xPix1506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[15] VREF PIX_IN[1506] NB2 NB1 CSA_VREF pixel
xPix1507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[15] VREF PIX_IN[1507] NB2 NB1 CSA_VREF pixel
xPix1508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[15] VREF PIX_IN[1508] NB2 NB1 CSA_VREF pixel
xPix1509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[15] VREF PIX_IN[1509] NB2 NB1 CSA_VREF pixel
xPix1510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[15] VREF PIX_IN[1510] NB2 NB1 CSA_VREF pixel
xPix1511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[15] VREF PIX_IN[1511] NB2 NB1 CSA_VREF pixel
xPix1512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[15] VREF PIX_IN[1512] NB2 NB1 CSA_VREF pixel
xPix1513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[15] VREF PIX_IN[1513] NB2 NB1 CSA_VREF pixel
xPix1514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[15] VREF PIX_IN[1514] NB2 NB1 CSA_VREF pixel
xPix1515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[15] VREF PIX_IN[1515] NB2 NB1 CSA_VREF pixel
xPix1516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[15] VREF PIX_IN[1516] NB2 NB1 CSA_VREF pixel
xPix1517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[15] VREF PIX_IN[1517] NB2 NB1 CSA_VREF pixel
xPix1518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[15] VREF PIX_IN[1518] NB2 NB1 CSA_VREF pixel
xPix1519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[15] VREF PIX_IN[1519] NB2 NB1 CSA_VREF pixel
xPix1520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[15] VREF PIX_IN[1520] NB2 NB1 CSA_VREF pixel
xPix1521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[15] VREF PIX_IN[1521] NB2 NB1 CSA_VREF pixel
xPix1522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[15] VREF PIX_IN[1522] NB2 NB1 CSA_VREF pixel
xPix1523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[15] VREF PIX_IN[1523] NB2 NB1 CSA_VREF pixel
xPix1524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[15] VREF PIX_IN[1524] NB2 NB1 CSA_VREF pixel
xPix1525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[15] VREF PIX_IN[1525] NB2 NB1 CSA_VREF pixel
xPix1526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[15] VREF PIX_IN[1526] NB2 NB1 CSA_VREF pixel
xPix1527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[15] VREF PIX_IN[1527] NB2 NB1 CSA_VREF pixel
xPix1528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[15] VREF PIX_IN[1528] NB2 NB1 CSA_VREF pixel
xPix1529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[15] VREF PIX_IN[1529] NB2 NB1 CSA_VREF pixel
xPix1530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[15] VREF PIX_IN[1530] NB2 NB1 CSA_VREF pixel
xPix1531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[15] VREF PIX_IN[1531] NB2 NB1 CSA_VREF pixel
xPix1532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[15] VREF PIX_IN[1532] NB2 NB1 CSA_VREF pixel
xPix1533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[15] VREF PIX_IN[1533] NB2 NB1 CSA_VREF pixel
xPix1534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[15] VREF PIX_IN[1534] NB2 NB1 CSA_VREF pixel
xPix1535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[15] VREF PIX_IN[1535] NB2 NB1 CSA_VREF pixel
xPix1536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[15] VREF PIX_IN[1536] NB2 NB1 CSA_VREF pixel
xPix1537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[15] VREF PIX_IN[1537] NB2 NB1 CSA_VREF pixel
xPix1538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[15] VREF PIX_IN[1538] NB2 NB1 CSA_VREF pixel
xPix1539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[15] VREF PIX_IN[1539] NB2 NB1 CSA_VREF pixel
xPix1540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[15] VREF PIX_IN[1540] NB2 NB1 CSA_VREF pixel
xPix1541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[15] VREF PIX_IN[1541] NB2 NB1 CSA_VREF pixel
xPix1542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[15] VREF PIX_IN[1542] NB2 NB1 CSA_VREF pixel
xPix1543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[15] VREF PIX_IN[1543] NB2 NB1 CSA_VREF pixel
xPix1544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[15] VREF PIX_IN[1544] NB2 NB1 CSA_VREF pixel
xPix1545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[15] VREF PIX_IN[1545] NB2 NB1 CSA_VREF pixel
xPix1546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[15] VREF PIX_IN[1546] NB2 NB1 CSA_VREF pixel
xPix1547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[15] VREF PIX_IN[1547] NB2 NB1 CSA_VREF pixel
xPix1548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[15] VREF PIX_IN[1548] NB2 NB1 CSA_VREF pixel
xPix1549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[15] VREF PIX_IN[1549] NB2 NB1 CSA_VREF pixel
xPix1550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[15] VREF PIX_IN[1550] NB2 NB1 CSA_VREF pixel
xPix1551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[15] VREF PIX_IN[1551] NB2 NB1 CSA_VREF pixel
xPix1552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[15] VREF PIX_IN[1552] NB2 NB1 CSA_VREF pixel
xPix1553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[15] VREF PIX_IN[1553] NB2 NB1 CSA_VREF pixel
xPix1554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[15] VREF PIX_IN[1554] NB2 NB1 CSA_VREF pixel
xPix1555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[15] VREF PIX_IN[1555] NB2 NB1 CSA_VREF pixel
xPix1556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[15] VREF PIX_IN[1556] NB2 NB1 CSA_VREF pixel
xPix1557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[15] VREF PIX_IN[1557] NB2 NB1 CSA_VREF pixel
xPix1558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[15] VREF PIX_IN[1558] NB2 NB1 CSA_VREF pixel
xPix1559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[15] VREF PIX_IN[1559] NB2 NB1 CSA_VREF pixel
xPix1560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[15] VREF PIX_IN[1560] NB2 NB1 CSA_VREF pixel
xPix1561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[15] VREF PIX_IN[1561] NB2 NB1 CSA_VREF pixel
xPix1562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[15] VREF PIX_IN[1562] NB2 NB1 CSA_VREF pixel
xPix1563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[15] VREF PIX_IN[1563] NB2 NB1 CSA_VREF pixel
xPix1564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[15] VREF PIX_IN[1564] NB2 NB1 CSA_VREF pixel
xPix1565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[15] VREF PIX_IN[1565] NB2 NB1 CSA_VREF pixel
xPix1566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[15] VREF PIX_IN[1566] NB2 NB1 CSA_VREF pixel
xPix1567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[15] VREF PIX_IN[1567] NB2 NB1 CSA_VREF pixel
xPix1568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[15] VREF PIX_IN[1568] NB2 NB1 CSA_VREF pixel
xPix1569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[15] VREF PIX_IN[1569] NB2 NB1 CSA_VREF pixel
xPix1570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[15] VREF PIX_IN[1570] NB2 NB1 CSA_VREF pixel
xPix1571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[15] VREF PIX_IN[1571] NB2 NB1 CSA_VREF pixel
xPix1572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[15] VREF PIX_IN[1572] NB2 NB1 CSA_VREF pixel
xPix1573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[15] VREF PIX_IN[1573] NB2 NB1 CSA_VREF pixel
xPix1574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[15] VREF PIX_IN[1574] NB2 NB1 CSA_VREF pixel
xPix1575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[15] VREF PIX_IN[1575] NB2 NB1 CSA_VREF pixel
xPix1576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[15] VREF PIX_IN[1576] NB2 NB1 CSA_VREF pixel
xPix1577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[15] VREF PIX_IN[1577] NB2 NB1 CSA_VREF pixel
xPix1578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[15] VREF PIX_IN[1578] NB2 NB1 CSA_VREF pixel
xPix1579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[15] VREF PIX_IN[1579] NB2 NB1 CSA_VREF pixel
xPix1580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[15] VREF PIX_IN[1580] NB2 NB1 CSA_VREF pixel
xPix1581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[15] VREF PIX_IN[1581] NB2 NB1 CSA_VREF pixel
xPix1582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[15] VREF PIX_IN[1582] NB2 NB1 CSA_VREF pixel
xPix1583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[15] VREF PIX_IN[1583] NB2 NB1 CSA_VREF pixel
xPix1584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[15] VREF PIX_IN[1584] NB2 NB1 CSA_VREF pixel
xPix1585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[15] VREF PIX_IN[1585] NB2 NB1 CSA_VREF pixel
xPix1586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[15] VREF PIX_IN[1586] NB2 NB1 CSA_VREF pixel
xPix1587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[15] VREF PIX_IN[1587] NB2 NB1 CSA_VREF pixel
xPix1588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[15] VREF PIX_IN[1588] NB2 NB1 CSA_VREF pixel
xPix1589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[15] VREF PIX_IN[1589] NB2 NB1 CSA_VREF pixel
xPix1590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[15] VREF PIX_IN[1590] NB2 NB1 CSA_VREF pixel
xPix1591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[15] VREF PIX_IN[1591] NB2 NB1 CSA_VREF pixel
xPix1592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[15] VREF PIX_IN[1592] NB2 NB1 CSA_VREF pixel
xPix1593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[15] VREF PIX_IN[1593] NB2 NB1 CSA_VREF pixel
xPix1594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[15] VREF PIX_IN[1594] NB2 NB1 CSA_VREF pixel
xPix1595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[15] VREF PIX_IN[1595] NB2 NB1 CSA_VREF pixel
xPix1596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[15] VREF PIX_IN[1596] NB2 NB1 CSA_VREF pixel
xPix1597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[15] VREF PIX_IN[1597] NB2 NB1 CSA_VREF pixel
xPix1598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[15] VREF PIX_IN[1598] NB2 NB1 CSA_VREF pixel
xPix1599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[15] VREF PIX_IN[1599] NB2 NB1 CSA_VREF pixel
xPix1600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[16] VREF PIX_IN[1600] NB2 NB1 CSA_VREF pixel
xPix1601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[16] VREF PIX_IN[1601] NB2 NB1 CSA_VREF pixel
xPix1602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[16] VREF PIX_IN[1602] NB2 NB1 CSA_VREF pixel
xPix1603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[16] VREF PIX_IN[1603] NB2 NB1 CSA_VREF pixel
xPix1604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[16] VREF PIX_IN[1604] NB2 NB1 CSA_VREF pixel
xPix1605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[16] VREF PIX_IN[1605] NB2 NB1 CSA_VREF pixel
xPix1606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[16] VREF PIX_IN[1606] NB2 NB1 CSA_VREF pixel
xPix1607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[16] VREF PIX_IN[1607] NB2 NB1 CSA_VREF pixel
xPix1608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[16] VREF PIX_IN[1608] NB2 NB1 CSA_VREF pixel
xPix1609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[16] VREF PIX_IN[1609] NB2 NB1 CSA_VREF pixel
xPix1610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[16] VREF PIX_IN[1610] NB2 NB1 CSA_VREF pixel
xPix1611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[16] VREF PIX_IN[1611] NB2 NB1 CSA_VREF pixel
xPix1612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[16] VREF PIX_IN[1612] NB2 NB1 CSA_VREF pixel
xPix1613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[16] VREF PIX_IN[1613] NB2 NB1 CSA_VREF pixel
xPix1614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[16] VREF PIX_IN[1614] NB2 NB1 CSA_VREF pixel
xPix1615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[16] VREF PIX_IN[1615] NB2 NB1 CSA_VREF pixel
xPix1616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[16] VREF PIX_IN[1616] NB2 NB1 CSA_VREF pixel
xPix1617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[16] VREF PIX_IN[1617] NB2 NB1 CSA_VREF pixel
xPix1618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[16] VREF PIX_IN[1618] NB2 NB1 CSA_VREF pixel
xPix1619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[16] VREF PIX_IN[1619] NB2 NB1 CSA_VREF pixel
xPix1620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[16] VREF PIX_IN[1620] NB2 NB1 CSA_VREF pixel
xPix1621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[16] VREF PIX_IN[1621] NB2 NB1 CSA_VREF pixel
xPix1622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[16] VREF PIX_IN[1622] NB2 NB1 CSA_VREF pixel
xPix1623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[16] VREF PIX_IN[1623] NB2 NB1 CSA_VREF pixel
xPix1624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[16] VREF PIX_IN[1624] NB2 NB1 CSA_VREF pixel
xPix1625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[16] VREF PIX_IN[1625] NB2 NB1 CSA_VREF pixel
xPix1626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[16] VREF PIX_IN[1626] NB2 NB1 CSA_VREF pixel
xPix1627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[16] VREF PIX_IN[1627] NB2 NB1 CSA_VREF pixel
xPix1628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[16] VREF PIX_IN[1628] NB2 NB1 CSA_VREF pixel
xPix1629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[16] VREF PIX_IN[1629] NB2 NB1 CSA_VREF pixel
xPix1630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[16] VREF PIX_IN[1630] NB2 NB1 CSA_VREF pixel
xPix1631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[16] VREF PIX_IN[1631] NB2 NB1 CSA_VREF pixel
xPix1632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[16] VREF PIX_IN[1632] NB2 NB1 CSA_VREF pixel
xPix1633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[16] VREF PIX_IN[1633] NB2 NB1 CSA_VREF pixel
xPix1634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[16] VREF PIX_IN[1634] NB2 NB1 CSA_VREF pixel
xPix1635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[16] VREF PIX_IN[1635] NB2 NB1 CSA_VREF pixel
xPix1636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[16] VREF PIX_IN[1636] NB2 NB1 CSA_VREF pixel
xPix1637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[16] VREF PIX_IN[1637] NB2 NB1 CSA_VREF pixel
xPix1638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[16] VREF PIX_IN[1638] NB2 NB1 CSA_VREF pixel
xPix1639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[16] VREF PIX_IN[1639] NB2 NB1 CSA_VREF pixel
xPix1640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[16] VREF PIX_IN[1640] NB2 NB1 CSA_VREF pixel
xPix1641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[16] VREF PIX_IN[1641] NB2 NB1 CSA_VREF pixel
xPix1642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[16] VREF PIX_IN[1642] NB2 NB1 CSA_VREF pixel
xPix1643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[16] VREF PIX_IN[1643] NB2 NB1 CSA_VREF pixel
xPix1644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[16] VREF PIX_IN[1644] NB2 NB1 CSA_VREF pixel
xPix1645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[16] VREF PIX_IN[1645] NB2 NB1 CSA_VREF pixel
xPix1646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[16] VREF PIX_IN[1646] NB2 NB1 CSA_VREF pixel
xPix1647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[16] VREF PIX_IN[1647] NB2 NB1 CSA_VREF pixel
xPix1648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[16] VREF PIX_IN[1648] NB2 NB1 CSA_VREF pixel
xPix1649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[16] VREF PIX_IN[1649] NB2 NB1 CSA_VREF pixel
xPix1650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[16] VREF PIX_IN[1650] NB2 NB1 CSA_VREF pixel
xPix1651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[16] VREF PIX_IN[1651] NB2 NB1 CSA_VREF pixel
xPix1652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[16] VREF PIX_IN[1652] NB2 NB1 CSA_VREF pixel
xPix1653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[16] VREF PIX_IN[1653] NB2 NB1 CSA_VREF pixel
xPix1654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[16] VREF PIX_IN[1654] NB2 NB1 CSA_VREF pixel
xPix1655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[16] VREF PIX_IN[1655] NB2 NB1 CSA_VREF pixel
xPix1656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[16] VREF PIX_IN[1656] NB2 NB1 CSA_VREF pixel
xPix1657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[16] VREF PIX_IN[1657] NB2 NB1 CSA_VREF pixel
xPix1658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[16] VREF PIX_IN[1658] NB2 NB1 CSA_VREF pixel
xPix1659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[16] VREF PIX_IN[1659] NB2 NB1 CSA_VREF pixel
xPix1660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[16] VREF PIX_IN[1660] NB2 NB1 CSA_VREF pixel
xPix1661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[16] VREF PIX_IN[1661] NB2 NB1 CSA_VREF pixel
xPix1662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[16] VREF PIX_IN[1662] NB2 NB1 CSA_VREF pixel
xPix1663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[16] VREF PIX_IN[1663] NB2 NB1 CSA_VREF pixel
xPix1664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[16] VREF PIX_IN[1664] NB2 NB1 CSA_VREF pixel
xPix1665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[16] VREF PIX_IN[1665] NB2 NB1 CSA_VREF pixel
xPix1666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[16] VREF PIX_IN[1666] NB2 NB1 CSA_VREF pixel
xPix1667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[16] VREF PIX_IN[1667] NB2 NB1 CSA_VREF pixel
xPix1668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[16] VREF PIX_IN[1668] NB2 NB1 CSA_VREF pixel
xPix1669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[16] VREF PIX_IN[1669] NB2 NB1 CSA_VREF pixel
xPix1670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[16] VREF PIX_IN[1670] NB2 NB1 CSA_VREF pixel
xPix1671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[16] VREF PIX_IN[1671] NB2 NB1 CSA_VREF pixel
xPix1672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[16] VREF PIX_IN[1672] NB2 NB1 CSA_VREF pixel
xPix1673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[16] VREF PIX_IN[1673] NB2 NB1 CSA_VREF pixel
xPix1674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[16] VREF PIX_IN[1674] NB2 NB1 CSA_VREF pixel
xPix1675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[16] VREF PIX_IN[1675] NB2 NB1 CSA_VREF pixel
xPix1676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[16] VREF PIX_IN[1676] NB2 NB1 CSA_VREF pixel
xPix1677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[16] VREF PIX_IN[1677] NB2 NB1 CSA_VREF pixel
xPix1678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[16] VREF PIX_IN[1678] NB2 NB1 CSA_VREF pixel
xPix1679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[16] VREF PIX_IN[1679] NB2 NB1 CSA_VREF pixel
xPix1680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[16] VREF PIX_IN[1680] NB2 NB1 CSA_VREF pixel
xPix1681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[16] VREF PIX_IN[1681] NB2 NB1 CSA_VREF pixel
xPix1682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[16] VREF PIX_IN[1682] NB2 NB1 CSA_VREF pixel
xPix1683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[16] VREF PIX_IN[1683] NB2 NB1 CSA_VREF pixel
xPix1684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[16] VREF PIX_IN[1684] NB2 NB1 CSA_VREF pixel
xPix1685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[16] VREF PIX_IN[1685] NB2 NB1 CSA_VREF pixel
xPix1686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[16] VREF PIX_IN[1686] NB2 NB1 CSA_VREF pixel
xPix1687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[16] VREF PIX_IN[1687] NB2 NB1 CSA_VREF pixel
xPix1688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[16] VREF PIX_IN[1688] NB2 NB1 CSA_VREF pixel
xPix1689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[16] VREF PIX_IN[1689] NB2 NB1 CSA_VREF pixel
xPix1690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[16] VREF PIX_IN[1690] NB2 NB1 CSA_VREF pixel
xPix1691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[16] VREF PIX_IN[1691] NB2 NB1 CSA_VREF pixel
xPix1692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[16] VREF PIX_IN[1692] NB2 NB1 CSA_VREF pixel
xPix1693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[16] VREF PIX_IN[1693] NB2 NB1 CSA_VREF pixel
xPix1694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[16] VREF PIX_IN[1694] NB2 NB1 CSA_VREF pixel
xPix1695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[16] VREF PIX_IN[1695] NB2 NB1 CSA_VREF pixel
xPix1696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[16] VREF PIX_IN[1696] NB2 NB1 CSA_VREF pixel
xPix1697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[16] VREF PIX_IN[1697] NB2 NB1 CSA_VREF pixel
xPix1698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[16] VREF PIX_IN[1698] NB2 NB1 CSA_VREF pixel
xPix1699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[16] VREF PIX_IN[1699] NB2 NB1 CSA_VREF pixel
xPix1700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[17] VREF PIX_IN[1700] NB2 NB1 CSA_VREF pixel
xPix1701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[17] VREF PIX_IN[1701] NB2 NB1 CSA_VREF pixel
xPix1702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[17] VREF PIX_IN[1702] NB2 NB1 CSA_VREF pixel
xPix1703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[17] VREF PIX_IN[1703] NB2 NB1 CSA_VREF pixel
xPix1704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[17] VREF PIX_IN[1704] NB2 NB1 CSA_VREF pixel
xPix1705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[17] VREF PIX_IN[1705] NB2 NB1 CSA_VREF pixel
xPix1706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[17] VREF PIX_IN[1706] NB2 NB1 CSA_VREF pixel
xPix1707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[17] VREF PIX_IN[1707] NB2 NB1 CSA_VREF pixel
xPix1708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[17] VREF PIX_IN[1708] NB2 NB1 CSA_VREF pixel
xPix1709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[17] VREF PIX_IN[1709] NB2 NB1 CSA_VREF pixel
xPix1710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[17] VREF PIX_IN[1710] NB2 NB1 CSA_VREF pixel
xPix1711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[17] VREF PIX_IN[1711] NB2 NB1 CSA_VREF pixel
xPix1712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[17] VREF PIX_IN[1712] NB2 NB1 CSA_VREF pixel
xPix1713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[17] VREF PIX_IN[1713] NB2 NB1 CSA_VREF pixel
xPix1714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[17] VREF PIX_IN[1714] NB2 NB1 CSA_VREF pixel
xPix1715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[17] VREF PIX_IN[1715] NB2 NB1 CSA_VREF pixel
xPix1716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[17] VREF PIX_IN[1716] NB2 NB1 CSA_VREF pixel
xPix1717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[17] VREF PIX_IN[1717] NB2 NB1 CSA_VREF pixel
xPix1718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[17] VREF PIX_IN[1718] NB2 NB1 CSA_VREF pixel
xPix1719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[17] VREF PIX_IN[1719] NB2 NB1 CSA_VREF pixel
xPix1720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[17] VREF PIX_IN[1720] NB2 NB1 CSA_VREF pixel
xPix1721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[17] VREF PIX_IN[1721] NB2 NB1 CSA_VREF pixel
xPix1722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[17] VREF PIX_IN[1722] NB2 NB1 CSA_VREF pixel
xPix1723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[17] VREF PIX_IN[1723] NB2 NB1 CSA_VREF pixel
xPix1724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[17] VREF PIX_IN[1724] NB2 NB1 CSA_VREF pixel
xPix1725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[17] VREF PIX_IN[1725] NB2 NB1 CSA_VREF pixel
xPix1726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[17] VREF PIX_IN[1726] NB2 NB1 CSA_VREF pixel
xPix1727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[17] VREF PIX_IN[1727] NB2 NB1 CSA_VREF pixel
xPix1728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[17] VREF PIX_IN[1728] NB2 NB1 CSA_VREF pixel
xPix1729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[17] VREF PIX_IN[1729] NB2 NB1 CSA_VREF pixel
xPix1730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[17] VREF PIX_IN[1730] NB2 NB1 CSA_VREF pixel
xPix1731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[17] VREF PIX_IN[1731] NB2 NB1 CSA_VREF pixel
xPix1732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[17] VREF PIX_IN[1732] NB2 NB1 CSA_VREF pixel
xPix1733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[17] VREF PIX_IN[1733] NB2 NB1 CSA_VREF pixel
xPix1734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[17] VREF PIX_IN[1734] NB2 NB1 CSA_VREF pixel
xPix1735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[17] VREF PIX_IN[1735] NB2 NB1 CSA_VREF pixel
xPix1736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[17] VREF PIX_IN[1736] NB2 NB1 CSA_VREF pixel
xPix1737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[17] VREF PIX_IN[1737] NB2 NB1 CSA_VREF pixel
xPix1738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[17] VREF PIX_IN[1738] NB2 NB1 CSA_VREF pixel
xPix1739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[17] VREF PIX_IN[1739] NB2 NB1 CSA_VREF pixel
xPix1740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[17] VREF PIX_IN[1740] NB2 NB1 CSA_VREF pixel
xPix1741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[17] VREF PIX_IN[1741] NB2 NB1 CSA_VREF pixel
xPix1742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[17] VREF PIX_IN[1742] NB2 NB1 CSA_VREF pixel
xPix1743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[17] VREF PIX_IN[1743] NB2 NB1 CSA_VREF pixel
xPix1744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[17] VREF PIX_IN[1744] NB2 NB1 CSA_VREF pixel
xPix1745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[17] VREF PIX_IN[1745] NB2 NB1 CSA_VREF pixel
xPix1746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[17] VREF PIX_IN[1746] NB2 NB1 CSA_VREF pixel
xPix1747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[17] VREF PIX_IN[1747] NB2 NB1 CSA_VREF pixel
xPix1748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[17] VREF PIX_IN[1748] NB2 NB1 CSA_VREF pixel
xPix1749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[17] VREF PIX_IN[1749] NB2 NB1 CSA_VREF pixel
xPix1750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[17] VREF PIX_IN[1750] NB2 NB1 CSA_VREF pixel
xPix1751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[17] VREF PIX_IN[1751] NB2 NB1 CSA_VREF pixel
xPix1752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[17] VREF PIX_IN[1752] NB2 NB1 CSA_VREF pixel
xPix1753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[17] VREF PIX_IN[1753] NB2 NB1 CSA_VREF pixel
xPix1754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[17] VREF PIX_IN[1754] NB2 NB1 CSA_VREF pixel
xPix1755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[17] VREF PIX_IN[1755] NB2 NB1 CSA_VREF pixel
xPix1756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[17] VREF PIX_IN[1756] NB2 NB1 CSA_VREF pixel
xPix1757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[17] VREF PIX_IN[1757] NB2 NB1 CSA_VREF pixel
xPix1758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[17] VREF PIX_IN[1758] NB2 NB1 CSA_VREF pixel
xPix1759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[17] VREF PIX_IN[1759] NB2 NB1 CSA_VREF pixel
xPix1760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[17] VREF PIX_IN[1760] NB2 NB1 CSA_VREF pixel
xPix1761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[17] VREF PIX_IN[1761] NB2 NB1 CSA_VREF pixel
xPix1762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[17] VREF PIX_IN[1762] NB2 NB1 CSA_VREF pixel
xPix1763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[17] VREF PIX_IN[1763] NB2 NB1 CSA_VREF pixel
xPix1764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[17] VREF PIX_IN[1764] NB2 NB1 CSA_VREF pixel
xPix1765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[17] VREF PIX_IN[1765] NB2 NB1 CSA_VREF pixel
xPix1766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[17] VREF PIX_IN[1766] NB2 NB1 CSA_VREF pixel
xPix1767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[17] VREF PIX_IN[1767] NB2 NB1 CSA_VREF pixel
xPix1768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[17] VREF PIX_IN[1768] NB2 NB1 CSA_VREF pixel
xPix1769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[17] VREF PIX_IN[1769] NB2 NB1 CSA_VREF pixel
xPix1770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[17] VREF PIX_IN[1770] NB2 NB1 CSA_VREF pixel
xPix1771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[17] VREF PIX_IN[1771] NB2 NB1 CSA_VREF pixel
xPix1772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[17] VREF PIX_IN[1772] NB2 NB1 CSA_VREF pixel
xPix1773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[17] VREF PIX_IN[1773] NB2 NB1 CSA_VREF pixel
xPix1774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[17] VREF PIX_IN[1774] NB2 NB1 CSA_VREF pixel
xPix1775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[17] VREF PIX_IN[1775] NB2 NB1 CSA_VREF pixel
xPix1776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[17] VREF PIX_IN[1776] NB2 NB1 CSA_VREF pixel
xPix1777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[17] VREF PIX_IN[1777] NB2 NB1 CSA_VREF pixel
xPix1778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[17] VREF PIX_IN[1778] NB2 NB1 CSA_VREF pixel
xPix1779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[17] VREF PIX_IN[1779] NB2 NB1 CSA_VREF pixel
xPix1780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[17] VREF PIX_IN[1780] NB2 NB1 CSA_VREF pixel
xPix1781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[17] VREF PIX_IN[1781] NB2 NB1 CSA_VREF pixel
xPix1782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[17] VREF PIX_IN[1782] NB2 NB1 CSA_VREF pixel
xPix1783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[17] VREF PIX_IN[1783] NB2 NB1 CSA_VREF pixel
xPix1784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[17] VREF PIX_IN[1784] NB2 NB1 CSA_VREF pixel
xPix1785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[17] VREF PIX_IN[1785] NB2 NB1 CSA_VREF pixel
xPix1786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[17] VREF PIX_IN[1786] NB2 NB1 CSA_VREF pixel
xPix1787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[17] VREF PIX_IN[1787] NB2 NB1 CSA_VREF pixel
xPix1788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[17] VREF PIX_IN[1788] NB2 NB1 CSA_VREF pixel
xPix1789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[17] VREF PIX_IN[1789] NB2 NB1 CSA_VREF pixel
xPix1790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[17] VREF PIX_IN[1790] NB2 NB1 CSA_VREF pixel
xPix1791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[17] VREF PIX_IN[1791] NB2 NB1 CSA_VREF pixel
xPix1792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[17] VREF PIX_IN[1792] NB2 NB1 CSA_VREF pixel
xPix1793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[17] VREF PIX_IN[1793] NB2 NB1 CSA_VREF pixel
xPix1794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[17] VREF PIX_IN[1794] NB2 NB1 CSA_VREF pixel
xPix1795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[17] VREF PIX_IN[1795] NB2 NB1 CSA_VREF pixel
xPix1796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[17] VREF PIX_IN[1796] NB2 NB1 CSA_VREF pixel
xPix1797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[17] VREF PIX_IN[1797] NB2 NB1 CSA_VREF pixel
xPix1798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[17] VREF PIX_IN[1798] NB2 NB1 CSA_VREF pixel
xPix1799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[17] VREF PIX_IN[1799] NB2 NB1 CSA_VREF pixel
xPix1800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[18] VREF PIX_IN[1800] NB2 NB1 CSA_VREF pixel
xPix1801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[18] VREF PIX_IN[1801] NB2 NB1 CSA_VREF pixel
xPix1802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[18] VREF PIX_IN[1802] NB2 NB1 CSA_VREF pixel
xPix1803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[18] VREF PIX_IN[1803] NB2 NB1 CSA_VREF pixel
xPix1804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[18] VREF PIX_IN[1804] NB2 NB1 CSA_VREF pixel
xPix1805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[18] VREF PIX_IN[1805] NB2 NB1 CSA_VREF pixel
xPix1806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[18] VREF PIX_IN[1806] NB2 NB1 CSA_VREF pixel
xPix1807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[18] VREF PIX_IN[1807] NB2 NB1 CSA_VREF pixel
xPix1808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[18] VREF PIX_IN[1808] NB2 NB1 CSA_VREF pixel
xPix1809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[18] VREF PIX_IN[1809] NB2 NB1 CSA_VREF pixel
xPix1810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[18] VREF PIX_IN[1810] NB2 NB1 CSA_VREF pixel
xPix1811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[18] VREF PIX_IN[1811] NB2 NB1 CSA_VREF pixel
xPix1812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[18] VREF PIX_IN[1812] NB2 NB1 CSA_VREF pixel
xPix1813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[18] VREF PIX_IN[1813] NB2 NB1 CSA_VREF pixel
xPix1814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[18] VREF PIX_IN[1814] NB2 NB1 CSA_VREF pixel
xPix1815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[18] VREF PIX_IN[1815] NB2 NB1 CSA_VREF pixel
xPix1816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[18] VREF PIX_IN[1816] NB2 NB1 CSA_VREF pixel
xPix1817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[18] VREF PIX_IN[1817] NB2 NB1 CSA_VREF pixel
xPix1818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[18] VREF PIX_IN[1818] NB2 NB1 CSA_VREF pixel
xPix1819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[18] VREF PIX_IN[1819] NB2 NB1 CSA_VREF pixel
xPix1820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[18] VREF PIX_IN[1820] NB2 NB1 CSA_VREF pixel
xPix1821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[18] VREF PIX_IN[1821] NB2 NB1 CSA_VREF pixel
xPix1822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[18] VREF PIX_IN[1822] NB2 NB1 CSA_VREF pixel
xPix1823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[18] VREF PIX_IN[1823] NB2 NB1 CSA_VREF pixel
xPix1824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[18] VREF PIX_IN[1824] NB2 NB1 CSA_VREF pixel
xPix1825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[18] VREF PIX_IN[1825] NB2 NB1 CSA_VREF pixel
xPix1826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[18] VREF PIX_IN[1826] NB2 NB1 CSA_VREF pixel
xPix1827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[18] VREF PIX_IN[1827] NB2 NB1 CSA_VREF pixel
xPix1828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[18] VREF PIX_IN[1828] NB2 NB1 CSA_VREF pixel
xPix1829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[18] VREF PIX_IN[1829] NB2 NB1 CSA_VREF pixel
xPix1830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[18] VREF PIX_IN[1830] NB2 NB1 CSA_VREF pixel
xPix1831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[18] VREF PIX_IN[1831] NB2 NB1 CSA_VREF pixel
xPix1832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[18] VREF PIX_IN[1832] NB2 NB1 CSA_VREF pixel
xPix1833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[18] VREF PIX_IN[1833] NB2 NB1 CSA_VREF pixel
xPix1834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[18] VREF PIX_IN[1834] NB2 NB1 CSA_VREF pixel
xPix1835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[18] VREF PIX_IN[1835] NB2 NB1 CSA_VREF pixel
xPix1836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[18] VREF PIX_IN[1836] NB2 NB1 CSA_VREF pixel
xPix1837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[18] VREF PIX_IN[1837] NB2 NB1 CSA_VREF pixel
xPix1838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[18] VREF PIX_IN[1838] NB2 NB1 CSA_VREF pixel
xPix1839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[18] VREF PIX_IN[1839] NB2 NB1 CSA_VREF pixel
xPix1840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[18] VREF PIX_IN[1840] NB2 NB1 CSA_VREF pixel
xPix1841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[18] VREF PIX_IN[1841] NB2 NB1 CSA_VREF pixel
xPix1842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[18] VREF PIX_IN[1842] NB2 NB1 CSA_VREF pixel
xPix1843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[18] VREF PIX_IN[1843] NB2 NB1 CSA_VREF pixel
xPix1844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[18] VREF PIX_IN[1844] NB2 NB1 CSA_VREF pixel
xPix1845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[18] VREF PIX_IN[1845] NB2 NB1 CSA_VREF pixel
xPix1846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[18] VREF PIX_IN[1846] NB2 NB1 CSA_VREF pixel
xPix1847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[18] VREF PIX_IN[1847] NB2 NB1 CSA_VREF pixel
xPix1848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[18] VREF PIX_IN[1848] NB2 NB1 CSA_VREF pixel
xPix1849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[18] VREF PIX_IN[1849] NB2 NB1 CSA_VREF pixel
xPix1850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[18] VREF PIX_IN[1850] NB2 NB1 CSA_VREF pixel
xPix1851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[18] VREF PIX_IN[1851] NB2 NB1 CSA_VREF pixel
xPix1852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[18] VREF PIX_IN[1852] NB2 NB1 CSA_VREF pixel
xPix1853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[18] VREF PIX_IN[1853] NB2 NB1 CSA_VREF pixel
xPix1854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[18] VREF PIX_IN[1854] NB2 NB1 CSA_VREF pixel
xPix1855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[18] VREF PIX_IN[1855] NB2 NB1 CSA_VREF pixel
xPix1856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[18] VREF PIX_IN[1856] NB2 NB1 CSA_VREF pixel
xPix1857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[18] VREF PIX_IN[1857] NB2 NB1 CSA_VREF pixel
xPix1858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[18] VREF PIX_IN[1858] NB2 NB1 CSA_VREF pixel
xPix1859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[18] VREF PIX_IN[1859] NB2 NB1 CSA_VREF pixel
xPix1860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[18] VREF PIX_IN[1860] NB2 NB1 CSA_VREF pixel
xPix1861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[18] VREF PIX_IN[1861] NB2 NB1 CSA_VREF pixel
xPix1862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[18] VREF PIX_IN[1862] NB2 NB1 CSA_VREF pixel
xPix1863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[18] VREF PIX_IN[1863] NB2 NB1 CSA_VREF pixel
xPix1864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[18] VREF PIX_IN[1864] NB2 NB1 CSA_VREF pixel
xPix1865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[18] VREF PIX_IN[1865] NB2 NB1 CSA_VREF pixel
xPix1866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[18] VREF PIX_IN[1866] NB2 NB1 CSA_VREF pixel
xPix1867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[18] VREF PIX_IN[1867] NB2 NB1 CSA_VREF pixel
xPix1868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[18] VREF PIX_IN[1868] NB2 NB1 CSA_VREF pixel
xPix1869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[18] VREF PIX_IN[1869] NB2 NB1 CSA_VREF pixel
xPix1870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[18] VREF PIX_IN[1870] NB2 NB1 CSA_VREF pixel
xPix1871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[18] VREF PIX_IN[1871] NB2 NB1 CSA_VREF pixel
xPix1872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[18] VREF PIX_IN[1872] NB2 NB1 CSA_VREF pixel
xPix1873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[18] VREF PIX_IN[1873] NB2 NB1 CSA_VREF pixel
xPix1874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[18] VREF PIX_IN[1874] NB2 NB1 CSA_VREF pixel
xPix1875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[18] VREF PIX_IN[1875] NB2 NB1 CSA_VREF pixel
xPix1876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[18] VREF PIX_IN[1876] NB2 NB1 CSA_VREF pixel
xPix1877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[18] VREF PIX_IN[1877] NB2 NB1 CSA_VREF pixel
xPix1878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[18] VREF PIX_IN[1878] NB2 NB1 CSA_VREF pixel
xPix1879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[18] VREF PIX_IN[1879] NB2 NB1 CSA_VREF pixel
xPix1880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[18] VREF PIX_IN[1880] NB2 NB1 CSA_VREF pixel
xPix1881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[18] VREF PIX_IN[1881] NB2 NB1 CSA_VREF pixel
xPix1882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[18] VREF PIX_IN[1882] NB2 NB1 CSA_VREF pixel
xPix1883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[18] VREF PIX_IN[1883] NB2 NB1 CSA_VREF pixel
xPix1884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[18] VREF PIX_IN[1884] NB2 NB1 CSA_VREF pixel
xPix1885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[18] VREF PIX_IN[1885] NB2 NB1 CSA_VREF pixel
xPix1886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[18] VREF PIX_IN[1886] NB2 NB1 CSA_VREF pixel
xPix1887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[18] VREF PIX_IN[1887] NB2 NB1 CSA_VREF pixel
xPix1888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[18] VREF PIX_IN[1888] NB2 NB1 CSA_VREF pixel
xPix1889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[18] VREF PIX_IN[1889] NB2 NB1 CSA_VREF pixel
xPix1890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[18] VREF PIX_IN[1890] NB2 NB1 CSA_VREF pixel
xPix1891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[18] VREF PIX_IN[1891] NB2 NB1 CSA_VREF pixel
xPix1892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[18] VREF PIX_IN[1892] NB2 NB1 CSA_VREF pixel
xPix1893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[18] VREF PIX_IN[1893] NB2 NB1 CSA_VREF pixel
xPix1894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[18] VREF PIX_IN[1894] NB2 NB1 CSA_VREF pixel
xPix1895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[18] VREF PIX_IN[1895] NB2 NB1 CSA_VREF pixel
xPix1896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[18] VREF PIX_IN[1896] NB2 NB1 CSA_VREF pixel
xPix1897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[18] VREF PIX_IN[1897] NB2 NB1 CSA_VREF pixel
xPix1898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[18] VREF PIX_IN[1898] NB2 NB1 CSA_VREF pixel
xPix1899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[18] VREF PIX_IN[1899] NB2 NB1 CSA_VREF pixel
xPix1900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[19] VREF PIX_IN[1900] NB2 NB1 CSA_VREF pixel
xPix1901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[19] VREF PIX_IN[1901] NB2 NB1 CSA_VREF pixel
xPix1902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[19] VREF PIX_IN[1902] NB2 NB1 CSA_VREF pixel
xPix1903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[19] VREF PIX_IN[1903] NB2 NB1 CSA_VREF pixel
xPix1904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[19] VREF PIX_IN[1904] NB2 NB1 CSA_VREF pixel
xPix1905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[19] VREF PIX_IN[1905] NB2 NB1 CSA_VREF pixel
xPix1906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[19] VREF PIX_IN[1906] NB2 NB1 CSA_VREF pixel
xPix1907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[19] VREF PIX_IN[1907] NB2 NB1 CSA_VREF pixel
xPix1908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[19] VREF PIX_IN[1908] NB2 NB1 CSA_VREF pixel
xPix1909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[19] VREF PIX_IN[1909] NB2 NB1 CSA_VREF pixel
xPix1910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[19] VREF PIX_IN[1910] NB2 NB1 CSA_VREF pixel
xPix1911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[19] VREF PIX_IN[1911] NB2 NB1 CSA_VREF pixel
xPix1912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[19] VREF PIX_IN[1912] NB2 NB1 CSA_VREF pixel
xPix1913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[19] VREF PIX_IN[1913] NB2 NB1 CSA_VREF pixel
xPix1914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[19] VREF PIX_IN[1914] NB2 NB1 CSA_VREF pixel
xPix1915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[19] VREF PIX_IN[1915] NB2 NB1 CSA_VREF pixel
xPix1916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[19] VREF PIX_IN[1916] NB2 NB1 CSA_VREF pixel
xPix1917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[19] VREF PIX_IN[1917] NB2 NB1 CSA_VREF pixel
xPix1918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[19] VREF PIX_IN[1918] NB2 NB1 CSA_VREF pixel
xPix1919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[19] VREF PIX_IN[1919] NB2 NB1 CSA_VREF pixel
xPix1920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[19] VREF PIX_IN[1920] NB2 NB1 CSA_VREF pixel
xPix1921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[19] VREF PIX_IN[1921] NB2 NB1 CSA_VREF pixel
xPix1922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[19] VREF PIX_IN[1922] NB2 NB1 CSA_VREF pixel
xPix1923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[19] VREF PIX_IN[1923] NB2 NB1 CSA_VREF pixel
xPix1924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[19] VREF PIX_IN[1924] NB2 NB1 CSA_VREF pixel
xPix1925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[19] VREF PIX_IN[1925] NB2 NB1 CSA_VREF pixel
xPix1926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[19] VREF PIX_IN[1926] NB2 NB1 CSA_VREF pixel
xPix1927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[19] VREF PIX_IN[1927] NB2 NB1 CSA_VREF pixel
xPix1928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[19] VREF PIX_IN[1928] NB2 NB1 CSA_VREF pixel
xPix1929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[19] VREF PIX_IN[1929] NB2 NB1 CSA_VREF pixel
xPix1930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[19] VREF PIX_IN[1930] NB2 NB1 CSA_VREF pixel
xPix1931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[19] VREF PIX_IN[1931] NB2 NB1 CSA_VREF pixel
xPix1932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[19] VREF PIX_IN[1932] NB2 NB1 CSA_VREF pixel
xPix1933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[19] VREF PIX_IN[1933] NB2 NB1 CSA_VREF pixel
xPix1934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[19] VREF PIX_IN[1934] NB2 NB1 CSA_VREF pixel
xPix1935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[19] VREF PIX_IN[1935] NB2 NB1 CSA_VREF pixel
xPix1936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[19] VREF PIX_IN[1936] NB2 NB1 CSA_VREF pixel
xPix1937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[19] VREF PIX_IN[1937] NB2 NB1 CSA_VREF pixel
xPix1938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[19] VREF PIX_IN[1938] NB2 NB1 CSA_VREF pixel
xPix1939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[19] VREF PIX_IN[1939] NB2 NB1 CSA_VREF pixel
xPix1940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[19] VREF PIX_IN[1940] NB2 NB1 CSA_VREF pixel
xPix1941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[19] VREF PIX_IN[1941] NB2 NB1 CSA_VREF pixel
xPix1942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[19] VREF PIX_IN[1942] NB2 NB1 CSA_VREF pixel
xPix1943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[19] VREF PIX_IN[1943] NB2 NB1 CSA_VREF pixel
xPix1944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[19] VREF PIX_IN[1944] NB2 NB1 CSA_VREF pixel
xPix1945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[19] VREF PIX_IN[1945] NB2 NB1 CSA_VREF pixel
xPix1946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[19] VREF PIX_IN[1946] NB2 NB1 CSA_VREF pixel
xPix1947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[19] VREF PIX_IN[1947] NB2 NB1 CSA_VREF pixel
xPix1948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[19] VREF PIX_IN[1948] NB2 NB1 CSA_VREF pixel
xPix1949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[19] VREF PIX_IN[1949] NB2 NB1 CSA_VREF pixel
xPix1950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[19] VREF PIX_IN[1950] NB2 NB1 CSA_VREF pixel
xPix1951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[19] VREF PIX_IN[1951] NB2 NB1 CSA_VREF pixel
xPix1952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[19] VREF PIX_IN[1952] NB2 NB1 CSA_VREF pixel
xPix1953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[19] VREF PIX_IN[1953] NB2 NB1 CSA_VREF pixel
xPix1954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[19] VREF PIX_IN[1954] NB2 NB1 CSA_VREF pixel
xPix1955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[19] VREF PIX_IN[1955] NB2 NB1 CSA_VREF pixel
xPix1956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[19] VREF PIX_IN[1956] NB2 NB1 CSA_VREF pixel
xPix1957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[19] VREF PIX_IN[1957] NB2 NB1 CSA_VREF pixel
xPix1958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[19] VREF PIX_IN[1958] NB2 NB1 CSA_VREF pixel
xPix1959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[19] VREF PIX_IN[1959] NB2 NB1 CSA_VREF pixel
xPix1960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[19] VREF PIX_IN[1960] NB2 NB1 CSA_VREF pixel
xPix1961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[19] VREF PIX_IN[1961] NB2 NB1 CSA_VREF pixel
xPix1962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[19] VREF PIX_IN[1962] NB2 NB1 CSA_VREF pixel
xPix1963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[19] VREF PIX_IN[1963] NB2 NB1 CSA_VREF pixel
xPix1964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[19] VREF PIX_IN[1964] NB2 NB1 CSA_VREF pixel
xPix1965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[19] VREF PIX_IN[1965] NB2 NB1 CSA_VREF pixel
xPix1966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[19] VREF PIX_IN[1966] NB2 NB1 CSA_VREF pixel
xPix1967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[19] VREF PIX_IN[1967] NB2 NB1 CSA_VREF pixel
xPix1968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[19] VREF PIX_IN[1968] NB2 NB1 CSA_VREF pixel
xPix1969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[19] VREF PIX_IN[1969] NB2 NB1 CSA_VREF pixel
xPix1970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[19] VREF PIX_IN[1970] NB2 NB1 CSA_VREF pixel
xPix1971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[19] VREF PIX_IN[1971] NB2 NB1 CSA_VREF pixel
xPix1972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[19] VREF PIX_IN[1972] NB2 NB1 CSA_VREF pixel
xPix1973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[19] VREF PIX_IN[1973] NB2 NB1 CSA_VREF pixel
xPix1974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[19] VREF PIX_IN[1974] NB2 NB1 CSA_VREF pixel
xPix1975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[19] VREF PIX_IN[1975] NB2 NB1 CSA_VREF pixel
xPix1976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[19] VREF PIX_IN[1976] NB2 NB1 CSA_VREF pixel
xPix1977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[19] VREF PIX_IN[1977] NB2 NB1 CSA_VREF pixel
xPix1978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[19] VREF PIX_IN[1978] NB2 NB1 CSA_VREF pixel
xPix1979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[19] VREF PIX_IN[1979] NB2 NB1 CSA_VREF pixel
xPix1980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[19] VREF PIX_IN[1980] NB2 NB1 CSA_VREF pixel
xPix1981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[19] VREF PIX_IN[1981] NB2 NB1 CSA_VREF pixel
xPix1982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[19] VREF PIX_IN[1982] NB2 NB1 CSA_VREF pixel
xPix1983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[19] VREF PIX_IN[1983] NB2 NB1 CSA_VREF pixel
xPix1984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[19] VREF PIX_IN[1984] NB2 NB1 CSA_VREF pixel
xPix1985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[19] VREF PIX_IN[1985] NB2 NB1 CSA_VREF pixel
xPix1986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[19] VREF PIX_IN[1986] NB2 NB1 CSA_VREF pixel
xPix1987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[19] VREF PIX_IN[1987] NB2 NB1 CSA_VREF pixel
xPix1988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[19] VREF PIX_IN[1988] NB2 NB1 CSA_VREF pixel
xPix1989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[19] VREF PIX_IN[1989] NB2 NB1 CSA_VREF pixel
xPix1990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[19] VREF PIX_IN[1990] NB2 NB1 CSA_VREF pixel
xPix1991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[19] VREF PIX_IN[1991] NB2 NB1 CSA_VREF pixel
xPix1992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[19] VREF PIX_IN[1992] NB2 NB1 CSA_VREF pixel
xPix1993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[19] VREF PIX_IN[1993] NB2 NB1 CSA_VREF pixel
xPix1994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[19] VREF PIX_IN[1994] NB2 NB1 CSA_VREF pixel
xPix1995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[19] VREF PIX_IN[1995] NB2 NB1 CSA_VREF pixel
xPix1996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[19] VREF PIX_IN[1996] NB2 NB1 CSA_VREF pixel
xPix1997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[19] VREF PIX_IN[1997] NB2 NB1 CSA_VREF pixel
xPix1998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[19] VREF PIX_IN[1998] NB2 NB1 CSA_VREF pixel
xPix1999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[19] VREF PIX_IN[1999] NB2 NB1 CSA_VREF pixel
xPix2000 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[20] VREF PIX_IN[2000] NB2 NB1 CSA_VREF pixel
xPix2001 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[20] VREF PIX_IN[2001] NB2 NB1 CSA_VREF pixel
xPix2002 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[20] VREF PIX_IN[2002] NB2 NB1 CSA_VREF pixel
xPix2003 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[20] VREF PIX_IN[2003] NB2 NB1 CSA_VREF pixel
xPix2004 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[20] VREF PIX_IN[2004] NB2 NB1 CSA_VREF pixel
xPix2005 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[20] VREF PIX_IN[2005] NB2 NB1 CSA_VREF pixel
xPix2006 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[20] VREF PIX_IN[2006] NB2 NB1 CSA_VREF pixel
xPix2007 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[20] VREF PIX_IN[2007] NB2 NB1 CSA_VREF pixel
xPix2008 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[20] VREF PIX_IN[2008] NB2 NB1 CSA_VREF pixel
xPix2009 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[20] VREF PIX_IN[2009] NB2 NB1 CSA_VREF pixel
xPix2010 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[20] VREF PIX_IN[2010] NB2 NB1 CSA_VREF pixel
xPix2011 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[20] VREF PIX_IN[2011] NB2 NB1 CSA_VREF pixel
xPix2012 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[20] VREF PIX_IN[2012] NB2 NB1 CSA_VREF pixel
xPix2013 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[20] VREF PIX_IN[2013] NB2 NB1 CSA_VREF pixel
xPix2014 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[20] VREF PIX_IN[2014] NB2 NB1 CSA_VREF pixel
xPix2015 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[20] VREF PIX_IN[2015] NB2 NB1 CSA_VREF pixel
xPix2016 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[20] VREF PIX_IN[2016] NB2 NB1 CSA_VREF pixel
xPix2017 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[20] VREF PIX_IN[2017] NB2 NB1 CSA_VREF pixel
xPix2018 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[20] VREF PIX_IN[2018] NB2 NB1 CSA_VREF pixel
xPix2019 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[20] VREF PIX_IN[2019] NB2 NB1 CSA_VREF pixel
xPix2020 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[20] VREF PIX_IN[2020] NB2 NB1 CSA_VREF pixel
xPix2021 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[20] VREF PIX_IN[2021] NB2 NB1 CSA_VREF pixel
xPix2022 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[20] VREF PIX_IN[2022] NB2 NB1 CSA_VREF pixel
xPix2023 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[20] VREF PIX_IN[2023] NB2 NB1 CSA_VREF pixel
xPix2024 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[20] VREF PIX_IN[2024] NB2 NB1 CSA_VREF pixel
xPix2025 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[20] VREF PIX_IN[2025] NB2 NB1 CSA_VREF pixel
xPix2026 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[20] VREF PIX_IN[2026] NB2 NB1 CSA_VREF pixel
xPix2027 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[20] VREF PIX_IN[2027] NB2 NB1 CSA_VREF pixel
xPix2028 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[20] VREF PIX_IN[2028] NB2 NB1 CSA_VREF pixel
xPix2029 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[20] VREF PIX_IN[2029] NB2 NB1 CSA_VREF pixel
xPix2030 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[20] VREF PIX_IN[2030] NB2 NB1 CSA_VREF pixel
xPix2031 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[20] VREF PIX_IN[2031] NB2 NB1 CSA_VREF pixel
xPix2032 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[20] VREF PIX_IN[2032] NB2 NB1 CSA_VREF pixel
xPix2033 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[20] VREF PIX_IN[2033] NB2 NB1 CSA_VREF pixel
xPix2034 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[20] VREF PIX_IN[2034] NB2 NB1 CSA_VREF pixel
xPix2035 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[20] VREF PIX_IN[2035] NB2 NB1 CSA_VREF pixel
xPix2036 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[20] VREF PIX_IN[2036] NB2 NB1 CSA_VREF pixel
xPix2037 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[20] VREF PIX_IN[2037] NB2 NB1 CSA_VREF pixel
xPix2038 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[20] VREF PIX_IN[2038] NB2 NB1 CSA_VREF pixel
xPix2039 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[20] VREF PIX_IN[2039] NB2 NB1 CSA_VREF pixel
xPix2040 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[20] VREF PIX_IN[2040] NB2 NB1 CSA_VREF pixel
xPix2041 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[20] VREF PIX_IN[2041] NB2 NB1 CSA_VREF pixel
xPix2042 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[20] VREF PIX_IN[2042] NB2 NB1 CSA_VREF pixel
xPix2043 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[20] VREF PIX_IN[2043] NB2 NB1 CSA_VREF pixel
xPix2044 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[20] VREF PIX_IN[2044] NB2 NB1 CSA_VREF pixel
xPix2045 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[20] VREF PIX_IN[2045] NB2 NB1 CSA_VREF pixel
xPix2046 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[20] VREF PIX_IN[2046] NB2 NB1 CSA_VREF pixel
xPix2047 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[20] VREF PIX_IN[2047] NB2 NB1 CSA_VREF pixel
xPix2048 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[20] VREF PIX_IN[2048] NB2 NB1 CSA_VREF pixel
xPix2049 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[20] VREF PIX_IN[2049] NB2 NB1 CSA_VREF pixel
xPix2050 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[20] VREF PIX_IN[2050] NB2 NB1 CSA_VREF pixel
xPix2051 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[20] VREF PIX_IN[2051] NB2 NB1 CSA_VREF pixel
xPix2052 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[20] VREF PIX_IN[2052] NB2 NB1 CSA_VREF pixel
xPix2053 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[20] VREF PIX_IN[2053] NB2 NB1 CSA_VREF pixel
xPix2054 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[20] VREF PIX_IN[2054] NB2 NB1 CSA_VREF pixel
xPix2055 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[20] VREF PIX_IN[2055] NB2 NB1 CSA_VREF pixel
xPix2056 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[20] VREF PIX_IN[2056] NB2 NB1 CSA_VREF pixel
xPix2057 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[20] VREF PIX_IN[2057] NB2 NB1 CSA_VREF pixel
xPix2058 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[20] VREF PIX_IN[2058] NB2 NB1 CSA_VREF pixel
xPix2059 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[20] VREF PIX_IN[2059] NB2 NB1 CSA_VREF pixel
xPix2060 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[20] VREF PIX_IN[2060] NB2 NB1 CSA_VREF pixel
xPix2061 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[20] VREF PIX_IN[2061] NB2 NB1 CSA_VREF pixel
xPix2062 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[20] VREF PIX_IN[2062] NB2 NB1 CSA_VREF pixel
xPix2063 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[20] VREF PIX_IN[2063] NB2 NB1 CSA_VREF pixel
xPix2064 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[20] VREF PIX_IN[2064] NB2 NB1 CSA_VREF pixel
xPix2065 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[20] VREF PIX_IN[2065] NB2 NB1 CSA_VREF pixel
xPix2066 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[20] VREF PIX_IN[2066] NB2 NB1 CSA_VREF pixel
xPix2067 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[20] VREF PIX_IN[2067] NB2 NB1 CSA_VREF pixel
xPix2068 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[20] VREF PIX_IN[2068] NB2 NB1 CSA_VREF pixel
xPix2069 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[20] VREF PIX_IN[2069] NB2 NB1 CSA_VREF pixel
xPix2070 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[20] VREF PIX_IN[2070] NB2 NB1 CSA_VREF pixel
xPix2071 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[20] VREF PIX_IN[2071] NB2 NB1 CSA_VREF pixel
xPix2072 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[20] VREF PIX_IN[2072] NB2 NB1 CSA_VREF pixel
xPix2073 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[20] VREF PIX_IN[2073] NB2 NB1 CSA_VREF pixel
xPix2074 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[20] VREF PIX_IN[2074] NB2 NB1 CSA_VREF pixel
xPix2075 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[20] VREF PIX_IN[2075] NB2 NB1 CSA_VREF pixel
xPix2076 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[20] VREF PIX_IN[2076] NB2 NB1 CSA_VREF pixel
xPix2077 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[20] VREF PIX_IN[2077] NB2 NB1 CSA_VREF pixel
xPix2078 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[20] VREF PIX_IN[2078] NB2 NB1 CSA_VREF pixel
xPix2079 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[20] VREF PIX_IN[2079] NB2 NB1 CSA_VREF pixel
xPix2080 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[20] VREF PIX_IN[2080] NB2 NB1 CSA_VREF pixel
xPix2081 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[20] VREF PIX_IN[2081] NB2 NB1 CSA_VREF pixel
xPix2082 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[20] VREF PIX_IN[2082] NB2 NB1 CSA_VREF pixel
xPix2083 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[20] VREF PIX_IN[2083] NB2 NB1 CSA_VREF pixel
xPix2084 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[20] VREF PIX_IN[2084] NB2 NB1 CSA_VREF pixel
xPix2085 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[20] VREF PIX_IN[2085] NB2 NB1 CSA_VREF pixel
xPix2086 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[20] VREF PIX_IN[2086] NB2 NB1 CSA_VREF pixel
xPix2087 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[20] VREF PIX_IN[2087] NB2 NB1 CSA_VREF pixel
xPix2088 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[20] VREF PIX_IN[2088] NB2 NB1 CSA_VREF pixel
xPix2089 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[20] VREF PIX_IN[2089] NB2 NB1 CSA_VREF pixel
xPix2090 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[20] VREF PIX_IN[2090] NB2 NB1 CSA_VREF pixel
xPix2091 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[20] VREF PIX_IN[2091] NB2 NB1 CSA_VREF pixel
xPix2092 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[20] VREF PIX_IN[2092] NB2 NB1 CSA_VREF pixel
xPix2093 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[20] VREF PIX_IN[2093] NB2 NB1 CSA_VREF pixel
xPix2094 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[20] VREF PIX_IN[2094] NB2 NB1 CSA_VREF pixel
xPix2095 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[20] VREF PIX_IN[2095] NB2 NB1 CSA_VREF pixel
xPix2096 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[20] VREF PIX_IN[2096] NB2 NB1 CSA_VREF pixel
xPix2097 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[20] VREF PIX_IN[2097] NB2 NB1 CSA_VREF pixel
xPix2098 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[20] VREF PIX_IN[2098] NB2 NB1 CSA_VREF pixel
xPix2099 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[20] VREF PIX_IN[2099] NB2 NB1 CSA_VREF pixel
xPix2100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[21] VREF PIX_IN[2100] NB2 NB1 CSA_VREF pixel
xPix2101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[21] VREF PIX_IN[2101] NB2 NB1 CSA_VREF pixel
xPix2102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[21] VREF PIX_IN[2102] NB2 NB1 CSA_VREF pixel
xPix2103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[21] VREF PIX_IN[2103] NB2 NB1 CSA_VREF pixel
xPix2104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[21] VREF PIX_IN[2104] NB2 NB1 CSA_VREF pixel
xPix2105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[21] VREF PIX_IN[2105] NB2 NB1 CSA_VREF pixel
xPix2106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[21] VREF PIX_IN[2106] NB2 NB1 CSA_VREF pixel
xPix2107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[21] VREF PIX_IN[2107] NB2 NB1 CSA_VREF pixel
xPix2108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[21] VREF PIX_IN[2108] NB2 NB1 CSA_VREF pixel
xPix2109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[21] VREF PIX_IN[2109] NB2 NB1 CSA_VREF pixel
xPix2110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[21] VREF PIX_IN[2110] NB2 NB1 CSA_VREF pixel
xPix2111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[21] VREF PIX_IN[2111] NB2 NB1 CSA_VREF pixel
xPix2112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[21] VREF PIX_IN[2112] NB2 NB1 CSA_VREF pixel
xPix2113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[21] VREF PIX_IN[2113] NB2 NB1 CSA_VREF pixel
xPix2114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[21] VREF PIX_IN[2114] NB2 NB1 CSA_VREF pixel
xPix2115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[21] VREF PIX_IN[2115] NB2 NB1 CSA_VREF pixel
xPix2116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[21] VREF PIX_IN[2116] NB2 NB1 CSA_VREF pixel
xPix2117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[21] VREF PIX_IN[2117] NB2 NB1 CSA_VREF pixel
xPix2118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[21] VREF PIX_IN[2118] NB2 NB1 CSA_VREF pixel
xPix2119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[21] VREF PIX_IN[2119] NB2 NB1 CSA_VREF pixel
xPix2120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[21] VREF PIX_IN[2120] NB2 NB1 CSA_VREF pixel
xPix2121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[21] VREF PIX_IN[2121] NB2 NB1 CSA_VREF pixel
xPix2122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[21] VREF PIX_IN[2122] NB2 NB1 CSA_VREF pixel
xPix2123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[21] VREF PIX_IN[2123] NB2 NB1 CSA_VREF pixel
xPix2124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[21] VREF PIX_IN[2124] NB2 NB1 CSA_VREF pixel
xPix2125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[21] VREF PIX_IN[2125] NB2 NB1 CSA_VREF pixel
xPix2126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[21] VREF PIX_IN[2126] NB2 NB1 CSA_VREF pixel
xPix2127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[21] VREF PIX_IN[2127] NB2 NB1 CSA_VREF pixel
xPix2128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[21] VREF PIX_IN[2128] NB2 NB1 CSA_VREF pixel
xPix2129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[21] VREF PIX_IN[2129] NB2 NB1 CSA_VREF pixel
xPix2130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[21] VREF PIX_IN[2130] NB2 NB1 CSA_VREF pixel
xPix2131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[21] VREF PIX_IN[2131] NB2 NB1 CSA_VREF pixel
xPix2132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[21] VREF PIX_IN[2132] NB2 NB1 CSA_VREF pixel
xPix2133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[21] VREF PIX_IN[2133] NB2 NB1 CSA_VREF pixel
xPix2134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[21] VREF PIX_IN[2134] NB2 NB1 CSA_VREF pixel
xPix2135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[21] VREF PIX_IN[2135] NB2 NB1 CSA_VREF pixel
xPix2136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[21] VREF PIX_IN[2136] NB2 NB1 CSA_VREF pixel
xPix2137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[21] VREF PIX_IN[2137] NB2 NB1 CSA_VREF pixel
xPix2138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[21] VREF PIX_IN[2138] NB2 NB1 CSA_VREF pixel
xPix2139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[21] VREF PIX_IN[2139] NB2 NB1 CSA_VREF pixel
xPix2140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[21] VREF PIX_IN[2140] NB2 NB1 CSA_VREF pixel
xPix2141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[21] VREF PIX_IN[2141] NB2 NB1 CSA_VREF pixel
xPix2142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[21] VREF PIX_IN[2142] NB2 NB1 CSA_VREF pixel
xPix2143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[21] VREF PIX_IN[2143] NB2 NB1 CSA_VREF pixel
xPix2144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[21] VREF PIX_IN[2144] NB2 NB1 CSA_VREF pixel
xPix2145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[21] VREF PIX_IN[2145] NB2 NB1 CSA_VREF pixel
xPix2146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[21] VREF PIX_IN[2146] NB2 NB1 CSA_VREF pixel
xPix2147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[21] VREF PIX_IN[2147] NB2 NB1 CSA_VREF pixel
xPix2148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[21] VREF PIX_IN[2148] NB2 NB1 CSA_VREF pixel
xPix2149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[21] VREF PIX_IN[2149] NB2 NB1 CSA_VREF pixel
xPix2150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[21] VREF PIX_IN[2150] NB2 NB1 CSA_VREF pixel
xPix2151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[21] VREF PIX_IN[2151] NB2 NB1 CSA_VREF pixel
xPix2152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[21] VREF PIX_IN[2152] NB2 NB1 CSA_VREF pixel
xPix2153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[21] VREF PIX_IN[2153] NB2 NB1 CSA_VREF pixel
xPix2154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[21] VREF PIX_IN[2154] NB2 NB1 CSA_VREF pixel
xPix2155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[21] VREF PIX_IN[2155] NB2 NB1 CSA_VREF pixel
xPix2156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[21] VREF PIX_IN[2156] NB2 NB1 CSA_VREF pixel
xPix2157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[21] VREF PIX_IN[2157] NB2 NB1 CSA_VREF pixel
xPix2158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[21] VREF PIX_IN[2158] NB2 NB1 CSA_VREF pixel
xPix2159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[21] VREF PIX_IN[2159] NB2 NB1 CSA_VREF pixel
xPix2160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[21] VREF PIX_IN[2160] NB2 NB1 CSA_VREF pixel
xPix2161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[21] VREF PIX_IN[2161] NB2 NB1 CSA_VREF pixel
xPix2162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[21] VREF PIX_IN[2162] NB2 NB1 CSA_VREF pixel
xPix2163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[21] VREF PIX_IN[2163] NB2 NB1 CSA_VREF pixel
xPix2164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[21] VREF PIX_IN[2164] NB2 NB1 CSA_VREF pixel
xPix2165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[21] VREF PIX_IN[2165] NB2 NB1 CSA_VREF pixel
xPix2166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[21] VREF PIX_IN[2166] NB2 NB1 CSA_VREF pixel
xPix2167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[21] VREF PIX_IN[2167] NB2 NB1 CSA_VREF pixel
xPix2168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[21] VREF PIX_IN[2168] NB2 NB1 CSA_VREF pixel
xPix2169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[21] VREF PIX_IN[2169] NB2 NB1 CSA_VREF pixel
xPix2170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[21] VREF PIX_IN[2170] NB2 NB1 CSA_VREF pixel
xPix2171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[21] VREF PIX_IN[2171] NB2 NB1 CSA_VREF pixel
xPix2172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[21] VREF PIX_IN[2172] NB2 NB1 CSA_VREF pixel
xPix2173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[21] VREF PIX_IN[2173] NB2 NB1 CSA_VREF pixel
xPix2174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[21] VREF PIX_IN[2174] NB2 NB1 CSA_VREF pixel
xPix2175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[21] VREF PIX_IN[2175] NB2 NB1 CSA_VREF pixel
xPix2176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[21] VREF PIX_IN[2176] NB2 NB1 CSA_VREF pixel
xPix2177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[21] VREF PIX_IN[2177] NB2 NB1 CSA_VREF pixel
xPix2178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[21] VREF PIX_IN[2178] NB2 NB1 CSA_VREF pixel
xPix2179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[21] VREF PIX_IN[2179] NB2 NB1 CSA_VREF pixel
xPix2180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[21] VREF PIX_IN[2180] NB2 NB1 CSA_VREF pixel
xPix2181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[21] VREF PIX_IN[2181] NB2 NB1 CSA_VREF pixel
xPix2182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[21] VREF PIX_IN[2182] NB2 NB1 CSA_VREF pixel
xPix2183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[21] VREF PIX_IN[2183] NB2 NB1 CSA_VREF pixel
xPix2184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[21] VREF PIX_IN[2184] NB2 NB1 CSA_VREF pixel
xPix2185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[21] VREF PIX_IN[2185] NB2 NB1 CSA_VREF pixel
xPix2186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[21] VREF PIX_IN[2186] NB2 NB1 CSA_VREF pixel
xPix2187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[21] VREF PIX_IN[2187] NB2 NB1 CSA_VREF pixel
xPix2188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[21] VREF PIX_IN[2188] NB2 NB1 CSA_VREF pixel
xPix2189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[21] VREF PIX_IN[2189] NB2 NB1 CSA_VREF pixel
xPix2190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[21] VREF PIX_IN[2190] NB2 NB1 CSA_VREF pixel
xPix2191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[21] VREF PIX_IN[2191] NB2 NB1 CSA_VREF pixel
xPix2192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[21] VREF PIX_IN[2192] NB2 NB1 CSA_VREF pixel
xPix2193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[21] VREF PIX_IN[2193] NB2 NB1 CSA_VREF pixel
xPix2194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[21] VREF PIX_IN[2194] NB2 NB1 CSA_VREF pixel
xPix2195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[21] VREF PIX_IN[2195] NB2 NB1 CSA_VREF pixel
xPix2196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[21] VREF PIX_IN[2196] NB2 NB1 CSA_VREF pixel
xPix2197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[21] VREF PIX_IN[2197] NB2 NB1 CSA_VREF pixel
xPix2198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[21] VREF PIX_IN[2198] NB2 NB1 CSA_VREF pixel
xPix2199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[21] VREF PIX_IN[2199] NB2 NB1 CSA_VREF pixel
xPix2200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[22] VREF PIX_IN[2200] NB2 NB1 CSA_VREF pixel
xPix2201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[22] VREF PIX_IN[2201] NB2 NB1 CSA_VREF pixel
xPix2202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[22] VREF PIX_IN[2202] NB2 NB1 CSA_VREF pixel
xPix2203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[22] VREF PIX_IN[2203] NB2 NB1 CSA_VREF pixel
xPix2204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[22] VREF PIX_IN[2204] NB2 NB1 CSA_VREF pixel
xPix2205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[22] VREF PIX_IN[2205] NB2 NB1 CSA_VREF pixel
xPix2206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[22] VREF PIX_IN[2206] NB2 NB1 CSA_VREF pixel
xPix2207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[22] VREF PIX_IN[2207] NB2 NB1 CSA_VREF pixel
xPix2208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[22] VREF PIX_IN[2208] NB2 NB1 CSA_VREF pixel
xPix2209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[22] VREF PIX_IN[2209] NB2 NB1 CSA_VREF pixel
xPix2210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[22] VREF PIX_IN[2210] NB2 NB1 CSA_VREF pixel
xPix2211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[22] VREF PIX_IN[2211] NB2 NB1 CSA_VREF pixel
xPix2212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[22] VREF PIX_IN[2212] NB2 NB1 CSA_VREF pixel
xPix2213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[22] VREF PIX_IN[2213] NB2 NB1 CSA_VREF pixel
xPix2214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[22] VREF PIX_IN[2214] NB2 NB1 CSA_VREF pixel
xPix2215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[22] VREF PIX_IN[2215] NB2 NB1 CSA_VREF pixel
xPix2216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[22] VREF PIX_IN[2216] NB2 NB1 CSA_VREF pixel
xPix2217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[22] VREF PIX_IN[2217] NB2 NB1 CSA_VREF pixel
xPix2218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[22] VREF PIX_IN[2218] NB2 NB1 CSA_VREF pixel
xPix2219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[22] VREF PIX_IN[2219] NB2 NB1 CSA_VREF pixel
xPix2220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[22] VREF PIX_IN[2220] NB2 NB1 CSA_VREF pixel
xPix2221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[22] VREF PIX_IN[2221] NB2 NB1 CSA_VREF pixel
xPix2222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[22] VREF PIX_IN[2222] NB2 NB1 CSA_VREF pixel
xPix2223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[22] VREF PIX_IN[2223] NB2 NB1 CSA_VREF pixel
xPix2224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[22] VREF PIX_IN[2224] NB2 NB1 CSA_VREF pixel
xPix2225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[22] VREF PIX_IN[2225] NB2 NB1 CSA_VREF pixel
xPix2226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[22] VREF PIX_IN[2226] NB2 NB1 CSA_VREF pixel
xPix2227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[22] VREF PIX_IN[2227] NB2 NB1 CSA_VREF pixel
xPix2228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[22] VREF PIX_IN[2228] NB2 NB1 CSA_VREF pixel
xPix2229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[22] VREF PIX_IN[2229] NB2 NB1 CSA_VREF pixel
xPix2230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[22] VREF PIX_IN[2230] NB2 NB1 CSA_VREF pixel
xPix2231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[22] VREF PIX_IN[2231] NB2 NB1 CSA_VREF pixel
xPix2232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[22] VREF PIX_IN[2232] NB2 NB1 CSA_VREF pixel
xPix2233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[22] VREF PIX_IN[2233] NB2 NB1 CSA_VREF pixel
xPix2234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[22] VREF PIX_IN[2234] NB2 NB1 CSA_VREF pixel
xPix2235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[22] VREF PIX_IN[2235] NB2 NB1 CSA_VREF pixel
xPix2236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[22] VREF PIX_IN[2236] NB2 NB1 CSA_VREF pixel
xPix2237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[22] VREF PIX_IN[2237] NB2 NB1 CSA_VREF pixel
xPix2238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[22] VREF PIX_IN[2238] NB2 NB1 CSA_VREF pixel
xPix2239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[22] VREF PIX_IN[2239] NB2 NB1 CSA_VREF pixel
xPix2240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[22] VREF PIX_IN[2240] NB2 NB1 CSA_VREF pixel
xPix2241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[22] VREF PIX_IN[2241] NB2 NB1 CSA_VREF pixel
xPix2242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[22] VREF PIX_IN[2242] NB2 NB1 CSA_VREF pixel
xPix2243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[22] VREF PIX_IN[2243] NB2 NB1 CSA_VREF pixel
xPix2244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[22] VREF PIX_IN[2244] NB2 NB1 CSA_VREF pixel
xPix2245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[22] VREF PIX_IN[2245] NB2 NB1 CSA_VREF pixel
xPix2246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[22] VREF PIX_IN[2246] NB2 NB1 CSA_VREF pixel
xPix2247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[22] VREF PIX_IN[2247] NB2 NB1 CSA_VREF pixel
xPix2248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[22] VREF PIX_IN[2248] NB2 NB1 CSA_VREF pixel
xPix2249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[22] VREF PIX_IN[2249] NB2 NB1 CSA_VREF pixel
xPix2250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[22] VREF PIX_IN[2250] NB2 NB1 CSA_VREF pixel
xPix2251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[22] VREF PIX_IN[2251] NB2 NB1 CSA_VREF pixel
xPix2252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[22] VREF PIX_IN[2252] NB2 NB1 CSA_VREF pixel
xPix2253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[22] VREF PIX_IN[2253] NB2 NB1 CSA_VREF pixel
xPix2254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[22] VREF PIX_IN[2254] NB2 NB1 CSA_VREF pixel
xPix2255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[22] VREF PIX_IN[2255] NB2 NB1 CSA_VREF pixel
xPix2256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[22] VREF PIX_IN[2256] NB2 NB1 CSA_VREF pixel
xPix2257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[22] VREF PIX_IN[2257] NB2 NB1 CSA_VREF pixel
xPix2258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[22] VREF PIX_IN[2258] NB2 NB1 CSA_VREF pixel
xPix2259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[22] VREF PIX_IN[2259] NB2 NB1 CSA_VREF pixel
xPix2260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[22] VREF PIX_IN[2260] NB2 NB1 CSA_VREF pixel
xPix2261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[22] VREF PIX_IN[2261] NB2 NB1 CSA_VREF pixel
xPix2262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[22] VREF PIX_IN[2262] NB2 NB1 CSA_VREF pixel
xPix2263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[22] VREF PIX_IN[2263] NB2 NB1 CSA_VREF pixel
xPix2264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[22] VREF PIX_IN[2264] NB2 NB1 CSA_VREF pixel
xPix2265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[22] VREF PIX_IN[2265] NB2 NB1 CSA_VREF pixel
xPix2266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[22] VREF PIX_IN[2266] NB2 NB1 CSA_VREF pixel
xPix2267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[22] VREF PIX_IN[2267] NB2 NB1 CSA_VREF pixel
xPix2268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[22] VREF PIX_IN[2268] NB2 NB1 CSA_VREF pixel
xPix2269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[22] VREF PIX_IN[2269] NB2 NB1 CSA_VREF pixel
xPix2270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[22] VREF PIX_IN[2270] NB2 NB1 CSA_VREF pixel
xPix2271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[22] VREF PIX_IN[2271] NB2 NB1 CSA_VREF pixel
xPix2272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[22] VREF PIX_IN[2272] NB2 NB1 CSA_VREF pixel
xPix2273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[22] VREF PIX_IN[2273] NB2 NB1 CSA_VREF pixel
xPix2274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[22] VREF PIX_IN[2274] NB2 NB1 CSA_VREF pixel
xPix2275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[22] VREF PIX_IN[2275] NB2 NB1 CSA_VREF pixel
xPix2276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[22] VREF PIX_IN[2276] NB2 NB1 CSA_VREF pixel
xPix2277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[22] VREF PIX_IN[2277] NB2 NB1 CSA_VREF pixel
xPix2278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[22] VREF PIX_IN[2278] NB2 NB1 CSA_VREF pixel
xPix2279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[22] VREF PIX_IN[2279] NB2 NB1 CSA_VREF pixel
xPix2280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[22] VREF PIX_IN[2280] NB2 NB1 CSA_VREF pixel
xPix2281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[22] VREF PIX_IN[2281] NB2 NB1 CSA_VREF pixel
xPix2282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[22] VREF PIX_IN[2282] NB2 NB1 CSA_VREF pixel
xPix2283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[22] VREF PIX_IN[2283] NB2 NB1 CSA_VREF pixel
xPix2284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[22] VREF PIX_IN[2284] NB2 NB1 CSA_VREF pixel
xPix2285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[22] VREF PIX_IN[2285] NB2 NB1 CSA_VREF pixel
xPix2286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[22] VREF PIX_IN[2286] NB2 NB1 CSA_VREF pixel
xPix2287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[22] VREF PIX_IN[2287] NB2 NB1 CSA_VREF pixel
xPix2288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[22] VREF PIX_IN[2288] NB2 NB1 CSA_VREF pixel
xPix2289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[22] VREF PIX_IN[2289] NB2 NB1 CSA_VREF pixel
xPix2290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[22] VREF PIX_IN[2290] NB2 NB1 CSA_VREF pixel
xPix2291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[22] VREF PIX_IN[2291] NB2 NB1 CSA_VREF pixel
xPix2292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[22] VREF PIX_IN[2292] NB2 NB1 CSA_VREF pixel
xPix2293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[22] VREF PIX_IN[2293] NB2 NB1 CSA_VREF pixel
xPix2294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[22] VREF PIX_IN[2294] NB2 NB1 CSA_VREF pixel
xPix2295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[22] VREF PIX_IN[2295] NB2 NB1 CSA_VREF pixel
xPix2296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[22] VREF PIX_IN[2296] NB2 NB1 CSA_VREF pixel
xPix2297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[22] VREF PIX_IN[2297] NB2 NB1 CSA_VREF pixel
xPix2298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[22] VREF PIX_IN[2298] NB2 NB1 CSA_VREF pixel
xPix2299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[22] VREF PIX_IN[2299] NB2 NB1 CSA_VREF pixel
xPix2300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[23] VREF PIX_IN[2300] NB2 NB1 CSA_VREF pixel
xPix2301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[23] VREF PIX_IN[2301] NB2 NB1 CSA_VREF pixel
xPix2302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[23] VREF PIX_IN[2302] NB2 NB1 CSA_VREF pixel
xPix2303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[23] VREF PIX_IN[2303] NB2 NB1 CSA_VREF pixel
xPix2304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[23] VREF PIX_IN[2304] NB2 NB1 CSA_VREF pixel
xPix2305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[23] VREF PIX_IN[2305] NB2 NB1 CSA_VREF pixel
xPix2306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[23] VREF PIX_IN[2306] NB2 NB1 CSA_VREF pixel
xPix2307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[23] VREF PIX_IN[2307] NB2 NB1 CSA_VREF pixel
xPix2308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[23] VREF PIX_IN[2308] NB2 NB1 CSA_VREF pixel
xPix2309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[23] VREF PIX_IN[2309] NB2 NB1 CSA_VREF pixel
xPix2310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[23] VREF PIX_IN[2310] NB2 NB1 CSA_VREF pixel
xPix2311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[23] VREF PIX_IN[2311] NB2 NB1 CSA_VREF pixel
xPix2312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[23] VREF PIX_IN[2312] NB2 NB1 CSA_VREF pixel
xPix2313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[23] VREF PIX_IN[2313] NB2 NB1 CSA_VREF pixel
xPix2314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[23] VREF PIX_IN[2314] NB2 NB1 CSA_VREF pixel
xPix2315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[23] VREF PIX_IN[2315] NB2 NB1 CSA_VREF pixel
xPix2316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[23] VREF PIX_IN[2316] NB2 NB1 CSA_VREF pixel
xPix2317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[23] VREF PIX_IN[2317] NB2 NB1 CSA_VREF pixel
xPix2318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[23] VREF PIX_IN[2318] NB2 NB1 CSA_VREF pixel
xPix2319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[23] VREF PIX_IN[2319] NB2 NB1 CSA_VREF pixel
xPix2320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[23] VREF PIX_IN[2320] NB2 NB1 CSA_VREF pixel
xPix2321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[23] VREF PIX_IN[2321] NB2 NB1 CSA_VREF pixel
xPix2322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[23] VREF PIX_IN[2322] NB2 NB1 CSA_VREF pixel
xPix2323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[23] VREF PIX_IN[2323] NB2 NB1 CSA_VREF pixel
xPix2324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[23] VREF PIX_IN[2324] NB2 NB1 CSA_VREF pixel
xPix2325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[23] VREF PIX_IN[2325] NB2 NB1 CSA_VREF pixel
xPix2326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[23] VREF PIX_IN[2326] NB2 NB1 CSA_VREF pixel
xPix2327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[23] VREF PIX_IN[2327] NB2 NB1 CSA_VREF pixel
xPix2328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[23] VREF PIX_IN[2328] NB2 NB1 CSA_VREF pixel
xPix2329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[23] VREF PIX_IN[2329] NB2 NB1 CSA_VREF pixel
xPix2330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[23] VREF PIX_IN[2330] NB2 NB1 CSA_VREF pixel
xPix2331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[23] VREF PIX_IN[2331] NB2 NB1 CSA_VREF pixel
xPix2332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[23] VREF PIX_IN[2332] NB2 NB1 CSA_VREF pixel
xPix2333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[23] VREF PIX_IN[2333] NB2 NB1 CSA_VREF pixel
xPix2334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[23] VREF PIX_IN[2334] NB2 NB1 CSA_VREF pixel
xPix2335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[23] VREF PIX_IN[2335] NB2 NB1 CSA_VREF pixel
xPix2336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[23] VREF PIX_IN[2336] NB2 NB1 CSA_VREF pixel
xPix2337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[23] VREF PIX_IN[2337] NB2 NB1 CSA_VREF pixel
xPix2338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[23] VREF PIX_IN[2338] NB2 NB1 CSA_VREF pixel
xPix2339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[23] VREF PIX_IN[2339] NB2 NB1 CSA_VREF pixel
xPix2340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[23] VREF PIX_IN[2340] NB2 NB1 CSA_VREF pixel
xPix2341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[23] VREF PIX_IN[2341] NB2 NB1 CSA_VREF pixel
xPix2342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[23] VREF PIX_IN[2342] NB2 NB1 CSA_VREF pixel
xPix2343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[23] VREF PIX_IN[2343] NB2 NB1 CSA_VREF pixel
xPix2344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[23] VREF PIX_IN[2344] NB2 NB1 CSA_VREF pixel
xPix2345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[23] VREF PIX_IN[2345] NB2 NB1 CSA_VREF pixel
xPix2346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[23] VREF PIX_IN[2346] NB2 NB1 CSA_VREF pixel
xPix2347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[23] VREF PIX_IN[2347] NB2 NB1 CSA_VREF pixel
xPix2348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[23] VREF PIX_IN[2348] NB2 NB1 CSA_VREF pixel
xPix2349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[23] VREF PIX_IN[2349] NB2 NB1 CSA_VREF pixel
xPix2350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[23] VREF PIX_IN[2350] NB2 NB1 CSA_VREF pixel
xPix2351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[23] VREF PIX_IN[2351] NB2 NB1 CSA_VREF pixel
xPix2352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[23] VREF PIX_IN[2352] NB2 NB1 CSA_VREF pixel
xPix2353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[23] VREF PIX_IN[2353] NB2 NB1 CSA_VREF pixel
xPix2354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[23] VREF PIX_IN[2354] NB2 NB1 CSA_VREF pixel
xPix2355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[23] VREF PIX_IN[2355] NB2 NB1 CSA_VREF pixel
xPix2356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[23] VREF PIX_IN[2356] NB2 NB1 CSA_VREF pixel
xPix2357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[23] VREF PIX_IN[2357] NB2 NB1 CSA_VREF pixel
xPix2358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[23] VREF PIX_IN[2358] NB2 NB1 CSA_VREF pixel
xPix2359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[23] VREF PIX_IN[2359] NB2 NB1 CSA_VREF pixel
xPix2360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[23] VREF PIX_IN[2360] NB2 NB1 CSA_VREF pixel
xPix2361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[23] VREF PIX_IN[2361] NB2 NB1 CSA_VREF pixel
xPix2362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[23] VREF PIX_IN[2362] NB2 NB1 CSA_VREF pixel
xPix2363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[23] VREF PIX_IN[2363] NB2 NB1 CSA_VREF pixel
xPix2364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[23] VREF PIX_IN[2364] NB2 NB1 CSA_VREF pixel
xPix2365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[23] VREF PIX_IN[2365] NB2 NB1 CSA_VREF pixel
xPix2366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[23] VREF PIX_IN[2366] NB2 NB1 CSA_VREF pixel
xPix2367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[23] VREF PIX_IN[2367] NB2 NB1 CSA_VREF pixel
xPix2368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[23] VREF PIX_IN[2368] NB2 NB1 CSA_VREF pixel
xPix2369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[23] VREF PIX_IN[2369] NB2 NB1 CSA_VREF pixel
xPix2370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[23] VREF PIX_IN[2370] NB2 NB1 CSA_VREF pixel
xPix2371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[23] VREF PIX_IN[2371] NB2 NB1 CSA_VREF pixel
xPix2372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[23] VREF PIX_IN[2372] NB2 NB1 CSA_VREF pixel
xPix2373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[23] VREF PIX_IN[2373] NB2 NB1 CSA_VREF pixel
xPix2374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[23] VREF PIX_IN[2374] NB2 NB1 CSA_VREF pixel
xPix2375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[23] VREF PIX_IN[2375] NB2 NB1 CSA_VREF pixel
xPix2376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[23] VREF PIX_IN[2376] NB2 NB1 CSA_VREF pixel
xPix2377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[23] VREF PIX_IN[2377] NB2 NB1 CSA_VREF pixel
xPix2378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[23] VREF PIX_IN[2378] NB2 NB1 CSA_VREF pixel
xPix2379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[23] VREF PIX_IN[2379] NB2 NB1 CSA_VREF pixel
xPix2380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[23] VREF PIX_IN[2380] NB2 NB1 CSA_VREF pixel
xPix2381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[23] VREF PIX_IN[2381] NB2 NB1 CSA_VREF pixel
xPix2382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[23] VREF PIX_IN[2382] NB2 NB1 CSA_VREF pixel
xPix2383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[23] VREF PIX_IN[2383] NB2 NB1 CSA_VREF pixel
xPix2384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[23] VREF PIX_IN[2384] NB2 NB1 CSA_VREF pixel
xPix2385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[23] VREF PIX_IN[2385] NB2 NB1 CSA_VREF pixel
xPix2386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[23] VREF PIX_IN[2386] NB2 NB1 CSA_VREF pixel
xPix2387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[23] VREF PIX_IN[2387] NB2 NB1 CSA_VREF pixel
xPix2388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[23] VREF PIX_IN[2388] NB2 NB1 CSA_VREF pixel
xPix2389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[23] VREF PIX_IN[2389] NB2 NB1 CSA_VREF pixel
xPix2390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[23] VREF PIX_IN[2390] NB2 NB1 CSA_VREF pixel
xPix2391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[23] VREF PIX_IN[2391] NB2 NB1 CSA_VREF pixel
xPix2392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[23] VREF PIX_IN[2392] NB2 NB1 CSA_VREF pixel
xPix2393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[23] VREF PIX_IN[2393] NB2 NB1 CSA_VREF pixel
xPix2394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[23] VREF PIX_IN[2394] NB2 NB1 CSA_VREF pixel
xPix2395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[23] VREF PIX_IN[2395] NB2 NB1 CSA_VREF pixel
xPix2396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[23] VREF PIX_IN[2396] NB2 NB1 CSA_VREF pixel
xPix2397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[23] VREF PIX_IN[2397] NB2 NB1 CSA_VREF pixel
xPix2398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[23] VREF PIX_IN[2398] NB2 NB1 CSA_VREF pixel
xPix2399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[23] VREF PIX_IN[2399] NB2 NB1 CSA_VREF pixel
xPix2400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[24] VREF PIX_IN[2400] NB2 NB1 CSA_VREF pixel
xPix2401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[24] VREF PIX_IN[2401] NB2 NB1 CSA_VREF pixel
xPix2402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[24] VREF PIX_IN[2402] NB2 NB1 CSA_VREF pixel
xPix2403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[24] VREF PIX_IN[2403] NB2 NB1 CSA_VREF pixel
xPix2404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[24] VREF PIX_IN[2404] NB2 NB1 CSA_VREF pixel
xPix2405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[24] VREF PIX_IN[2405] NB2 NB1 CSA_VREF pixel
xPix2406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[24] VREF PIX_IN[2406] NB2 NB1 CSA_VREF pixel
xPix2407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[24] VREF PIX_IN[2407] NB2 NB1 CSA_VREF pixel
xPix2408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[24] VREF PIX_IN[2408] NB2 NB1 CSA_VREF pixel
xPix2409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[24] VREF PIX_IN[2409] NB2 NB1 CSA_VREF pixel
xPix2410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[24] VREF PIX_IN[2410] NB2 NB1 CSA_VREF pixel
xPix2411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[24] VREF PIX_IN[2411] NB2 NB1 CSA_VREF pixel
xPix2412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[24] VREF PIX_IN[2412] NB2 NB1 CSA_VREF pixel
xPix2413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[24] VREF PIX_IN[2413] NB2 NB1 CSA_VREF pixel
xPix2414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[24] VREF PIX_IN[2414] NB2 NB1 CSA_VREF pixel
xPix2415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[24] VREF PIX_IN[2415] NB2 NB1 CSA_VREF pixel
xPix2416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[24] VREF PIX_IN[2416] NB2 NB1 CSA_VREF pixel
xPix2417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[24] VREF PIX_IN[2417] NB2 NB1 CSA_VREF pixel
xPix2418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[24] VREF PIX_IN[2418] NB2 NB1 CSA_VREF pixel
xPix2419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[24] VREF PIX_IN[2419] NB2 NB1 CSA_VREF pixel
xPix2420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[24] VREF PIX_IN[2420] NB2 NB1 CSA_VREF pixel
xPix2421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[24] VREF PIX_IN[2421] NB2 NB1 CSA_VREF pixel
xPix2422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[24] VREF PIX_IN[2422] NB2 NB1 CSA_VREF pixel
xPix2423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[24] VREF PIX_IN[2423] NB2 NB1 CSA_VREF pixel
xPix2424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[24] VREF PIX_IN[2424] NB2 NB1 CSA_VREF pixel
xPix2425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[24] VREF PIX_IN[2425] NB2 NB1 CSA_VREF pixel
xPix2426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[24] VREF PIX_IN[2426] NB2 NB1 CSA_VREF pixel
xPix2427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[24] VREF PIX_IN[2427] NB2 NB1 CSA_VREF pixel
xPix2428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[24] VREF PIX_IN[2428] NB2 NB1 CSA_VREF pixel
xPix2429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[24] VREF PIX_IN[2429] NB2 NB1 CSA_VREF pixel
xPix2430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[24] VREF PIX_IN[2430] NB2 NB1 CSA_VREF pixel
xPix2431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[24] VREF PIX_IN[2431] NB2 NB1 CSA_VREF pixel
xPix2432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[24] VREF PIX_IN[2432] NB2 NB1 CSA_VREF pixel
xPix2433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[24] VREF PIX_IN[2433] NB2 NB1 CSA_VREF pixel
xPix2434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[24] VREF PIX_IN[2434] NB2 NB1 CSA_VREF pixel
xPix2435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[24] VREF PIX_IN[2435] NB2 NB1 CSA_VREF pixel
xPix2436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[24] VREF PIX_IN[2436] NB2 NB1 CSA_VREF pixel
xPix2437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[24] VREF PIX_IN[2437] NB2 NB1 CSA_VREF pixel
xPix2438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[24] VREF PIX_IN[2438] NB2 NB1 CSA_VREF pixel
xPix2439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[24] VREF PIX_IN[2439] NB2 NB1 CSA_VREF pixel
xPix2440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[24] VREF PIX_IN[2440] NB2 NB1 CSA_VREF pixel
xPix2441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[24] VREF PIX_IN[2441] NB2 NB1 CSA_VREF pixel
xPix2442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[24] VREF PIX_IN[2442] NB2 NB1 CSA_VREF pixel
xPix2443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[24] VREF PIX_IN[2443] NB2 NB1 CSA_VREF pixel
xPix2444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[24] VREF PIX_IN[2444] NB2 NB1 CSA_VREF pixel
xPix2445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[24] VREF PIX_IN[2445] NB2 NB1 CSA_VREF pixel
xPix2446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[24] VREF PIX_IN[2446] NB2 NB1 CSA_VREF pixel
xPix2447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[24] VREF PIX_IN[2447] NB2 NB1 CSA_VREF pixel
xPix2448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[24] VREF PIX_IN[2448] NB2 NB1 CSA_VREF pixel
xPix2449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[24] VREF PIX_IN[2449] NB2 NB1 CSA_VREF pixel
xPix2450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[24] VREF PIX_IN[2450] NB2 NB1 CSA_VREF pixel
xPix2451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[24] VREF PIX_IN[2451] NB2 NB1 CSA_VREF pixel
xPix2452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[24] VREF PIX_IN[2452] NB2 NB1 CSA_VREF pixel
xPix2453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[24] VREF PIX_IN[2453] NB2 NB1 CSA_VREF pixel
xPix2454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[24] VREF PIX_IN[2454] NB2 NB1 CSA_VREF pixel
xPix2455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[24] VREF PIX_IN[2455] NB2 NB1 CSA_VREF pixel
xPix2456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[24] VREF PIX_IN[2456] NB2 NB1 CSA_VREF pixel
xPix2457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[24] VREF PIX_IN[2457] NB2 NB1 CSA_VREF pixel
xPix2458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[24] VREF PIX_IN[2458] NB2 NB1 CSA_VREF pixel
xPix2459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[24] VREF PIX_IN[2459] NB2 NB1 CSA_VREF pixel
xPix2460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[24] VREF PIX_IN[2460] NB2 NB1 CSA_VREF pixel
xPix2461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[24] VREF PIX_IN[2461] NB2 NB1 CSA_VREF pixel
xPix2462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[24] VREF PIX_IN[2462] NB2 NB1 CSA_VREF pixel
xPix2463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[24] VREF PIX_IN[2463] NB2 NB1 CSA_VREF pixel
xPix2464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[24] VREF PIX_IN[2464] NB2 NB1 CSA_VREF pixel
xPix2465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[24] VREF PIX_IN[2465] NB2 NB1 CSA_VREF pixel
xPix2466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[24] VREF PIX_IN[2466] NB2 NB1 CSA_VREF pixel
xPix2467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[24] VREF PIX_IN[2467] NB2 NB1 CSA_VREF pixel
xPix2468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[24] VREF PIX_IN[2468] NB2 NB1 CSA_VREF pixel
xPix2469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[24] VREF PIX_IN[2469] NB2 NB1 CSA_VREF pixel
xPix2470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[24] VREF PIX_IN[2470] NB2 NB1 CSA_VREF pixel
xPix2471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[24] VREF PIX_IN[2471] NB2 NB1 CSA_VREF pixel
xPix2472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[24] VREF PIX_IN[2472] NB2 NB1 CSA_VREF pixel
xPix2473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[24] VREF PIX_IN[2473] NB2 NB1 CSA_VREF pixel
xPix2474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[24] VREF PIX_IN[2474] NB2 NB1 CSA_VREF pixel
xPix2475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[24] VREF PIX_IN[2475] NB2 NB1 CSA_VREF pixel
xPix2476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[24] VREF PIX_IN[2476] NB2 NB1 CSA_VREF pixel
xPix2477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[24] VREF PIX_IN[2477] NB2 NB1 CSA_VREF pixel
xPix2478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[24] VREF PIX_IN[2478] NB2 NB1 CSA_VREF pixel
xPix2479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[24] VREF PIX_IN[2479] NB2 NB1 CSA_VREF pixel
xPix2480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[24] VREF PIX_IN[2480] NB2 NB1 CSA_VREF pixel
xPix2481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[24] VREF PIX_IN[2481] NB2 NB1 CSA_VREF pixel
xPix2482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[24] VREF PIX_IN[2482] NB2 NB1 CSA_VREF pixel
xPix2483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[24] VREF PIX_IN[2483] NB2 NB1 CSA_VREF pixel
xPix2484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[24] VREF PIX_IN[2484] NB2 NB1 CSA_VREF pixel
xPix2485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[24] VREF PIX_IN[2485] NB2 NB1 CSA_VREF pixel
xPix2486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[24] VREF PIX_IN[2486] NB2 NB1 CSA_VREF pixel
xPix2487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[24] VREF PIX_IN[2487] NB2 NB1 CSA_VREF pixel
xPix2488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[24] VREF PIX_IN[2488] NB2 NB1 CSA_VREF pixel
xPix2489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[24] VREF PIX_IN[2489] NB2 NB1 CSA_VREF pixel
xPix2490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[24] VREF PIX_IN[2490] NB2 NB1 CSA_VREF pixel
xPix2491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[24] VREF PIX_IN[2491] NB2 NB1 CSA_VREF pixel
xPix2492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[24] VREF PIX_IN[2492] NB2 NB1 CSA_VREF pixel
xPix2493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[24] VREF PIX_IN[2493] NB2 NB1 CSA_VREF pixel
xPix2494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[24] VREF PIX_IN[2494] NB2 NB1 CSA_VREF pixel
xPix2495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[24] VREF PIX_IN[2495] NB2 NB1 CSA_VREF pixel
xPix2496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[24] VREF PIX_IN[2496] NB2 NB1 CSA_VREF pixel
xPix2497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[24] VREF PIX_IN[2497] NB2 NB1 CSA_VREF pixel
xPix2498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[24] VREF PIX_IN[2498] NB2 NB1 CSA_VREF pixel
xPix2499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[24] VREF PIX_IN[2499] NB2 NB1 CSA_VREF pixel
xPix2500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[25] VREF PIX_IN[2500] NB2 NB1 CSA_VREF pixel
xPix2501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[25] VREF PIX_IN[2501] NB2 NB1 CSA_VREF pixel
xPix2502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[25] VREF PIX_IN[2502] NB2 NB1 CSA_VREF pixel
xPix2503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[25] VREF PIX_IN[2503] NB2 NB1 CSA_VREF pixel
xPix2504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[25] VREF PIX_IN[2504] NB2 NB1 CSA_VREF pixel
xPix2505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[25] VREF PIX_IN[2505] NB2 NB1 CSA_VREF pixel
xPix2506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[25] VREF PIX_IN[2506] NB2 NB1 CSA_VREF pixel
xPix2507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[25] VREF PIX_IN[2507] NB2 NB1 CSA_VREF pixel
xPix2508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[25] VREF PIX_IN[2508] NB2 NB1 CSA_VREF pixel
xPix2509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[25] VREF PIX_IN[2509] NB2 NB1 CSA_VREF pixel
xPix2510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[25] VREF PIX_IN[2510] NB2 NB1 CSA_VREF pixel
xPix2511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[25] VREF PIX_IN[2511] NB2 NB1 CSA_VREF pixel
xPix2512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[25] VREF PIX_IN[2512] NB2 NB1 CSA_VREF pixel
xPix2513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[25] VREF PIX_IN[2513] NB2 NB1 CSA_VREF pixel
xPix2514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[25] VREF PIX_IN[2514] NB2 NB1 CSA_VREF pixel
xPix2515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[25] VREF PIX_IN[2515] NB2 NB1 CSA_VREF pixel
xPix2516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[25] VREF PIX_IN[2516] NB2 NB1 CSA_VREF pixel
xPix2517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[25] VREF PIX_IN[2517] NB2 NB1 CSA_VREF pixel
xPix2518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[25] VREF PIX_IN[2518] NB2 NB1 CSA_VREF pixel
xPix2519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[25] VREF PIX_IN[2519] NB2 NB1 CSA_VREF pixel
xPix2520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[25] VREF PIX_IN[2520] NB2 NB1 CSA_VREF pixel
xPix2521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[25] VREF PIX_IN[2521] NB2 NB1 CSA_VREF pixel
xPix2522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[25] VREF PIX_IN[2522] NB2 NB1 CSA_VREF pixel
xPix2523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[25] VREF PIX_IN[2523] NB2 NB1 CSA_VREF pixel
xPix2524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[25] VREF PIX_IN[2524] NB2 NB1 CSA_VREF pixel
xPix2525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[25] VREF PIX_IN[2525] NB2 NB1 CSA_VREF pixel
xPix2526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[25] VREF PIX_IN[2526] NB2 NB1 CSA_VREF pixel
xPix2527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[25] VREF PIX_IN[2527] NB2 NB1 CSA_VREF pixel
xPix2528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[25] VREF PIX_IN[2528] NB2 NB1 CSA_VREF pixel
xPix2529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[25] VREF PIX_IN[2529] NB2 NB1 CSA_VREF pixel
xPix2530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[25] VREF PIX_IN[2530] NB2 NB1 CSA_VREF pixel
xPix2531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[25] VREF PIX_IN[2531] NB2 NB1 CSA_VREF pixel
xPix2532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[25] VREF PIX_IN[2532] NB2 NB1 CSA_VREF pixel
xPix2533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[25] VREF PIX_IN[2533] NB2 NB1 CSA_VREF pixel
xPix2534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[25] VREF PIX_IN[2534] NB2 NB1 CSA_VREF pixel
xPix2535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[25] VREF PIX_IN[2535] NB2 NB1 CSA_VREF pixel
xPix2536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[25] VREF PIX_IN[2536] NB2 NB1 CSA_VREF pixel
xPix2537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[25] VREF PIX_IN[2537] NB2 NB1 CSA_VREF pixel
xPix2538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[25] VREF PIX_IN[2538] NB2 NB1 CSA_VREF pixel
xPix2539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[25] VREF PIX_IN[2539] NB2 NB1 CSA_VREF pixel
xPix2540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[25] VREF PIX_IN[2540] NB2 NB1 CSA_VREF pixel
xPix2541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[25] VREF PIX_IN[2541] NB2 NB1 CSA_VREF pixel
xPix2542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[25] VREF PIX_IN[2542] NB2 NB1 CSA_VREF pixel
xPix2543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[25] VREF PIX_IN[2543] NB2 NB1 CSA_VREF pixel
xPix2544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[25] VREF PIX_IN[2544] NB2 NB1 CSA_VREF pixel
xPix2545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[25] VREF PIX_IN[2545] NB2 NB1 CSA_VREF pixel
xPix2546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[25] VREF PIX_IN[2546] NB2 NB1 CSA_VREF pixel
xPix2547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[25] VREF PIX_IN[2547] NB2 NB1 CSA_VREF pixel
xPix2548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[25] VREF PIX_IN[2548] NB2 NB1 CSA_VREF pixel
xPix2549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[25] VREF PIX_IN[2549] NB2 NB1 CSA_VREF pixel
xPix2550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[25] VREF PIX_IN[2550] NB2 NB1 CSA_VREF pixel
xPix2551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[25] VREF PIX_IN[2551] NB2 NB1 CSA_VREF pixel
xPix2552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[25] VREF PIX_IN[2552] NB2 NB1 CSA_VREF pixel
xPix2553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[25] VREF PIX_IN[2553] NB2 NB1 CSA_VREF pixel
xPix2554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[25] VREF PIX_IN[2554] NB2 NB1 CSA_VREF pixel
xPix2555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[25] VREF PIX_IN[2555] NB2 NB1 CSA_VREF pixel
xPix2556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[25] VREF PIX_IN[2556] NB2 NB1 CSA_VREF pixel
xPix2557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[25] VREF PIX_IN[2557] NB2 NB1 CSA_VREF pixel
xPix2558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[25] VREF PIX_IN[2558] NB2 NB1 CSA_VREF pixel
xPix2559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[25] VREF PIX_IN[2559] NB2 NB1 CSA_VREF pixel
xPix2560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[25] VREF PIX_IN[2560] NB2 NB1 CSA_VREF pixel
xPix2561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[25] VREF PIX_IN[2561] NB2 NB1 CSA_VREF pixel
xPix2562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[25] VREF PIX_IN[2562] NB2 NB1 CSA_VREF pixel
xPix2563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[25] VREF PIX_IN[2563] NB2 NB1 CSA_VREF pixel
xPix2564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[25] VREF PIX_IN[2564] NB2 NB1 CSA_VREF pixel
xPix2565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[25] VREF PIX_IN[2565] NB2 NB1 CSA_VREF pixel
xPix2566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[25] VREF PIX_IN[2566] NB2 NB1 CSA_VREF pixel
xPix2567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[25] VREF PIX_IN[2567] NB2 NB1 CSA_VREF pixel
xPix2568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[25] VREF PIX_IN[2568] NB2 NB1 CSA_VREF pixel
xPix2569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[25] VREF PIX_IN[2569] NB2 NB1 CSA_VREF pixel
xPix2570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[25] VREF PIX_IN[2570] NB2 NB1 CSA_VREF pixel
xPix2571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[25] VREF PIX_IN[2571] NB2 NB1 CSA_VREF pixel
xPix2572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[25] VREF PIX_IN[2572] NB2 NB1 CSA_VREF pixel
xPix2573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[25] VREF PIX_IN[2573] NB2 NB1 CSA_VREF pixel
xPix2574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[25] VREF PIX_IN[2574] NB2 NB1 CSA_VREF pixel
xPix2575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[25] VREF PIX_IN[2575] NB2 NB1 CSA_VREF pixel
xPix2576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[25] VREF PIX_IN[2576] NB2 NB1 CSA_VREF pixel
xPix2577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[25] VREF PIX_IN[2577] NB2 NB1 CSA_VREF pixel
xPix2578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[25] VREF PIX_IN[2578] NB2 NB1 CSA_VREF pixel
xPix2579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[25] VREF PIX_IN[2579] NB2 NB1 CSA_VREF pixel
xPix2580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[25] VREF PIX_IN[2580] NB2 NB1 CSA_VREF pixel
xPix2581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[25] VREF PIX_IN[2581] NB2 NB1 CSA_VREF pixel
xPix2582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[25] VREF PIX_IN[2582] NB2 NB1 CSA_VREF pixel
xPix2583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[25] VREF PIX_IN[2583] NB2 NB1 CSA_VREF pixel
xPix2584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[25] VREF PIX_IN[2584] NB2 NB1 CSA_VREF pixel
xPix2585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[25] VREF PIX_IN[2585] NB2 NB1 CSA_VREF pixel
xPix2586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[25] VREF PIX_IN[2586] NB2 NB1 CSA_VREF pixel
xPix2587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[25] VREF PIX_IN[2587] NB2 NB1 CSA_VREF pixel
xPix2588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[25] VREF PIX_IN[2588] NB2 NB1 CSA_VREF pixel
xPix2589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[25] VREF PIX_IN[2589] NB2 NB1 CSA_VREF pixel
xPix2590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[25] VREF PIX_IN[2590] NB2 NB1 CSA_VREF pixel
xPix2591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[25] VREF PIX_IN[2591] NB2 NB1 CSA_VREF pixel
xPix2592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[25] VREF PIX_IN[2592] NB2 NB1 CSA_VREF pixel
xPix2593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[25] VREF PIX_IN[2593] NB2 NB1 CSA_VREF pixel
xPix2594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[25] VREF PIX_IN[2594] NB2 NB1 CSA_VREF pixel
xPix2595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[25] VREF PIX_IN[2595] NB2 NB1 CSA_VREF pixel
xPix2596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[25] VREF PIX_IN[2596] NB2 NB1 CSA_VREF pixel
xPix2597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[25] VREF PIX_IN[2597] NB2 NB1 CSA_VREF pixel
xPix2598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[25] VREF PIX_IN[2598] NB2 NB1 CSA_VREF pixel
xPix2599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[25] VREF PIX_IN[2599] NB2 NB1 CSA_VREF pixel
xPix2600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[26] VREF PIX_IN[2600] NB2 NB1 CSA_VREF pixel
xPix2601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[26] VREF PIX_IN[2601] NB2 NB1 CSA_VREF pixel
xPix2602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[26] VREF PIX_IN[2602] NB2 NB1 CSA_VREF pixel
xPix2603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[26] VREF PIX_IN[2603] NB2 NB1 CSA_VREF pixel
xPix2604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[26] VREF PIX_IN[2604] NB2 NB1 CSA_VREF pixel
xPix2605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[26] VREF PIX_IN[2605] NB2 NB1 CSA_VREF pixel
xPix2606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[26] VREF PIX_IN[2606] NB2 NB1 CSA_VREF pixel
xPix2607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[26] VREF PIX_IN[2607] NB2 NB1 CSA_VREF pixel
xPix2608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[26] VREF PIX_IN[2608] NB2 NB1 CSA_VREF pixel
xPix2609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[26] VREF PIX_IN[2609] NB2 NB1 CSA_VREF pixel
xPix2610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[26] VREF PIX_IN[2610] NB2 NB1 CSA_VREF pixel
xPix2611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[26] VREF PIX_IN[2611] NB2 NB1 CSA_VREF pixel
xPix2612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[26] VREF PIX_IN[2612] NB2 NB1 CSA_VREF pixel
xPix2613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[26] VREF PIX_IN[2613] NB2 NB1 CSA_VREF pixel
xPix2614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[26] VREF PIX_IN[2614] NB2 NB1 CSA_VREF pixel
xPix2615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[26] VREF PIX_IN[2615] NB2 NB1 CSA_VREF pixel
xPix2616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[26] VREF PIX_IN[2616] NB2 NB1 CSA_VREF pixel
xPix2617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[26] VREF PIX_IN[2617] NB2 NB1 CSA_VREF pixel
xPix2618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[26] VREF PIX_IN[2618] NB2 NB1 CSA_VREF pixel
xPix2619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[26] VREF PIX_IN[2619] NB2 NB1 CSA_VREF pixel
xPix2620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[26] VREF PIX_IN[2620] NB2 NB1 CSA_VREF pixel
xPix2621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[26] VREF PIX_IN[2621] NB2 NB1 CSA_VREF pixel
xPix2622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[26] VREF PIX_IN[2622] NB2 NB1 CSA_VREF pixel
xPix2623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[26] VREF PIX_IN[2623] NB2 NB1 CSA_VREF pixel
xPix2624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[26] VREF PIX_IN[2624] NB2 NB1 CSA_VREF pixel
xPix2625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[26] VREF PIX_IN[2625] NB2 NB1 CSA_VREF pixel
xPix2626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[26] VREF PIX_IN[2626] NB2 NB1 CSA_VREF pixel
xPix2627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[26] VREF PIX_IN[2627] NB2 NB1 CSA_VREF pixel
xPix2628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[26] VREF PIX_IN[2628] NB2 NB1 CSA_VREF pixel
xPix2629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[26] VREF PIX_IN[2629] NB2 NB1 CSA_VREF pixel
xPix2630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[26] VREF PIX_IN[2630] NB2 NB1 CSA_VREF pixel
xPix2631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[26] VREF PIX_IN[2631] NB2 NB1 CSA_VREF pixel
xPix2632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[26] VREF PIX_IN[2632] NB2 NB1 CSA_VREF pixel
xPix2633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[26] VREF PIX_IN[2633] NB2 NB1 CSA_VREF pixel
xPix2634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[26] VREF PIX_IN[2634] NB2 NB1 CSA_VREF pixel
xPix2635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[26] VREF PIX_IN[2635] NB2 NB1 CSA_VREF pixel
xPix2636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[26] VREF PIX_IN[2636] NB2 NB1 CSA_VREF pixel
xPix2637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[26] VREF PIX_IN[2637] NB2 NB1 CSA_VREF pixel
xPix2638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[26] VREF PIX_IN[2638] NB2 NB1 CSA_VREF pixel
xPix2639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[26] VREF PIX_IN[2639] NB2 NB1 CSA_VREF pixel
xPix2640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[26] VREF PIX_IN[2640] NB2 NB1 CSA_VREF pixel
xPix2641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[26] VREF PIX_IN[2641] NB2 NB1 CSA_VREF pixel
xPix2642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[26] VREF PIX_IN[2642] NB2 NB1 CSA_VREF pixel
xPix2643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[26] VREF PIX_IN[2643] NB2 NB1 CSA_VREF pixel
xPix2644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[26] VREF PIX_IN[2644] NB2 NB1 CSA_VREF pixel
xPix2645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[26] VREF PIX_IN[2645] NB2 NB1 CSA_VREF pixel
xPix2646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[26] VREF PIX_IN[2646] NB2 NB1 CSA_VREF pixel
xPix2647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[26] VREF PIX_IN[2647] NB2 NB1 CSA_VREF pixel
xPix2648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[26] VREF PIX_IN[2648] NB2 NB1 CSA_VREF pixel
xPix2649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[26] VREF PIX_IN[2649] NB2 NB1 CSA_VREF pixel
xPix2650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[26] VREF PIX_IN[2650] NB2 NB1 CSA_VREF pixel
xPix2651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[26] VREF PIX_IN[2651] NB2 NB1 CSA_VREF pixel
xPix2652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[26] VREF PIX_IN[2652] NB2 NB1 CSA_VREF pixel
xPix2653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[26] VREF PIX_IN[2653] NB2 NB1 CSA_VREF pixel
xPix2654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[26] VREF PIX_IN[2654] NB2 NB1 CSA_VREF pixel
xPix2655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[26] VREF PIX_IN[2655] NB2 NB1 CSA_VREF pixel
xPix2656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[26] VREF PIX_IN[2656] NB2 NB1 CSA_VREF pixel
xPix2657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[26] VREF PIX_IN[2657] NB2 NB1 CSA_VREF pixel
xPix2658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[26] VREF PIX_IN[2658] NB2 NB1 CSA_VREF pixel
xPix2659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[26] VREF PIX_IN[2659] NB2 NB1 CSA_VREF pixel
xPix2660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[26] VREF PIX_IN[2660] NB2 NB1 CSA_VREF pixel
xPix2661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[26] VREF PIX_IN[2661] NB2 NB1 CSA_VREF pixel
xPix2662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[26] VREF PIX_IN[2662] NB2 NB1 CSA_VREF pixel
xPix2663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[26] VREF PIX_IN[2663] NB2 NB1 CSA_VREF pixel
xPix2664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[26] VREF PIX_IN[2664] NB2 NB1 CSA_VREF pixel
xPix2665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[26] VREF PIX_IN[2665] NB2 NB1 CSA_VREF pixel
xPix2666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[26] VREF PIX_IN[2666] NB2 NB1 CSA_VREF pixel
xPix2667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[26] VREF PIX_IN[2667] NB2 NB1 CSA_VREF pixel
xPix2668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[26] VREF PIX_IN[2668] NB2 NB1 CSA_VREF pixel
xPix2669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[26] VREF PIX_IN[2669] NB2 NB1 CSA_VREF pixel
xPix2670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[26] VREF PIX_IN[2670] NB2 NB1 CSA_VREF pixel
xPix2671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[26] VREF PIX_IN[2671] NB2 NB1 CSA_VREF pixel
xPix2672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[26] VREF PIX_IN[2672] NB2 NB1 CSA_VREF pixel
xPix2673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[26] VREF PIX_IN[2673] NB2 NB1 CSA_VREF pixel
xPix2674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[26] VREF PIX_IN[2674] NB2 NB1 CSA_VREF pixel
xPix2675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[26] VREF PIX_IN[2675] NB2 NB1 CSA_VREF pixel
xPix2676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[26] VREF PIX_IN[2676] NB2 NB1 CSA_VREF pixel
xPix2677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[26] VREF PIX_IN[2677] NB2 NB1 CSA_VREF pixel
xPix2678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[26] VREF PIX_IN[2678] NB2 NB1 CSA_VREF pixel
xPix2679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[26] VREF PIX_IN[2679] NB2 NB1 CSA_VREF pixel
xPix2680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[26] VREF PIX_IN[2680] NB2 NB1 CSA_VREF pixel
xPix2681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[26] VREF PIX_IN[2681] NB2 NB1 CSA_VREF pixel
xPix2682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[26] VREF PIX_IN[2682] NB2 NB1 CSA_VREF pixel
xPix2683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[26] VREF PIX_IN[2683] NB2 NB1 CSA_VREF pixel
xPix2684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[26] VREF PIX_IN[2684] NB2 NB1 CSA_VREF pixel
xPix2685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[26] VREF PIX_IN[2685] NB2 NB1 CSA_VREF pixel
xPix2686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[26] VREF PIX_IN[2686] NB2 NB1 CSA_VREF pixel
xPix2687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[26] VREF PIX_IN[2687] NB2 NB1 CSA_VREF pixel
xPix2688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[26] VREF PIX_IN[2688] NB2 NB1 CSA_VREF pixel
xPix2689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[26] VREF PIX_IN[2689] NB2 NB1 CSA_VREF pixel
xPix2690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[26] VREF PIX_IN[2690] NB2 NB1 CSA_VREF pixel
xPix2691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[26] VREF PIX_IN[2691] NB2 NB1 CSA_VREF pixel
xPix2692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[26] VREF PIX_IN[2692] NB2 NB1 CSA_VREF pixel
xPix2693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[26] VREF PIX_IN[2693] NB2 NB1 CSA_VREF pixel
xPix2694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[26] VREF PIX_IN[2694] NB2 NB1 CSA_VREF pixel
xPix2695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[26] VREF PIX_IN[2695] NB2 NB1 CSA_VREF pixel
xPix2696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[26] VREF PIX_IN[2696] NB2 NB1 CSA_VREF pixel
xPix2697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[26] VREF PIX_IN[2697] NB2 NB1 CSA_VREF pixel
xPix2698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[26] VREF PIX_IN[2698] NB2 NB1 CSA_VREF pixel
xPix2699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[26] VREF PIX_IN[2699] NB2 NB1 CSA_VREF pixel
xPix2700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[27] VREF PIX_IN[2700] NB2 NB1 CSA_VREF pixel
xPix2701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[27] VREF PIX_IN[2701] NB2 NB1 CSA_VREF pixel
xPix2702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[27] VREF PIX_IN[2702] NB2 NB1 CSA_VREF pixel
xPix2703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[27] VREF PIX_IN[2703] NB2 NB1 CSA_VREF pixel
xPix2704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[27] VREF PIX_IN[2704] NB2 NB1 CSA_VREF pixel
xPix2705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[27] VREF PIX_IN[2705] NB2 NB1 CSA_VREF pixel
xPix2706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[27] VREF PIX_IN[2706] NB2 NB1 CSA_VREF pixel
xPix2707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[27] VREF PIX_IN[2707] NB2 NB1 CSA_VREF pixel
xPix2708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[27] VREF PIX_IN[2708] NB2 NB1 CSA_VREF pixel
xPix2709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[27] VREF PIX_IN[2709] NB2 NB1 CSA_VREF pixel
xPix2710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[27] VREF PIX_IN[2710] NB2 NB1 CSA_VREF pixel
xPix2711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[27] VREF PIX_IN[2711] NB2 NB1 CSA_VREF pixel
xPix2712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[27] VREF PIX_IN[2712] NB2 NB1 CSA_VREF pixel
xPix2713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[27] VREF PIX_IN[2713] NB2 NB1 CSA_VREF pixel
xPix2714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[27] VREF PIX_IN[2714] NB2 NB1 CSA_VREF pixel
xPix2715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[27] VREF PIX_IN[2715] NB2 NB1 CSA_VREF pixel
xPix2716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[27] VREF PIX_IN[2716] NB2 NB1 CSA_VREF pixel
xPix2717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[27] VREF PIX_IN[2717] NB2 NB1 CSA_VREF pixel
xPix2718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[27] VREF PIX_IN[2718] NB2 NB1 CSA_VREF pixel
xPix2719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[27] VREF PIX_IN[2719] NB2 NB1 CSA_VREF pixel
xPix2720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[27] VREF PIX_IN[2720] NB2 NB1 CSA_VREF pixel
xPix2721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[27] VREF PIX_IN[2721] NB2 NB1 CSA_VREF pixel
xPix2722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[27] VREF PIX_IN[2722] NB2 NB1 CSA_VREF pixel
xPix2723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[27] VREF PIX_IN[2723] NB2 NB1 CSA_VREF pixel
xPix2724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[27] VREF PIX_IN[2724] NB2 NB1 CSA_VREF pixel
xPix2725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[27] VREF PIX_IN[2725] NB2 NB1 CSA_VREF pixel
xPix2726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[27] VREF PIX_IN[2726] NB2 NB1 CSA_VREF pixel
xPix2727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[27] VREF PIX_IN[2727] NB2 NB1 CSA_VREF pixel
xPix2728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[27] VREF PIX_IN[2728] NB2 NB1 CSA_VREF pixel
xPix2729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[27] VREF PIX_IN[2729] NB2 NB1 CSA_VREF pixel
xPix2730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[27] VREF PIX_IN[2730] NB2 NB1 CSA_VREF pixel
xPix2731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[27] VREF PIX_IN[2731] NB2 NB1 CSA_VREF pixel
xPix2732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[27] VREF PIX_IN[2732] NB2 NB1 CSA_VREF pixel
xPix2733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[27] VREF PIX_IN[2733] NB2 NB1 CSA_VREF pixel
xPix2734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[27] VREF PIX_IN[2734] NB2 NB1 CSA_VREF pixel
xPix2735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[27] VREF PIX_IN[2735] NB2 NB1 CSA_VREF pixel
xPix2736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[27] VREF PIX_IN[2736] NB2 NB1 CSA_VREF pixel
xPix2737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[27] VREF PIX_IN[2737] NB2 NB1 CSA_VREF pixel
xPix2738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[27] VREF PIX_IN[2738] NB2 NB1 CSA_VREF pixel
xPix2739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[27] VREF PIX_IN[2739] NB2 NB1 CSA_VREF pixel
xPix2740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[27] VREF PIX_IN[2740] NB2 NB1 CSA_VREF pixel
xPix2741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[27] VREF PIX_IN[2741] NB2 NB1 CSA_VREF pixel
xPix2742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[27] VREF PIX_IN[2742] NB2 NB1 CSA_VREF pixel
xPix2743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[27] VREF PIX_IN[2743] NB2 NB1 CSA_VREF pixel
xPix2744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[27] VREF PIX_IN[2744] NB2 NB1 CSA_VREF pixel
xPix2745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[27] VREF PIX_IN[2745] NB2 NB1 CSA_VREF pixel
xPix2746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[27] VREF PIX_IN[2746] NB2 NB1 CSA_VREF pixel
xPix2747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[27] VREF PIX_IN[2747] NB2 NB1 CSA_VREF pixel
xPix2748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[27] VREF PIX_IN[2748] NB2 NB1 CSA_VREF pixel
xPix2749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[27] VREF PIX_IN[2749] NB2 NB1 CSA_VREF pixel
xPix2750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[27] VREF PIX_IN[2750] NB2 NB1 CSA_VREF pixel
xPix2751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[27] VREF PIX_IN[2751] NB2 NB1 CSA_VREF pixel
xPix2752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[27] VREF PIX_IN[2752] NB2 NB1 CSA_VREF pixel
xPix2753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[27] VREF PIX_IN[2753] NB2 NB1 CSA_VREF pixel
xPix2754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[27] VREF PIX_IN[2754] NB2 NB1 CSA_VREF pixel
xPix2755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[27] VREF PIX_IN[2755] NB2 NB1 CSA_VREF pixel
xPix2756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[27] VREF PIX_IN[2756] NB2 NB1 CSA_VREF pixel
xPix2757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[27] VREF PIX_IN[2757] NB2 NB1 CSA_VREF pixel
xPix2758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[27] VREF PIX_IN[2758] NB2 NB1 CSA_VREF pixel
xPix2759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[27] VREF PIX_IN[2759] NB2 NB1 CSA_VREF pixel
xPix2760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[27] VREF PIX_IN[2760] NB2 NB1 CSA_VREF pixel
xPix2761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[27] VREF PIX_IN[2761] NB2 NB1 CSA_VREF pixel
xPix2762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[27] VREF PIX_IN[2762] NB2 NB1 CSA_VREF pixel
xPix2763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[27] VREF PIX_IN[2763] NB2 NB1 CSA_VREF pixel
xPix2764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[27] VREF PIX_IN[2764] NB2 NB1 CSA_VREF pixel
xPix2765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[27] VREF PIX_IN[2765] NB2 NB1 CSA_VREF pixel
xPix2766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[27] VREF PIX_IN[2766] NB2 NB1 CSA_VREF pixel
xPix2767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[27] VREF PIX_IN[2767] NB2 NB1 CSA_VREF pixel
xPix2768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[27] VREF PIX_IN[2768] NB2 NB1 CSA_VREF pixel
xPix2769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[27] VREF PIX_IN[2769] NB2 NB1 CSA_VREF pixel
xPix2770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[27] VREF PIX_IN[2770] NB2 NB1 CSA_VREF pixel
xPix2771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[27] VREF PIX_IN[2771] NB2 NB1 CSA_VREF pixel
xPix2772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[27] VREF PIX_IN[2772] NB2 NB1 CSA_VREF pixel
xPix2773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[27] VREF PIX_IN[2773] NB2 NB1 CSA_VREF pixel
xPix2774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[27] VREF PIX_IN[2774] NB2 NB1 CSA_VREF pixel
xPix2775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[27] VREF PIX_IN[2775] NB2 NB1 CSA_VREF pixel
xPix2776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[27] VREF PIX_IN[2776] NB2 NB1 CSA_VREF pixel
xPix2777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[27] VREF PIX_IN[2777] NB2 NB1 CSA_VREF pixel
xPix2778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[27] VREF PIX_IN[2778] NB2 NB1 CSA_VREF pixel
xPix2779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[27] VREF PIX_IN[2779] NB2 NB1 CSA_VREF pixel
xPix2780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[27] VREF PIX_IN[2780] NB2 NB1 CSA_VREF pixel
xPix2781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[27] VREF PIX_IN[2781] NB2 NB1 CSA_VREF pixel
xPix2782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[27] VREF PIX_IN[2782] NB2 NB1 CSA_VREF pixel
xPix2783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[27] VREF PIX_IN[2783] NB2 NB1 CSA_VREF pixel
xPix2784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[27] VREF PIX_IN[2784] NB2 NB1 CSA_VREF pixel
xPix2785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[27] VREF PIX_IN[2785] NB2 NB1 CSA_VREF pixel
xPix2786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[27] VREF PIX_IN[2786] NB2 NB1 CSA_VREF pixel
xPix2787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[27] VREF PIX_IN[2787] NB2 NB1 CSA_VREF pixel
xPix2788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[27] VREF PIX_IN[2788] NB2 NB1 CSA_VREF pixel
xPix2789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[27] VREF PIX_IN[2789] NB2 NB1 CSA_VREF pixel
xPix2790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[27] VREF PIX_IN[2790] NB2 NB1 CSA_VREF pixel
xPix2791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[27] VREF PIX_IN[2791] NB2 NB1 CSA_VREF pixel
xPix2792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[27] VREF PIX_IN[2792] NB2 NB1 CSA_VREF pixel
xPix2793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[27] VREF PIX_IN[2793] NB2 NB1 CSA_VREF pixel
xPix2794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[27] VREF PIX_IN[2794] NB2 NB1 CSA_VREF pixel
xPix2795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[27] VREF PIX_IN[2795] NB2 NB1 CSA_VREF pixel
xPix2796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[27] VREF PIX_IN[2796] NB2 NB1 CSA_VREF pixel
xPix2797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[27] VREF PIX_IN[2797] NB2 NB1 CSA_VREF pixel
xPix2798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[27] VREF PIX_IN[2798] NB2 NB1 CSA_VREF pixel
xPix2799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[27] VREF PIX_IN[2799] NB2 NB1 CSA_VREF pixel
xPix2800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[28] VREF PIX_IN[2800] NB2 NB1 CSA_VREF pixel
xPix2801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[28] VREF PIX_IN[2801] NB2 NB1 CSA_VREF pixel
xPix2802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[28] VREF PIX_IN[2802] NB2 NB1 CSA_VREF pixel
xPix2803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[28] VREF PIX_IN[2803] NB2 NB1 CSA_VREF pixel
xPix2804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[28] VREF PIX_IN[2804] NB2 NB1 CSA_VREF pixel
xPix2805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[28] VREF PIX_IN[2805] NB2 NB1 CSA_VREF pixel
xPix2806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[28] VREF PIX_IN[2806] NB2 NB1 CSA_VREF pixel
xPix2807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[28] VREF PIX_IN[2807] NB2 NB1 CSA_VREF pixel
xPix2808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[28] VREF PIX_IN[2808] NB2 NB1 CSA_VREF pixel
xPix2809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[28] VREF PIX_IN[2809] NB2 NB1 CSA_VREF pixel
xPix2810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[28] VREF PIX_IN[2810] NB2 NB1 CSA_VREF pixel
xPix2811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[28] VREF PIX_IN[2811] NB2 NB1 CSA_VREF pixel
xPix2812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[28] VREF PIX_IN[2812] NB2 NB1 CSA_VREF pixel
xPix2813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[28] VREF PIX_IN[2813] NB2 NB1 CSA_VREF pixel
xPix2814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[28] VREF PIX_IN[2814] NB2 NB1 CSA_VREF pixel
xPix2815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[28] VREF PIX_IN[2815] NB2 NB1 CSA_VREF pixel
xPix2816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[28] VREF PIX_IN[2816] NB2 NB1 CSA_VREF pixel
xPix2817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[28] VREF PIX_IN[2817] NB2 NB1 CSA_VREF pixel
xPix2818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[28] VREF PIX_IN[2818] NB2 NB1 CSA_VREF pixel
xPix2819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[28] VREF PIX_IN[2819] NB2 NB1 CSA_VREF pixel
xPix2820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[28] VREF PIX_IN[2820] NB2 NB1 CSA_VREF pixel
xPix2821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[28] VREF PIX_IN[2821] NB2 NB1 CSA_VREF pixel
xPix2822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[28] VREF PIX_IN[2822] NB2 NB1 CSA_VREF pixel
xPix2823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[28] VREF PIX_IN[2823] NB2 NB1 CSA_VREF pixel
xPix2824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[28] VREF PIX_IN[2824] NB2 NB1 CSA_VREF pixel
xPix2825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[28] VREF PIX_IN[2825] NB2 NB1 CSA_VREF pixel
xPix2826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[28] VREF PIX_IN[2826] NB2 NB1 CSA_VREF pixel
xPix2827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[28] VREF PIX_IN[2827] NB2 NB1 CSA_VREF pixel
xPix2828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[28] VREF PIX_IN[2828] NB2 NB1 CSA_VREF pixel
xPix2829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[28] VREF PIX_IN[2829] NB2 NB1 CSA_VREF pixel
xPix2830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[28] VREF PIX_IN[2830] NB2 NB1 CSA_VREF pixel
xPix2831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[28] VREF PIX_IN[2831] NB2 NB1 CSA_VREF pixel
xPix2832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[28] VREF PIX_IN[2832] NB2 NB1 CSA_VREF pixel
xPix2833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[28] VREF PIX_IN[2833] NB2 NB1 CSA_VREF pixel
xPix2834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[28] VREF PIX_IN[2834] NB2 NB1 CSA_VREF pixel
xPix2835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[28] VREF PIX_IN[2835] NB2 NB1 CSA_VREF pixel
xPix2836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[28] VREF PIX_IN[2836] NB2 NB1 CSA_VREF pixel
xPix2837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[28] VREF PIX_IN[2837] NB2 NB1 CSA_VREF pixel
xPix2838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[28] VREF PIX_IN[2838] NB2 NB1 CSA_VREF pixel
xPix2839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[28] VREF PIX_IN[2839] NB2 NB1 CSA_VREF pixel
xPix2840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[28] VREF PIX_IN[2840] NB2 NB1 CSA_VREF pixel
xPix2841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[28] VREF PIX_IN[2841] NB2 NB1 CSA_VREF pixel
xPix2842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[28] VREF PIX_IN[2842] NB2 NB1 CSA_VREF pixel
xPix2843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[28] VREF PIX_IN[2843] NB2 NB1 CSA_VREF pixel
xPix2844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[28] VREF PIX_IN[2844] NB2 NB1 CSA_VREF pixel
xPix2845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[28] VREF PIX_IN[2845] NB2 NB1 CSA_VREF pixel
xPix2846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[28] VREF PIX_IN[2846] NB2 NB1 CSA_VREF pixel
xPix2847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[28] VREF PIX_IN[2847] NB2 NB1 CSA_VREF pixel
xPix2848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[28] VREF PIX_IN[2848] NB2 NB1 CSA_VREF pixel
xPix2849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[28] VREF PIX_IN[2849] NB2 NB1 CSA_VREF pixel
xPix2850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[28] VREF PIX_IN[2850] NB2 NB1 CSA_VREF pixel
xPix2851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[28] VREF PIX_IN[2851] NB2 NB1 CSA_VREF pixel
xPix2852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[28] VREF PIX_IN[2852] NB2 NB1 CSA_VREF pixel
xPix2853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[28] VREF PIX_IN[2853] NB2 NB1 CSA_VREF pixel
xPix2854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[28] VREF PIX_IN[2854] NB2 NB1 CSA_VREF pixel
xPix2855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[28] VREF PIX_IN[2855] NB2 NB1 CSA_VREF pixel
xPix2856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[28] VREF PIX_IN[2856] NB2 NB1 CSA_VREF pixel
xPix2857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[28] VREF PIX_IN[2857] NB2 NB1 CSA_VREF pixel
xPix2858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[28] VREF PIX_IN[2858] NB2 NB1 CSA_VREF pixel
xPix2859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[28] VREF PIX_IN[2859] NB2 NB1 CSA_VREF pixel
xPix2860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[28] VREF PIX_IN[2860] NB2 NB1 CSA_VREF pixel
xPix2861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[28] VREF PIX_IN[2861] NB2 NB1 CSA_VREF pixel
xPix2862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[28] VREF PIX_IN[2862] NB2 NB1 CSA_VREF pixel
xPix2863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[28] VREF PIX_IN[2863] NB2 NB1 CSA_VREF pixel
xPix2864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[28] VREF PIX_IN[2864] NB2 NB1 CSA_VREF pixel
xPix2865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[28] VREF PIX_IN[2865] NB2 NB1 CSA_VREF pixel
xPix2866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[28] VREF PIX_IN[2866] NB2 NB1 CSA_VREF pixel
xPix2867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[28] VREF PIX_IN[2867] NB2 NB1 CSA_VREF pixel
xPix2868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[28] VREF PIX_IN[2868] NB2 NB1 CSA_VREF pixel
xPix2869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[28] VREF PIX_IN[2869] NB2 NB1 CSA_VREF pixel
xPix2870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[28] VREF PIX_IN[2870] NB2 NB1 CSA_VREF pixel
xPix2871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[28] VREF PIX_IN[2871] NB2 NB1 CSA_VREF pixel
xPix2872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[28] VREF PIX_IN[2872] NB2 NB1 CSA_VREF pixel
xPix2873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[28] VREF PIX_IN[2873] NB2 NB1 CSA_VREF pixel
xPix2874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[28] VREF PIX_IN[2874] NB2 NB1 CSA_VREF pixel
xPix2875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[28] VREF PIX_IN[2875] NB2 NB1 CSA_VREF pixel
xPix2876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[28] VREF PIX_IN[2876] NB2 NB1 CSA_VREF pixel
xPix2877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[28] VREF PIX_IN[2877] NB2 NB1 CSA_VREF pixel
xPix2878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[28] VREF PIX_IN[2878] NB2 NB1 CSA_VREF pixel
xPix2879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[28] VREF PIX_IN[2879] NB2 NB1 CSA_VREF pixel
xPix2880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[28] VREF PIX_IN[2880] NB2 NB1 CSA_VREF pixel
xPix2881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[28] VREF PIX_IN[2881] NB2 NB1 CSA_VREF pixel
xPix2882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[28] VREF PIX_IN[2882] NB2 NB1 CSA_VREF pixel
xPix2883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[28] VREF PIX_IN[2883] NB2 NB1 CSA_VREF pixel
xPix2884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[28] VREF PIX_IN[2884] NB2 NB1 CSA_VREF pixel
xPix2885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[28] VREF PIX_IN[2885] NB2 NB1 CSA_VREF pixel
xPix2886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[28] VREF PIX_IN[2886] NB2 NB1 CSA_VREF pixel
xPix2887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[28] VREF PIX_IN[2887] NB2 NB1 CSA_VREF pixel
xPix2888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[28] VREF PIX_IN[2888] NB2 NB1 CSA_VREF pixel
xPix2889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[28] VREF PIX_IN[2889] NB2 NB1 CSA_VREF pixel
xPix2890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[28] VREF PIX_IN[2890] NB2 NB1 CSA_VREF pixel
xPix2891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[28] VREF PIX_IN[2891] NB2 NB1 CSA_VREF pixel
xPix2892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[28] VREF PIX_IN[2892] NB2 NB1 CSA_VREF pixel
xPix2893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[28] VREF PIX_IN[2893] NB2 NB1 CSA_VREF pixel
xPix2894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[28] VREF PIX_IN[2894] NB2 NB1 CSA_VREF pixel
xPix2895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[28] VREF PIX_IN[2895] NB2 NB1 CSA_VREF pixel
xPix2896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[28] VREF PIX_IN[2896] NB2 NB1 CSA_VREF pixel
xPix2897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[28] VREF PIX_IN[2897] NB2 NB1 CSA_VREF pixel
xPix2898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[28] VREF PIX_IN[2898] NB2 NB1 CSA_VREF pixel
xPix2899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[28] VREF PIX_IN[2899] NB2 NB1 CSA_VREF pixel
xPix2900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[29] VREF PIX_IN[2900] NB2 NB1 CSA_VREF pixel
xPix2901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[29] VREF PIX_IN[2901] NB2 NB1 CSA_VREF pixel
xPix2902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[29] VREF PIX_IN[2902] NB2 NB1 CSA_VREF pixel
xPix2903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[29] VREF PIX_IN[2903] NB2 NB1 CSA_VREF pixel
xPix2904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[29] VREF PIX_IN[2904] NB2 NB1 CSA_VREF pixel
xPix2905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[29] VREF PIX_IN[2905] NB2 NB1 CSA_VREF pixel
xPix2906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[29] VREF PIX_IN[2906] NB2 NB1 CSA_VREF pixel
xPix2907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[29] VREF PIX_IN[2907] NB2 NB1 CSA_VREF pixel
xPix2908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[29] VREF PIX_IN[2908] NB2 NB1 CSA_VREF pixel
xPix2909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[29] VREF PIX_IN[2909] NB2 NB1 CSA_VREF pixel
xPix2910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[29] VREF PIX_IN[2910] NB2 NB1 CSA_VREF pixel
xPix2911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[29] VREF PIX_IN[2911] NB2 NB1 CSA_VREF pixel
xPix2912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[29] VREF PIX_IN[2912] NB2 NB1 CSA_VREF pixel
xPix2913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[29] VREF PIX_IN[2913] NB2 NB1 CSA_VREF pixel
xPix2914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[29] VREF PIX_IN[2914] NB2 NB1 CSA_VREF pixel
xPix2915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[29] VREF PIX_IN[2915] NB2 NB1 CSA_VREF pixel
xPix2916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[29] VREF PIX_IN[2916] NB2 NB1 CSA_VREF pixel
xPix2917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[29] VREF PIX_IN[2917] NB2 NB1 CSA_VREF pixel
xPix2918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[29] VREF PIX_IN[2918] NB2 NB1 CSA_VREF pixel
xPix2919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[29] VREF PIX_IN[2919] NB2 NB1 CSA_VREF pixel
xPix2920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[29] VREF PIX_IN[2920] NB2 NB1 CSA_VREF pixel
xPix2921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[29] VREF PIX_IN[2921] NB2 NB1 CSA_VREF pixel
xPix2922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[29] VREF PIX_IN[2922] NB2 NB1 CSA_VREF pixel
xPix2923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[29] VREF PIX_IN[2923] NB2 NB1 CSA_VREF pixel
xPix2924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[29] VREF PIX_IN[2924] NB2 NB1 CSA_VREF pixel
xPix2925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[29] VREF PIX_IN[2925] NB2 NB1 CSA_VREF pixel
xPix2926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[29] VREF PIX_IN[2926] NB2 NB1 CSA_VREF pixel
xPix2927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[29] VREF PIX_IN[2927] NB2 NB1 CSA_VREF pixel
xPix2928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[29] VREF PIX_IN[2928] NB2 NB1 CSA_VREF pixel
xPix2929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[29] VREF PIX_IN[2929] NB2 NB1 CSA_VREF pixel
xPix2930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[29] VREF PIX_IN[2930] NB2 NB1 CSA_VREF pixel
xPix2931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[29] VREF PIX_IN[2931] NB2 NB1 CSA_VREF pixel
xPix2932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[29] VREF PIX_IN[2932] NB2 NB1 CSA_VREF pixel
xPix2933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[29] VREF PIX_IN[2933] NB2 NB1 CSA_VREF pixel
xPix2934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[29] VREF PIX_IN[2934] NB2 NB1 CSA_VREF pixel
xPix2935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[29] VREF PIX_IN[2935] NB2 NB1 CSA_VREF pixel
xPix2936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[29] VREF PIX_IN[2936] NB2 NB1 CSA_VREF pixel
xPix2937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[29] VREF PIX_IN[2937] NB2 NB1 CSA_VREF pixel
xPix2938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[29] VREF PIX_IN[2938] NB2 NB1 CSA_VREF pixel
xPix2939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[29] VREF PIX_IN[2939] NB2 NB1 CSA_VREF pixel
xPix2940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[29] VREF PIX_IN[2940] NB2 NB1 CSA_VREF pixel
xPix2941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[29] VREF PIX_IN[2941] NB2 NB1 CSA_VREF pixel
xPix2942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[29] VREF PIX_IN[2942] NB2 NB1 CSA_VREF pixel
xPix2943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[29] VREF PIX_IN[2943] NB2 NB1 CSA_VREF pixel
xPix2944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[29] VREF PIX_IN[2944] NB2 NB1 CSA_VREF pixel
xPix2945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[29] VREF PIX_IN[2945] NB2 NB1 CSA_VREF pixel
xPix2946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[29] VREF PIX_IN[2946] NB2 NB1 CSA_VREF pixel
xPix2947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[29] VREF PIX_IN[2947] NB2 NB1 CSA_VREF pixel
xPix2948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[29] VREF PIX_IN[2948] NB2 NB1 CSA_VREF pixel
xPix2949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[29] VREF PIX_IN[2949] NB2 NB1 CSA_VREF pixel
xPix2950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[29] VREF PIX_IN[2950] NB2 NB1 CSA_VREF pixel
xPix2951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[29] VREF PIX_IN[2951] NB2 NB1 CSA_VREF pixel
xPix2952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[29] VREF PIX_IN[2952] NB2 NB1 CSA_VREF pixel
xPix2953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[29] VREF PIX_IN[2953] NB2 NB1 CSA_VREF pixel
xPix2954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[29] VREF PIX_IN[2954] NB2 NB1 CSA_VREF pixel
xPix2955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[29] VREF PIX_IN[2955] NB2 NB1 CSA_VREF pixel
xPix2956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[29] VREF PIX_IN[2956] NB2 NB1 CSA_VREF pixel
xPix2957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[29] VREF PIX_IN[2957] NB2 NB1 CSA_VREF pixel
xPix2958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[29] VREF PIX_IN[2958] NB2 NB1 CSA_VREF pixel
xPix2959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[29] VREF PIX_IN[2959] NB2 NB1 CSA_VREF pixel
xPix2960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[29] VREF PIX_IN[2960] NB2 NB1 CSA_VREF pixel
xPix2961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[29] VREF PIX_IN[2961] NB2 NB1 CSA_VREF pixel
xPix2962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[29] VREF PIX_IN[2962] NB2 NB1 CSA_VREF pixel
xPix2963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[29] VREF PIX_IN[2963] NB2 NB1 CSA_VREF pixel
xPix2964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[29] VREF PIX_IN[2964] NB2 NB1 CSA_VREF pixel
xPix2965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[29] VREF PIX_IN[2965] NB2 NB1 CSA_VREF pixel
xPix2966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[29] VREF PIX_IN[2966] NB2 NB1 CSA_VREF pixel
xPix2967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[29] VREF PIX_IN[2967] NB2 NB1 CSA_VREF pixel
xPix2968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[29] VREF PIX_IN[2968] NB2 NB1 CSA_VREF pixel
xPix2969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[29] VREF PIX_IN[2969] NB2 NB1 CSA_VREF pixel
xPix2970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[29] VREF PIX_IN[2970] NB2 NB1 CSA_VREF pixel
xPix2971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[29] VREF PIX_IN[2971] NB2 NB1 CSA_VREF pixel
xPix2972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[29] VREF PIX_IN[2972] NB2 NB1 CSA_VREF pixel
xPix2973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[29] VREF PIX_IN[2973] NB2 NB1 CSA_VREF pixel
xPix2974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[29] VREF PIX_IN[2974] NB2 NB1 CSA_VREF pixel
xPix2975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[29] VREF PIX_IN[2975] NB2 NB1 CSA_VREF pixel
xPix2976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[29] VREF PIX_IN[2976] NB2 NB1 CSA_VREF pixel
xPix2977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[29] VREF PIX_IN[2977] NB2 NB1 CSA_VREF pixel
xPix2978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[29] VREF PIX_IN[2978] NB2 NB1 CSA_VREF pixel
xPix2979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[29] VREF PIX_IN[2979] NB2 NB1 CSA_VREF pixel
xPix2980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[29] VREF PIX_IN[2980] NB2 NB1 CSA_VREF pixel
xPix2981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[29] VREF PIX_IN[2981] NB2 NB1 CSA_VREF pixel
xPix2982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[29] VREF PIX_IN[2982] NB2 NB1 CSA_VREF pixel
xPix2983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[29] VREF PIX_IN[2983] NB2 NB1 CSA_VREF pixel
xPix2984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[29] VREF PIX_IN[2984] NB2 NB1 CSA_VREF pixel
xPix2985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[29] VREF PIX_IN[2985] NB2 NB1 CSA_VREF pixel
xPix2986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[29] VREF PIX_IN[2986] NB2 NB1 CSA_VREF pixel
xPix2987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[29] VREF PIX_IN[2987] NB2 NB1 CSA_VREF pixel
xPix2988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[29] VREF PIX_IN[2988] NB2 NB1 CSA_VREF pixel
xPix2989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[29] VREF PIX_IN[2989] NB2 NB1 CSA_VREF pixel
xPix2990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[29] VREF PIX_IN[2990] NB2 NB1 CSA_VREF pixel
xPix2991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[29] VREF PIX_IN[2991] NB2 NB1 CSA_VREF pixel
xPix2992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[29] VREF PIX_IN[2992] NB2 NB1 CSA_VREF pixel
xPix2993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[29] VREF PIX_IN[2993] NB2 NB1 CSA_VREF pixel
xPix2994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[29] VREF PIX_IN[2994] NB2 NB1 CSA_VREF pixel
xPix2995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[29] VREF PIX_IN[2995] NB2 NB1 CSA_VREF pixel
xPix2996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[29] VREF PIX_IN[2996] NB2 NB1 CSA_VREF pixel
xPix2997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[29] VREF PIX_IN[2997] NB2 NB1 CSA_VREF pixel
xPix2998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[29] VREF PIX_IN[2998] NB2 NB1 CSA_VREF pixel
xPix2999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[29] VREF PIX_IN[2999] NB2 NB1 CSA_VREF pixel
xPix3000 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[30] VREF PIX_IN[3000] NB2 NB1 CSA_VREF pixel
xPix3001 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[30] VREF PIX_IN[3001] NB2 NB1 CSA_VREF pixel
xPix3002 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[30] VREF PIX_IN[3002] NB2 NB1 CSA_VREF pixel
xPix3003 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[30] VREF PIX_IN[3003] NB2 NB1 CSA_VREF pixel
xPix3004 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[30] VREF PIX_IN[3004] NB2 NB1 CSA_VREF pixel
xPix3005 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[30] VREF PIX_IN[3005] NB2 NB1 CSA_VREF pixel
xPix3006 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[30] VREF PIX_IN[3006] NB2 NB1 CSA_VREF pixel
xPix3007 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[30] VREF PIX_IN[3007] NB2 NB1 CSA_VREF pixel
xPix3008 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[30] VREF PIX_IN[3008] NB2 NB1 CSA_VREF pixel
xPix3009 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[30] VREF PIX_IN[3009] NB2 NB1 CSA_VREF pixel
xPix3010 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[30] VREF PIX_IN[3010] NB2 NB1 CSA_VREF pixel
xPix3011 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[30] VREF PIX_IN[3011] NB2 NB1 CSA_VREF pixel
xPix3012 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[30] VREF PIX_IN[3012] NB2 NB1 CSA_VREF pixel
xPix3013 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[30] VREF PIX_IN[3013] NB2 NB1 CSA_VREF pixel
xPix3014 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[30] VREF PIX_IN[3014] NB2 NB1 CSA_VREF pixel
xPix3015 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[30] VREF PIX_IN[3015] NB2 NB1 CSA_VREF pixel
xPix3016 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[30] VREF PIX_IN[3016] NB2 NB1 CSA_VREF pixel
xPix3017 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[30] VREF PIX_IN[3017] NB2 NB1 CSA_VREF pixel
xPix3018 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[30] VREF PIX_IN[3018] NB2 NB1 CSA_VREF pixel
xPix3019 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[30] VREF PIX_IN[3019] NB2 NB1 CSA_VREF pixel
xPix3020 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[30] VREF PIX_IN[3020] NB2 NB1 CSA_VREF pixel
xPix3021 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[30] VREF PIX_IN[3021] NB2 NB1 CSA_VREF pixel
xPix3022 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[30] VREF PIX_IN[3022] NB2 NB1 CSA_VREF pixel
xPix3023 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[30] VREF PIX_IN[3023] NB2 NB1 CSA_VREF pixel
xPix3024 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[30] VREF PIX_IN[3024] NB2 NB1 CSA_VREF pixel
xPix3025 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[30] VREF PIX_IN[3025] NB2 NB1 CSA_VREF pixel
xPix3026 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[30] VREF PIX_IN[3026] NB2 NB1 CSA_VREF pixel
xPix3027 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[30] VREF PIX_IN[3027] NB2 NB1 CSA_VREF pixel
xPix3028 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[30] VREF PIX_IN[3028] NB2 NB1 CSA_VREF pixel
xPix3029 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[30] VREF PIX_IN[3029] NB2 NB1 CSA_VREF pixel
xPix3030 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[30] VREF PIX_IN[3030] NB2 NB1 CSA_VREF pixel
xPix3031 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[30] VREF PIX_IN[3031] NB2 NB1 CSA_VREF pixel
xPix3032 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[30] VREF PIX_IN[3032] NB2 NB1 CSA_VREF pixel
xPix3033 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[30] VREF PIX_IN[3033] NB2 NB1 CSA_VREF pixel
xPix3034 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[30] VREF PIX_IN[3034] NB2 NB1 CSA_VREF pixel
xPix3035 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[30] VREF PIX_IN[3035] NB2 NB1 CSA_VREF pixel
xPix3036 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[30] VREF PIX_IN[3036] NB2 NB1 CSA_VREF pixel
xPix3037 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[30] VREF PIX_IN[3037] NB2 NB1 CSA_VREF pixel
xPix3038 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[30] VREF PIX_IN[3038] NB2 NB1 CSA_VREF pixel
xPix3039 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[30] VREF PIX_IN[3039] NB2 NB1 CSA_VREF pixel
xPix3040 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[30] VREF PIX_IN[3040] NB2 NB1 CSA_VREF pixel
xPix3041 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[30] VREF PIX_IN[3041] NB2 NB1 CSA_VREF pixel
xPix3042 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[30] VREF PIX_IN[3042] NB2 NB1 CSA_VREF pixel
xPix3043 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[30] VREF PIX_IN[3043] NB2 NB1 CSA_VREF pixel
xPix3044 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[30] VREF PIX_IN[3044] NB2 NB1 CSA_VREF pixel
xPix3045 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[30] VREF PIX_IN[3045] NB2 NB1 CSA_VREF pixel
xPix3046 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[30] VREF PIX_IN[3046] NB2 NB1 CSA_VREF pixel
xPix3047 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[30] VREF PIX_IN[3047] NB2 NB1 CSA_VREF pixel
xPix3048 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[30] VREF PIX_IN[3048] NB2 NB1 CSA_VREF pixel
xPix3049 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[30] VREF PIX_IN[3049] NB2 NB1 CSA_VREF pixel
xPix3050 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[30] VREF PIX_IN[3050] NB2 NB1 CSA_VREF pixel
xPix3051 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[30] VREF PIX_IN[3051] NB2 NB1 CSA_VREF pixel
xPix3052 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[30] VREF PIX_IN[3052] NB2 NB1 CSA_VREF pixel
xPix3053 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[30] VREF PIX_IN[3053] NB2 NB1 CSA_VREF pixel
xPix3054 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[30] VREF PIX_IN[3054] NB2 NB1 CSA_VREF pixel
xPix3055 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[30] VREF PIX_IN[3055] NB2 NB1 CSA_VREF pixel
xPix3056 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[30] VREF PIX_IN[3056] NB2 NB1 CSA_VREF pixel
xPix3057 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[30] VREF PIX_IN[3057] NB2 NB1 CSA_VREF pixel
xPix3058 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[30] VREF PIX_IN[3058] NB2 NB1 CSA_VREF pixel
xPix3059 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[30] VREF PIX_IN[3059] NB2 NB1 CSA_VREF pixel
xPix3060 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[30] VREF PIX_IN[3060] NB2 NB1 CSA_VREF pixel
xPix3061 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[30] VREF PIX_IN[3061] NB2 NB1 CSA_VREF pixel
xPix3062 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[30] VREF PIX_IN[3062] NB2 NB1 CSA_VREF pixel
xPix3063 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[30] VREF PIX_IN[3063] NB2 NB1 CSA_VREF pixel
xPix3064 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[30] VREF PIX_IN[3064] NB2 NB1 CSA_VREF pixel
xPix3065 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[30] VREF PIX_IN[3065] NB2 NB1 CSA_VREF pixel
xPix3066 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[30] VREF PIX_IN[3066] NB2 NB1 CSA_VREF pixel
xPix3067 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[30] VREF PIX_IN[3067] NB2 NB1 CSA_VREF pixel
xPix3068 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[30] VREF PIX_IN[3068] NB2 NB1 CSA_VREF pixel
xPix3069 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[30] VREF PIX_IN[3069] NB2 NB1 CSA_VREF pixel
xPix3070 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[30] VREF PIX_IN[3070] NB2 NB1 CSA_VREF pixel
xPix3071 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[30] VREF PIX_IN[3071] NB2 NB1 CSA_VREF pixel
xPix3072 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[30] VREF PIX_IN[3072] NB2 NB1 CSA_VREF pixel
xPix3073 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[30] VREF PIX_IN[3073] NB2 NB1 CSA_VREF pixel
xPix3074 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[30] VREF PIX_IN[3074] NB2 NB1 CSA_VREF pixel
xPix3075 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[30] VREF PIX_IN[3075] NB2 NB1 CSA_VREF pixel
xPix3076 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[30] VREF PIX_IN[3076] NB2 NB1 CSA_VREF pixel
xPix3077 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[30] VREF PIX_IN[3077] NB2 NB1 CSA_VREF pixel
xPix3078 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[30] VREF PIX_IN[3078] NB2 NB1 CSA_VREF pixel
xPix3079 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[30] VREF PIX_IN[3079] NB2 NB1 CSA_VREF pixel
xPix3080 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[30] VREF PIX_IN[3080] NB2 NB1 CSA_VREF pixel
xPix3081 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[30] VREF PIX_IN[3081] NB2 NB1 CSA_VREF pixel
xPix3082 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[30] VREF PIX_IN[3082] NB2 NB1 CSA_VREF pixel
xPix3083 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[30] VREF PIX_IN[3083] NB2 NB1 CSA_VREF pixel
xPix3084 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[30] VREF PIX_IN[3084] NB2 NB1 CSA_VREF pixel
xPix3085 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[30] VREF PIX_IN[3085] NB2 NB1 CSA_VREF pixel
xPix3086 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[30] VREF PIX_IN[3086] NB2 NB1 CSA_VREF pixel
xPix3087 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[30] VREF PIX_IN[3087] NB2 NB1 CSA_VREF pixel
xPix3088 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[30] VREF PIX_IN[3088] NB2 NB1 CSA_VREF pixel
xPix3089 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[30] VREF PIX_IN[3089] NB2 NB1 CSA_VREF pixel
xPix3090 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[30] VREF PIX_IN[3090] NB2 NB1 CSA_VREF pixel
xPix3091 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[30] VREF PIX_IN[3091] NB2 NB1 CSA_VREF pixel
xPix3092 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[30] VREF PIX_IN[3092] NB2 NB1 CSA_VREF pixel
xPix3093 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[30] VREF PIX_IN[3093] NB2 NB1 CSA_VREF pixel
xPix3094 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[30] VREF PIX_IN[3094] NB2 NB1 CSA_VREF pixel
xPix3095 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[30] VREF PIX_IN[3095] NB2 NB1 CSA_VREF pixel
xPix3096 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[30] VREF PIX_IN[3096] NB2 NB1 CSA_VREF pixel
xPix3097 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[30] VREF PIX_IN[3097] NB2 NB1 CSA_VREF pixel
xPix3098 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[30] VREF PIX_IN[3098] NB2 NB1 CSA_VREF pixel
xPix3099 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[30] VREF PIX_IN[3099] NB2 NB1 CSA_VREF pixel
xPix3100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[31] VREF PIX_IN[3100] NB2 NB1 CSA_VREF pixel
xPix3101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[31] VREF PIX_IN[3101] NB2 NB1 CSA_VREF pixel
xPix3102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[31] VREF PIX_IN[3102] NB2 NB1 CSA_VREF pixel
xPix3103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[31] VREF PIX_IN[3103] NB2 NB1 CSA_VREF pixel
xPix3104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[31] VREF PIX_IN[3104] NB2 NB1 CSA_VREF pixel
xPix3105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[31] VREF PIX_IN[3105] NB2 NB1 CSA_VREF pixel
xPix3106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[31] VREF PIX_IN[3106] NB2 NB1 CSA_VREF pixel
xPix3107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[31] VREF PIX_IN[3107] NB2 NB1 CSA_VREF pixel
xPix3108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[31] VREF PIX_IN[3108] NB2 NB1 CSA_VREF pixel
xPix3109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[31] VREF PIX_IN[3109] NB2 NB1 CSA_VREF pixel
xPix3110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[31] VREF PIX_IN[3110] NB2 NB1 CSA_VREF pixel
xPix3111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[31] VREF PIX_IN[3111] NB2 NB1 CSA_VREF pixel
xPix3112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[31] VREF PIX_IN[3112] NB2 NB1 CSA_VREF pixel
xPix3113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[31] VREF PIX_IN[3113] NB2 NB1 CSA_VREF pixel
xPix3114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[31] VREF PIX_IN[3114] NB2 NB1 CSA_VREF pixel
xPix3115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[31] VREF PIX_IN[3115] NB2 NB1 CSA_VREF pixel
xPix3116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[31] VREF PIX_IN[3116] NB2 NB1 CSA_VREF pixel
xPix3117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[31] VREF PIX_IN[3117] NB2 NB1 CSA_VREF pixel
xPix3118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[31] VREF PIX_IN[3118] NB2 NB1 CSA_VREF pixel
xPix3119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[31] VREF PIX_IN[3119] NB2 NB1 CSA_VREF pixel
xPix3120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[31] VREF PIX_IN[3120] NB2 NB1 CSA_VREF pixel
xPix3121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[31] VREF PIX_IN[3121] NB2 NB1 CSA_VREF pixel
xPix3122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[31] VREF PIX_IN[3122] NB2 NB1 CSA_VREF pixel
xPix3123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[31] VREF PIX_IN[3123] NB2 NB1 CSA_VREF pixel
xPix3124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[31] VREF PIX_IN[3124] NB2 NB1 CSA_VREF pixel
xPix3125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[31] VREF PIX_IN[3125] NB2 NB1 CSA_VREF pixel
xPix3126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[31] VREF PIX_IN[3126] NB2 NB1 CSA_VREF pixel
xPix3127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[31] VREF PIX_IN[3127] NB2 NB1 CSA_VREF pixel
xPix3128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[31] VREF PIX_IN[3128] NB2 NB1 CSA_VREF pixel
xPix3129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[31] VREF PIX_IN[3129] NB2 NB1 CSA_VREF pixel
xPix3130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[31] VREF PIX_IN[3130] NB2 NB1 CSA_VREF pixel
xPix3131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[31] VREF PIX_IN[3131] NB2 NB1 CSA_VREF pixel
xPix3132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[31] VREF PIX_IN[3132] NB2 NB1 CSA_VREF pixel
xPix3133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[31] VREF PIX_IN[3133] NB2 NB1 CSA_VREF pixel
xPix3134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[31] VREF PIX_IN[3134] NB2 NB1 CSA_VREF pixel
xPix3135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[31] VREF PIX_IN[3135] NB2 NB1 CSA_VREF pixel
xPix3136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[31] VREF PIX_IN[3136] NB2 NB1 CSA_VREF pixel
xPix3137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[31] VREF PIX_IN[3137] NB2 NB1 CSA_VREF pixel
xPix3138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[31] VREF PIX_IN[3138] NB2 NB1 CSA_VREF pixel
xPix3139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[31] VREF PIX_IN[3139] NB2 NB1 CSA_VREF pixel
xPix3140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[31] VREF PIX_IN[3140] NB2 NB1 CSA_VREF pixel
xPix3141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[31] VREF PIX_IN[3141] NB2 NB1 CSA_VREF pixel
xPix3142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[31] VREF PIX_IN[3142] NB2 NB1 CSA_VREF pixel
xPix3143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[31] VREF PIX_IN[3143] NB2 NB1 CSA_VREF pixel
xPix3144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[31] VREF PIX_IN[3144] NB2 NB1 CSA_VREF pixel
xPix3145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[31] VREF PIX_IN[3145] NB2 NB1 CSA_VREF pixel
xPix3146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[31] VREF PIX_IN[3146] NB2 NB1 CSA_VREF pixel
xPix3147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[31] VREF PIX_IN[3147] NB2 NB1 CSA_VREF pixel
xPix3148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[31] VREF PIX_IN[3148] NB2 NB1 CSA_VREF pixel
xPix3149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[31] VREF PIX_IN[3149] NB2 NB1 CSA_VREF pixel
xPix3150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[31] VREF PIX_IN[3150] NB2 NB1 CSA_VREF pixel
xPix3151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[31] VREF PIX_IN[3151] NB2 NB1 CSA_VREF pixel
xPix3152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[31] VREF PIX_IN[3152] NB2 NB1 CSA_VREF pixel
xPix3153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[31] VREF PIX_IN[3153] NB2 NB1 CSA_VREF pixel
xPix3154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[31] VREF PIX_IN[3154] NB2 NB1 CSA_VREF pixel
xPix3155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[31] VREF PIX_IN[3155] NB2 NB1 CSA_VREF pixel
xPix3156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[31] VREF PIX_IN[3156] NB2 NB1 CSA_VREF pixel
xPix3157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[31] VREF PIX_IN[3157] NB2 NB1 CSA_VREF pixel
xPix3158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[31] VREF PIX_IN[3158] NB2 NB1 CSA_VREF pixel
xPix3159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[31] VREF PIX_IN[3159] NB2 NB1 CSA_VREF pixel
xPix3160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[31] VREF PIX_IN[3160] NB2 NB1 CSA_VREF pixel
xPix3161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[31] VREF PIX_IN[3161] NB2 NB1 CSA_VREF pixel
xPix3162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[31] VREF PIX_IN[3162] NB2 NB1 CSA_VREF pixel
xPix3163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[31] VREF PIX_IN[3163] NB2 NB1 CSA_VREF pixel
xPix3164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[31] VREF PIX_IN[3164] NB2 NB1 CSA_VREF pixel
xPix3165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[31] VREF PIX_IN[3165] NB2 NB1 CSA_VREF pixel
xPix3166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[31] VREF PIX_IN[3166] NB2 NB1 CSA_VREF pixel
xPix3167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[31] VREF PIX_IN[3167] NB2 NB1 CSA_VREF pixel
xPix3168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[31] VREF PIX_IN[3168] NB2 NB1 CSA_VREF pixel
xPix3169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[31] VREF PIX_IN[3169] NB2 NB1 CSA_VREF pixel
xPix3170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[31] VREF PIX_IN[3170] NB2 NB1 CSA_VREF pixel
xPix3171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[31] VREF PIX_IN[3171] NB2 NB1 CSA_VREF pixel
xPix3172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[31] VREF PIX_IN[3172] NB2 NB1 CSA_VREF pixel
xPix3173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[31] VREF PIX_IN[3173] NB2 NB1 CSA_VREF pixel
xPix3174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[31] VREF PIX_IN[3174] NB2 NB1 CSA_VREF pixel
xPix3175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[31] VREF PIX_IN[3175] NB2 NB1 CSA_VREF pixel
xPix3176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[31] VREF PIX_IN[3176] NB2 NB1 CSA_VREF pixel
xPix3177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[31] VREF PIX_IN[3177] NB2 NB1 CSA_VREF pixel
xPix3178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[31] VREF PIX_IN[3178] NB2 NB1 CSA_VREF pixel
xPix3179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[31] VREF PIX_IN[3179] NB2 NB1 CSA_VREF pixel
xPix3180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[31] VREF PIX_IN[3180] NB2 NB1 CSA_VREF pixel
xPix3181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[31] VREF PIX_IN[3181] NB2 NB1 CSA_VREF pixel
xPix3182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[31] VREF PIX_IN[3182] NB2 NB1 CSA_VREF pixel
xPix3183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[31] VREF PIX_IN[3183] NB2 NB1 CSA_VREF pixel
xPix3184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[31] VREF PIX_IN[3184] NB2 NB1 CSA_VREF pixel
xPix3185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[31] VREF PIX_IN[3185] NB2 NB1 CSA_VREF pixel
xPix3186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[31] VREF PIX_IN[3186] NB2 NB1 CSA_VREF pixel
xPix3187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[31] VREF PIX_IN[3187] NB2 NB1 CSA_VREF pixel
xPix3188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[31] VREF PIX_IN[3188] NB2 NB1 CSA_VREF pixel
xPix3189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[31] VREF PIX_IN[3189] NB2 NB1 CSA_VREF pixel
xPix3190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[31] VREF PIX_IN[3190] NB2 NB1 CSA_VREF pixel
xPix3191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[31] VREF PIX_IN[3191] NB2 NB1 CSA_VREF pixel
xPix3192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[31] VREF PIX_IN[3192] NB2 NB1 CSA_VREF pixel
xPix3193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[31] VREF PIX_IN[3193] NB2 NB1 CSA_VREF pixel
xPix3194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[31] VREF PIX_IN[3194] NB2 NB1 CSA_VREF pixel
xPix3195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[31] VREF PIX_IN[3195] NB2 NB1 CSA_VREF pixel
xPix3196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[31] VREF PIX_IN[3196] NB2 NB1 CSA_VREF pixel
xPix3197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[31] VREF PIX_IN[3197] NB2 NB1 CSA_VREF pixel
xPix3198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[31] VREF PIX_IN[3198] NB2 NB1 CSA_VREF pixel
xPix3199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[31] VREF PIX_IN[3199] NB2 NB1 CSA_VREF pixel
xPix3200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[32] VREF PIX_IN[3200] NB2 NB1 CSA_VREF pixel
xPix3201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[32] VREF PIX_IN[3201] NB2 NB1 CSA_VREF pixel
xPix3202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[32] VREF PIX_IN[3202] NB2 NB1 CSA_VREF pixel
xPix3203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[32] VREF PIX_IN[3203] NB2 NB1 CSA_VREF pixel
xPix3204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[32] VREF PIX_IN[3204] NB2 NB1 CSA_VREF pixel
xPix3205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[32] VREF PIX_IN[3205] NB2 NB1 CSA_VREF pixel
xPix3206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[32] VREF PIX_IN[3206] NB2 NB1 CSA_VREF pixel
xPix3207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[32] VREF PIX_IN[3207] NB2 NB1 CSA_VREF pixel
xPix3208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[32] VREF PIX_IN[3208] NB2 NB1 CSA_VREF pixel
xPix3209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[32] VREF PIX_IN[3209] NB2 NB1 CSA_VREF pixel
xPix3210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[32] VREF PIX_IN[3210] NB2 NB1 CSA_VREF pixel
xPix3211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[32] VREF PIX_IN[3211] NB2 NB1 CSA_VREF pixel
xPix3212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[32] VREF PIX_IN[3212] NB2 NB1 CSA_VREF pixel
xPix3213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[32] VREF PIX_IN[3213] NB2 NB1 CSA_VREF pixel
xPix3214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[32] VREF PIX_IN[3214] NB2 NB1 CSA_VREF pixel
xPix3215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[32] VREF PIX_IN[3215] NB2 NB1 CSA_VREF pixel
xPix3216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[32] VREF PIX_IN[3216] NB2 NB1 CSA_VREF pixel
xPix3217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[32] VREF PIX_IN[3217] NB2 NB1 CSA_VREF pixel
xPix3218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[32] VREF PIX_IN[3218] NB2 NB1 CSA_VREF pixel
xPix3219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[32] VREF PIX_IN[3219] NB2 NB1 CSA_VREF pixel
xPix3220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[32] VREF PIX_IN[3220] NB2 NB1 CSA_VREF pixel
xPix3221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[32] VREF PIX_IN[3221] NB2 NB1 CSA_VREF pixel
xPix3222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[32] VREF PIX_IN[3222] NB2 NB1 CSA_VREF pixel
xPix3223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[32] VREF PIX_IN[3223] NB2 NB1 CSA_VREF pixel
xPix3224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[32] VREF PIX_IN[3224] NB2 NB1 CSA_VREF pixel
xPix3225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[32] VREF PIX_IN[3225] NB2 NB1 CSA_VREF pixel
xPix3226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[32] VREF PIX_IN[3226] NB2 NB1 CSA_VREF pixel
xPix3227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[32] VREF PIX_IN[3227] NB2 NB1 CSA_VREF pixel
xPix3228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[32] VREF PIX_IN[3228] NB2 NB1 CSA_VREF pixel
xPix3229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[32] VREF PIX_IN[3229] NB2 NB1 CSA_VREF pixel
xPix3230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[32] VREF PIX_IN[3230] NB2 NB1 CSA_VREF pixel
xPix3231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[32] VREF PIX_IN[3231] NB2 NB1 CSA_VREF pixel
xPix3232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[32] VREF PIX_IN[3232] NB2 NB1 CSA_VREF pixel
xPix3233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[32] VREF PIX_IN[3233] NB2 NB1 CSA_VREF pixel
xPix3234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[32] VREF PIX_IN[3234] NB2 NB1 CSA_VREF pixel
xPix3235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[32] VREF PIX_IN[3235] NB2 NB1 CSA_VREF pixel
xPix3236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[32] VREF PIX_IN[3236] NB2 NB1 CSA_VREF pixel
xPix3237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[32] VREF PIX_IN[3237] NB2 NB1 CSA_VREF pixel
xPix3238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[32] VREF PIX_IN[3238] NB2 NB1 CSA_VREF pixel
xPix3239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[32] VREF PIX_IN[3239] NB2 NB1 CSA_VREF pixel
xPix3240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[32] VREF PIX_IN[3240] NB2 NB1 CSA_VREF pixel
xPix3241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[32] VREF PIX_IN[3241] NB2 NB1 CSA_VREF pixel
xPix3242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[32] VREF PIX_IN[3242] NB2 NB1 CSA_VREF pixel
xPix3243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[32] VREF PIX_IN[3243] NB2 NB1 CSA_VREF pixel
xPix3244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[32] VREF PIX_IN[3244] NB2 NB1 CSA_VREF pixel
xPix3245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[32] VREF PIX_IN[3245] NB2 NB1 CSA_VREF pixel
xPix3246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[32] VREF PIX_IN[3246] NB2 NB1 CSA_VREF pixel
xPix3247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[32] VREF PIX_IN[3247] NB2 NB1 CSA_VREF pixel
xPix3248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[32] VREF PIX_IN[3248] NB2 NB1 CSA_VREF pixel
xPix3249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[32] VREF PIX_IN[3249] NB2 NB1 CSA_VREF pixel
xPix3250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[32] VREF PIX_IN[3250] NB2 NB1 CSA_VREF pixel
xPix3251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[32] VREF PIX_IN[3251] NB2 NB1 CSA_VREF pixel
xPix3252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[32] VREF PIX_IN[3252] NB2 NB1 CSA_VREF pixel
xPix3253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[32] VREF PIX_IN[3253] NB2 NB1 CSA_VREF pixel
xPix3254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[32] VREF PIX_IN[3254] NB2 NB1 CSA_VREF pixel
xPix3255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[32] VREF PIX_IN[3255] NB2 NB1 CSA_VREF pixel
xPix3256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[32] VREF PIX_IN[3256] NB2 NB1 CSA_VREF pixel
xPix3257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[32] VREF PIX_IN[3257] NB2 NB1 CSA_VREF pixel
xPix3258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[32] VREF PIX_IN[3258] NB2 NB1 CSA_VREF pixel
xPix3259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[32] VREF PIX_IN[3259] NB2 NB1 CSA_VREF pixel
xPix3260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[32] VREF PIX_IN[3260] NB2 NB1 CSA_VREF pixel
xPix3261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[32] VREF PIX_IN[3261] NB2 NB1 CSA_VREF pixel
xPix3262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[32] VREF PIX_IN[3262] NB2 NB1 CSA_VREF pixel
xPix3263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[32] VREF PIX_IN[3263] NB2 NB1 CSA_VREF pixel
xPix3264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[32] VREF PIX_IN[3264] NB2 NB1 CSA_VREF pixel
xPix3265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[32] VREF PIX_IN[3265] NB2 NB1 CSA_VREF pixel
xPix3266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[32] VREF PIX_IN[3266] NB2 NB1 CSA_VREF pixel
xPix3267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[32] VREF PIX_IN[3267] NB2 NB1 CSA_VREF pixel
xPix3268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[32] VREF PIX_IN[3268] NB2 NB1 CSA_VREF pixel
xPix3269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[32] VREF PIX_IN[3269] NB2 NB1 CSA_VREF pixel
xPix3270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[32] VREF PIX_IN[3270] NB2 NB1 CSA_VREF pixel
xPix3271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[32] VREF PIX_IN[3271] NB2 NB1 CSA_VREF pixel
xPix3272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[32] VREF PIX_IN[3272] NB2 NB1 CSA_VREF pixel
xPix3273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[32] VREF PIX_IN[3273] NB2 NB1 CSA_VREF pixel
xPix3274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[32] VREF PIX_IN[3274] NB2 NB1 CSA_VREF pixel
xPix3275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[32] VREF PIX_IN[3275] NB2 NB1 CSA_VREF pixel
xPix3276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[32] VREF PIX_IN[3276] NB2 NB1 CSA_VREF pixel
xPix3277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[32] VREF PIX_IN[3277] NB2 NB1 CSA_VREF pixel
xPix3278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[32] VREF PIX_IN[3278] NB2 NB1 CSA_VREF pixel
xPix3279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[32] VREF PIX_IN[3279] NB2 NB1 CSA_VREF pixel
xPix3280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[32] VREF PIX_IN[3280] NB2 NB1 CSA_VREF pixel
xPix3281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[32] VREF PIX_IN[3281] NB2 NB1 CSA_VREF pixel
xPix3282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[32] VREF PIX_IN[3282] NB2 NB1 CSA_VREF pixel
xPix3283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[32] VREF PIX_IN[3283] NB2 NB1 CSA_VREF pixel
xPix3284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[32] VREF PIX_IN[3284] NB2 NB1 CSA_VREF pixel
xPix3285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[32] VREF PIX_IN[3285] NB2 NB1 CSA_VREF pixel
xPix3286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[32] VREF PIX_IN[3286] NB2 NB1 CSA_VREF pixel
xPix3287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[32] VREF PIX_IN[3287] NB2 NB1 CSA_VREF pixel
xPix3288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[32] VREF PIX_IN[3288] NB2 NB1 CSA_VREF pixel
xPix3289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[32] VREF PIX_IN[3289] NB2 NB1 CSA_VREF pixel
xPix3290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[32] VREF PIX_IN[3290] NB2 NB1 CSA_VREF pixel
xPix3291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[32] VREF PIX_IN[3291] NB2 NB1 CSA_VREF pixel
xPix3292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[32] VREF PIX_IN[3292] NB2 NB1 CSA_VREF pixel
xPix3293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[32] VREF PIX_IN[3293] NB2 NB1 CSA_VREF pixel
xPix3294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[32] VREF PIX_IN[3294] NB2 NB1 CSA_VREF pixel
xPix3295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[32] VREF PIX_IN[3295] NB2 NB1 CSA_VREF pixel
xPix3296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[32] VREF PIX_IN[3296] NB2 NB1 CSA_VREF pixel
xPix3297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[32] VREF PIX_IN[3297] NB2 NB1 CSA_VREF pixel
xPix3298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[32] VREF PIX_IN[3298] NB2 NB1 CSA_VREF pixel
xPix3299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[32] VREF PIX_IN[3299] NB2 NB1 CSA_VREF pixel
xPix3300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[33] VREF PIX_IN[3300] NB2 NB1 CSA_VREF pixel
xPix3301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[33] VREF PIX_IN[3301] NB2 NB1 CSA_VREF pixel
xPix3302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[33] VREF PIX_IN[3302] NB2 NB1 CSA_VREF pixel
xPix3303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[33] VREF PIX_IN[3303] NB2 NB1 CSA_VREF pixel
xPix3304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[33] VREF PIX_IN[3304] NB2 NB1 CSA_VREF pixel
xPix3305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[33] VREF PIX_IN[3305] NB2 NB1 CSA_VREF pixel
xPix3306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[33] VREF PIX_IN[3306] NB2 NB1 CSA_VREF pixel
xPix3307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[33] VREF PIX_IN[3307] NB2 NB1 CSA_VREF pixel
xPix3308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[33] VREF PIX_IN[3308] NB2 NB1 CSA_VREF pixel
xPix3309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[33] VREF PIX_IN[3309] NB2 NB1 CSA_VREF pixel
xPix3310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[33] VREF PIX_IN[3310] NB2 NB1 CSA_VREF pixel
xPix3311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[33] VREF PIX_IN[3311] NB2 NB1 CSA_VREF pixel
xPix3312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[33] VREF PIX_IN[3312] NB2 NB1 CSA_VREF pixel
xPix3313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[33] VREF PIX_IN[3313] NB2 NB1 CSA_VREF pixel
xPix3314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[33] VREF PIX_IN[3314] NB2 NB1 CSA_VREF pixel
xPix3315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[33] VREF PIX_IN[3315] NB2 NB1 CSA_VREF pixel
xPix3316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[33] VREF PIX_IN[3316] NB2 NB1 CSA_VREF pixel
xPix3317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[33] VREF PIX_IN[3317] NB2 NB1 CSA_VREF pixel
xPix3318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[33] VREF PIX_IN[3318] NB2 NB1 CSA_VREF pixel
xPix3319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[33] VREF PIX_IN[3319] NB2 NB1 CSA_VREF pixel
xPix3320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[33] VREF PIX_IN[3320] NB2 NB1 CSA_VREF pixel
xPix3321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[33] VREF PIX_IN[3321] NB2 NB1 CSA_VREF pixel
xPix3322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[33] VREF PIX_IN[3322] NB2 NB1 CSA_VREF pixel
xPix3323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[33] VREF PIX_IN[3323] NB2 NB1 CSA_VREF pixel
xPix3324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[33] VREF PIX_IN[3324] NB2 NB1 CSA_VREF pixel
xPix3325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[33] VREF PIX_IN[3325] NB2 NB1 CSA_VREF pixel
xPix3326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[33] VREF PIX_IN[3326] NB2 NB1 CSA_VREF pixel
xPix3327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[33] VREF PIX_IN[3327] NB2 NB1 CSA_VREF pixel
xPix3328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[33] VREF PIX_IN[3328] NB2 NB1 CSA_VREF pixel
xPix3329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[33] VREF PIX_IN[3329] NB2 NB1 CSA_VREF pixel
xPix3330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[33] VREF PIX_IN[3330] NB2 NB1 CSA_VREF pixel
xPix3331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[33] VREF PIX_IN[3331] NB2 NB1 CSA_VREF pixel
xPix3332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[33] VREF PIX_IN[3332] NB2 NB1 CSA_VREF pixel
xPix3333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[33] VREF PIX_IN[3333] NB2 NB1 CSA_VREF pixel
xPix3334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[33] VREF PIX_IN[3334] NB2 NB1 CSA_VREF pixel
xPix3335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[33] VREF PIX_IN[3335] NB2 NB1 CSA_VREF pixel
xPix3336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[33] VREF PIX_IN[3336] NB2 NB1 CSA_VREF pixel
xPix3337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[33] VREF PIX_IN[3337] NB2 NB1 CSA_VREF pixel
xPix3338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[33] VREF PIX_IN[3338] NB2 NB1 CSA_VREF pixel
xPix3339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[33] VREF PIX_IN[3339] NB2 NB1 CSA_VREF pixel
xPix3340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[33] VREF PIX_IN[3340] NB2 NB1 CSA_VREF pixel
xPix3341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[33] VREF PIX_IN[3341] NB2 NB1 CSA_VREF pixel
xPix3342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[33] VREF PIX_IN[3342] NB2 NB1 CSA_VREF pixel
xPix3343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[33] VREF PIX_IN[3343] NB2 NB1 CSA_VREF pixel
xPix3344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[33] VREF PIX_IN[3344] NB2 NB1 CSA_VREF pixel
xPix3345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[33] VREF PIX_IN[3345] NB2 NB1 CSA_VREF pixel
xPix3346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[33] VREF PIX_IN[3346] NB2 NB1 CSA_VREF pixel
xPix3347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[33] VREF PIX_IN[3347] NB2 NB1 CSA_VREF pixel
xPix3348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[33] VREF PIX_IN[3348] NB2 NB1 CSA_VREF pixel
xPix3349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[33] VREF PIX_IN[3349] NB2 NB1 CSA_VREF pixel
xPix3350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[33] VREF PIX_IN[3350] NB2 NB1 CSA_VREF pixel
xPix3351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[33] VREF PIX_IN[3351] NB2 NB1 CSA_VREF pixel
xPix3352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[33] VREF PIX_IN[3352] NB2 NB1 CSA_VREF pixel
xPix3353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[33] VREF PIX_IN[3353] NB2 NB1 CSA_VREF pixel
xPix3354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[33] VREF PIX_IN[3354] NB2 NB1 CSA_VREF pixel
xPix3355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[33] VREF PIX_IN[3355] NB2 NB1 CSA_VREF pixel
xPix3356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[33] VREF PIX_IN[3356] NB2 NB1 CSA_VREF pixel
xPix3357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[33] VREF PIX_IN[3357] NB2 NB1 CSA_VREF pixel
xPix3358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[33] VREF PIX_IN[3358] NB2 NB1 CSA_VREF pixel
xPix3359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[33] VREF PIX_IN[3359] NB2 NB1 CSA_VREF pixel
xPix3360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[33] VREF PIX_IN[3360] NB2 NB1 CSA_VREF pixel
xPix3361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[33] VREF PIX_IN[3361] NB2 NB1 CSA_VREF pixel
xPix3362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[33] VREF PIX_IN[3362] NB2 NB1 CSA_VREF pixel
xPix3363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[33] VREF PIX_IN[3363] NB2 NB1 CSA_VREF pixel
xPix3364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[33] VREF PIX_IN[3364] NB2 NB1 CSA_VREF pixel
xPix3365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[33] VREF PIX_IN[3365] NB2 NB1 CSA_VREF pixel
xPix3366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[33] VREF PIX_IN[3366] NB2 NB1 CSA_VREF pixel
xPix3367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[33] VREF PIX_IN[3367] NB2 NB1 CSA_VREF pixel
xPix3368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[33] VREF PIX_IN[3368] NB2 NB1 CSA_VREF pixel
xPix3369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[33] VREF PIX_IN[3369] NB2 NB1 CSA_VREF pixel
xPix3370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[33] VREF PIX_IN[3370] NB2 NB1 CSA_VREF pixel
xPix3371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[33] VREF PIX_IN[3371] NB2 NB1 CSA_VREF pixel
xPix3372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[33] VREF PIX_IN[3372] NB2 NB1 CSA_VREF pixel
xPix3373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[33] VREF PIX_IN[3373] NB2 NB1 CSA_VREF pixel
xPix3374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[33] VREF PIX_IN[3374] NB2 NB1 CSA_VREF pixel
xPix3375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[33] VREF PIX_IN[3375] NB2 NB1 CSA_VREF pixel
xPix3376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[33] VREF PIX_IN[3376] NB2 NB1 CSA_VREF pixel
xPix3377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[33] VREF PIX_IN[3377] NB2 NB1 CSA_VREF pixel
xPix3378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[33] VREF PIX_IN[3378] NB2 NB1 CSA_VREF pixel
xPix3379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[33] VREF PIX_IN[3379] NB2 NB1 CSA_VREF pixel
xPix3380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[33] VREF PIX_IN[3380] NB2 NB1 CSA_VREF pixel
xPix3381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[33] VREF PIX_IN[3381] NB2 NB1 CSA_VREF pixel
xPix3382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[33] VREF PIX_IN[3382] NB2 NB1 CSA_VREF pixel
xPix3383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[33] VREF PIX_IN[3383] NB2 NB1 CSA_VREF pixel
xPix3384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[33] VREF PIX_IN[3384] NB2 NB1 CSA_VREF pixel
xPix3385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[33] VREF PIX_IN[3385] NB2 NB1 CSA_VREF pixel
xPix3386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[33] VREF PIX_IN[3386] NB2 NB1 CSA_VREF pixel
xPix3387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[33] VREF PIX_IN[3387] NB2 NB1 CSA_VREF pixel
xPix3388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[33] VREF PIX_IN[3388] NB2 NB1 CSA_VREF pixel
xPix3389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[33] VREF PIX_IN[3389] NB2 NB1 CSA_VREF pixel
xPix3390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[33] VREF PIX_IN[3390] NB2 NB1 CSA_VREF pixel
xPix3391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[33] VREF PIX_IN[3391] NB2 NB1 CSA_VREF pixel
xPix3392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[33] VREF PIX_IN[3392] NB2 NB1 CSA_VREF pixel
xPix3393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[33] VREF PIX_IN[3393] NB2 NB1 CSA_VREF pixel
xPix3394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[33] VREF PIX_IN[3394] NB2 NB1 CSA_VREF pixel
xPix3395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[33] VREF PIX_IN[3395] NB2 NB1 CSA_VREF pixel
xPix3396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[33] VREF PIX_IN[3396] NB2 NB1 CSA_VREF pixel
xPix3397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[33] VREF PIX_IN[3397] NB2 NB1 CSA_VREF pixel
xPix3398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[33] VREF PIX_IN[3398] NB2 NB1 CSA_VREF pixel
xPix3399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[33] VREF PIX_IN[3399] NB2 NB1 CSA_VREF pixel
xPix3400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[34] VREF PIX_IN[3400] NB2 NB1 CSA_VREF pixel
xPix3401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[34] VREF PIX_IN[3401] NB2 NB1 CSA_VREF pixel
xPix3402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[34] VREF PIX_IN[3402] NB2 NB1 CSA_VREF pixel
xPix3403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[34] VREF PIX_IN[3403] NB2 NB1 CSA_VREF pixel
xPix3404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[34] VREF PIX_IN[3404] NB2 NB1 CSA_VREF pixel
xPix3405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[34] VREF PIX_IN[3405] NB2 NB1 CSA_VREF pixel
xPix3406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[34] VREF PIX_IN[3406] NB2 NB1 CSA_VREF pixel
xPix3407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[34] VREF PIX_IN[3407] NB2 NB1 CSA_VREF pixel
xPix3408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[34] VREF PIX_IN[3408] NB2 NB1 CSA_VREF pixel
xPix3409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[34] VREF PIX_IN[3409] NB2 NB1 CSA_VREF pixel
xPix3410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[34] VREF PIX_IN[3410] NB2 NB1 CSA_VREF pixel
xPix3411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[34] VREF PIX_IN[3411] NB2 NB1 CSA_VREF pixel
xPix3412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[34] VREF PIX_IN[3412] NB2 NB1 CSA_VREF pixel
xPix3413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[34] VREF PIX_IN[3413] NB2 NB1 CSA_VREF pixel
xPix3414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[34] VREF PIX_IN[3414] NB2 NB1 CSA_VREF pixel
xPix3415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[34] VREF PIX_IN[3415] NB2 NB1 CSA_VREF pixel
xPix3416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[34] VREF PIX_IN[3416] NB2 NB1 CSA_VREF pixel
xPix3417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[34] VREF PIX_IN[3417] NB2 NB1 CSA_VREF pixel
xPix3418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[34] VREF PIX_IN[3418] NB2 NB1 CSA_VREF pixel
xPix3419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[34] VREF PIX_IN[3419] NB2 NB1 CSA_VREF pixel
xPix3420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[34] VREF PIX_IN[3420] NB2 NB1 CSA_VREF pixel
xPix3421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[34] VREF PIX_IN[3421] NB2 NB1 CSA_VREF pixel
xPix3422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[34] VREF PIX_IN[3422] NB2 NB1 CSA_VREF pixel
xPix3423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[34] VREF PIX_IN[3423] NB2 NB1 CSA_VREF pixel
xPix3424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[34] VREF PIX_IN[3424] NB2 NB1 CSA_VREF pixel
xPix3425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[34] VREF PIX_IN[3425] NB2 NB1 CSA_VREF pixel
xPix3426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[34] VREF PIX_IN[3426] NB2 NB1 CSA_VREF pixel
xPix3427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[34] VREF PIX_IN[3427] NB2 NB1 CSA_VREF pixel
xPix3428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[34] VREF PIX_IN[3428] NB2 NB1 CSA_VREF pixel
xPix3429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[34] VREF PIX_IN[3429] NB2 NB1 CSA_VREF pixel
xPix3430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[34] VREF PIX_IN[3430] NB2 NB1 CSA_VREF pixel
xPix3431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[34] VREF PIX_IN[3431] NB2 NB1 CSA_VREF pixel
xPix3432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[34] VREF PIX_IN[3432] NB2 NB1 CSA_VREF pixel
xPix3433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[34] VREF PIX_IN[3433] NB2 NB1 CSA_VREF pixel
xPix3434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[34] VREF PIX_IN[3434] NB2 NB1 CSA_VREF pixel
xPix3435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[34] VREF PIX_IN[3435] NB2 NB1 CSA_VREF pixel
xPix3436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[34] VREF PIX_IN[3436] NB2 NB1 CSA_VREF pixel
xPix3437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[34] VREF PIX_IN[3437] NB2 NB1 CSA_VREF pixel
xPix3438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[34] VREF PIX_IN[3438] NB2 NB1 CSA_VREF pixel
xPix3439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[34] VREF PIX_IN[3439] NB2 NB1 CSA_VREF pixel
xPix3440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[34] VREF PIX_IN[3440] NB2 NB1 CSA_VREF pixel
xPix3441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[34] VREF PIX_IN[3441] NB2 NB1 CSA_VREF pixel
xPix3442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[34] VREF PIX_IN[3442] NB2 NB1 CSA_VREF pixel
xPix3443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[34] VREF PIX_IN[3443] NB2 NB1 CSA_VREF pixel
xPix3444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[34] VREF PIX_IN[3444] NB2 NB1 CSA_VREF pixel
xPix3445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[34] VREF PIX_IN[3445] NB2 NB1 CSA_VREF pixel
xPix3446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[34] VREF PIX_IN[3446] NB2 NB1 CSA_VREF pixel
xPix3447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[34] VREF PIX_IN[3447] NB2 NB1 CSA_VREF pixel
xPix3448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[34] VREF PIX_IN[3448] NB2 NB1 CSA_VREF pixel
xPix3449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[34] VREF PIX_IN[3449] NB2 NB1 CSA_VREF pixel
xPix3450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[34] VREF PIX_IN[3450] NB2 NB1 CSA_VREF pixel
xPix3451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[34] VREF PIX_IN[3451] NB2 NB1 CSA_VREF pixel
xPix3452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[34] VREF PIX_IN[3452] NB2 NB1 CSA_VREF pixel
xPix3453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[34] VREF PIX_IN[3453] NB2 NB1 CSA_VREF pixel
xPix3454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[34] VREF PIX_IN[3454] NB2 NB1 CSA_VREF pixel
xPix3455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[34] VREF PIX_IN[3455] NB2 NB1 CSA_VREF pixel
xPix3456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[34] VREF PIX_IN[3456] NB2 NB1 CSA_VREF pixel
xPix3457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[34] VREF PIX_IN[3457] NB2 NB1 CSA_VREF pixel
xPix3458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[34] VREF PIX_IN[3458] NB2 NB1 CSA_VREF pixel
xPix3459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[34] VREF PIX_IN[3459] NB2 NB1 CSA_VREF pixel
xPix3460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[34] VREF PIX_IN[3460] NB2 NB1 CSA_VREF pixel
xPix3461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[34] VREF PIX_IN[3461] NB2 NB1 CSA_VREF pixel
xPix3462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[34] VREF PIX_IN[3462] NB2 NB1 CSA_VREF pixel
xPix3463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[34] VREF PIX_IN[3463] NB2 NB1 CSA_VREF pixel
xPix3464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[34] VREF PIX_IN[3464] NB2 NB1 CSA_VREF pixel
xPix3465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[34] VREF PIX_IN[3465] NB2 NB1 CSA_VREF pixel
xPix3466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[34] VREF PIX_IN[3466] NB2 NB1 CSA_VREF pixel
xPix3467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[34] VREF PIX_IN[3467] NB2 NB1 CSA_VREF pixel
xPix3468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[34] VREF PIX_IN[3468] NB2 NB1 CSA_VREF pixel
xPix3469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[34] VREF PIX_IN[3469] NB2 NB1 CSA_VREF pixel
xPix3470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[34] VREF PIX_IN[3470] NB2 NB1 CSA_VREF pixel
xPix3471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[34] VREF PIX_IN[3471] NB2 NB1 CSA_VREF pixel
xPix3472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[34] VREF PIX_IN[3472] NB2 NB1 CSA_VREF pixel
xPix3473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[34] VREF PIX_IN[3473] NB2 NB1 CSA_VREF pixel
xPix3474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[34] VREF PIX_IN[3474] NB2 NB1 CSA_VREF pixel
xPix3475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[34] VREF PIX_IN[3475] NB2 NB1 CSA_VREF pixel
xPix3476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[34] VREF PIX_IN[3476] NB2 NB1 CSA_VREF pixel
xPix3477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[34] VREF PIX_IN[3477] NB2 NB1 CSA_VREF pixel
xPix3478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[34] VREF PIX_IN[3478] NB2 NB1 CSA_VREF pixel
xPix3479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[34] VREF PIX_IN[3479] NB2 NB1 CSA_VREF pixel
xPix3480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[34] VREF PIX_IN[3480] NB2 NB1 CSA_VREF pixel
xPix3481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[34] VREF PIX_IN[3481] NB2 NB1 CSA_VREF pixel
xPix3482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[34] VREF PIX_IN[3482] NB2 NB1 CSA_VREF pixel
xPix3483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[34] VREF PIX_IN[3483] NB2 NB1 CSA_VREF pixel
xPix3484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[34] VREF PIX_IN[3484] NB2 NB1 CSA_VREF pixel
xPix3485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[34] VREF PIX_IN[3485] NB2 NB1 CSA_VREF pixel
xPix3486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[34] VREF PIX_IN[3486] NB2 NB1 CSA_VREF pixel
xPix3487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[34] VREF PIX_IN[3487] NB2 NB1 CSA_VREF pixel
xPix3488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[34] VREF PIX_IN[3488] NB2 NB1 CSA_VREF pixel
xPix3489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[34] VREF PIX_IN[3489] NB2 NB1 CSA_VREF pixel
xPix3490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[34] VREF PIX_IN[3490] NB2 NB1 CSA_VREF pixel
xPix3491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[34] VREF PIX_IN[3491] NB2 NB1 CSA_VREF pixel
xPix3492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[34] VREF PIX_IN[3492] NB2 NB1 CSA_VREF pixel
xPix3493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[34] VREF PIX_IN[3493] NB2 NB1 CSA_VREF pixel
xPix3494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[34] VREF PIX_IN[3494] NB2 NB1 CSA_VREF pixel
xPix3495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[34] VREF PIX_IN[3495] NB2 NB1 CSA_VREF pixel
xPix3496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[34] VREF PIX_IN[3496] NB2 NB1 CSA_VREF pixel
xPix3497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[34] VREF PIX_IN[3497] NB2 NB1 CSA_VREF pixel
xPix3498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[34] VREF PIX_IN[3498] NB2 NB1 CSA_VREF pixel
xPix3499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[34] VREF PIX_IN[3499] NB2 NB1 CSA_VREF pixel
xPix3500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[35] VREF PIX_IN[3500] NB2 NB1 CSA_VREF pixel
xPix3501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[35] VREF PIX_IN[3501] NB2 NB1 CSA_VREF pixel
xPix3502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[35] VREF PIX_IN[3502] NB2 NB1 CSA_VREF pixel
xPix3503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[35] VREF PIX_IN[3503] NB2 NB1 CSA_VREF pixel
xPix3504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[35] VREF PIX_IN[3504] NB2 NB1 CSA_VREF pixel
xPix3505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[35] VREF PIX_IN[3505] NB2 NB1 CSA_VREF pixel
xPix3506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[35] VREF PIX_IN[3506] NB2 NB1 CSA_VREF pixel
xPix3507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[35] VREF PIX_IN[3507] NB2 NB1 CSA_VREF pixel
xPix3508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[35] VREF PIX_IN[3508] NB2 NB1 CSA_VREF pixel
xPix3509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[35] VREF PIX_IN[3509] NB2 NB1 CSA_VREF pixel
xPix3510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[35] VREF PIX_IN[3510] NB2 NB1 CSA_VREF pixel
xPix3511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[35] VREF PIX_IN[3511] NB2 NB1 CSA_VREF pixel
xPix3512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[35] VREF PIX_IN[3512] NB2 NB1 CSA_VREF pixel
xPix3513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[35] VREF PIX_IN[3513] NB2 NB1 CSA_VREF pixel
xPix3514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[35] VREF PIX_IN[3514] NB2 NB1 CSA_VREF pixel
xPix3515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[35] VREF PIX_IN[3515] NB2 NB1 CSA_VREF pixel
xPix3516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[35] VREF PIX_IN[3516] NB2 NB1 CSA_VREF pixel
xPix3517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[35] VREF PIX_IN[3517] NB2 NB1 CSA_VREF pixel
xPix3518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[35] VREF PIX_IN[3518] NB2 NB1 CSA_VREF pixel
xPix3519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[35] VREF PIX_IN[3519] NB2 NB1 CSA_VREF pixel
xPix3520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[35] VREF PIX_IN[3520] NB2 NB1 CSA_VREF pixel
xPix3521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[35] VREF PIX_IN[3521] NB2 NB1 CSA_VREF pixel
xPix3522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[35] VREF PIX_IN[3522] NB2 NB1 CSA_VREF pixel
xPix3523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[35] VREF PIX_IN[3523] NB2 NB1 CSA_VREF pixel
xPix3524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[35] VREF PIX_IN[3524] NB2 NB1 CSA_VREF pixel
xPix3525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[35] VREF PIX_IN[3525] NB2 NB1 CSA_VREF pixel
xPix3526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[35] VREF PIX_IN[3526] NB2 NB1 CSA_VREF pixel
xPix3527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[35] VREF PIX_IN[3527] NB2 NB1 CSA_VREF pixel
xPix3528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[35] VREF PIX_IN[3528] NB2 NB1 CSA_VREF pixel
xPix3529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[35] VREF PIX_IN[3529] NB2 NB1 CSA_VREF pixel
xPix3530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[35] VREF PIX_IN[3530] NB2 NB1 CSA_VREF pixel
xPix3531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[35] VREF PIX_IN[3531] NB2 NB1 CSA_VREF pixel
xPix3532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[35] VREF PIX_IN[3532] NB2 NB1 CSA_VREF pixel
xPix3533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[35] VREF PIX_IN[3533] NB2 NB1 CSA_VREF pixel
xPix3534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[35] VREF PIX_IN[3534] NB2 NB1 CSA_VREF pixel
xPix3535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[35] VREF PIX_IN[3535] NB2 NB1 CSA_VREF pixel
xPix3536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[35] VREF PIX_IN[3536] NB2 NB1 CSA_VREF pixel
xPix3537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[35] VREF PIX_IN[3537] NB2 NB1 CSA_VREF pixel
xPix3538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[35] VREF PIX_IN[3538] NB2 NB1 CSA_VREF pixel
xPix3539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[35] VREF PIX_IN[3539] NB2 NB1 CSA_VREF pixel
xPix3540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[35] VREF PIX_IN[3540] NB2 NB1 CSA_VREF pixel
xPix3541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[35] VREF PIX_IN[3541] NB2 NB1 CSA_VREF pixel
xPix3542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[35] VREF PIX_IN[3542] NB2 NB1 CSA_VREF pixel
xPix3543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[35] VREF PIX_IN[3543] NB2 NB1 CSA_VREF pixel
xPix3544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[35] VREF PIX_IN[3544] NB2 NB1 CSA_VREF pixel
xPix3545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[35] VREF PIX_IN[3545] NB2 NB1 CSA_VREF pixel
xPix3546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[35] VREF PIX_IN[3546] NB2 NB1 CSA_VREF pixel
xPix3547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[35] VREF PIX_IN[3547] NB2 NB1 CSA_VREF pixel
xPix3548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[35] VREF PIX_IN[3548] NB2 NB1 CSA_VREF pixel
xPix3549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[35] VREF PIX_IN[3549] NB2 NB1 CSA_VREF pixel
xPix3550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[35] VREF PIX_IN[3550] NB2 NB1 CSA_VREF pixel
xPix3551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[35] VREF PIX_IN[3551] NB2 NB1 CSA_VREF pixel
xPix3552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[35] VREF PIX_IN[3552] NB2 NB1 CSA_VREF pixel
xPix3553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[35] VREF PIX_IN[3553] NB2 NB1 CSA_VREF pixel
xPix3554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[35] VREF PIX_IN[3554] NB2 NB1 CSA_VREF pixel
xPix3555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[35] VREF PIX_IN[3555] NB2 NB1 CSA_VREF pixel
xPix3556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[35] VREF PIX_IN[3556] NB2 NB1 CSA_VREF pixel
xPix3557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[35] VREF PIX_IN[3557] NB2 NB1 CSA_VREF pixel
xPix3558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[35] VREF PIX_IN[3558] NB2 NB1 CSA_VREF pixel
xPix3559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[35] VREF PIX_IN[3559] NB2 NB1 CSA_VREF pixel
xPix3560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[35] VREF PIX_IN[3560] NB2 NB1 CSA_VREF pixel
xPix3561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[35] VREF PIX_IN[3561] NB2 NB1 CSA_VREF pixel
xPix3562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[35] VREF PIX_IN[3562] NB2 NB1 CSA_VREF pixel
xPix3563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[35] VREF PIX_IN[3563] NB2 NB1 CSA_VREF pixel
xPix3564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[35] VREF PIX_IN[3564] NB2 NB1 CSA_VREF pixel
xPix3565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[35] VREF PIX_IN[3565] NB2 NB1 CSA_VREF pixel
xPix3566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[35] VREF PIX_IN[3566] NB2 NB1 CSA_VREF pixel
xPix3567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[35] VREF PIX_IN[3567] NB2 NB1 CSA_VREF pixel
xPix3568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[35] VREF PIX_IN[3568] NB2 NB1 CSA_VREF pixel
xPix3569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[35] VREF PIX_IN[3569] NB2 NB1 CSA_VREF pixel
xPix3570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[35] VREF PIX_IN[3570] NB2 NB1 CSA_VREF pixel
xPix3571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[35] VREF PIX_IN[3571] NB2 NB1 CSA_VREF pixel
xPix3572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[35] VREF PIX_IN[3572] NB2 NB1 CSA_VREF pixel
xPix3573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[35] VREF PIX_IN[3573] NB2 NB1 CSA_VREF pixel
xPix3574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[35] VREF PIX_IN[3574] NB2 NB1 CSA_VREF pixel
xPix3575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[35] VREF PIX_IN[3575] NB2 NB1 CSA_VREF pixel
xPix3576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[35] VREF PIX_IN[3576] NB2 NB1 CSA_VREF pixel
xPix3577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[35] VREF PIX_IN[3577] NB2 NB1 CSA_VREF pixel
xPix3578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[35] VREF PIX_IN[3578] NB2 NB1 CSA_VREF pixel
xPix3579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[35] VREF PIX_IN[3579] NB2 NB1 CSA_VREF pixel
xPix3580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[35] VREF PIX_IN[3580] NB2 NB1 CSA_VREF pixel
xPix3581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[35] VREF PIX_IN[3581] NB2 NB1 CSA_VREF pixel
xPix3582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[35] VREF PIX_IN[3582] NB2 NB1 CSA_VREF pixel
xPix3583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[35] VREF PIX_IN[3583] NB2 NB1 CSA_VREF pixel
xPix3584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[35] VREF PIX_IN[3584] NB2 NB1 CSA_VREF pixel
xPix3585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[35] VREF PIX_IN[3585] NB2 NB1 CSA_VREF pixel
xPix3586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[35] VREF PIX_IN[3586] NB2 NB1 CSA_VREF pixel
xPix3587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[35] VREF PIX_IN[3587] NB2 NB1 CSA_VREF pixel
xPix3588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[35] VREF PIX_IN[3588] NB2 NB1 CSA_VREF pixel
xPix3589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[35] VREF PIX_IN[3589] NB2 NB1 CSA_VREF pixel
xPix3590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[35] VREF PIX_IN[3590] NB2 NB1 CSA_VREF pixel
xPix3591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[35] VREF PIX_IN[3591] NB2 NB1 CSA_VREF pixel
xPix3592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[35] VREF PIX_IN[3592] NB2 NB1 CSA_VREF pixel
xPix3593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[35] VREF PIX_IN[3593] NB2 NB1 CSA_VREF pixel
xPix3594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[35] VREF PIX_IN[3594] NB2 NB1 CSA_VREF pixel
xPix3595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[35] VREF PIX_IN[3595] NB2 NB1 CSA_VREF pixel
xPix3596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[35] VREF PIX_IN[3596] NB2 NB1 CSA_VREF pixel
xPix3597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[35] VREF PIX_IN[3597] NB2 NB1 CSA_VREF pixel
xPix3598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[35] VREF PIX_IN[3598] NB2 NB1 CSA_VREF pixel
xPix3599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[35] VREF PIX_IN[3599] NB2 NB1 CSA_VREF pixel
xPix3600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[36] VREF PIX_IN[3600] NB2 NB1 CSA_VREF pixel
xPix3601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[36] VREF PIX_IN[3601] NB2 NB1 CSA_VREF pixel
xPix3602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[36] VREF PIX_IN[3602] NB2 NB1 CSA_VREF pixel
xPix3603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[36] VREF PIX_IN[3603] NB2 NB1 CSA_VREF pixel
xPix3604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[36] VREF PIX_IN[3604] NB2 NB1 CSA_VREF pixel
xPix3605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[36] VREF PIX_IN[3605] NB2 NB1 CSA_VREF pixel
xPix3606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[36] VREF PIX_IN[3606] NB2 NB1 CSA_VREF pixel
xPix3607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[36] VREF PIX_IN[3607] NB2 NB1 CSA_VREF pixel
xPix3608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[36] VREF PIX_IN[3608] NB2 NB1 CSA_VREF pixel
xPix3609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[36] VREF PIX_IN[3609] NB2 NB1 CSA_VREF pixel
xPix3610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[36] VREF PIX_IN[3610] NB2 NB1 CSA_VREF pixel
xPix3611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[36] VREF PIX_IN[3611] NB2 NB1 CSA_VREF pixel
xPix3612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[36] VREF PIX_IN[3612] NB2 NB1 CSA_VREF pixel
xPix3613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[36] VREF PIX_IN[3613] NB2 NB1 CSA_VREF pixel
xPix3614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[36] VREF PIX_IN[3614] NB2 NB1 CSA_VREF pixel
xPix3615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[36] VREF PIX_IN[3615] NB2 NB1 CSA_VREF pixel
xPix3616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[36] VREF PIX_IN[3616] NB2 NB1 CSA_VREF pixel
xPix3617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[36] VREF PIX_IN[3617] NB2 NB1 CSA_VREF pixel
xPix3618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[36] VREF PIX_IN[3618] NB2 NB1 CSA_VREF pixel
xPix3619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[36] VREF PIX_IN[3619] NB2 NB1 CSA_VREF pixel
xPix3620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[36] VREF PIX_IN[3620] NB2 NB1 CSA_VREF pixel
xPix3621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[36] VREF PIX_IN[3621] NB2 NB1 CSA_VREF pixel
xPix3622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[36] VREF PIX_IN[3622] NB2 NB1 CSA_VREF pixel
xPix3623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[36] VREF PIX_IN[3623] NB2 NB1 CSA_VREF pixel
xPix3624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[36] VREF PIX_IN[3624] NB2 NB1 CSA_VREF pixel
xPix3625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[36] VREF PIX_IN[3625] NB2 NB1 CSA_VREF pixel
xPix3626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[36] VREF PIX_IN[3626] NB2 NB1 CSA_VREF pixel
xPix3627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[36] VREF PIX_IN[3627] NB2 NB1 CSA_VREF pixel
xPix3628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[36] VREF PIX_IN[3628] NB2 NB1 CSA_VREF pixel
xPix3629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[36] VREF PIX_IN[3629] NB2 NB1 CSA_VREF pixel
xPix3630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[36] VREF PIX_IN[3630] NB2 NB1 CSA_VREF pixel
xPix3631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[36] VREF PIX_IN[3631] NB2 NB1 CSA_VREF pixel
xPix3632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[36] VREF PIX_IN[3632] NB2 NB1 CSA_VREF pixel
xPix3633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[36] VREF PIX_IN[3633] NB2 NB1 CSA_VREF pixel
xPix3634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[36] VREF PIX_IN[3634] NB2 NB1 CSA_VREF pixel
xPix3635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[36] VREF PIX_IN[3635] NB2 NB1 CSA_VREF pixel
xPix3636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[36] VREF PIX_IN[3636] NB2 NB1 CSA_VREF pixel
xPix3637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[36] VREF PIX_IN[3637] NB2 NB1 CSA_VREF pixel
xPix3638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[36] VREF PIX_IN[3638] NB2 NB1 CSA_VREF pixel
xPix3639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[36] VREF PIX_IN[3639] NB2 NB1 CSA_VREF pixel
xPix3640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[36] VREF PIX_IN[3640] NB2 NB1 CSA_VREF pixel
xPix3641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[36] VREF PIX_IN[3641] NB2 NB1 CSA_VREF pixel
xPix3642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[36] VREF PIX_IN[3642] NB2 NB1 CSA_VREF pixel
xPix3643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[36] VREF PIX_IN[3643] NB2 NB1 CSA_VREF pixel
xPix3644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[36] VREF PIX_IN[3644] NB2 NB1 CSA_VREF pixel
xPix3645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[36] VREF PIX_IN[3645] NB2 NB1 CSA_VREF pixel
xPix3646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[36] VREF PIX_IN[3646] NB2 NB1 CSA_VREF pixel
xPix3647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[36] VREF PIX_IN[3647] NB2 NB1 CSA_VREF pixel
xPix3648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[36] VREF PIX_IN[3648] NB2 NB1 CSA_VREF pixel
xPix3649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[36] VREF PIX_IN[3649] NB2 NB1 CSA_VREF pixel
xPix3650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[36] VREF PIX_IN[3650] NB2 NB1 CSA_VREF pixel
xPix3651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[36] VREF PIX_IN[3651] NB2 NB1 CSA_VREF pixel
xPix3652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[36] VREF PIX_IN[3652] NB2 NB1 CSA_VREF pixel
xPix3653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[36] VREF PIX_IN[3653] NB2 NB1 CSA_VREF pixel
xPix3654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[36] VREF PIX_IN[3654] NB2 NB1 CSA_VREF pixel
xPix3655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[36] VREF PIX_IN[3655] NB2 NB1 CSA_VREF pixel
xPix3656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[36] VREF PIX_IN[3656] NB2 NB1 CSA_VREF pixel
xPix3657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[36] VREF PIX_IN[3657] NB2 NB1 CSA_VREF pixel
xPix3658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[36] VREF PIX_IN[3658] NB2 NB1 CSA_VREF pixel
xPix3659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[36] VREF PIX_IN[3659] NB2 NB1 CSA_VREF pixel
xPix3660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[36] VREF PIX_IN[3660] NB2 NB1 CSA_VREF pixel
xPix3661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[36] VREF PIX_IN[3661] NB2 NB1 CSA_VREF pixel
xPix3662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[36] VREF PIX_IN[3662] NB2 NB1 CSA_VREF pixel
xPix3663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[36] VREF PIX_IN[3663] NB2 NB1 CSA_VREF pixel
xPix3664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[36] VREF PIX_IN[3664] NB2 NB1 CSA_VREF pixel
xPix3665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[36] VREF PIX_IN[3665] NB2 NB1 CSA_VREF pixel
xPix3666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[36] VREF PIX_IN[3666] NB2 NB1 CSA_VREF pixel
xPix3667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[36] VREF PIX_IN[3667] NB2 NB1 CSA_VREF pixel
xPix3668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[36] VREF PIX_IN[3668] NB2 NB1 CSA_VREF pixel
xPix3669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[36] VREF PIX_IN[3669] NB2 NB1 CSA_VREF pixel
xPix3670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[36] VREF PIX_IN[3670] NB2 NB1 CSA_VREF pixel
xPix3671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[36] VREF PIX_IN[3671] NB2 NB1 CSA_VREF pixel
xPix3672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[36] VREF PIX_IN[3672] NB2 NB1 CSA_VREF pixel
xPix3673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[36] VREF PIX_IN[3673] NB2 NB1 CSA_VREF pixel
xPix3674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[36] VREF PIX_IN[3674] NB2 NB1 CSA_VREF pixel
xPix3675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[36] VREF PIX_IN[3675] NB2 NB1 CSA_VREF pixel
xPix3676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[36] VREF PIX_IN[3676] NB2 NB1 CSA_VREF pixel
xPix3677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[36] VREF PIX_IN[3677] NB2 NB1 CSA_VREF pixel
xPix3678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[36] VREF PIX_IN[3678] NB2 NB1 CSA_VREF pixel
xPix3679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[36] VREF PIX_IN[3679] NB2 NB1 CSA_VREF pixel
xPix3680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[36] VREF PIX_IN[3680] NB2 NB1 CSA_VREF pixel
xPix3681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[36] VREF PIX_IN[3681] NB2 NB1 CSA_VREF pixel
xPix3682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[36] VREF PIX_IN[3682] NB2 NB1 CSA_VREF pixel
xPix3683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[36] VREF PIX_IN[3683] NB2 NB1 CSA_VREF pixel
xPix3684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[36] VREF PIX_IN[3684] NB2 NB1 CSA_VREF pixel
xPix3685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[36] VREF PIX_IN[3685] NB2 NB1 CSA_VREF pixel
xPix3686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[36] VREF PIX_IN[3686] NB2 NB1 CSA_VREF pixel
xPix3687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[36] VREF PIX_IN[3687] NB2 NB1 CSA_VREF pixel
xPix3688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[36] VREF PIX_IN[3688] NB2 NB1 CSA_VREF pixel
xPix3689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[36] VREF PIX_IN[3689] NB2 NB1 CSA_VREF pixel
xPix3690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[36] VREF PIX_IN[3690] NB2 NB1 CSA_VREF pixel
xPix3691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[36] VREF PIX_IN[3691] NB2 NB1 CSA_VREF pixel
xPix3692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[36] VREF PIX_IN[3692] NB2 NB1 CSA_VREF pixel
xPix3693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[36] VREF PIX_IN[3693] NB2 NB1 CSA_VREF pixel
xPix3694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[36] VREF PIX_IN[3694] NB2 NB1 CSA_VREF pixel
xPix3695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[36] VREF PIX_IN[3695] NB2 NB1 CSA_VREF pixel
xPix3696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[36] VREF PIX_IN[3696] NB2 NB1 CSA_VREF pixel
xPix3697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[36] VREF PIX_IN[3697] NB2 NB1 CSA_VREF pixel
xPix3698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[36] VREF PIX_IN[3698] NB2 NB1 CSA_VREF pixel
xPix3699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[36] VREF PIX_IN[3699] NB2 NB1 CSA_VREF pixel
xPix3700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[37] VREF PIX_IN[3700] NB2 NB1 CSA_VREF pixel
xPix3701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[37] VREF PIX_IN[3701] NB2 NB1 CSA_VREF pixel
xPix3702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[37] VREF PIX_IN[3702] NB2 NB1 CSA_VREF pixel
xPix3703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[37] VREF PIX_IN[3703] NB2 NB1 CSA_VREF pixel
xPix3704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[37] VREF PIX_IN[3704] NB2 NB1 CSA_VREF pixel
xPix3705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[37] VREF PIX_IN[3705] NB2 NB1 CSA_VREF pixel
xPix3706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[37] VREF PIX_IN[3706] NB2 NB1 CSA_VREF pixel
xPix3707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[37] VREF PIX_IN[3707] NB2 NB1 CSA_VREF pixel
xPix3708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[37] VREF PIX_IN[3708] NB2 NB1 CSA_VREF pixel
xPix3709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[37] VREF PIX_IN[3709] NB2 NB1 CSA_VREF pixel
xPix3710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[37] VREF PIX_IN[3710] NB2 NB1 CSA_VREF pixel
xPix3711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[37] VREF PIX_IN[3711] NB2 NB1 CSA_VREF pixel
xPix3712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[37] VREF PIX_IN[3712] NB2 NB1 CSA_VREF pixel
xPix3713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[37] VREF PIX_IN[3713] NB2 NB1 CSA_VREF pixel
xPix3714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[37] VREF PIX_IN[3714] NB2 NB1 CSA_VREF pixel
xPix3715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[37] VREF PIX_IN[3715] NB2 NB1 CSA_VREF pixel
xPix3716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[37] VREF PIX_IN[3716] NB2 NB1 CSA_VREF pixel
xPix3717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[37] VREF PIX_IN[3717] NB2 NB1 CSA_VREF pixel
xPix3718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[37] VREF PIX_IN[3718] NB2 NB1 CSA_VREF pixel
xPix3719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[37] VREF PIX_IN[3719] NB2 NB1 CSA_VREF pixel
xPix3720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[37] VREF PIX_IN[3720] NB2 NB1 CSA_VREF pixel
xPix3721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[37] VREF PIX_IN[3721] NB2 NB1 CSA_VREF pixel
xPix3722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[37] VREF PIX_IN[3722] NB2 NB1 CSA_VREF pixel
xPix3723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[37] VREF PIX_IN[3723] NB2 NB1 CSA_VREF pixel
xPix3724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[37] VREF PIX_IN[3724] NB2 NB1 CSA_VREF pixel
xPix3725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[37] VREF PIX_IN[3725] NB2 NB1 CSA_VREF pixel
xPix3726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[37] VREF PIX_IN[3726] NB2 NB1 CSA_VREF pixel
xPix3727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[37] VREF PIX_IN[3727] NB2 NB1 CSA_VREF pixel
xPix3728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[37] VREF PIX_IN[3728] NB2 NB1 CSA_VREF pixel
xPix3729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[37] VREF PIX_IN[3729] NB2 NB1 CSA_VREF pixel
xPix3730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[37] VREF PIX_IN[3730] NB2 NB1 CSA_VREF pixel
xPix3731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[37] VREF PIX_IN[3731] NB2 NB1 CSA_VREF pixel
xPix3732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[37] VREF PIX_IN[3732] NB2 NB1 CSA_VREF pixel
xPix3733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[37] VREF PIX_IN[3733] NB2 NB1 CSA_VREF pixel
xPix3734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[37] VREF PIX_IN[3734] NB2 NB1 CSA_VREF pixel
xPix3735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[37] VREF PIX_IN[3735] NB2 NB1 CSA_VREF pixel
xPix3736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[37] VREF PIX_IN[3736] NB2 NB1 CSA_VREF pixel
xPix3737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[37] VREF PIX_IN[3737] NB2 NB1 CSA_VREF pixel
xPix3738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[37] VREF PIX_IN[3738] NB2 NB1 CSA_VREF pixel
xPix3739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[37] VREF PIX_IN[3739] NB2 NB1 CSA_VREF pixel
xPix3740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[37] VREF PIX_IN[3740] NB2 NB1 CSA_VREF pixel
xPix3741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[37] VREF PIX_IN[3741] NB2 NB1 CSA_VREF pixel
xPix3742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[37] VREF PIX_IN[3742] NB2 NB1 CSA_VREF pixel
xPix3743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[37] VREF PIX_IN[3743] NB2 NB1 CSA_VREF pixel
xPix3744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[37] VREF PIX_IN[3744] NB2 NB1 CSA_VREF pixel
xPix3745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[37] VREF PIX_IN[3745] NB2 NB1 CSA_VREF pixel
xPix3746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[37] VREF PIX_IN[3746] NB2 NB1 CSA_VREF pixel
xPix3747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[37] VREF PIX_IN[3747] NB2 NB1 CSA_VREF pixel
xPix3748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[37] VREF PIX_IN[3748] NB2 NB1 CSA_VREF pixel
xPix3749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[37] VREF PIX_IN[3749] NB2 NB1 CSA_VREF pixel
xPix3750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[37] VREF PIX_IN[3750] NB2 NB1 CSA_VREF pixel
xPix3751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[37] VREF PIX_IN[3751] NB2 NB1 CSA_VREF pixel
xPix3752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[37] VREF PIX_IN[3752] NB2 NB1 CSA_VREF pixel
xPix3753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[37] VREF PIX_IN[3753] NB2 NB1 CSA_VREF pixel
xPix3754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[37] VREF PIX_IN[3754] NB2 NB1 CSA_VREF pixel
xPix3755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[37] VREF PIX_IN[3755] NB2 NB1 CSA_VREF pixel
xPix3756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[37] VREF PIX_IN[3756] NB2 NB1 CSA_VREF pixel
xPix3757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[37] VREF PIX_IN[3757] NB2 NB1 CSA_VREF pixel
xPix3758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[37] VREF PIX_IN[3758] NB2 NB1 CSA_VREF pixel
xPix3759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[37] VREF PIX_IN[3759] NB2 NB1 CSA_VREF pixel
xPix3760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[37] VREF PIX_IN[3760] NB2 NB1 CSA_VREF pixel
xPix3761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[37] VREF PIX_IN[3761] NB2 NB1 CSA_VREF pixel
xPix3762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[37] VREF PIX_IN[3762] NB2 NB1 CSA_VREF pixel
xPix3763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[37] VREF PIX_IN[3763] NB2 NB1 CSA_VREF pixel
xPix3764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[37] VREF PIX_IN[3764] NB2 NB1 CSA_VREF pixel
xPix3765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[37] VREF PIX_IN[3765] NB2 NB1 CSA_VREF pixel
xPix3766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[37] VREF PIX_IN[3766] NB2 NB1 CSA_VREF pixel
xPix3767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[37] VREF PIX_IN[3767] NB2 NB1 CSA_VREF pixel
xPix3768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[37] VREF PIX_IN[3768] NB2 NB1 CSA_VREF pixel
xPix3769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[37] VREF PIX_IN[3769] NB2 NB1 CSA_VREF pixel
xPix3770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[37] VREF PIX_IN[3770] NB2 NB1 CSA_VREF pixel
xPix3771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[37] VREF PIX_IN[3771] NB2 NB1 CSA_VREF pixel
xPix3772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[37] VREF PIX_IN[3772] NB2 NB1 CSA_VREF pixel
xPix3773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[37] VREF PIX_IN[3773] NB2 NB1 CSA_VREF pixel
xPix3774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[37] VREF PIX_IN[3774] NB2 NB1 CSA_VREF pixel
xPix3775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[37] VREF PIX_IN[3775] NB2 NB1 CSA_VREF pixel
xPix3776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[37] VREF PIX_IN[3776] NB2 NB1 CSA_VREF pixel
xPix3777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[37] VREF PIX_IN[3777] NB2 NB1 CSA_VREF pixel
xPix3778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[37] VREF PIX_IN[3778] NB2 NB1 CSA_VREF pixel
xPix3779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[37] VREF PIX_IN[3779] NB2 NB1 CSA_VREF pixel
xPix3780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[37] VREF PIX_IN[3780] NB2 NB1 CSA_VREF pixel
xPix3781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[37] VREF PIX_IN[3781] NB2 NB1 CSA_VREF pixel
xPix3782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[37] VREF PIX_IN[3782] NB2 NB1 CSA_VREF pixel
xPix3783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[37] VREF PIX_IN[3783] NB2 NB1 CSA_VREF pixel
xPix3784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[37] VREF PIX_IN[3784] NB2 NB1 CSA_VREF pixel
xPix3785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[37] VREF PIX_IN[3785] NB2 NB1 CSA_VREF pixel
xPix3786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[37] VREF PIX_IN[3786] NB2 NB1 CSA_VREF pixel
xPix3787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[37] VREF PIX_IN[3787] NB2 NB1 CSA_VREF pixel
xPix3788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[37] VREF PIX_IN[3788] NB2 NB1 CSA_VREF pixel
xPix3789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[37] VREF PIX_IN[3789] NB2 NB1 CSA_VREF pixel
xPix3790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[37] VREF PIX_IN[3790] NB2 NB1 CSA_VREF pixel
xPix3791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[37] VREF PIX_IN[3791] NB2 NB1 CSA_VREF pixel
xPix3792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[37] VREF PIX_IN[3792] NB2 NB1 CSA_VREF pixel
xPix3793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[37] VREF PIX_IN[3793] NB2 NB1 CSA_VREF pixel
xPix3794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[37] VREF PIX_IN[3794] NB2 NB1 CSA_VREF pixel
xPix3795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[37] VREF PIX_IN[3795] NB2 NB1 CSA_VREF pixel
xPix3796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[37] VREF PIX_IN[3796] NB2 NB1 CSA_VREF pixel
xPix3797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[37] VREF PIX_IN[3797] NB2 NB1 CSA_VREF pixel
xPix3798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[37] VREF PIX_IN[3798] NB2 NB1 CSA_VREF pixel
xPix3799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[37] VREF PIX_IN[3799] NB2 NB1 CSA_VREF pixel
xPix3800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[38] VREF PIX_IN[3800] NB2 NB1 CSA_VREF pixel
xPix3801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[38] VREF PIX_IN[3801] NB2 NB1 CSA_VREF pixel
xPix3802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[38] VREF PIX_IN[3802] NB2 NB1 CSA_VREF pixel
xPix3803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[38] VREF PIX_IN[3803] NB2 NB1 CSA_VREF pixel
xPix3804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[38] VREF PIX_IN[3804] NB2 NB1 CSA_VREF pixel
xPix3805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[38] VREF PIX_IN[3805] NB2 NB1 CSA_VREF pixel
xPix3806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[38] VREF PIX_IN[3806] NB2 NB1 CSA_VREF pixel
xPix3807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[38] VREF PIX_IN[3807] NB2 NB1 CSA_VREF pixel
xPix3808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[38] VREF PIX_IN[3808] NB2 NB1 CSA_VREF pixel
xPix3809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[38] VREF PIX_IN[3809] NB2 NB1 CSA_VREF pixel
xPix3810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[38] VREF PIX_IN[3810] NB2 NB1 CSA_VREF pixel
xPix3811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[38] VREF PIX_IN[3811] NB2 NB1 CSA_VREF pixel
xPix3812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[38] VREF PIX_IN[3812] NB2 NB1 CSA_VREF pixel
xPix3813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[38] VREF PIX_IN[3813] NB2 NB1 CSA_VREF pixel
xPix3814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[38] VREF PIX_IN[3814] NB2 NB1 CSA_VREF pixel
xPix3815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[38] VREF PIX_IN[3815] NB2 NB1 CSA_VREF pixel
xPix3816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[38] VREF PIX_IN[3816] NB2 NB1 CSA_VREF pixel
xPix3817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[38] VREF PIX_IN[3817] NB2 NB1 CSA_VREF pixel
xPix3818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[38] VREF PIX_IN[3818] NB2 NB1 CSA_VREF pixel
xPix3819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[38] VREF PIX_IN[3819] NB2 NB1 CSA_VREF pixel
xPix3820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[38] VREF PIX_IN[3820] NB2 NB1 CSA_VREF pixel
xPix3821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[38] VREF PIX_IN[3821] NB2 NB1 CSA_VREF pixel
xPix3822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[38] VREF PIX_IN[3822] NB2 NB1 CSA_VREF pixel
xPix3823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[38] VREF PIX_IN[3823] NB2 NB1 CSA_VREF pixel
xPix3824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[38] VREF PIX_IN[3824] NB2 NB1 CSA_VREF pixel
xPix3825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[38] VREF PIX_IN[3825] NB2 NB1 CSA_VREF pixel
xPix3826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[38] VREF PIX_IN[3826] NB2 NB1 CSA_VREF pixel
xPix3827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[38] VREF PIX_IN[3827] NB2 NB1 CSA_VREF pixel
xPix3828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[38] VREF PIX_IN[3828] NB2 NB1 CSA_VREF pixel
xPix3829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[38] VREF PIX_IN[3829] NB2 NB1 CSA_VREF pixel
xPix3830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[38] VREF PIX_IN[3830] NB2 NB1 CSA_VREF pixel
xPix3831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[38] VREF PIX_IN[3831] NB2 NB1 CSA_VREF pixel
xPix3832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[38] VREF PIX_IN[3832] NB2 NB1 CSA_VREF pixel
xPix3833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[38] VREF PIX_IN[3833] NB2 NB1 CSA_VREF pixel
xPix3834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[38] VREF PIX_IN[3834] NB2 NB1 CSA_VREF pixel
xPix3835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[38] VREF PIX_IN[3835] NB2 NB1 CSA_VREF pixel
xPix3836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[38] VREF PIX_IN[3836] NB2 NB1 CSA_VREF pixel
xPix3837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[38] VREF PIX_IN[3837] NB2 NB1 CSA_VREF pixel
xPix3838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[38] VREF PIX_IN[3838] NB2 NB1 CSA_VREF pixel
xPix3839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[38] VREF PIX_IN[3839] NB2 NB1 CSA_VREF pixel
xPix3840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[38] VREF PIX_IN[3840] NB2 NB1 CSA_VREF pixel
xPix3841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[38] VREF PIX_IN[3841] NB2 NB1 CSA_VREF pixel
xPix3842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[38] VREF PIX_IN[3842] NB2 NB1 CSA_VREF pixel
xPix3843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[38] VREF PIX_IN[3843] NB2 NB1 CSA_VREF pixel
xPix3844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[38] VREF PIX_IN[3844] NB2 NB1 CSA_VREF pixel
xPix3845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[38] VREF PIX_IN[3845] NB2 NB1 CSA_VREF pixel
xPix3846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[38] VREF PIX_IN[3846] NB2 NB1 CSA_VREF pixel
xPix3847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[38] VREF PIX_IN[3847] NB2 NB1 CSA_VREF pixel
xPix3848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[38] VREF PIX_IN[3848] NB2 NB1 CSA_VREF pixel
xPix3849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[38] VREF PIX_IN[3849] NB2 NB1 CSA_VREF pixel
xPix3850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[38] VREF PIX_IN[3850] NB2 NB1 CSA_VREF pixel
xPix3851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[38] VREF PIX_IN[3851] NB2 NB1 CSA_VREF pixel
xPix3852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[38] VREF PIX_IN[3852] NB2 NB1 CSA_VREF pixel
xPix3853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[38] VREF PIX_IN[3853] NB2 NB1 CSA_VREF pixel
xPix3854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[38] VREF PIX_IN[3854] NB2 NB1 CSA_VREF pixel
xPix3855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[38] VREF PIX_IN[3855] NB2 NB1 CSA_VREF pixel
xPix3856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[38] VREF PIX_IN[3856] NB2 NB1 CSA_VREF pixel
xPix3857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[38] VREF PIX_IN[3857] NB2 NB1 CSA_VREF pixel
xPix3858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[38] VREF PIX_IN[3858] NB2 NB1 CSA_VREF pixel
xPix3859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[38] VREF PIX_IN[3859] NB2 NB1 CSA_VREF pixel
xPix3860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[38] VREF PIX_IN[3860] NB2 NB1 CSA_VREF pixel
xPix3861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[38] VREF PIX_IN[3861] NB2 NB1 CSA_VREF pixel
xPix3862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[38] VREF PIX_IN[3862] NB2 NB1 CSA_VREF pixel
xPix3863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[38] VREF PIX_IN[3863] NB2 NB1 CSA_VREF pixel
xPix3864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[38] VREF PIX_IN[3864] NB2 NB1 CSA_VREF pixel
xPix3865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[38] VREF PIX_IN[3865] NB2 NB1 CSA_VREF pixel
xPix3866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[38] VREF PIX_IN[3866] NB2 NB1 CSA_VREF pixel
xPix3867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[38] VREF PIX_IN[3867] NB2 NB1 CSA_VREF pixel
xPix3868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[38] VREF PIX_IN[3868] NB2 NB1 CSA_VREF pixel
xPix3869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[38] VREF PIX_IN[3869] NB2 NB1 CSA_VREF pixel
xPix3870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[38] VREF PIX_IN[3870] NB2 NB1 CSA_VREF pixel
xPix3871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[38] VREF PIX_IN[3871] NB2 NB1 CSA_VREF pixel
xPix3872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[38] VREF PIX_IN[3872] NB2 NB1 CSA_VREF pixel
xPix3873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[38] VREF PIX_IN[3873] NB2 NB1 CSA_VREF pixel
xPix3874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[38] VREF PIX_IN[3874] NB2 NB1 CSA_VREF pixel
xPix3875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[38] VREF PIX_IN[3875] NB2 NB1 CSA_VREF pixel
xPix3876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[38] VREF PIX_IN[3876] NB2 NB1 CSA_VREF pixel
xPix3877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[38] VREF PIX_IN[3877] NB2 NB1 CSA_VREF pixel
xPix3878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[38] VREF PIX_IN[3878] NB2 NB1 CSA_VREF pixel
xPix3879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[38] VREF PIX_IN[3879] NB2 NB1 CSA_VREF pixel
xPix3880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[38] VREF PIX_IN[3880] NB2 NB1 CSA_VREF pixel
xPix3881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[38] VREF PIX_IN[3881] NB2 NB1 CSA_VREF pixel
xPix3882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[38] VREF PIX_IN[3882] NB2 NB1 CSA_VREF pixel
xPix3883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[38] VREF PIX_IN[3883] NB2 NB1 CSA_VREF pixel
xPix3884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[38] VREF PIX_IN[3884] NB2 NB1 CSA_VREF pixel
xPix3885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[38] VREF PIX_IN[3885] NB2 NB1 CSA_VREF pixel
xPix3886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[38] VREF PIX_IN[3886] NB2 NB1 CSA_VREF pixel
xPix3887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[38] VREF PIX_IN[3887] NB2 NB1 CSA_VREF pixel
xPix3888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[38] VREF PIX_IN[3888] NB2 NB1 CSA_VREF pixel
xPix3889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[38] VREF PIX_IN[3889] NB2 NB1 CSA_VREF pixel
xPix3890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[38] VREF PIX_IN[3890] NB2 NB1 CSA_VREF pixel
xPix3891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[38] VREF PIX_IN[3891] NB2 NB1 CSA_VREF pixel
xPix3892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[38] VREF PIX_IN[3892] NB2 NB1 CSA_VREF pixel
xPix3893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[38] VREF PIX_IN[3893] NB2 NB1 CSA_VREF pixel
xPix3894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[38] VREF PIX_IN[3894] NB2 NB1 CSA_VREF pixel
xPix3895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[38] VREF PIX_IN[3895] NB2 NB1 CSA_VREF pixel
xPix3896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[38] VREF PIX_IN[3896] NB2 NB1 CSA_VREF pixel
xPix3897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[38] VREF PIX_IN[3897] NB2 NB1 CSA_VREF pixel
xPix3898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[38] VREF PIX_IN[3898] NB2 NB1 CSA_VREF pixel
xPix3899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[38] VREF PIX_IN[3899] NB2 NB1 CSA_VREF pixel
xPix3900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[39] VREF PIX_IN[3900] NB2 NB1 CSA_VREF pixel
xPix3901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[39] VREF PIX_IN[3901] NB2 NB1 CSA_VREF pixel
xPix3902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[39] VREF PIX_IN[3902] NB2 NB1 CSA_VREF pixel
xPix3903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[39] VREF PIX_IN[3903] NB2 NB1 CSA_VREF pixel
xPix3904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[39] VREF PIX_IN[3904] NB2 NB1 CSA_VREF pixel
xPix3905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[39] VREF PIX_IN[3905] NB2 NB1 CSA_VREF pixel
xPix3906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[39] VREF PIX_IN[3906] NB2 NB1 CSA_VREF pixel
xPix3907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[39] VREF PIX_IN[3907] NB2 NB1 CSA_VREF pixel
xPix3908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[39] VREF PIX_IN[3908] NB2 NB1 CSA_VREF pixel
xPix3909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[39] VREF PIX_IN[3909] NB2 NB1 CSA_VREF pixel
xPix3910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[39] VREF PIX_IN[3910] NB2 NB1 CSA_VREF pixel
xPix3911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[39] VREF PIX_IN[3911] NB2 NB1 CSA_VREF pixel
xPix3912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[39] VREF PIX_IN[3912] NB2 NB1 CSA_VREF pixel
xPix3913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[39] VREF PIX_IN[3913] NB2 NB1 CSA_VREF pixel
xPix3914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[39] VREF PIX_IN[3914] NB2 NB1 CSA_VREF pixel
xPix3915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[39] VREF PIX_IN[3915] NB2 NB1 CSA_VREF pixel
xPix3916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[39] VREF PIX_IN[3916] NB2 NB1 CSA_VREF pixel
xPix3917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[39] VREF PIX_IN[3917] NB2 NB1 CSA_VREF pixel
xPix3918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[39] VREF PIX_IN[3918] NB2 NB1 CSA_VREF pixel
xPix3919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[39] VREF PIX_IN[3919] NB2 NB1 CSA_VREF pixel
xPix3920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[39] VREF PIX_IN[3920] NB2 NB1 CSA_VREF pixel
xPix3921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[39] VREF PIX_IN[3921] NB2 NB1 CSA_VREF pixel
xPix3922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[39] VREF PIX_IN[3922] NB2 NB1 CSA_VREF pixel
xPix3923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[39] VREF PIX_IN[3923] NB2 NB1 CSA_VREF pixel
xPix3924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[39] VREF PIX_IN[3924] NB2 NB1 CSA_VREF pixel
xPix3925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[39] VREF PIX_IN[3925] NB2 NB1 CSA_VREF pixel
xPix3926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[39] VREF PIX_IN[3926] NB2 NB1 CSA_VREF pixel
xPix3927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[39] VREF PIX_IN[3927] NB2 NB1 CSA_VREF pixel
xPix3928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[39] VREF PIX_IN[3928] NB2 NB1 CSA_VREF pixel
xPix3929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[39] VREF PIX_IN[3929] NB2 NB1 CSA_VREF pixel
xPix3930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[39] VREF PIX_IN[3930] NB2 NB1 CSA_VREF pixel
xPix3931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[39] VREF PIX_IN[3931] NB2 NB1 CSA_VREF pixel
xPix3932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[39] VREF PIX_IN[3932] NB2 NB1 CSA_VREF pixel
xPix3933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[39] VREF PIX_IN[3933] NB2 NB1 CSA_VREF pixel
xPix3934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[39] VREF PIX_IN[3934] NB2 NB1 CSA_VREF pixel
xPix3935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[39] VREF PIX_IN[3935] NB2 NB1 CSA_VREF pixel
xPix3936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[39] VREF PIX_IN[3936] NB2 NB1 CSA_VREF pixel
xPix3937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[39] VREF PIX_IN[3937] NB2 NB1 CSA_VREF pixel
xPix3938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[39] VREF PIX_IN[3938] NB2 NB1 CSA_VREF pixel
xPix3939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[39] VREF PIX_IN[3939] NB2 NB1 CSA_VREF pixel
xPix3940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[39] VREF PIX_IN[3940] NB2 NB1 CSA_VREF pixel
xPix3941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[39] VREF PIX_IN[3941] NB2 NB1 CSA_VREF pixel
xPix3942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[39] VREF PIX_IN[3942] NB2 NB1 CSA_VREF pixel
xPix3943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[39] VREF PIX_IN[3943] NB2 NB1 CSA_VREF pixel
xPix3944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[39] VREF PIX_IN[3944] NB2 NB1 CSA_VREF pixel
xPix3945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[39] VREF PIX_IN[3945] NB2 NB1 CSA_VREF pixel
xPix3946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[39] VREF PIX_IN[3946] NB2 NB1 CSA_VREF pixel
xPix3947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[39] VREF PIX_IN[3947] NB2 NB1 CSA_VREF pixel
xPix3948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[39] VREF PIX_IN[3948] NB2 NB1 CSA_VREF pixel
xPix3949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[39] VREF PIX_IN[3949] NB2 NB1 CSA_VREF pixel
xPix3950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[39] VREF PIX_IN[3950] NB2 NB1 CSA_VREF pixel
xPix3951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[39] VREF PIX_IN[3951] NB2 NB1 CSA_VREF pixel
xPix3952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[39] VREF PIX_IN[3952] NB2 NB1 CSA_VREF pixel
xPix3953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[39] VREF PIX_IN[3953] NB2 NB1 CSA_VREF pixel
xPix3954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[39] VREF PIX_IN[3954] NB2 NB1 CSA_VREF pixel
xPix3955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[39] VREF PIX_IN[3955] NB2 NB1 CSA_VREF pixel
xPix3956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[39] VREF PIX_IN[3956] NB2 NB1 CSA_VREF pixel
xPix3957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[39] VREF PIX_IN[3957] NB2 NB1 CSA_VREF pixel
xPix3958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[39] VREF PIX_IN[3958] NB2 NB1 CSA_VREF pixel
xPix3959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[39] VREF PIX_IN[3959] NB2 NB1 CSA_VREF pixel
xPix3960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[39] VREF PIX_IN[3960] NB2 NB1 CSA_VREF pixel
xPix3961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[39] VREF PIX_IN[3961] NB2 NB1 CSA_VREF pixel
xPix3962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[39] VREF PIX_IN[3962] NB2 NB1 CSA_VREF pixel
xPix3963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[39] VREF PIX_IN[3963] NB2 NB1 CSA_VREF pixel
xPix3964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[39] VREF PIX_IN[3964] NB2 NB1 CSA_VREF pixel
xPix3965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[39] VREF PIX_IN[3965] NB2 NB1 CSA_VREF pixel
xPix3966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[39] VREF PIX_IN[3966] NB2 NB1 CSA_VREF pixel
xPix3967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[39] VREF PIX_IN[3967] NB2 NB1 CSA_VREF pixel
xPix3968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[39] VREF PIX_IN[3968] NB2 NB1 CSA_VREF pixel
xPix3969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[39] VREF PIX_IN[3969] NB2 NB1 CSA_VREF pixel
xPix3970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[39] VREF PIX_IN[3970] NB2 NB1 CSA_VREF pixel
xPix3971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[39] VREF PIX_IN[3971] NB2 NB1 CSA_VREF pixel
xPix3972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[39] VREF PIX_IN[3972] NB2 NB1 CSA_VREF pixel
xPix3973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[39] VREF PIX_IN[3973] NB2 NB1 CSA_VREF pixel
xPix3974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[39] VREF PIX_IN[3974] NB2 NB1 CSA_VREF pixel
xPix3975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[39] VREF PIX_IN[3975] NB2 NB1 CSA_VREF pixel
xPix3976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[39] VREF PIX_IN[3976] NB2 NB1 CSA_VREF pixel
xPix3977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[39] VREF PIX_IN[3977] NB2 NB1 CSA_VREF pixel
xPix3978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[39] VREF PIX_IN[3978] NB2 NB1 CSA_VREF pixel
xPix3979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[39] VREF PIX_IN[3979] NB2 NB1 CSA_VREF pixel
xPix3980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[39] VREF PIX_IN[3980] NB2 NB1 CSA_VREF pixel
xPix3981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[39] VREF PIX_IN[3981] NB2 NB1 CSA_VREF pixel
xPix3982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[39] VREF PIX_IN[3982] NB2 NB1 CSA_VREF pixel
xPix3983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[39] VREF PIX_IN[3983] NB2 NB1 CSA_VREF pixel
xPix3984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[39] VREF PIX_IN[3984] NB2 NB1 CSA_VREF pixel
xPix3985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[39] VREF PIX_IN[3985] NB2 NB1 CSA_VREF pixel
xPix3986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[39] VREF PIX_IN[3986] NB2 NB1 CSA_VREF pixel
xPix3987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[39] VREF PIX_IN[3987] NB2 NB1 CSA_VREF pixel
xPix3988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[39] VREF PIX_IN[3988] NB2 NB1 CSA_VREF pixel
xPix3989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[39] VREF PIX_IN[3989] NB2 NB1 CSA_VREF pixel
xPix3990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[39] VREF PIX_IN[3990] NB2 NB1 CSA_VREF pixel
xPix3991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[39] VREF PIX_IN[3991] NB2 NB1 CSA_VREF pixel
xPix3992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[39] VREF PIX_IN[3992] NB2 NB1 CSA_VREF pixel
xPix3993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[39] VREF PIX_IN[3993] NB2 NB1 CSA_VREF pixel
xPix3994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[39] VREF PIX_IN[3994] NB2 NB1 CSA_VREF pixel
xPix3995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[39] VREF PIX_IN[3995] NB2 NB1 CSA_VREF pixel
xPix3996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[39] VREF PIX_IN[3996] NB2 NB1 CSA_VREF pixel
xPix3997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[39] VREF PIX_IN[3997] NB2 NB1 CSA_VREF pixel
xPix3998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[39] VREF PIX_IN[3998] NB2 NB1 CSA_VREF pixel
xPix3999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[39] VREF PIX_IN[3999] NB2 NB1 CSA_VREF pixel
xPix4000 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[40] VREF PIX_IN[4000] NB2 NB1 CSA_VREF pixel
xPix4001 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[40] VREF PIX_IN[4001] NB2 NB1 CSA_VREF pixel
xPix4002 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[40] VREF PIX_IN[4002] NB2 NB1 CSA_VREF pixel
xPix4003 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[40] VREF PIX_IN[4003] NB2 NB1 CSA_VREF pixel
xPix4004 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[40] VREF PIX_IN[4004] NB2 NB1 CSA_VREF pixel
xPix4005 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[40] VREF PIX_IN[4005] NB2 NB1 CSA_VREF pixel
xPix4006 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[40] VREF PIX_IN[4006] NB2 NB1 CSA_VREF pixel
xPix4007 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[40] VREF PIX_IN[4007] NB2 NB1 CSA_VREF pixel
xPix4008 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[40] VREF PIX_IN[4008] NB2 NB1 CSA_VREF pixel
xPix4009 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[40] VREF PIX_IN[4009] NB2 NB1 CSA_VREF pixel
xPix4010 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[40] VREF PIX_IN[4010] NB2 NB1 CSA_VREF pixel
xPix4011 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[40] VREF PIX_IN[4011] NB2 NB1 CSA_VREF pixel
xPix4012 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[40] VREF PIX_IN[4012] NB2 NB1 CSA_VREF pixel
xPix4013 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[40] VREF PIX_IN[4013] NB2 NB1 CSA_VREF pixel
xPix4014 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[40] VREF PIX_IN[4014] NB2 NB1 CSA_VREF pixel
xPix4015 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[40] VREF PIX_IN[4015] NB2 NB1 CSA_VREF pixel
xPix4016 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[40] VREF PIX_IN[4016] NB2 NB1 CSA_VREF pixel
xPix4017 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[40] VREF PIX_IN[4017] NB2 NB1 CSA_VREF pixel
xPix4018 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[40] VREF PIX_IN[4018] NB2 NB1 CSA_VREF pixel
xPix4019 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[40] VREF PIX_IN[4019] NB2 NB1 CSA_VREF pixel
xPix4020 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[40] VREF PIX_IN[4020] NB2 NB1 CSA_VREF pixel
xPix4021 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[40] VREF PIX_IN[4021] NB2 NB1 CSA_VREF pixel
xPix4022 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[40] VREF PIX_IN[4022] NB2 NB1 CSA_VREF pixel
xPix4023 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[40] VREF PIX_IN[4023] NB2 NB1 CSA_VREF pixel
xPix4024 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[40] VREF PIX_IN[4024] NB2 NB1 CSA_VREF pixel
xPix4025 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[40] VREF PIX_IN[4025] NB2 NB1 CSA_VREF pixel
xPix4026 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[40] VREF PIX_IN[4026] NB2 NB1 CSA_VREF pixel
xPix4027 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[40] VREF PIX_IN[4027] NB2 NB1 CSA_VREF pixel
xPix4028 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[40] VREF PIX_IN[4028] NB2 NB1 CSA_VREF pixel
xPix4029 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[40] VREF PIX_IN[4029] NB2 NB1 CSA_VREF pixel
xPix4030 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[40] VREF PIX_IN[4030] NB2 NB1 CSA_VREF pixel
xPix4031 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[40] VREF PIX_IN[4031] NB2 NB1 CSA_VREF pixel
xPix4032 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[40] VREF PIX_IN[4032] NB2 NB1 CSA_VREF pixel
xPix4033 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[40] VREF PIX_IN[4033] NB2 NB1 CSA_VREF pixel
xPix4034 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[40] VREF PIX_IN[4034] NB2 NB1 CSA_VREF pixel
xPix4035 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[40] VREF PIX_IN[4035] NB2 NB1 CSA_VREF pixel
xPix4036 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[40] VREF PIX_IN[4036] NB2 NB1 CSA_VREF pixel
xPix4037 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[40] VREF PIX_IN[4037] NB2 NB1 CSA_VREF pixel
xPix4038 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[40] VREF PIX_IN[4038] NB2 NB1 CSA_VREF pixel
xPix4039 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[40] VREF PIX_IN[4039] NB2 NB1 CSA_VREF pixel
xPix4040 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[40] VREF PIX_IN[4040] NB2 NB1 CSA_VREF pixel
xPix4041 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[40] VREF PIX_IN[4041] NB2 NB1 CSA_VREF pixel
xPix4042 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[40] VREF PIX_IN[4042] NB2 NB1 CSA_VREF pixel
xPix4043 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[40] VREF PIX_IN[4043] NB2 NB1 CSA_VREF pixel
xPix4044 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[40] VREF PIX_IN[4044] NB2 NB1 CSA_VREF pixel
xPix4045 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[40] VREF PIX_IN[4045] NB2 NB1 CSA_VREF pixel
xPix4046 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[40] VREF PIX_IN[4046] NB2 NB1 CSA_VREF pixel
xPix4047 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[40] VREF PIX_IN[4047] NB2 NB1 CSA_VREF pixel
xPix4048 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[40] VREF PIX_IN[4048] NB2 NB1 CSA_VREF pixel
xPix4049 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[40] VREF PIX_IN[4049] NB2 NB1 CSA_VREF pixel
xPix4050 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[40] VREF PIX_IN[4050] NB2 NB1 CSA_VREF pixel
xPix4051 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[40] VREF PIX_IN[4051] NB2 NB1 CSA_VREF pixel
xPix4052 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[40] VREF PIX_IN[4052] NB2 NB1 CSA_VREF pixel
xPix4053 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[40] VREF PIX_IN[4053] NB2 NB1 CSA_VREF pixel
xPix4054 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[40] VREF PIX_IN[4054] NB2 NB1 CSA_VREF pixel
xPix4055 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[40] VREF PIX_IN[4055] NB2 NB1 CSA_VREF pixel
xPix4056 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[40] VREF PIX_IN[4056] NB2 NB1 CSA_VREF pixel
xPix4057 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[40] VREF PIX_IN[4057] NB2 NB1 CSA_VREF pixel
xPix4058 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[40] VREF PIX_IN[4058] NB2 NB1 CSA_VREF pixel
xPix4059 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[40] VREF PIX_IN[4059] NB2 NB1 CSA_VREF pixel
xPix4060 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[40] VREF PIX_IN[4060] NB2 NB1 CSA_VREF pixel
xPix4061 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[40] VREF PIX_IN[4061] NB2 NB1 CSA_VREF pixel
xPix4062 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[40] VREF PIX_IN[4062] NB2 NB1 CSA_VREF pixel
xPix4063 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[40] VREF PIX_IN[4063] NB2 NB1 CSA_VREF pixel
xPix4064 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[40] VREF PIX_IN[4064] NB2 NB1 CSA_VREF pixel
xPix4065 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[40] VREF PIX_IN[4065] NB2 NB1 CSA_VREF pixel
xPix4066 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[40] VREF PIX_IN[4066] NB2 NB1 CSA_VREF pixel
xPix4067 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[40] VREF PIX_IN[4067] NB2 NB1 CSA_VREF pixel
xPix4068 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[40] VREF PIX_IN[4068] NB2 NB1 CSA_VREF pixel
xPix4069 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[40] VREF PIX_IN[4069] NB2 NB1 CSA_VREF pixel
xPix4070 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[40] VREF PIX_IN[4070] NB2 NB1 CSA_VREF pixel
xPix4071 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[40] VREF PIX_IN[4071] NB2 NB1 CSA_VREF pixel
xPix4072 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[40] VREF PIX_IN[4072] NB2 NB1 CSA_VREF pixel
xPix4073 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[40] VREF PIX_IN[4073] NB2 NB1 CSA_VREF pixel
xPix4074 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[40] VREF PIX_IN[4074] NB2 NB1 CSA_VREF pixel
xPix4075 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[40] VREF PIX_IN[4075] NB2 NB1 CSA_VREF pixel
xPix4076 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[40] VREF PIX_IN[4076] NB2 NB1 CSA_VREF pixel
xPix4077 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[40] VREF PIX_IN[4077] NB2 NB1 CSA_VREF pixel
xPix4078 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[40] VREF PIX_IN[4078] NB2 NB1 CSA_VREF pixel
xPix4079 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[40] VREF PIX_IN[4079] NB2 NB1 CSA_VREF pixel
xPix4080 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[40] VREF PIX_IN[4080] NB2 NB1 CSA_VREF pixel
xPix4081 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[40] VREF PIX_IN[4081] NB2 NB1 CSA_VREF pixel
xPix4082 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[40] VREF PIX_IN[4082] NB2 NB1 CSA_VREF pixel
xPix4083 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[40] VREF PIX_IN[4083] NB2 NB1 CSA_VREF pixel
xPix4084 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[40] VREF PIX_IN[4084] NB2 NB1 CSA_VREF pixel
xPix4085 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[40] VREF PIX_IN[4085] NB2 NB1 CSA_VREF pixel
xPix4086 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[40] VREF PIX_IN[4086] NB2 NB1 CSA_VREF pixel
xPix4087 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[40] VREF PIX_IN[4087] NB2 NB1 CSA_VREF pixel
xPix4088 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[40] VREF PIX_IN[4088] NB2 NB1 CSA_VREF pixel
xPix4089 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[40] VREF PIX_IN[4089] NB2 NB1 CSA_VREF pixel
xPix4090 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[40] VREF PIX_IN[4090] NB2 NB1 CSA_VREF pixel
xPix4091 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[40] VREF PIX_IN[4091] NB2 NB1 CSA_VREF pixel
xPix4092 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[40] VREF PIX_IN[4092] NB2 NB1 CSA_VREF pixel
xPix4093 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[40] VREF PIX_IN[4093] NB2 NB1 CSA_VREF pixel
xPix4094 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[40] VREF PIX_IN[4094] NB2 NB1 CSA_VREF pixel
xPix4095 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[40] VREF PIX_IN[4095] NB2 NB1 CSA_VREF pixel
xPix4096 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[40] VREF PIX_IN[4096] NB2 NB1 CSA_VREF pixel
xPix4097 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[40] VREF PIX_IN[4097] NB2 NB1 CSA_VREF pixel
xPix4098 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[40] VREF PIX_IN[4098] NB2 NB1 CSA_VREF pixel
xPix4099 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[40] VREF PIX_IN[4099] NB2 NB1 CSA_VREF pixel
xPix4100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[41] VREF PIX_IN[4100] NB2 NB1 CSA_VREF pixel
xPix4101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[41] VREF PIX_IN[4101] NB2 NB1 CSA_VREF pixel
xPix4102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[41] VREF PIX_IN[4102] NB2 NB1 CSA_VREF pixel
xPix4103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[41] VREF PIX_IN[4103] NB2 NB1 CSA_VREF pixel
xPix4104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[41] VREF PIX_IN[4104] NB2 NB1 CSA_VREF pixel
xPix4105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[41] VREF PIX_IN[4105] NB2 NB1 CSA_VREF pixel
xPix4106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[41] VREF PIX_IN[4106] NB2 NB1 CSA_VREF pixel
xPix4107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[41] VREF PIX_IN[4107] NB2 NB1 CSA_VREF pixel
xPix4108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[41] VREF PIX_IN[4108] NB2 NB1 CSA_VREF pixel
xPix4109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[41] VREF PIX_IN[4109] NB2 NB1 CSA_VREF pixel
xPix4110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[41] VREF PIX_IN[4110] NB2 NB1 CSA_VREF pixel
xPix4111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[41] VREF PIX_IN[4111] NB2 NB1 CSA_VREF pixel
xPix4112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[41] VREF PIX_IN[4112] NB2 NB1 CSA_VREF pixel
xPix4113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[41] VREF PIX_IN[4113] NB2 NB1 CSA_VREF pixel
xPix4114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[41] VREF PIX_IN[4114] NB2 NB1 CSA_VREF pixel
xPix4115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[41] VREF PIX_IN[4115] NB2 NB1 CSA_VREF pixel
xPix4116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[41] VREF PIX_IN[4116] NB2 NB1 CSA_VREF pixel
xPix4117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[41] VREF PIX_IN[4117] NB2 NB1 CSA_VREF pixel
xPix4118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[41] VREF PIX_IN[4118] NB2 NB1 CSA_VREF pixel
xPix4119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[41] VREF PIX_IN[4119] NB2 NB1 CSA_VREF pixel
xPix4120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[41] VREF PIX_IN[4120] NB2 NB1 CSA_VREF pixel
xPix4121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[41] VREF PIX_IN[4121] NB2 NB1 CSA_VREF pixel
xPix4122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[41] VREF PIX_IN[4122] NB2 NB1 CSA_VREF pixel
xPix4123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[41] VREF PIX_IN[4123] NB2 NB1 CSA_VREF pixel
xPix4124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[41] VREF PIX_IN[4124] NB2 NB1 CSA_VREF pixel
xPix4125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[41] VREF PIX_IN[4125] NB2 NB1 CSA_VREF pixel
xPix4126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[41] VREF PIX_IN[4126] NB2 NB1 CSA_VREF pixel
xPix4127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[41] VREF PIX_IN[4127] NB2 NB1 CSA_VREF pixel
xPix4128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[41] VREF PIX_IN[4128] NB2 NB1 CSA_VREF pixel
xPix4129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[41] VREF PIX_IN[4129] NB2 NB1 CSA_VREF pixel
xPix4130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[41] VREF PIX_IN[4130] NB2 NB1 CSA_VREF pixel
xPix4131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[41] VREF PIX_IN[4131] NB2 NB1 CSA_VREF pixel
xPix4132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[41] VREF PIX_IN[4132] NB2 NB1 CSA_VREF pixel
xPix4133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[41] VREF PIX_IN[4133] NB2 NB1 CSA_VREF pixel
xPix4134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[41] VREF PIX_IN[4134] NB2 NB1 CSA_VREF pixel
xPix4135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[41] VREF PIX_IN[4135] NB2 NB1 CSA_VREF pixel
xPix4136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[41] VREF PIX_IN[4136] NB2 NB1 CSA_VREF pixel
xPix4137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[41] VREF PIX_IN[4137] NB2 NB1 CSA_VREF pixel
xPix4138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[41] VREF PIX_IN[4138] NB2 NB1 CSA_VREF pixel
xPix4139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[41] VREF PIX_IN[4139] NB2 NB1 CSA_VREF pixel
xPix4140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[41] VREF PIX_IN[4140] NB2 NB1 CSA_VREF pixel
xPix4141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[41] VREF PIX_IN[4141] NB2 NB1 CSA_VREF pixel
xPix4142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[41] VREF PIX_IN[4142] NB2 NB1 CSA_VREF pixel
xPix4143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[41] VREF PIX_IN[4143] NB2 NB1 CSA_VREF pixel
xPix4144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[41] VREF PIX_IN[4144] NB2 NB1 CSA_VREF pixel
xPix4145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[41] VREF PIX_IN[4145] NB2 NB1 CSA_VREF pixel
xPix4146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[41] VREF PIX_IN[4146] NB2 NB1 CSA_VREF pixel
xPix4147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[41] VREF PIX_IN[4147] NB2 NB1 CSA_VREF pixel
xPix4148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[41] VREF PIX_IN[4148] NB2 NB1 CSA_VREF pixel
xPix4149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[41] VREF PIX_IN[4149] NB2 NB1 CSA_VREF pixel
xPix4150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[41] VREF PIX_IN[4150] NB2 NB1 CSA_VREF pixel
xPix4151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[41] VREF PIX_IN[4151] NB2 NB1 CSA_VREF pixel
xPix4152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[41] VREF PIX_IN[4152] NB2 NB1 CSA_VREF pixel
xPix4153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[41] VREF PIX_IN[4153] NB2 NB1 CSA_VREF pixel
xPix4154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[41] VREF PIX_IN[4154] NB2 NB1 CSA_VREF pixel
xPix4155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[41] VREF PIX_IN[4155] NB2 NB1 CSA_VREF pixel
xPix4156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[41] VREF PIX_IN[4156] NB2 NB1 CSA_VREF pixel
xPix4157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[41] VREF PIX_IN[4157] NB2 NB1 CSA_VREF pixel
xPix4158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[41] VREF PIX_IN[4158] NB2 NB1 CSA_VREF pixel
xPix4159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[41] VREF PIX_IN[4159] NB2 NB1 CSA_VREF pixel
xPix4160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[41] VREF PIX_IN[4160] NB2 NB1 CSA_VREF pixel
xPix4161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[41] VREF PIX_IN[4161] NB2 NB1 CSA_VREF pixel
xPix4162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[41] VREF PIX_IN[4162] NB2 NB1 CSA_VREF pixel
xPix4163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[41] VREF PIX_IN[4163] NB2 NB1 CSA_VREF pixel
xPix4164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[41] VREF PIX_IN[4164] NB2 NB1 CSA_VREF pixel
xPix4165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[41] VREF PIX_IN[4165] NB2 NB1 CSA_VREF pixel
xPix4166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[41] VREF PIX_IN[4166] NB2 NB1 CSA_VREF pixel
xPix4167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[41] VREF PIX_IN[4167] NB2 NB1 CSA_VREF pixel
xPix4168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[41] VREF PIX_IN[4168] NB2 NB1 CSA_VREF pixel
xPix4169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[41] VREF PIX_IN[4169] NB2 NB1 CSA_VREF pixel
xPix4170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[41] VREF PIX_IN[4170] NB2 NB1 CSA_VREF pixel
xPix4171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[41] VREF PIX_IN[4171] NB2 NB1 CSA_VREF pixel
xPix4172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[41] VREF PIX_IN[4172] NB2 NB1 CSA_VREF pixel
xPix4173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[41] VREF PIX_IN[4173] NB2 NB1 CSA_VREF pixel
xPix4174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[41] VREF PIX_IN[4174] NB2 NB1 CSA_VREF pixel
xPix4175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[41] VREF PIX_IN[4175] NB2 NB1 CSA_VREF pixel
xPix4176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[41] VREF PIX_IN[4176] NB2 NB1 CSA_VREF pixel
xPix4177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[41] VREF PIX_IN[4177] NB2 NB1 CSA_VREF pixel
xPix4178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[41] VREF PIX_IN[4178] NB2 NB1 CSA_VREF pixel
xPix4179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[41] VREF PIX_IN[4179] NB2 NB1 CSA_VREF pixel
xPix4180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[41] VREF PIX_IN[4180] NB2 NB1 CSA_VREF pixel
xPix4181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[41] VREF PIX_IN[4181] NB2 NB1 CSA_VREF pixel
xPix4182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[41] VREF PIX_IN[4182] NB2 NB1 CSA_VREF pixel
xPix4183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[41] VREF PIX_IN[4183] NB2 NB1 CSA_VREF pixel
xPix4184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[41] VREF PIX_IN[4184] NB2 NB1 CSA_VREF pixel
xPix4185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[41] VREF PIX_IN[4185] NB2 NB1 CSA_VREF pixel
xPix4186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[41] VREF PIX_IN[4186] NB2 NB1 CSA_VREF pixel
xPix4187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[41] VREF PIX_IN[4187] NB2 NB1 CSA_VREF pixel
xPix4188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[41] VREF PIX_IN[4188] NB2 NB1 CSA_VREF pixel
xPix4189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[41] VREF PIX_IN[4189] NB2 NB1 CSA_VREF pixel
xPix4190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[41] VREF PIX_IN[4190] NB2 NB1 CSA_VREF pixel
xPix4191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[41] VREF PIX_IN[4191] NB2 NB1 CSA_VREF pixel
xPix4192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[41] VREF PIX_IN[4192] NB2 NB1 CSA_VREF pixel
xPix4193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[41] VREF PIX_IN[4193] NB2 NB1 CSA_VREF pixel
xPix4194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[41] VREF PIX_IN[4194] NB2 NB1 CSA_VREF pixel
xPix4195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[41] VREF PIX_IN[4195] NB2 NB1 CSA_VREF pixel
xPix4196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[41] VREF PIX_IN[4196] NB2 NB1 CSA_VREF pixel
xPix4197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[41] VREF PIX_IN[4197] NB2 NB1 CSA_VREF pixel
xPix4198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[41] VREF PIX_IN[4198] NB2 NB1 CSA_VREF pixel
xPix4199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[41] VREF PIX_IN[4199] NB2 NB1 CSA_VREF pixel
xPix4200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[42] VREF PIX_IN[4200] NB2 NB1 CSA_VREF pixel
xPix4201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[42] VREF PIX_IN[4201] NB2 NB1 CSA_VREF pixel
xPix4202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[42] VREF PIX_IN[4202] NB2 NB1 CSA_VREF pixel
xPix4203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[42] VREF PIX_IN[4203] NB2 NB1 CSA_VREF pixel
xPix4204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[42] VREF PIX_IN[4204] NB2 NB1 CSA_VREF pixel
xPix4205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[42] VREF PIX_IN[4205] NB2 NB1 CSA_VREF pixel
xPix4206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[42] VREF PIX_IN[4206] NB2 NB1 CSA_VREF pixel
xPix4207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[42] VREF PIX_IN[4207] NB2 NB1 CSA_VREF pixel
xPix4208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[42] VREF PIX_IN[4208] NB2 NB1 CSA_VREF pixel
xPix4209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[42] VREF PIX_IN[4209] NB2 NB1 CSA_VREF pixel
xPix4210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[42] VREF PIX_IN[4210] NB2 NB1 CSA_VREF pixel
xPix4211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[42] VREF PIX_IN[4211] NB2 NB1 CSA_VREF pixel
xPix4212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[42] VREF PIX_IN[4212] NB2 NB1 CSA_VREF pixel
xPix4213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[42] VREF PIX_IN[4213] NB2 NB1 CSA_VREF pixel
xPix4214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[42] VREF PIX_IN[4214] NB2 NB1 CSA_VREF pixel
xPix4215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[42] VREF PIX_IN[4215] NB2 NB1 CSA_VREF pixel
xPix4216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[42] VREF PIX_IN[4216] NB2 NB1 CSA_VREF pixel
xPix4217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[42] VREF PIX_IN[4217] NB2 NB1 CSA_VREF pixel
xPix4218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[42] VREF PIX_IN[4218] NB2 NB1 CSA_VREF pixel
xPix4219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[42] VREF PIX_IN[4219] NB2 NB1 CSA_VREF pixel
xPix4220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[42] VREF PIX_IN[4220] NB2 NB1 CSA_VREF pixel
xPix4221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[42] VREF PIX_IN[4221] NB2 NB1 CSA_VREF pixel
xPix4222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[42] VREF PIX_IN[4222] NB2 NB1 CSA_VREF pixel
xPix4223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[42] VREF PIX_IN[4223] NB2 NB1 CSA_VREF pixel
xPix4224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[42] VREF PIX_IN[4224] NB2 NB1 CSA_VREF pixel
xPix4225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[42] VREF PIX_IN[4225] NB2 NB1 CSA_VREF pixel
xPix4226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[42] VREF PIX_IN[4226] NB2 NB1 CSA_VREF pixel
xPix4227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[42] VREF PIX_IN[4227] NB2 NB1 CSA_VREF pixel
xPix4228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[42] VREF PIX_IN[4228] NB2 NB1 CSA_VREF pixel
xPix4229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[42] VREF PIX_IN[4229] NB2 NB1 CSA_VREF pixel
xPix4230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[42] VREF PIX_IN[4230] NB2 NB1 CSA_VREF pixel
xPix4231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[42] VREF PIX_IN[4231] NB2 NB1 CSA_VREF pixel
xPix4232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[42] VREF PIX_IN[4232] NB2 NB1 CSA_VREF pixel
xPix4233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[42] VREF PIX_IN[4233] NB2 NB1 CSA_VREF pixel
xPix4234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[42] VREF PIX_IN[4234] NB2 NB1 CSA_VREF pixel
xPix4235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[42] VREF PIX_IN[4235] NB2 NB1 CSA_VREF pixel
xPix4236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[42] VREF PIX_IN[4236] NB2 NB1 CSA_VREF pixel
xPix4237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[42] VREF PIX_IN[4237] NB2 NB1 CSA_VREF pixel
xPix4238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[42] VREF PIX_IN[4238] NB2 NB1 CSA_VREF pixel
xPix4239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[42] VREF PIX_IN[4239] NB2 NB1 CSA_VREF pixel
xPix4240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[42] VREF PIX_IN[4240] NB2 NB1 CSA_VREF pixel
xPix4241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[42] VREF PIX_IN[4241] NB2 NB1 CSA_VREF pixel
xPix4242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[42] VREF PIX_IN[4242] NB2 NB1 CSA_VREF pixel
xPix4243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[42] VREF PIX_IN[4243] NB2 NB1 CSA_VREF pixel
xPix4244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[42] VREF PIX_IN[4244] NB2 NB1 CSA_VREF pixel
xPix4245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[42] VREF PIX_IN[4245] NB2 NB1 CSA_VREF pixel
xPix4246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[42] VREF PIX_IN[4246] NB2 NB1 CSA_VREF pixel
xPix4247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[42] VREF PIX_IN[4247] NB2 NB1 CSA_VREF pixel
xPix4248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[42] VREF PIX_IN[4248] NB2 NB1 CSA_VREF pixel
xPix4249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[42] VREF PIX_IN[4249] NB2 NB1 CSA_VREF pixel
xPix4250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[42] VREF PIX_IN[4250] NB2 NB1 CSA_VREF pixel
xPix4251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[42] VREF PIX_IN[4251] NB2 NB1 CSA_VREF pixel
xPix4252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[42] VREF PIX_IN[4252] NB2 NB1 CSA_VREF pixel
xPix4253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[42] VREF PIX_IN[4253] NB2 NB1 CSA_VREF pixel
xPix4254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[42] VREF PIX_IN[4254] NB2 NB1 CSA_VREF pixel
xPix4255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[42] VREF PIX_IN[4255] NB2 NB1 CSA_VREF pixel
xPix4256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[42] VREF PIX_IN[4256] NB2 NB1 CSA_VREF pixel
xPix4257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[42] VREF PIX_IN[4257] NB2 NB1 CSA_VREF pixel
xPix4258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[42] VREF PIX_IN[4258] NB2 NB1 CSA_VREF pixel
xPix4259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[42] VREF PIX_IN[4259] NB2 NB1 CSA_VREF pixel
xPix4260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[42] VREF PIX_IN[4260] NB2 NB1 CSA_VREF pixel
xPix4261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[42] VREF PIX_IN[4261] NB2 NB1 CSA_VREF pixel
xPix4262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[42] VREF PIX_IN[4262] NB2 NB1 CSA_VREF pixel
xPix4263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[42] VREF PIX_IN[4263] NB2 NB1 CSA_VREF pixel
xPix4264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[42] VREF PIX_IN[4264] NB2 NB1 CSA_VREF pixel
xPix4265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[42] VREF PIX_IN[4265] NB2 NB1 CSA_VREF pixel
xPix4266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[42] VREF PIX_IN[4266] NB2 NB1 CSA_VREF pixel
xPix4267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[42] VREF PIX_IN[4267] NB2 NB1 CSA_VREF pixel
xPix4268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[42] VREF PIX_IN[4268] NB2 NB1 CSA_VREF pixel
xPix4269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[42] VREF PIX_IN[4269] NB2 NB1 CSA_VREF pixel
xPix4270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[42] VREF PIX_IN[4270] NB2 NB1 CSA_VREF pixel
xPix4271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[42] VREF PIX_IN[4271] NB2 NB1 CSA_VREF pixel
xPix4272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[42] VREF PIX_IN[4272] NB2 NB1 CSA_VREF pixel
xPix4273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[42] VREF PIX_IN[4273] NB2 NB1 CSA_VREF pixel
xPix4274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[42] VREF PIX_IN[4274] NB2 NB1 CSA_VREF pixel
xPix4275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[42] VREF PIX_IN[4275] NB2 NB1 CSA_VREF pixel
xPix4276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[42] VREF PIX_IN[4276] NB2 NB1 CSA_VREF pixel
xPix4277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[42] VREF PIX_IN[4277] NB2 NB1 CSA_VREF pixel
xPix4278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[42] VREF PIX_IN[4278] NB2 NB1 CSA_VREF pixel
xPix4279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[42] VREF PIX_IN[4279] NB2 NB1 CSA_VREF pixel
xPix4280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[42] VREF PIX_IN[4280] NB2 NB1 CSA_VREF pixel
xPix4281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[42] VREF PIX_IN[4281] NB2 NB1 CSA_VREF pixel
xPix4282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[42] VREF PIX_IN[4282] NB2 NB1 CSA_VREF pixel
xPix4283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[42] VREF PIX_IN[4283] NB2 NB1 CSA_VREF pixel
xPix4284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[42] VREF PIX_IN[4284] NB2 NB1 CSA_VREF pixel
xPix4285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[42] VREF PIX_IN[4285] NB2 NB1 CSA_VREF pixel
xPix4286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[42] VREF PIX_IN[4286] NB2 NB1 CSA_VREF pixel
xPix4287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[42] VREF PIX_IN[4287] NB2 NB1 CSA_VREF pixel
xPix4288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[42] VREF PIX_IN[4288] NB2 NB1 CSA_VREF pixel
xPix4289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[42] VREF PIX_IN[4289] NB2 NB1 CSA_VREF pixel
xPix4290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[42] VREF PIX_IN[4290] NB2 NB1 CSA_VREF pixel
xPix4291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[42] VREF PIX_IN[4291] NB2 NB1 CSA_VREF pixel
xPix4292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[42] VREF PIX_IN[4292] NB2 NB1 CSA_VREF pixel
xPix4293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[42] VREF PIX_IN[4293] NB2 NB1 CSA_VREF pixel
xPix4294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[42] VREF PIX_IN[4294] NB2 NB1 CSA_VREF pixel
xPix4295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[42] VREF PIX_IN[4295] NB2 NB1 CSA_VREF pixel
xPix4296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[42] VREF PIX_IN[4296] NB2 NB1 CSA_VREF pixel
xPix4297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[42] VREF PIX_IN[4297] NB2 NB1 CSA_VREF pixel
xPix4298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[42] VREF PIX_IN[4298] NB2 NB1 CSA_VREF pixel
xPix4299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[42] VREF PIX_IN[4299] NB2 NB1 CSA_VREF pixel
xPix4300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[43] VREF PIX_IN[4300] NB2 NB1 CSA_VREF pixel
xPix4301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[43] VREF PIX_IN[4301] NB2 NB1 CSA_VREF pixel
xPix4302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[43] VREF PIX_IN[4302] NB2 NB1 CSA_VREF pixel
xPix4303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[43] VREF PIX_IN[4303] NB2 NB1 CSA_VREF pixel
xPix4304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[43] VREF PIX_IN[4304] NB2 NB1 CSA_VREF pixel
xPix4305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[43] VREF PIX_IN[4305] NB2 NB1 CSA_VREF pixel
xPix4306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[43] VREF PIX_IN[4306] NB2 NB1 CSA_VREF pixel
xPix4307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[43] VREF PIX_IN[4307] NB2 NB1 CSA_VREF pixel
xPix4308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[43] VREF PIX_IN[4308] NB2 NB1 CSA_VREF pixel
xPix4309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[43] VREF PIX_IN[4309] NB2 NB1 CSA_VREF pixel
xPix4310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[43] VREF PIX_IN[4310] NB2 NB1 CSA_VREF pixel
xPix4311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[43] VREF PIX_IN[4311] NB2 NB1 CSA_VREF pixel
xPix4312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[43] VREF PIX_IN[4312] NB2 NB1 CSA_VREF pixel
xPix4313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[43] VREF PIX_IN[4313] NB2 NB1 CSA_VREF pixel
xPix4314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[43] VREF PIX_IN[4314] NB2 NB1 CSA_VREF pixel
xPix4315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[43] VREF PIX_IN[4315] NB2 NB1 CSA_VREF pixel
xPix4316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[43] VREF PIX_IN[4316] NB2 NB1 CSA_VREF pixel
xPix4317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[43] VREF PIX_IN[4317] NB2 NB1 CSA_VREF pixel
xPix4318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[43] VREF PIX_IN[4318] NB2 NB1 CSA_VREF pixel
xPix4319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[43] VREF PIX_IN[4319] NB2 NB1 CSA_VREF pixel
xPix4320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[43] VREF PIX_IN[4320] NB2 NB1 CSA_VREF pixel
xPix4321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[43] VREF PIX_IN[4321] NB2 NB1 CSA_VREF pixel
xPix4322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[43] VREF PIX_IN[4322] NB2 NB1 CSA_VREF pixel
xPix4323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[43] VREF PIX_IN[4323] NB2 NB1 CSA_VREF pixel
xPix4324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[43] VREF PIX_IN[4324] NB2 NB1 CSA_VREF pixel
xPix4325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[43] VREF PIX_IN[4325] NB2 NB1 CSA_VREF pixel
xPix4326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[43] VREF PIX_IN[4326] NB2 NB1 CSA_VREF pixel
xPix4327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[43] VREF PIX_IN[4327] NB2 NB1 CSA_VREF pixel
xPix4328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[43] VREF PIX_IN[4328] NB2 NB1 CSA_VREF pixel
xPix4329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[43] VREF PIX_IN[4329] NB2 NB1 CSA_VREF pixel
xPix4330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[43] VREF PIX_IN[4330] NB2 NB1 CSA_VREF pixel
xPix4331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[43] VREF PIX_IN[4331] NB2 NB1 CSA_VREF pixel
xPix4332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[43] VREF PIX_IN[4332] NB2 NB1 CSA_VREF pixel
xPix4333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[43] VREF PIX_IN[4333] NB2 NB1 CSA_VREF pixel
xPix4334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[43] VREF PIX_IN[4334] NB2 NB1 CSA_VREF pixel
xPix4335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[43] VREF PIX_IN[4335] NB2 NB1 CSA_VREF pixel
xPix4336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[43] VREF PIX_IN[4336] NB2 NB1 CSA_VREF pixel
xPix4337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[43] VREF PIX_IN[4337] NB2 NB1 CSA_VREF pixel
xPix4338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[43] VREF PIX_IN[4338] NB2 NB1 CSA_VREF pixel
xPix4339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[43] VREF PIX_IN[4339] NB2 NB1 CSA_VREF pixel
xPix4340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[43] VREF PIX_IN[4340] NB2 NB1 CSA_VREF pixel
xPix4341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[43] VREF PIX_IN[4341] NB2 NB1 CSA_VREF pixel
xPix4342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[43] VREF PIX_IN[4342] NB2 NB1 CSA_VREF pixel
xPix4343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[43] VREF PIX_IN[4343] NB2 NB1 CSA_VREF pixel
xPix4344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[43] VREF PIX_IN[4344] NB2 NB1 CSA_VREF pixel
xPix4345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[43] VREF PIX_IN[4345] NB2 NB1 CSA_VREF pixel
xPix4346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[43] VREF PIX_IN[4346] NB2 NB1 CSA_VREF pixel
xPix4347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[43] VREF PIX_IN[4347] NB2 NB1 CSA_VREF pixel
xPix4348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[43] VREF PIX_IN[4348] NB2 NB1 CSA_VREF pixel
xPix4349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[43] VREF PIX_IN[4349] NB2 NB1 CSA_VREF pixel
xPix4350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[43] VREF PIX_IN[4350] NB2 NB1 CSA_VREF pixel
xPix4351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[43] VREF PIX_IN[4351] NB2 NB1 CSA_VREF pixel
xPix4352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[43] VREF PIX_IN[4352] NB2 NB1 CSA_VREF pixel
xPix4353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[43] VREF PIX_IN[4353] NB2 NB1 CSA_VREF pixel
xPix4354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[43] VREF PIX_IN[4354] NB2 NB1 CSA_VREF pixel
xPix4355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[43] VREF PIX_IN[4355] NB2 NB1 CSA_VREF pixel
xPix4356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[43] VREF PIX_IN[4356] NB2 NB1 CSA_VREF pixel
xPix4357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[43] VREF PIX_IN[4357] NB2 NB1 CSA_VREF pixel
xPix4358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[43] VREF PIX_IN[4358] NB2 NB1 CSA_VREF pixel
xPix4359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[43] VREF PIX_IN[4359] NB2 NB1 CSA_VREF pixel
xPix4360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[43] VREF PIX_IN[4360] NB2 NB1 CSA_VREF pixel
xPix4361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[43] VREF PIX_IN[4361] NB2 NB1 CSA_VREF pixel
xPix4362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[43] VREF PIX_IN[4362] NB2 NB1 CSA_VREF pixel
xPix4363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[43] VREF PIX_IN[4363] NB2 NB1 CSA_VREF pixel
xPix4364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[43] VREF PIX_IN[4364] NB2 NB1 CSA_VREF pixel
xPix4365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[43] VREF PIX_IN[4365] NB2 NB1 CSA_VREF pixel
xPix4366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[43] VREF PIX_IN[4366] NB2 NB1 CSA_VREF pixel
xPix4367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[43] VREF PIX_IN[4367] NB2 NB1 CSA_VREF pixel
xPix4368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[43] VREF PIX_IN[4368] NB2 NB1 CSA_VREF pixel
xPix4369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[43] VREF PIX_IN[4369] NB2 NB1 CSA_VREF pixel
xPix4370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[43] VREF PIX_IN[4370] NB2 NB1 CSA_VREF pixel
xPix4371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[43] VREF PIX_IN[4371] NB2 NB1 CSA_VREF pixel
xPix4372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[43] VREF PIX_IN[4372] NB2 NB1 CSA_VREF pixel
xPix4373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[43] VREF PIX_IN[4373] NB2 NB1 CSA_VREF pixel
xPix4374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[43] VREF PIX_IN[4374] NB2 NB1 CSA_VREF pixel
xPix4375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[43] VREF PIX_IN[4375] NB2 NB1 CSA_VREF pixel
xPix4376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[43] VREF PIX_IN[4376] NB2 NB1 CSA_VREF pixel
xPix4377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[43] VREF PIX_IN[4377] NB2 NB1 CSA_VREF pixel
xPix4378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[43] VREF PIX_IN[4378] NB2 NB1 CSA_VREF pixel
xPix4379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[43] VREF PIX_IN[4379] NB2 NB1 CSA_VREF pixel
xPix4380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[43] VREF PIX_IN[4380] NB2 NB1 CSA_VREF pixel
xPix4381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[43] VREF PIX_IN[4381] NB2 NB1 CSA_VREF pixel
xPix4382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[43] VREF PIX_IN[4382] NB2 NB1 CSA_VREF pixel
xPix4383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[43] VREF PIX_IN[4383] NB2 NB1 CSA_VREF pixel
xPix4384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[43] VREF PIX_IN[4384] NB2 NB1 CSA_VREF pixel
xPix4385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[43] VREF PIX_IN[4385] NB2 NB1 CSA_VREF pixel
xPix4386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[43] VREF PIX_IN[4386] NB2 NB1 CSA_VREF pixel
xPix4387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[43] VREF PIX_IN[4387] NB2 NB1 CSA_VREF pixel
xPix4388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[43] VREF PIX_IN[4388] NB2 NB1 CSA_VREF pixel
xPix4389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[43] VREF PIX_IN[4389] NB2 NB1 CSA_VREF pixel
xPix4390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[43] VREF PIX_IN[4390] NB2 NB1 CSA_VREF pixel
xPix4391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[43] VREF PIX_IN[4391] NB2 NB1 CSA_VREF pixel
xPix4392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[43] VREF PIX_IN[4392] NB2 NB1 CSA_VREF pixel
xPix4393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[43] VREF PIX_IN[4393] NB2 NB1 CSA_VREF pixel
xPix4394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[43] VREF PIX_IN[4394] NB2 NB1 CSA_VREF pixel
xPix4395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[43] VREF PIX_IN[4395] NB2 NB1 CSA_VREF pixel
xPix4396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[43] VREF PIX_IN[4396] NB2 NB1 CSA_VREF pixel
xPix4397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[43] VREF PIX_IN[4397] NB2 NB1 CSA_VREF pixel
xPix4398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[43] VREF PIX_IN[4398] NB2 NB1 CSA_VREF pixel
xPix4399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[43] VREF PIX_IN[4399] NB2 NB1 CSA_VREF pixel
xPix4400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[44] VREF PIX_IN[4400] NB2 NB1 CSA_VREF pixel
xPix4401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[44] VREF PIX_IN[4401] NB2 NB1 CSA_VREF pixel
xPix4402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[44] VREF PIX_IN[4402] NB2 NB1 CSA_VREF pixel
xPix4403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[44] VREF PIX_IN[4403] NB2 NB1 CSA_VREF pixel
xPix4404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[44] VREF PIX_IN[4404] NB2 NB1 CSA_VREF pixel
xPix4405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[44] VREF PIX_IN[4405] NB2 NB1 CSA_VREF pixel
xPix4406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[44] VREF PIX_IN[4406] NB2 NB1 CSA_VREF pixel
xPix4407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[44] VREF PIX_IN[4407] NB2 NB1 CSA_VREF pixel
xPix4408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[44] VREF PIX_IN[4408] NB2 NB1 CSA_VREF pixel
xPix4409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[44] VREF PIX_IN[4409] NB2 NB1 CSA_VREF pixel
xPix4410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[44] VREF PIX_IN[4410] NB2 NB1 CSA_VREF pixel
xPix4411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[44] VREF PIX_IN[4411] NB2 NB1 CSA_VREF pixel
xPix4412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[44] VREF PIX_IN[4412] NB2 NB1 CSA_VREF pixel
xPix4413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[44] VREF PIX_IN[4413] NB2 NB1 CSA_VREF pixel
xPix4414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[44] VREF PIX_IN[4414] NB2 NB1 CSA_VREF pixel
xPix4415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[44] VREF PIX_IN[4415] NB2 NB1 CSA_VREF pixel
xPix4416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[44] VREF PIX_IN[4416] NB2 NB1 CSA_VREF pixel
xPix4417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[44] VREF PIX_IN[4417] NB2 NB1 CSA_VREF pixel
xPix4418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[44] VREF PIX_IN[4418] NB2 NB1 CSA_VREF pixel
xPix4419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[44] VREF PIX_IN[4419] NB2 NB1 CSA_VREF pixel
xPix4420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[44] VREF PIX_IN[4420] NB2 NB1 CSA_VREF pixel
xPix4421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[44] VREF PIX_IN[4421] NB2 NB1 CSA_VREF pixel
xPix4422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[44] VREF PIX_IN[4422] NB2 NB1 CSA_VREF pixel
xPix4423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[44] VREF PIX_IN[4423] NB2 NB1 CSA_VREF pixel
xPix4424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[44] VREF PIX_IN[4424] NB2 NB1 CSA_VREF pixel
xPix4425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[44] VREF PIX_IN[4425] NB2 NB1 CSA_VREF pixel
xPix4426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[44] VREF PIX_IN[4426] NB2 NB1 CSA_VREF pixel
xPix4427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[44] VREF PIX_IN[4427] NB2 NB1 CSA_VREF pixel
xPix4428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[44] VREF PIX_IN[4428] NB2 NB1 CSA_VREF pixel
xPix4429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[44] VREF PIX_IN[4429] NB2 NB1 CSA_VREF pixel
xPix4430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[44] VREF PIX_IN[4430] NB2 NB1 CSA_VREF pixel
xPix4431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[44] VREF PIX_IN[4431] NB2 NB1 CSA_VREF pixel
xPix4432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[44] VREF PIX_IN[4432] NB2 NB1 CSA_VREF pixel
xPix4433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[44] VREF PIX_IN[4433] NB2 NB1 CSA_VREF pixel
xPix4434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[44] VREF PIX_IN[4434] NB2 NB1 CSA_VREF pixel
xPix4435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[44] VREF PIX_IN[4435] NB2 NB1 CSA_VREF pixel
xPix4436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[44] VREF PIX_IN[4436] NB2 NB1 CSA_VREF pixel
xPix4437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[44] VREF PIX_IN[4437] NB2 NB1 CSA_VREF pixel
xPix4438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[44] VREF PIX_IN[4438] NB2 NB1 CSA_VREF pixel
xPix4439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[44] VREF PIX_IN[4439] NB2 NB1 CSA_VREF pixel
xPix4440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[44] VREF PIX_IN[4440] NB2 NB1 CSA_VREF pixel
xPix4441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[44] VREF PIX_IN[4441] NB2 NB1 CSA_VREF pixel
xPix4442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[44] VREF PIX_IN[4442] NB2 NB1 CSA_VREF pixel
xPix4443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[44] VREF PIX_IN[4443] NB2 NB1 CSA_VREF pixel
xPix4444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[44] VREF PIX_IN[4444] NB2 NB1 CSA_VREF pixel
xPix4445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[44] VREF PIX_IN[4445] NB2 NB1 CSA_VREF pixel
xPix4446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[44] VREF PIX_IN[4446] NB2 NB1 CSA_VREF pixel
xPix4447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[44] VREF PIX_IN[4447] NB2 NB1 CSA_VREF pixel
xPix4448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[44] VREF PIX_IN[4448] NB2 NB1 CSA_VREF pixel
xPix4449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[44] VREF PIX_IN[4449] NB2 NB1 CSA_VREF pixel
xPix4450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[44] VREF PIX_IN[4450] NB2 NB1 CSA_VREF pixel
xPix4451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[44] VREF PIX_IN[4451] NB2 NB1 CSA_VREF pixel
xPix4452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[44] VREF PIX_IN[4452] NB2 NB1 CSA_VREF pixel
xPix4453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[44] VREF PIX_IN[4453] NB2 NB1 CSA_VREF pixel
xPix4454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[44] VREF PIX_IN[4454] NB2 NB1 CSA_VREF pixel
xPix4455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[44] VREF PIX_IN[4455] NB2 NB1 CSA_VREF pixel
xPix4456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[44] VREF PIX_IN[4456] NB2 NB1 CSA_VREF pixel
xPix4457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[44] VREF PIX_IN[4457] NB2 NB1 CSA_VREF pixel
xPix4458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[44] VREF PIX_IN[4458] NB2 NB1 CSA_VREF pixel
xPix4459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[44] VREF PIX_IN[4459] NB2 NB1 CSA_VREF pixel
xPix4460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[44] VREF PIX_IN[4460] NB2 NB1 CSA_VREF pixel
xPix4461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[44] VREF PIX_IN[4461] NB2 NB1 CSA_VREF pixel
xPix4462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[44] VREF PIX_IN[4462] NB2 NB1 CSA_VREF pixel
xPix4463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[44] VREF PIX_IN[4463] NB2 NB1 CSA_VREF pixel
xPix4464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[44] VREF PIX_IN[4464] NB2 NB1 CSA_VREF pixel
xPix4465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[44] VREF PIX_IN[4465] NB2 NB1 CSA_VREF pixel
xPix4466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[44] VREF PIX_IN[4466] NB2 NB1 CSA_VREF pixel
xPix4467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[44] VREF PIX_IN[4467] NB2 NB1 CSA_VREF pixel
xPix4468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[44] VREF PIX_IN[4468] NB2 NB1 CSA_VREF pixel
xPix4469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[44] VREF PIX_IN[4469] NB2 NB1 CSA_VREF pixel
xPix4470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[44] VREF PIX_IN[4470] NB2 NB1 CSA_VREF pixel
xPix4471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[44] VREF PIX_IN[4471] NB2 NB1 CSA_VREF pixel
xPix4472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[44] VREF PIX_IN[4472] NB2 NB1 CSA_VREF pixel
xPix4473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[44] VREF PIX_IN[4473] NB2 NB1 CSA_VREF pixel
xPix4474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[44] VREF PIX_IN[4474] NB2 NB1 CSA_VREF pixel
xPix4475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[44] VREF PIX_IN[4475] NB2 NB1 CSA_VREF pixel
xPix4476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[44] VREF PIX_IN[4476] NB2 NB1 CSA_VREF pixel
xPix4477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[44] VREF PIX_IN[4477] NB2 NB1 CSA_VREF pixel
xPix4478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[44] VREF PIX_IN[4478] NB2 NB1 CSA_VREF pixel
xPix4479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[44] VREF PIX_IN[4479] NB2 NB1 CSA_VREF pixel
xPix4480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[44] VREF PIX_IN[4480] NB2 NB1 CSA_VREF pixel
xPix4481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[44] VREF PIX_IN[4481] NB2 NB1 CSA_VREF pixel
xPix4482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[44] VREF PIX_IN[4482] NB2 NB1 CSA_VREF pixel
xPix4483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[44] VREF PIX_IN[4483] NB2 NB1 CSA_VREF pixel
xPix4484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[44] VREF PIX_IN[4484] NB2 NB1 CSA_VREF pixel
xPix4485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[44] VREF PIX_IN[4485] NB2 NB1 CSA_VREF pixel
xPix4486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[44] VREF PIX_IN[4486] NB2 NB1 CSA_VREF pixel
xPix4487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[44] VREF PIX_IN[4487] NB2 NB1 CSA_VREF pixel
xPix4488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[44] VREF PIX_IN[4488] NB2 NB1 CSA_VREF pixel
xPix4489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[44] VREF PIX_IN[4489] NB2 NB1 CSA_VREF pixel
xPix4490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[44] VREF PIX_IN[4490] NB2 NB1 CSA_VREF pixel
xPix4491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[44] VREF PIX_IN[4491] NB2 NB1 CSA_VREF pixel
xPix4492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[44] VREF PIX_IN[4492] NB2 NB1 CSA_VREF pixel
xPix4493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[44] VREF PIX_IN[4493] NB2 NB1 CSA_VREF pixel
xPix4494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[44] VREF PIX_IN[4494] NB2 NB1 CSA_VREF pixel
xPix4495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[44] VREF PIX_IN[4495] NB2 NB1 CSA_VREF pixel
xPix4496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[44] VREF PIX_IN[4496] NB2 NB1 CSA_VREF pixel
xPix4497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[44] VREF PIX_IN[4497] NB2 NB1 CSA_VREF pixel
xPix4498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[44] VREF PIX_IN[4498] NB2 NB1 CSA_VREF pixel
xPix4499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[44] VREF PIX_IN[4499] NB2 NB1 CSA_VREF pixel
xPix4500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[45] VREF PIX_IN[4500] NB2 NB1 CSA_VREF pixel
xPix4501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[45] VREF PIX_IN[4501] NB2 NB1 CSA_VREF pixel
xPix4502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[45] VREF PIX_IN[4502] NB2 NB1 CSA_VREF pixel
xPix4503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[45] VREF PIX_IN[4503] NB2 NB1 CSA_VREF pixel
xPix4504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[45] VREF PIX_IN[4504] NB2 NB1 CSA_VREF pixel
xPix4505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[45] VREF PIX_IN[4505] NB2 NB1 CSA_VREF pixel
xPix4506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[45] VREF PIX_IN[4506] NB2 NB1 CSA_VREF pixel
xPix4507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[45] VREF PIX_IN[4507] NB2 NB1 CSA_VREF pixel
xPix4508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[45] VREF PIX_IN[4508] NB2 NB1 CSA_VREF pixel
xPix4509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[45] VREF PIX_IN[4509] NB2 NB1 CSA_VREF pixel
xPix4510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[45] VREF PIX_IN[4510] NB2 NB1 CSA_VREF pixel
xPix4511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[45] VREF PIX_IN[4511] NB2 NB1 CSA_VREF pixel
xPix4512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[45] VREF PIX_IN[4512] NB2 NB1 CSA_VREF pixel
xPix4513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[45] VREF PIX_IN[4513] NB2 NB1 CSA_VREF pixel
xPix4514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[45] VREF PIX_IN[4514] NB2 NB1 CSA_VREF pixel
xPix4515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[45] VREF PIX_IN[4515] NB2 NB1 CSA_VREF pixel
xPix4516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[45] VREF PIX_IN[4516] NB2 NB1 CSA_VREF pixel
xPix4517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[45] VREF PIX_IN[4517] NB2 NB1 CSA_VREF pixel
xPix4518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[45] VREF PIX_IN[4518] NB2 NB1 CSA_VREF pixel
xPix4519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[45] VREF PIX_IN[4519] NB2 NB1 CSA_VREF pixel
xPix4520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[45] VREF PIX_IN[4520] NB2 NB1 CSA_VREF pixel
xPix4521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[45] VREF PIX_IN[4521] NB2 NB1 CSA_VREF pixel
xPix4522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[45] VREF PIX_IN[4522] NB2 NB1 CSA_VREF pixel
xPix4523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[45] VREF PIX_IN[4523] NB2 NB1 CSA_VREF pixel
xPix4524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[45] VREF PIX_IN[4524] NB2 NB1 CSA_VREF pixel
xPix4525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[45] VREF PIX_IN[4525] NB2 NB1 CSA_VREF pixel
xPix4526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[45] VREF PIX_IN[4526] NB2 NB1 CSA_VREF pixel
xPix4527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[45] VREF PIX_IN[4527] NB2 NB1 CSA_VREF pixel
xPix4528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[45] VREF PIX_IN[4528] NB2 NB1 CSA_VREF pixel
xPix4529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[45] VREF PIX_IN[4529] NB2 NB1 CSA_VREF pixel
xPix4530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[45] VREF PIX_IN[4530] NB2 NB1 CSA_VREF pixel
xPix4531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[45] VREF PIX_IN[4531] NB2 NB1 CSA_VREF pixel
xPix4532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[45] VREF PIX_IN[4532] NB2 NB1 CSA_VREF pixel
xPix4533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[45] VREF PIX_IN[4533] NB2 NB1 CSA_VREF pixel
xPix4534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[45] VREF PIX_IN[4534] NB2 NB1 CSA_VREF pixel
xPix4535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[45] VREF PIX_IN[4535] NB2 NB1 CSA_VREF pixel
xPix4536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[45] VREF PIX_IN[4536] NB2 NB1 CSA_VREF pixel
xPix4537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[45] VREF PIX_IN[4537] NB2 NB1 CSA_VREF pixel
xPix4538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[45] VREF PIX_IN[4538] NB2 NB1 CSA_VREF pixel
xPix4539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[45] VREF PIX_IN[4539] NB2 NB1 CSA_VREF pixel
xPix4540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[45] VREF PIX_IN[4540] NB2 NB1 CSA_VREF pixel
xPix4541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[45] VREF PIX_IN[4541] NB2 NB1 CSA_VREF pixel
xPix4542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[45] VREF PIX_IN[4542] NB2 NB1 CSA_VREF pixel
xPix4543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[45] VREF PIX_IN[4543] NB2 NB1 CSA_VREF pixel
xPix4544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[45] VREF PIX_IN[4544] NB2 NB1 CSA_VREF pixel
xPix4545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[45] VREF PIX_IN[4545] NB2 NB1 CSA_VREF pixel
xPix4546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[45] VREF PIX_IN[4546] NB2 NB1 CSA_VREF pixel
xPix4547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[45] VREF PIX_IN[4547] NB2 NB1 CSA_VREF pixel
xPix4548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[45] VREF PIX_IN[4548] NB2 NB1 CSA_VREF pixel
xPix4549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[45] VREF PIX_IN[4549] NB2 NB1 CSA_VREF pixel
xPix4550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[45] VREF PIX_IN[4550] NB2 NB1 CSA_VREF pixel
xPix4551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[45] VREF PIX_IN[4551] NB2 NB1 CSA_VREF pixel
xPix4552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[45] VREF PIX_IN[4552] NB2 NB1 CSA_VREF pixel
xPix4553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[45] VREF PIX_IN[4553] NB2 NB1 CSA_VREF pixel
xPix4554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[45] VREF PIX_IN[4554] NB2 NB1 CSA_VREF pixel
xPix4555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[45] VREF PIX_IN[4555] NB2 NB1 CSA_VREF pixel
xPix4556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[45] VREF PIX_IN[4556] NB2 NB1 CSA_VREF pixel
xPix4557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[45] VREF PIX_IN[4557] NB2 NB1 CSA_VREF pixel
xPix4558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[45] VREF PIX_IN[4558] NB2 NB1 CSA_VREF pixel
xPix4559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[45] VREF PIX_IN[4559] NB2 NB1 CSA_VREF pixel
xPix4560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[45] VREF PIX_IN[4560] NB2 NB1 CSA_VREF pixel
xPix4561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[45] VREF PIX_IN[4561] NB2 NB1 CSA_VREF pixel
xPix4562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[45] VREF PIX_IN[4562] NB2 NB1 CSA_VREF pixel
xPix4563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[45] VREF PIX_IN[4563] NB2 NB1 CSA_VREF pixel
xPix4564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[45] VREF PIX_IN[4564] NB2 NB1 CSA_VREF pixel
xPix4565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[45] VREF PIX_IN[4565] NB2 NB1 CSA_VREF pixel
xPix4566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[45] VREF PIX_IN[4566] NB2 NB1 CSA_VREF pixel
xPix4567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[45] VREF PIX_IN[4567] NB2 NB1 CSA_VREF pixel
xPix4568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[45] VREF PIX_IN[4568] NB2 NB1 CSA_VREF pixel
xPix4569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[45] VREF PIX_IN[4569] NB2 NB1 CSA_VREF pixel
xPix4570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[45] VREF PIX_IN[4570] NB2 NB1 CSA_VREF pixel
xPix4571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[45] VREF PIX_IN[4571] NB2 NB1 CSA_VREF pixel
xPix4572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[45] VREF PIX_IN[4572] NB2 NB1 CSA_VREF pixel
xPix4573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[45] VREF PIX_IN[4573] NB2 NB1 CSA_VREF pixel
xPix4574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[45] VREF PIX_IN[4574] NB2 NB1 CSA_VREF pixel
xPix4575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[45] VREF PIX_IN[4575] NB2 NB1 CSA_VREF pixel
xPix4576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[45] VREF PIX_IN[4576] NB2 NB1 CSA_VREF pixel
xPix4577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[45] VREF PIX_IN[4577] NB2 NB1 CSA_VREF pixel
xPix4578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[45] VREF PIX_IN[4578] NB2 NB1 CSA_VREF pixel
xPix4579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[45] VREF PIX_IN[4579] NB2 NB1 CSA_VREF pixel
xPix4580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[45] VREF PIX_IN[4580] NB2 NB1 CSA_VREF pixel
xPix4581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[45] VREF PIX_IN[4581] NB2 NB1 CSA_VREF pixel
xPix4582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[45] VREF PIX_IN[4582] NB2 NB1 CSA_VREF pixel
xPix4583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[45] VREF PIX_IN[4583] NB2 NB1 CSA_VREF pixel
xPix4584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[45] VREF PIX_IN[4584] NB2 NB1 CSA_VREF pixel
xPix4585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[45] VREF PIX_IN[4585] NB2 NB1 CSA_VREF pixel
xPix4586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[45] VREF PIX_IN[4586] NB2 NB1 CSA_VREF pixel
xPix4587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[45] VREF PIX_IN[4587] NB2 NB1 CSA_VREF pixel
xPix4588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[45] VREF PIX_IN[4588] NB2 NB1 CSA_VREF pixel
xPix4589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[45] VREF PIX_IN[4589] NB2 NB1 CSA_VREF pixel
xPix4590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[45] VREF PIX_IN[4590] NB2 NB1 CSA_VREF pixel
xPix4591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[45] VREF PIX_IN[4591] NB2 NB1 CSA_VREF pixel
xPix4592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[45] VREF PIX_IN[4592] NB2 NB1 CSA_VREF pixel
xPix4593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[45] VREF PIX_IN[4593] NB2 NB1 CSA_VREF pixel
xPix4594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[45] VREF PIX_IN[4594] NB2 NB1 CSA_VREF pixel
xPix4595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[45] VREF PIX_IN[4595] NB2 NB1 CSA_VREF pixel
xPix4596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[45] VREF PIX_IN[4596] NB2 NB1 CSA_VREF pixel
xPix4597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[45] VREF PIX_IN[4597] NB2 NB1 CSA_VREF pixel
xPix4598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[45] VREF PIX_IN[4598] NB2 NB1 CSA_VREF pixel
xPix4599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[45] VREF PIX_IN[4599] NB2 NB1 CSA_VREF pixel
xPix4600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[46] VREF PIX_IN[4600] NB2 NB1 CSA_VREF pixel
xPix4601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[46] VREF PIX_IN[4601] NB2 NB1 CSA_VREF pixel
xPix4602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[46] VREF PIX_IN[4602] NB2 NB1 CSA_VREF pixel
xPix4603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[46] VREF PIX_IN[4603] NB2 NB1 CSA_VREF pixel
xPix4604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[46] VREF PIX_IN[4604] NB2 NB1 CSA_VREF pixel
xPix4605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[46] VREF PIX_IN[4605] NB2 NB1 CSA_VREF pixel
xPix4606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[46] VREF PIX_IN[4606] NB2 NB1 CSA_VREF pixel
xPix4607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[46] VREF PIX_IN[4607] NB2 NB1 CSA_VREF pixel
xPix4608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[46] VREF PIX_IN[4608] NB2 NB1 CSA_VREF pixel
xPix4609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[46] VREF PIX_IN[4609] NB2 NB1 CSA_VREF pixel
xPix4610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[46] VREF PIX_IN[4610] NB2 NB1 CSA_VREF pixel
xPix4611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[46] VREF PIX_IN[4611] NB2 NB1 CSA_VREF pixel
xPix4612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[46] VREF PIX_IN[4612] NB2 NB1 CSA_VREF pixel
xPix4613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[46] VREF PIX_IN[4613] NB2 NB1 CSA_VREF pixel
xPix4614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[46] VREF PIX_IN[4614] NB2 NB1 CSA_VREF pixel
xPix4615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[46] VREF PIX_IN[4615] NB2 NB1 CSA_VREF pixel
xPix4616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[46] VREF PIX_IN[4616] NB2 NB1 CSA_VREF pixel
xPix4617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[46] VREF PIX_IN[4617] NB2 NB1 CSA_VREF pixel
xPix4618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[46] VREF PIX_IN[4618] NB2 NB1 CSA_VREF pixel
xPix4619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[46] VREF PIX_IN[4619] NB2 NB1 CSA_VREF pixel
xPix4620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[46] VREF PIX_IN[4620] NB2 NB1 CSA_VREF pixel
xPix4621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[46] VREF PIX_IN[4621] NB2 NB1 CSA_VREF pixel
xPix4622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[46] VREF PIX_IN[4622] NB2 NB1 CSA_VREF pixel
xPix4623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[46] VREF PIX_IN[4623] NB2 NB1 CSA_VREF pixel
xPix4624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[46] VREF PIX_IN[4624] NB2 NB1 CSA_VREF pixel
xPix4625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[46] VREF PIX_IN[4625] NB2 NB1 CSA_VREF pixel
xPix4626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[46] VREF PIX_IN[4626] NB2 NB1 CSA_VREF pixel
xPix4627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[46] VREF PIX_IN[4627] NB2 NB1 CSA_VREF pixel
xPix4628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[46] VREF PIX_IN[4628] NB2 NB1 CSA_VREF pixel
xPix4629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[46] VREF PIX_IN[4629] NB2 NB1 CSA_VREF pixel
xPix4630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[46] VREF PIX_IN[4630] NB2 NB1 CSA_VREF pixel
xPix4631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[46] VREF PIX_IN[4631] NB2 NB1 CSA_VREF pixel
xPix4632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[46] VREF PIX_IN[4632] NB2 NB1 CSA_VREF pixel
xPix4633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[46] VREF PIX_IN[4633] NB2 NB1 CSA_VREF pixel
xPix4634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[46] VREF PIX_IN[4634] NB2 NB1 CSA_VREF pixel
xPix4635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[46] VREF PIX_IN[4635] NB2 NB1 CSA_VREF pixel
xPix4636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[46] VREF PIX_IN[4636] NB2 NB1 CSA_VREF pixel
xPix4637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[46] VREF PIX_IN[4637] NB2 NB1 CSA_VREF pixel
xPix4638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[46] VREF PIX_IN[4638] NB2 NB1 CSA_VREF pixel
xPix4639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[46] VREF PIX_IN[4639] NB2 NB1 CSA_VREF pixel
xPix4640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[46] VREF PIX_IN[4640] NB2 NB1 CSA_VREF pixel
xPix4641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[46] VREF PIX_IN[4641] NB2 NB1 CSA_VREF pixel
xPix4642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[46] VREF PIX_IN[4642] NB2 NB1 CSA_VREF pixel
xPix4643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[46] VREF PIX_IN[4643] NB2 NB1 CSA_VREF pixel
xPix4644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[46] VREF PIX_IN[4644] NB2 NB1 CSA_VREF pixel
xPix4645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[46] VREF PIX_IN[4645] NB2 NB1 CSA_VREF pixel
xPix4646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[46] VREF PIX_IN[4646] NB2 NB1 CSA_VREF pixel
xPix4647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[46] VREF PIX_IN[4647] NB2 NB1 CSA_VREF pixel
xPix4648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[46] VREF PIX_IN[4648] NB2 NB1 CSA_VREF pixel
xPix4649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[46] VREF PIX_IN[4649] NB2 NB1 CSA_VREF pixel
xPix4650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[46] VREF PIX_IN[4650] NB2 NB1 CSA_VREF pixel
xPix4651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[46] VREF PIX_IN[4651] NB2 NB1 CSA_VREF pixel
xPix4652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[46] VREF PIX_IN[4652] NB2 NB1 CSA_VREF pixel
xPix4653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[46] VREF PIX_IN[4653] NB2 NB1 CSA_VREF pixel
xPix4654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[46] VREF PIX_IN[4654] NB2 NB1 CSA_VREF pixel
xPix4655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[46] VREF PIX_IN[4655] NB2 NB1 CSA_VREF pixel
xPix4656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[46] VREF PIX_IN[4656] NB2 NB1 CSA_VREF pixel
xPix4657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[46] VREF PIX_IN[4657] NB2 NB1 CSA_VREF pixel
xPix4658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[46] VREF PIX_IN[4658] NB2 NB1 CSA_VREF pixel
xPix4659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[46] VREF PIX_IN[4659] NB2 NB1 CSA_VREF pixel
xPix4660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[46] VREF PIX_IN[4660] NB2 NB1 CSA_VREF pixel
xPix4661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[46] VREF PIX_IN[4661] NB2 NB1 CSA_VREF pixel
xPix4662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[46] VREF PIX_IN[4662] NB2 NB1 CSA_VREF pixel
xPix4663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[46] VREF PIX_IN[4663] NB2 NB1 CSA_VREF pixel
xPix4664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[46] VREF PIX_IN[4664] NB2 NB1 CSA_VREF pixel
xPix4665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[46] VREF PIX_IN[4665] NB2 NB1 CSA_VREF pixel
xPix4666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[46] VREF PIX_IN[4666] NB2 NB1 CSA_VREF pixel
xPix4667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[46] VREF PIX_IN[4667] NB2 NB1 CSA_VREF pixel
xPix4668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[46] VREF PIX_IN[4668] NB2 NB1 CSA_VREF pixel
xPix4669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[46] VREF PIX_IN[4669] NB2 NB1 CSA_VREF pixel
xPix4670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[46] VREF PIX_IN[4670] NB2 NB1 CSA_VREF pixel
xPix4671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[46] VREF PIX_IN[4671] NB2 NB1 CSA_VREF pixel
xPix4672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[46] VREF PIX_IN[4672] NB2 NB1 CSA_VREF pixel
xPix4673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[46] VREF PIX_IN[4673] NB2 NB1 CSA_VREF pixel
xPix4674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[46] VREF PIX_IN[4674] NB2 NB1 CSA_VREF pixel
xPix4675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[46] VREF PIX_IN[4675] NB2 NB1 CSA_VREF pixel
xPix4676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[46] VREF PIX_IN[4676] NB2 NB1 CSA_VREF pixel
xPix4677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[46] VREF PIX_IN[4677] NB2 NB1 CSA_VREF pixel
xPix4678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[46] VREF PIX_IN[4678] NB2 NB1 CSA_VREF pixel
xPix4679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[46] VREF PIX_IN[4679] NB2 NB1 CSA_VREF pixel
xPix4680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[46] VREF PIX_IN[4680] NB2 NB1 CSA_VREF pixel
xPix4681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[46] VREF PIX_IN[4681] NB2 NB1 CSA_VREF pixel
xPix4682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[46] VREF PIX_IN[4682] NB2 NB1 CSA_VREF pixel
xPix4683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[46] VREF PIX_IN[4683] NB2 NB1 CSA_VREF pixel
xPix4684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[46] VREF PIX_IN[4684] NB2 NB1 CSA_VREF pixel
xPix4685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[46] VREF PIX_IN[4685] NB2 NB1 CSA_VREF pixel
xPix4686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[46] VREF PIX_IN[4686] NB2 NB1 CSA_VREF pixel
xPix4687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[46] VREF PIX_IN[4687] NB2 NB1 CSA_VREF pixel
xPix4688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[46] VREF PIX_IN[4688] NB2 NB1 CSA_VREF pixel
xPix4689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[46] VREF PIX_IN[4689] NB2 NB1 CSA_VREF pixel
xPix4690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[46] VREF PIX_IN[4690] NB2 NB1 CSA_VREF pixel
xPix4691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[46] VREF PIX_IN[4691] NB2 NB1 CSA_VREF pixel
xPix4692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[46] VREF PIX_IN[4692] NB2 NB1 CSA_VREF pixel
xPix4693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[46] VREF PIX_IN[4693] NB2 NB1 CSA_VREF pixel
xPix4694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[46] VREF PIX_IN[4694] NB2 NB1 CSA_VREF pixel
xPix4695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[46] VREF PIX_IN[4695] NB2 NB1 CSA_VREF pixel
xPix4696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[46] VREF PIX_IN[4696] NB2 NB1 CSA_VREF pixel
xPix4697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[46] VREF PIX_IN[4697] NB2 NB1 CSA_VREF pixel
xPix4698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[46] VREF PIX_IN[4698] NB2 NB1 CSA_VREF pixel
xPix4699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[46] VREF PIX_IN[4699] NB2 NB1 CSA_VREF pixel
xPix4700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[47] VREF PIX_IN[4700] NB2 NB1 CSA_VREF pixel
xPix4701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[47] VREF PIX_IN[4701] NB2 NB1 CSA_VREF pixel
xPix4702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[47] VREF PIX_IN[4702] NB2 NB1 CSA_VREF pixel
xPix4703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[47] VREF PIX_IN[4703] NB2 NB1 CSA_VREF pixel
xPix4704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[47] VREF PIX_IN[4704] NB2 NB1 CSA_VREF pixel
xPix4705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[47] VREF PIX_IN[4705] NB2 NB1 CSA_VREF pixel
xPix4706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[47] VREF PIX_IN[4706] NB2 NB1 CSA_VREF pixel
xPix4707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[47] VREF PIX_IN[4707] NB2 NB1 CSA_VREF pixel
xPix4708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[47] VREF PIX_IN[4708] NB2 NB1 CSA_VREF pixel
xPix4709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[47] VREF PIX_IN[4709] NB2 NB1 CSA_VREF pixel
xPix4710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[47] VREF PIX_IN[4710] NB2 NB1 CSA_VREF pixel
xPix4711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[47] VREF PIX_IN[4711] NB2 NB1 CSA_VREF pixel
xPix4712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[47] VREF PIX_IN[4712] NB2 NB1 CSA_VREF pixel
xPix4713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[47] VREF PIX_IN[4713] NB2 NB1 CSA_VREF pixel
xPix4714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[47] VREF PIX_IN[4714] NB2 NB1 CSA_VREF pixel
xPix4715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[47] VREF PIX_IN[4715] NB2 NB1 CSA_VREF pixel
xPix4716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[47] VREF PIX_IN[4716] NB2 NB1 CSA_VREF pixel
xPix4717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[47] VREF PIX_IN[4717] NB2 NB1 CSA_VREF pixel
xPix4718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[47] VREF PIX_IN[4718] NB2 NB1 CSA_VREF pixel
xPix4719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[47] VREF PIX_IN[4719] NB2 NB1 CSA_VREF pixel
xPix4720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[47] VREF PIX_IN[4720] NB2 NB1 CSA_VREF pixel
xPix4721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[47] VREF PIX_IN[4721] NB2 NB1 CSA_VREF pixel
xPix4722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[47] VREF PIX_IN[4722] NB2 NB1 CSA_VREF pixel
xPix4723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[47] VREF PIX_IN[4723] NB2 NB1 CSA_VREF pixel
xPix4724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[47] VREF PIX_IN[4724] NB2 NB1 CSA_VREF pixel
xPix4725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[47] VREF PIX_IN[4725] NB2 NB1 CSA_VREF pixel
xPix4726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[47] VREF PIX_IN[4726] NB2 NB1 CSA_VREF pixel
xPix4727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[47] VREF PIX_IN[4727] NB2 NB1 CSA_VREF pixel
xPix4728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[47] VREF PIX_IN[4728] NB2 NB1 CSA_VREF pixel
xPix4729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[47] VREF PIX_IN[4729] NB2 NB1 CSA_VREF pixel
xPix4730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[47] VREF PIX_IN[4730] NB2 NB1 CSA_VREF pixel
xPix4731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[47] VREF PIX_IN[4731] NB2 NB1 CSA_VREF pixel
xPix4732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[47] VREF PIX_IN[4732] NB2 NB1 CSA_VREF pixel
xPix4733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[47] VREF PIX_IN[4733] NB2 NB1 CSA_VREF pixel
xPix4734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[47] VREF PIX_IN[4734] NB2 NB1 CSA_VREF pixel
xPix4735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[47] VREF PIX_IN[4735] NB2 NB1 CSA_VREF pixel
xPix4736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[47] VREF PIX_IN[4736] NB2 NB1 CSA_VREF pixel
xPix4737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[47] VREF PIX_IN[4737] NB2 NB1 CSA_VREF pixel
xPix4738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[47] VREF PIX_IN[4738] NB2 NB1 CSA_VREF pixel
xPix4739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[47] VREF PIX_IN[4739] NB2 NB1 CSA_VREF pixel
xPix4740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[47] VREF PIX_IN[4740] NB2 NB1 CSA_VREF pixel
xPix4741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[47] VREF PIX_IN[4741] NB2 NB1 CSA_VREF pixel
xPix4742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[47] VREF PIX_IN[4742] NB2 NB1 CSA_VREF pixel
xPix4743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[47] VREF PIX_IN[4743] NB2 NB1 CSA_VREF pixel
xPix4744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[47] VREF PIX_IN[4744] NB2 NB1 CSA_VREF pixel
xPix4745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[47] VREF PIX_IN[4745] NB2 NB1 CSA_VREF pixel
xPix4746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[47] VREF PIX_IN[4746] NB2 NB1 CSA_VREF pixel
xPix4747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[47] VREF PIX_IN[4747] NB2 NB1 CSA_VREF pixel
xPix4748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[47] VREF PIX_IN[4748] NB2 NB1 CSA_VREF pixel
xPix4749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[47] VREF PIX_IN[4749] NB2 NB1 CSA_VREF pixel
xPix4750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[47] VREF PIX_IN[4750] NB2 NB1 CSA_VREF pixel
xPix4751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[47] VREF PIX_IN[4751] NB2 NB1 CSA_VREF pixel
xPix4752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[47] VREF PIX_IN[4752] NB2 NB1 CSA_VREF pixel
xPix4753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[47] VREF PIX_IN[4753] NB2 NB1 CSA_VREF pixel
xPix4754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[47] VREF PIX_IN[4754] NB2 NB1 CSA_VREF pixel
xPix4755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[47] VREF PIX_IN[4755] NB2 NB1 CSA_VREF pixel
xPix4756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[47] VREF PIX_IN[4756] NB2 NB1 CSA_VREF pixel
xPix4757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[47] VREF PIX_IN[4757] NB2 NB1 CSA_VREF pixel
xPix4758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[47] VREF PIX_IN[4758] NB2 NB1 CSA_VREF pixel
xPix4759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[47] VREF PIX_IN[4759] NB2 NB1 CSA_VREF pixel
xPix4760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[47] VREF PIX_IN[4760] NB2 NB1 CSA_VREF pixel
xPix4761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[47] VREF PIX_IN[4761] NB2 NB1 CSA_VREF pixel
xPix4762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[47] VREF PIX_IN[4762] NB2 NB1 CSA_VREF pixel
xPix4763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[47] VREF PIX_IN[4763] NB2 NB1 CSA_VREF pixel
xPix4764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[47] VREF PIX_IN[4764] NB2 NB1 CSA_VREF pixel
xPix4765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[47] VREF PIX_IN[4765] NB2 NB1 CSA_VREF pixel
xPix4766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[47] VREF PIX_IN[4766] NB2 NB1 CSA_VREF pixel
xPix4767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[47] VREF PIX_IN[4767] NB2 NB1 CSA_VREF pixel
xPix4768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[47] VREF PIX_IN[4768] NB2 NB1 CSA_VREF pixel
xPix4769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[47] VREF PIX_IN[4769] NB2 NB1 CSA_VREF pixel
xPix4770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[47] VREF PIX_IN[4770] NB2 NB1 CSA_VREF pixel
xPix4771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[47] VREF PIX_IN[4771] NB2 NB1 CSA_VREF pixel
xPix4772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[47] VREF PIX_IN[4772] NB2 NB1 CSA_VREF pixel
xPix4773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[47] VREF PIX_IN[4773] NB2 NB1 CSA_VREF pixel
xPix4774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[47] VREF PIX_IN[4774] NB2 NB1 CSA_VREF pixel
xPix4775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[47] VREF PIX_IN[4775] NB2 NB1 CSA_VREF pixel
xPix4776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[47] VREF PIX_IN[4776] NB2 NB1 CSA_VREF pixel
xPix4777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[47] VREF PIX_IN[4777] NB2 NB1 CSA_VREF pixel
xPix4778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[47] VREF PIX_IN[4778] NB2 NB1 CSA_VREF pixel
xPix4779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[47] VREF PIX_IN[4779] NB2 NB1 CSA_VREF pixel
xPix4780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[47] VREF PIX_IN[4780] NB2 NB1 CSA_VREF pixel
xPix4781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[47] VREF PIX_IN[4781] NB2 NB1 CSA_VREF pixel
xPix4782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[47] VREF PIX_IN[4782] NB2 NB1 CSA_VREF pixel
xPix4783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[47] VREF PIX_IN[4783] NB2 NB1 CSA_VREF pixel
xPix4784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[47] VREF PIX_IN[4784] NB2 NB1 CSA_VREF pixel
xPix4785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[47] VREF PIX_IN[4785] NB2 NB1 CSA_VREF pixel
xPix4786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[47] VREF PIX_IN[4786] NB2 NB1 CSA_VREF pixel
xPix4787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[47] VREF PIX_IN[4787] NB2 NB1 CSA_VREF pixel
xPix4788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[47] VREF PIX_IN[4788] NB2 NB1 CSA_VREF pixel
xPix4789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[47] VREF PIX_IN[4789] NB2 NB1 CSA_VREF pixel
xPix4790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[47] VREF PIX_IN[4790] NB2 NB1 CSA_VREF pixel
xPix4791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[47] VREF PIX_IN[4791] NB2 NB1 CSA_VREF pixel
xPix4792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[47] VREF PIX_IN[4792] NB2 NB1 CSA_VREF pixel
xPix4793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[47] VREF PIX_IN[4793] NB2 NB1 CSA_VREF pixel
xPix4794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[47] VREF PIX_IN[4794] NB2 NB1 CSA_VREF pixel
xPix4795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[47] VREF PIX_IN[4795] NB2 NB1 CSA_VREF pixel
xPix4796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[47] VREF PIX_IN[4796] NB2 NB1 CSA_VREF pixel
xPix4797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[47] VREF PIX_IN[4797] NB2 NB1 CSA_VREF pixel
xPix4798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[47] VREF PIX_IN[4798] NB2 NB1 CSA_VREF pixel
xPix4799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[47] VREF PIX_IN[4799] NB2 NB1 CSA_VREF pixel
xPix4800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[48] VREF PIX_IN[4800] NB2 NB1 CSA_VREF pixel
xPix4801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[48] VREF PIX_IN[4801] NB2 NB1 CSA_VREF pixel
xPix4802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[48] VREF PIX_IN[4802] NB2 NB1 CSA_VREF pixel
xPix4803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[48] VREF PIX_IN[4803] NB2 NB1 CSA_VREF pixel
xPix4804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[48] VREF PIX_IN[4804] NB2 NB1 CSA_VREF pixel
xPix4805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[48] VREF PIX_IN[4805] NB2 NB1 CSA_VREF pixel
xPix4806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[48] VREF PIX_IN[4806] NB2 NB1 CSA_VREF pixel
xPix4807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[48] VREF PIX_IN[4807] NB2 NB1 CSA_VREF pixel
xPix4808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[48] VREF PIX_IN[4808] NB2 NB1 CSA_VREF pixel
xPix4809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[48] VREF PIX_IN[4809] NB2 NB1 CSA_VREF pixel
xPix4810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[48] VREF PIX_IN[4810] NB2 NB1 CSA_VREF pixel
xPix4811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[48] VREF PIX_IN[4811] NB2 NB1 CSA_VREF pixel
xPix4812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[48] VREF PIX_IN[4812] NB2 NB1 CSA_VREF pixel
xPix4813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[48] VREF PIX_IN[4813] NB2 NB1 CSA_VREF pixel
xPix4814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[48] VREF PIX_IN[4814] NB2 NB1 CSA_VREF pixel
xPix4815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[48] VREF PIX_IN[4815] NB2 NB1 CSA_VREF pixel
xPix4816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[48] VREF PIX_IN[4816] NB2 NB1 CSA_VREF pixel
xPix4817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[48] VREF PIX_IN[4817] NB2 NB1 CSA_VREF pixel
xPix4818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[48] VREF PIX_IN[4818] NB2 NB1 CSA_VREF pixel
xPix4819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[48] VREF PIX_IN[4819] NB2 NB1 CSA_VREF pixel
xPix4820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[48] VREF PIX_IN[4820] NB2 NB1 CSA_VREF pixel
xPix4821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[48] VREF PIX_IN[4821] NB2 NB1 CSA_VREF pixel
xPix4822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[48] VREF PIX_IN[4822] NB2 NB1 CSA_VREF pixel
xPix4823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[48] VREF PIX_IN[4823] NB2 NB1 CSA_VREF pixel
xPix4824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[48] VREF PIX_IN[4824] NB2 NB1 CSA_VREF pixel
xPix4825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[48] VREF PIX_IN[4825] NB2 NB1 CSA_VREF pixel
xPix4826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[48] VREF PIX_IN[4826] NB2 NB1 CSA_VREF pixel
xPix4827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[48] VREF PIX_IN[4827] NB2 NB1 CSA_VREF pixel
xPix4828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[48] VREF PIX_IN[4828] NB2 NB1 CSA_VREF pixel
xPix4829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[48] VREF PIX_IN[4829] NB2 NB1 CSA_VREF pixel
xPix4830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[48] VREF PIX_IN[4830] NB2 NB1 CSA_VREF pixel
xPix4831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[48] VREF PIX_IN[4831] NB2 NB1 CSA_VREF pixel
xPix4832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[48] VREF PIX_IN[4832] NB2 NB1 CSA_VREF pixel
xPix4833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[48] VREF PIX_IN[4833] NB2 NB1 CSA_VREF pixel
xPix4834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[48] VREF PIX_IN[4834] NB2 NB1 CSA_VREF pixel
xPix4835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[48] VREF PIX_IN[4835] NB2 NB1 CSA_VREF pixel
xPix4836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[48] VREF PIX_IN[4836] NB2 NB1 CSA_VREF pixel
xPix4837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[48] VREF PIX_IN[4837] NB2 NB1 CSA_VREF pixel
xPix4838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[48] VREF PIX_IN[4838] NB2 NB1 CSA_VREF pixel
xPix4839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[48] VREF PIX_IN[4839] NB2 NB1 CSA_VREF pixel
xPix4840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[48] VREF PIX_IN[4840] NB2 NB1 CSA_VREF pixel
xPix4841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[48] VREF PIX_IN[4841] NB2 NB1 CSA_VREF pixel
xPix4842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[48] VREF PIX_IN[4842] NB2 NB1 CSA_VREF pixel
xPix4843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[48] VREF PIX_IN[4843] NB2 NB1 CSA_VREF pixel
xPix4844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[48] VREF PIX_IN[4844] NB2 NB1 CSA_VREF pixel
xPix4845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[48] VREF PIX_IN[4845] NB2 NB1 CSA_VREF pixel
xPix4846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[48] VREF PIX_IN[4846] NB2 NB1 CSA_VREF pixel
xPix4847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[48] VREF PIX_IN[4847] NB2 NB1 CSA_VREF pixel
xPix4848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[48] VREF PIX_IN[4848] NB2 NB1 CSA_VREF pixel
xPix4849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[48] VREF PIX_IN[4849] NB2 NB1 CSA_VREF pixel
xPix4850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[48] VREF PIX_IN[4850] NB2 NB1 CSA_VREF pixel
xPix4851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[48] VREF PIX_IN[4851] NB2 NB1 CSA_VREF pixel
xPix4852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[48] VREF PIX_IN[4852] NB2 NB1 CSA_VREF pixel
xPix4853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[48] VREF PIX_IN[4853] NB2 NB1 CSA_VREF pixel
xPix4854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[48] VREF PIX_IN[4854] NB2 NB1 CSA_VREF pixel
xPix4855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[48] VREF PIX_IN[4855] NB2 NB1 CSA_VREF pixel
xPix4856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[48] VREF PIX_IN[4856] NB2 NB1 CSA_VREF pixel
xPix4857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[48] VREF PIX_IN[4857] NB2 NB1 CSA_VREF pixel
xPix4858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[48] VREF PIX_IN[4858] NB2 NB1 CSA_VREF pixel
xPix4859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[48] VREF PIX_IN[4859] NB2 NB1 CSA_VREF pixel
xPix4860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[48] VREF PIX_IN[4860] NB2 NB1 CSA_VREF pixel
xPix4861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[48] VREF PIX_IN[4861] NB2 NB1 CSA_VREF pixel
xPix4862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[48] VREF PIX_IN[4862] NB2 NB1 CSA_VREF pixel
xPix4863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[48] VREF PIX_IN[4863] NB2 NB1 CSA_VREF pixel
xPix4864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[48] VREF PIX_IN[4864] NB2 NB1 CSA_VREF pixel
xPix4865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[48] VREF PIX_IN[4865] NB2 NB1 CSA_VREF pixel
xPix4866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[48] VREF PIX_IN[4866] NB2 NB1 CSA_VREF pixel
xPix4867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[48] VREF PIX_IN[4867] NB2 NB1 CSA_VREF pixel
xPix4868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[48] VREF PIX_IN[4868] NB2 NB1 CSA_VREF pixel
xPix4869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[48] VREF PIX_IN[4869] NB2 NB1 CSA_VREF pixel
xPix4870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[48] VREF PIX_IN[4870] NB2 NB1 CSA_VREF pixel
xPix4871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[48] VREF PIX_IN[4871] NB2 NB1 CSA_VREF pixel
xPix4872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[48] VREF PIX_IN[4872] NB2 NB1 CSA_VREF pixel
xPix4873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[48] VREF PIX_IN[4873] NB2 NB1 CSA_VREF pixel
xPix4874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[48] VREF PIX_IN[4874] NB2 NB1 CSA_VREF pixel
xPix4875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[48] VREF PIX_IN[4875] NB2 NB1 CSA_VREF pixel
xPix4876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[48] VREF PIX_IN[4876] NB2 NB1 CSA_VREF pixel
xPix4877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[48] VREF PIX_IN[4877] NB2 NB1 CSA_VREF pixel
xPix4878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[48] VREF PIX_IN[4878] NB2 NB1 CSA_VREF pixel
xPix4879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[48] VREF PIX_IN[4879] NB2 NB1 CSA_VREF pixel
xPix4880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[48] VREF PIX_IN[4880] NB2 NB1 CSA_VREF pixel
xPix4881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[48] VREF PIX_IN[4881] NB2 NB1 CSA_VREF pixel
xPix4882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[48] VREF PIX_IN[4882] NB2 NB1 CSA_VREF pixel
xPix4883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[48] VREF PIX_IN[4883] NB2 NB1 CSA_VREF pixel
xPix4884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[48] VREF PIX_IN[4884] NB2 NB1 CSA_VREF pixel
xPix4885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[48] VREF PIX_IN[4885] NB2 NB1 CSA_VREF pixel
xPix4886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[48] VREF PIX_IN[4886] NB2 NB1 CSA_VREF pixel
xPix4887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[48] VREF PIX_IN[4887] NB2 NB1 CSA_VREF pixel
xPix4888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[48] VREF PIX_IN[4888] NB2 NB1 CSA_VREF pixel
xPix4889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[48] VREF PIX_IN[4889] NB2 NB1 CSA_VREF pixel
xPix4890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[48] VREF PIX_IN[4890] NB2 NB1 CSA_VREF pixel
xPix4891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[48] VREF PIX_IN[4891] NB2 NB1 CSA_VREF pixel
xPix4892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[48] VREF PIX_IN[4892] NB2 NB1 CSA_VREF pixel
xPix4893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[48] VREF PIX_IN[4893] NB2 NB1 CSA_VREF pixel
xPix4894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[48] VREF PIX_IN[4894] NB2 NB1 CSA_VREF pixel
xPix4895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[48] VREF PIX_IN[4895] NB2 NB1 CSA_VREF pixel
xPix4896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[48] VREF PIX_IN[4896] NB2 NB1 CSA_VREF pixel
xPix4897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[48] VREF PIX_IN[4897] NB2 NB1 CSA_VREF pixel
xPix4898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[48] VREF PIX_IN[4898] NB2 NB1 CSA_VREF pixel
xPix4899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[48] VREF PIX_IN[4899] NB2 NB1 CSA_VREF pixel
xPix4900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[49] VREF PIX_IN[4900] NB2 NB1 CSA_VREF pixel
xPix4901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[49] VREF PIX_IN[4901] NB2 NB1 CSA_VREF pixel
xPix4902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[49] VREF PIX_IN[4902] NB2 NB1 CSA_VREF pixel
xPix4903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[49] VREF PIX_IN[4903] NB2 NB1 CSA_VREF pixel
xPix4904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[49] VREF PIX_IN[4904] NB2 NB1 CSA_VREF pixel
xPix4905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[49] VREF PIX_IN[4905] NB2 NB1 CSA_VREF pixel
xPix4906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[49] VREF PIX_IN[4906] NB2 NB1 CSA_VREF pixel
xPix4907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[49] VREF PIX_IN[4907] NB2 NB1 CSA_VREF pixel
xPix4908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[49] VREF PIX_IN[4908] NB2 NB1 CSA_VREF pixel
xPix4909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[49] VREF PIX_IN[4909] NB2 NB1 CSA_VREF pixel
xPix4910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[49] VREF PIX_IN[4910] NB2 NB1 CSA_VREF pixel
xPix4911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[49] VREF PIX_IN[4911] NB2 NB1 CSA_VREF pixel
xPix4912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[49] VREF PIX_IN[4912] NB2 NB1 CSA_VREF pixel
xPix4913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[49] VREF PIX_IN[4913] NB2 NB1 CSA_VREF pixel
xPix4914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[49] VREF PIX_IN[4914] NB2 NB1 CSA_VREF pixel
xPix4915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[49] VREF PIX_IN[4915] NB2 NB1 CSA_VREF pixel
xPix4916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[49] VREF PIX_IN[4916] NB2 NB1 CSA_VREF pixel
xPix4917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[49] VREF PIX_IN[4917] NB2 NB1 CSA_VREF pixel
xPix4918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[49] VREF PIX_IN[4918] NB2 NB1 CSA_VREF pixel
xPix4919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[49] VREF PIX_IN[4919] NB2 NB1 CSA_VREF pixel
xPix4920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[49] VREF PIX_IN[4920] NB2 NB1 CSA_VREF pixel
xPix4921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[49] VREF PIX_IN[4921] NB2 NB1 CSA_VREF pixel
xPix4922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[49] VREF PIX_IN[4922] NB2 NB1 CSA_VREF pixel
xPix4923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[49] VREF PIX_IN[4923] NB2 NB1 CSA_VREF pixel
xPix4924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[49] VREF PIX_IN[4924] NB2 NB1 CSA_VREF pixel
xPix4925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[49] VREF PIX_IN[4925] NB2 NB1 CSA_VREF pixel
xPix4926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[49] VREF PIX_IN[4926] NB2 NB1 CSA_VREF pixel
xPix4927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[49] VREF PIX_IN[4927] NB2 NB1 CSA_VREF pixel
xPix4928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[49] VREF PIX_IN[4928] NB2 NB1 CSA_VREF pixel
xPix4929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[49] VREF PIX_IN[4929] NB2 NB1 CSA_VREF pixel
xPix4930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[49] VREF PIX_IN[4930] NB2 NB1 CSA_VREF pixel
xPix4931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[49] VREF PIX_IN[4931] NB2 NB1 CSA_VREF pixel
xPix4932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[49] VREF PIX_IN[4932] NB2 NB1 CSA_VREF pixel
xPix4933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[49] VREF PIX_IN[4933] NB2 NB1 CSA_VREF pixel
xPix4934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[49] VREF PIX_IN[4934] NB2 NB1 CSA_VREF pixel
xPix4935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[49] VREF PIX_IN[4935] NB2 NB1 CSA_VREF pixel
xPix4936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[49] VREF PIX_IN[4936] NB2 NB1 CSA_VREF pixel
xPix4937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[49] VREF PIX_IN[4937] NB2 NB1 CSA_VREF pixel
xPix4938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[49] VREF PIX_IN[4938] NB2 NB1 CSA_VREF pixel
xPix4939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[49] VREF PIX_IN[4939] NB2 NB1 CSA_VREF pixel
xPix4940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[49] VREF PIX_IN[4940] NB2 NB1 CSA_VREF pixel
xPix4941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[49] VREF PIX_IN[4941] NB2 NB1 CSA_VREF pixel
xPix4942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[49] VREF PIX_IN[4942] NB2 NB1 CSA_VREF pixel
xPix4943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[49] VREF PIX_IN[4943] NB2 NB1 CSA_VREF pixel
xPix4944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[49] VREF PIX_IN[4944] NB2 NB1 CSA_VREF pixel
xPix4945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[49] VREF PIX_IN[4945] NB2 NB1 CSA_VREF pixel
xPix4946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[49] VREF PIX_IN[4946] NB2 NB1 CSA_VREF pixel
xPix4947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[49] VREF PIX_IN[4947] NB2 NB1 CSA_VREF pixel
xPix4948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[49] VREF PIX_IN[4948] NB2 NB1 CSA_VREF pixel
xPix4949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[49] VREF PIX_IN[4949] NB2 NB1 CSA_VREF pixel
xPix4950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[49] VREF PIX_IN[4950] NB2 NB1 CSA_VREF pixel
xPix4951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[49] VREF PIX_IN[4951] NB2 NB1 CSA_VREF pixel
xPix4952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[49] VREF PIX_IN[4952] NB2 NB1 CSA_VREF pixel
xPix4953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[49] VREF PIX_IN[4953] NB2 NB1 CSA_VREF pixel
xPix4954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[49] VREF PIX_IN[4954] NB2 NB1 CSA_VREF pixel
xPix4955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[49] VREF PIX_IN[4955] NB2 NB1 CSA_VREF pixel
xPix4956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[49] VREF PIX_IN[4956] NB2 NB1 CSA_VREF pixel
xPix4957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[49] VREF PIX_IN[4957] NB2 NB1 CSA_VREF pixel
xPix4958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[49] VREF PIX_IN[4958] NB2 NB1 CSA_VREF pixel
xPix4959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[49] VREF PIX_IN[4959] NB2 NB1 CSA_VREF pixel
xPix4960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[49] VREF PIX_IN[4960] NB2 NB1 CSA_VREF pixel
xPix4961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[49] VREF PIX_IN[4961] NB2 NB1 CSA_VREF pixel
xPix4962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[49] VREF PIX_IN[4962] NB2 NB1 CSA_VREF pixel
xPix4963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[49] VREF PIX_IN[4963] NB2 NB1 CSA_VREF pixel
xPix4964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[49] VREF PIX_IN[4964] NB2 NB1 CSA_VREF pixel
xPix4965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[49] VREF PIX_IN[4965] NB2 NB1 CSA_VREF pixel
xPix4966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[49] VREF PIX_IN[4966] NB2 NB1 CSA_VREF pixel
xPix4967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[49] VREF PIX_IN[4967] NB2 NB1 CSA_VREF pixel
xPix4968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[49] VREF PIX_IN[4968] NB2 NB1 CSA_VREF pixel
xPix4969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[49] VREF PIX_IN[4969] NB2 NB1 CSA_VREF pixel
xPix4970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[49] VREF PIX_IN[4970] NB2 NB1 CSA_VREF pixel
xPix4971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[49] VREF PIX_IN[4971] NB2 NB1 CSA_VREF pixel
xPix4972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[49] VREF PIX_IN[4972] NB2 NB1 CSA_VREF pixel
xPix4973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[49] VREF PIX_IN[4973] NB2 NB1 CSA_VREF pixel
xPix4974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[49] VREF PIX_IN[4974] NB2 NB1 CSA_VREF pixel
xPix4975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[49] VREF PIX_IN[4975] NB2 NB1 CSA_VREF pixel
xPix4976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[49] VREF PIX_IN[4976] NB2 NB1 CSA_VREF pixel
xPix4977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[49] VREF PIX_IN[4977] NB2 NB1 CSA_VREF pixel
xPix4978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[49] VREF PIX_IN[4978] NB2 NB1 CSA_VREF pixel
xPix4979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[49] VREF PIX_IN[4979] NB2 NB1 CSA_VREF pixel
xPix4980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[49] VREF PIX_IN[4980] NB2 NB1 CSA_VREF pixel
xPix4981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[49] VREF PIX_IN[4981] NB2 NB1 CSA_VREF pixel
xPix4982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[49] VREF PIX_IN[4982] NB2 NB1 CSA_VREF pixel
xPix4983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[49] VREF PIX_IN[4983] NB2 NB1 CSA_VREF pixel
xPix4984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[49] VREF PIX_IN[4984] NB2 NB1 CSA_VREF pixel
xPix4985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[49] VREF PIX_IN[4985] NB2 NB1 CSA_VREF pixel
xPix4986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[49] VREF PIX_IN[4986] NB2 NB1 CSA_VREF pixel
xPix4987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[49] VREF PIX_IN[4987] NB2 NB1 CSA_VREF pixel
xPix4988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[49] VREF PIX_IN[4988] NB2 NB1 CSA_VREF pixel
xPix4989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[49] VREF PIX_IN[4989] NB2 NB1 CSA_VREF pixel
xPix4990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[49] VREF PIX_IN[4990] NB2 NB1 CSA_VREF pixel
xPix4991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[49] VREF PIX_IN[4991] NB2 NB1 CSA_VREF pixel
xPix4992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[49] VREF PIX_IN[4992] NB2 NB1 CSA_VREF pixel
xPix4993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[49] VREF PIX_IN[4993] NB2 NB1 CSA_VREF pixel
xPix4994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[49] VREF PIX_IN[4994] NB2 NB1 CSA_VREF pixel
xPix4995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[49] VREF PIX_IN[4995] NB2 NB1 CSA_VREF pixel
xPix4996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[49] VREF PIX_IN[4996] NB2 NB1 CSA_VREF pixel
xPix4997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[49] VREF PIX_IN[4997] NB2 NB1 CSA_VREF pixel
xPix4998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[49] VREF PIX_IN[4998] NB2 NB1 CSA_VREF pixel
xPix4999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[49] VREF PIX_IN[4999] NB2 NB1 CSA_VREF pixel
xPix5000 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[50] VREF PIX_IN[5000] NB2 NB1 CSA_VREF pixel
xPix5001 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[50] VREF PIX_IN[5001] NB2 NB1 CSA_VREF pixel
xPix5002 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[50] VREF PIX_IN[5002] NB2 NB1 CSA_VREF pixel
xPix5003 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[50] VREF PIX_IN[5003] NB2 NB1 CSA_VREF pixel
xPix5004 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[50] VREF PIX_IN[5004] NB2 NB1 CSA_VREF pixel
xPix5005 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[50] VREF PIX_IN[5005] NB2 NB1 CSA_VREF pixel
xPix5006 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[50] VREF PIX_IN[5006] NB2 NB1 CSA_VREF pixel
xPix5007 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[50] VREF PIX_IN[5007] NB2 NB1 CSA_VREF pixel
xPix5008 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[50] VREF PIX_IN[5008] NB2 NB1 CSA_VREF pixel
xPix5009 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[50] VREF PIX_IN[5009] NB2 NB1 CSA_VREF pixel
xPix5010 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[50] VREF PIX_IN[5010] NB2 NB1 CSA_VREF pixel
xPix5011 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[50] VREF PIX_IN[5011] NB2 NB1 CSA_VREF pixel
xPix5012 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[50] VREF PIX_IN[5012] NB2 NB1 CSA_VREF pixel
xPix5013 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[50] VREF PIX_IN[5013] NB2 NB1 CSA_VREF pixel
xPix5014 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[50] VREF PIX_IN[5014] NB2 NB1 CSA_VREF pixel
xPix5015 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[50] VREF PIX_IN[5015] NB2 NB1 CSA_VREF pixel
xPix5016 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[50] VREF PIX_IN[5016] NB2 NB1 CSA_VREF pixel
xPix5017 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[50] VREF PIX_IN[5017] NB2 NB1 CSA_VREF pixel
xPix5018 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[50] VREF PIX_IN[5018] NB2 NB1 CSA_VREF pixel
xPix5019 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[50] VREF PIX_IN[5019] NB2 NB1 CSA_VREF pixel
xPix5020 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[50] VREF PIX_IN[5020] NB2 NB1 CSA_VREF pixel
xPix5021 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[50] VREF PIX_IN[5021] NB2 NB1 CSA_VREF pixel
xPix5022 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[50] VREF PIX_IN[5022] NB2 NB1 CSA_VREF pixel
xPix5023 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[50] VREF PIX_IN[5023] NB2 NB1 CSA_VREF pixel
xPix5024 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[50] VREF PIX_IN[5024] NB2 NB1 CSA_VREF pixel
xPix5025 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[50] VREF PIX_IN[5025] NB2 NB1 CSA_VREF pixel
xPix5026 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[50] VREF PIX_IN[5026] NB2 NB1 CSA_VREF pixel
xPix5027 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[50] VREF PIX_IN[5027] NB2 NB1 CSA_VREF pixel
xPix5028 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[50] VREF PIX_IN[5028] NB2 NB1 CSA_VREF pixel
xPix5029 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[50] VREF PIX_IN[5029] NB2 NB1 CSA_VREF pixel
xPix5030 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[50] VREF PIX_IN[5030] NB2 NB1 CSA_VREF pixel
xPix5031 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[50] VREF PIX_IN[5031] NB2 NB1 CSA_VREF pixel
xPix5032 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[50] VREF PIX_IN[5032] NB2 NB1 CSA_VREF pixel
xPix5033 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[50] VREF PIX_IN[5033] NB2 NB1 CSA_VREF pixel
xPix5034 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[50] VREF PIX_IN[5034] NB2 NB1 CSA_VREF pixel
xPix5035 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[50] VREF PIX_IN[5035] NB2 NB1 CSA_VREF pixel
xPix5036 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[50] VREF PIX_IN[5036] NB2 NB1 CSA_VREF pixel
xPix5037 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[50] VREF PIX_IN[5037] NB2 NB1 CSA_VREF pixel
xPix5038 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[50] VREF PIX_IN[5038] NB2 NB1 CSA_VREF pixel
xPix5039 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[50] VREF PIX_IN[5039] NB2 NB1 CSA_VREF pixel
xPix5040 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[50] VREF PIX_IN[5040] NB2 NB1 CSA_VREF pixel
xPix5041 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[50] VREF PIX_IN[5041] NB2 NB1 CSA_VREF pixel
xPix5042 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[50] VREF PIX_IN[5042] NB2 NB1 CSA_VREF pixel
xPix5043 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[50] VREF PIX_IN[5043] NB2 NB1 CSA_VREF pixel
xPix5044 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[50] VREF PIX_IN[5044] NB2 NB1 CSA_VREF pixel
xPix5045 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[50] VREF PIX_IN[5045] NB2 NB1 CSA_VREF pixel
xPix5046 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[50] VREF PIX_IN[5046] NB2 NB1 CSA_VREF pixel
xPix5047 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[50] VREF PIX_IN[5047] NB2 NB1 CSA_VREF pixel
xPix5048 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[50] VREF PIX_IN[5048] NB2 NB1 CSA_VREF pixel
xPix5049 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[50] VREF PIX_IN[5049] NB2 NB1 CSA_VREF pixel
xPix5050 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[50] VREF PIX_IN[5050] NB2 NB1 CSA_VREF pixel
xPix5051 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[50] VREF PIX_IN[5051] NB2 NB1 CSA_VREF pixel
xPix5052 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[50] VREF PIX_IN[5052] NB2 NB1 CSA_VREF pixel
xPix5053 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[50] VREF PIX_IN[5053] NB2 NB1 CSA_VREF pixel
xPix5054 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[50] VREF PIX_IN[5054] NB2 NB1 CSA_VREF pixel
xPix5055 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[50] VREF PIX_IN[5055] NB2 NB1 CSA_VREF pixel
xPix5056 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[50] VREF PIX_IN[5056] NB2 NB1 CSA_VREF pixel
xPix5057 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[50] VREF PIX_IN[5057] NB2 NB1 CSA_VREF pixel
xPix5058 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[50] VREF PIX_IN[5058] NB2 NB1 CSA_VREF pixel
xPix5059 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[50] VREF PIX_IN[5059] NB2 NB1 CSA_VREF pixel
xPix5060 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[50] VREF PIX_IN[5060] NB2 NB1 CSA_VREF pixel
xPix5061 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[50] VREF PIX_IN[5061] NB2 NB1 CSA_VREF pixel
xPix5062 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[50] VREF PIX_IN[5062] NB2 NB1 CSA_VREF pixel
xPix5063 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[50] VREF PIX_IN[5063] NB2 NB1 CSA_VREF pixel
xPix5064 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[50] VREF PIX_IN[5064] NB2 NB1 CSA_VREF pixel
xPix5065 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[50] VREF PIX_IN[5065] NB2 NB1 CSA_VREF pixel
xPix5066 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[50] VREF PIX_IN[5066] NB2 NB1 CSA_VREF pixel
xPix5067 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[50] VREF PIX_IN[5067] NB2 NB1 CSA_VREF pixel
xPix5068 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[50] VREF PIX_IN[5068] NB2 NB1 CSA_VREF pixel
xPix5069 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[50] VREF PIX_IN[5069] NB2 NB1 CSA_VREF pixel
xPix5070 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[50] VREF PIX_IN[5070] NB2 NB1 CSA_VREF pixel
xPix5071 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[50] VREF PIX_IN[5071] NB2 NB1 CSA_VREF pixel
xPix5072 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[50] VREF PIX_IN[5072] NB2 NB1 CSA_VREF pixel
xPix5073 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[50] VREF PIX_IN[5073] NB2 NB1 CSA_VREF pixel
xPix5074 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[50] VREF PIX_IN[5074] NB2 NB1 CSA_VREF pixel
xPix5075 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[50] VREF PIX_IN[5075] NB2 NB1 CSA_VREF pixel
xPix5076 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[50] VREF PIX_IN[5076] NB2 NB1 CSA_VREF pixel
xPix5077 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[50] VREF PIX_IN[5077] NB2 NB1 CSA_VREF pixel
xPix5078 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[50] VREF PIX_IN[5078] NB2 NB1 CSA_VREF pixel
xPix5079 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[50] VREF PIX_IN[5079] NB2 NB1 CSA_VREF pixel
xPix5080 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[50] VREF PIX_IN[5080] NB2 NB1 CSA_VREF pixel
xPix5081 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[50] VREF PIX_IN[5081] NB2 NB1 CSA_VREF pixel
xPix5082 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[50] VREF PIX_IN[5082] NB2 NB1 CSA_VREF pixel
xPix5083 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[50] VREF PIX_IN[5083] NB2 NB1 CSA_VREF pixel
xPix5084 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[50] VREF PIX_IN[5084] NB2 NB1 CSA_VREF pixel
xPix5085 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[50] VREF PIX_IN[5085] NB2 NB1 CSA_VREF pixel
xPix5086 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[50] VREF PIX_IN[5086] NB2 NB1 CSA_VREF pixel
xPix5087 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[50] VREF PIX_IN[5087] NB2 NB1 CSA_VREF pixel
xPix5088 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[50] VREF PIX_IN[5088] NB2 NB1 CSA_VREF pixel
xPix5089 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[50] VREF PIX_IN[5089] NB2 NB1 CSA_VREF pixel
xPix5090 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[50] VREF PIX_IN[5090] NB2 NB1 CSA_VREF pixel
xPix5091 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[50] VREF PIX_IN[5091] NB2 NB1 CSA_VREF pixel
xPix5092 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[50] VREF PIX_IN[5092] NB2 NB1 CSA_VREF pixel
xPix5093 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[50] VREF PIX_IN[5093] NB2 NB1 CSA_VREF pixel
xPix5094 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[50] VREF PIX_IN[5094] NB2 NB1 CSA_VREF pixel
xPix5095 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[50] VREF PIX_IN[5095] NB2 NB1 CSA_VREF pixel
xPix5096 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[50] VREF PIX_IN[5096] NB2 NB1 CSA_VREF pixel
xPix5097 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[50] VREF PIX_IN[5097] NB2 NB1 CSA_VREF pixel
xPix5098 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[50] VREF PIX_IN[5098] NB2 NB1 CSA_VREF pixel
xPix5099 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[50] VREF PIX_IN[5099] NB2 NB1 CSA_VREF pixel
xPix5100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[51] VREF PIX_IN[5100] NB2 NB1 CSA_VREF pixel
xPix5101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[51] VREF PIX_IN[5101] NB2 NB1 CSA_VREF pixel
xPix5102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[51] VREF PIX_IN[5102] NB2 NB1 CSA_VREF pixel
xPix5103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[51] VREF PIX_IN[5103] NB2 NB1 CSA_VREF pixel
xPix5104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[51] VREF PIX_IN[5104] NB2 NB1 CSA_VREF pixel
xPix5105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[51] VREF PIX_IN[5105] NB2 NB1 CSA_VREF pixel
xPix5106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[51] VREF PIX_IN[5106] NB2 NB1 CSA_VREF pixel
xPix5107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[51] VREF PIX_IN[5107] NB2 NB1 CSA_VREF pixel
xPix5108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[51] VREF PIX_IN[5108] NB2 NB1 CSA_VREF pixel
xPix5109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[51] VREF PIX_IN[5109] NB2 NB1 CSA_VREF pixel
xPix5110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[51] VREF PIX_IN[5110] NB2 NB1 CSA_VREF pixel
xPix5111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[51] VREF PIX_IN[5111] NB2 NB1 CSA_VREF pixel
xPix5112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[51] VREF PIX_IN[5112] NB2 NB1 CSA_VREF pixel
xPix5113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[51] VREF PIX_IN[5113] NB2 NB1 CSA_VREF pixel
xPix5114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[51] VREF PIX_IN[5114] NB2 NB1 CSA_VREF pixel
xPix5115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[51] VREF PIX_IN[5115] NB2 NB1 CSA_VREF pixel
xPix5116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[51] VREF PIX_IN[5116] NB2 NB1 CSA_VREF pixel
xPix5117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[51] VREF PIX_IN[5117] NB2 NB1 CSA_VREF pixel
xPix5118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[51] VREF PIX_IN[5118] NB2 NB1 CSA_VREF pixel
xPix5119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[51] VREF PIX_IN[5119] NB2 NB1 CSA_VREF pixel
xPix5120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[51] VREF PIX_IN[5120] NB2 NB1 CSA_VREF pixel
xPix5121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[51] VREF PIX_IN[5121] NB2 NB1 CSA_VREF pixel
xPix5122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[51] VREF PIX_IN[5122] NB2 NB1 CSA_VREF pixel
xPix5123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[51] VREF PIX_IN[5123] NB2 NB1 CSA_VREF pixel
xPix5124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[51] VREF PIX_IN[5124] NB2 NB1 CSA_VREF pixel
xPix5125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[51] VREF PIX_IN[5125] NB2 NB1 CSA_VREF pixel
xPix5126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[51] VREF PIX_IN[5126] NB2 NB1 CSA_VREF pixel
xPix5127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[51] VREF PIX_IN[5127] NB2 NB1 CSA_VREF pixel
xPix5128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[51] VREF PIX_IN[5128] NB2 NB1 CSA_VREF pixel
xPix5129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[51] VREF PIX_IN[5129] NB2 NB1 CSA_VREF pixel
xPix5130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[51] VREF PIX_IN[5130] NB2 NB1 CSA_VREF pixel
xPix5131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[51] VREF PIX_IN[5131] NB2 NB1 CSA_VREF pixel
xPix5132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[51] VREF PIX_IN[5132] NB2 NB1 CSA_VREF pixel
xPix5133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[51] VREF PIX_IN[5133] NB2 NB1 CSA_VREF pixel
xPix5134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[51] VREF PIX_IN[5134] NB2 NB1 CSA_VREF pixel
xPix5135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[51] VREF PIX_IN[5135] NB2 NB1 CSA_VREF pixel
xPix5136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[51] VREF PIX_IN[5136] NB2 NB1 CSA_VREF pixel
xPix5137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[51] VREF PIX_IN[5137] NB2 NB1 CSA_VREF pixel
xPix5138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[51] VREF PIX_IN[5138] NB2 NB1 CSA_VREF pixel
xPix5139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[51] VREF PIX_IN[5139] NB2 NB1 CSA_VREF pixel
xPix5140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[51] VREF PIX_IN[5140] NB2 NB1 CSA_VREF pixel
xPix5141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[51] VREF PIX_IN[5141] NB2 NB1 CSA_VREF pixel
xPix5142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[51] VREF PIX_IN[5142] NB2 NB1 CSA_VREF pixel
xPix5143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[51] VREF PIX_IN[5143] NB2 NB1 CSA_VREF pixel
xPix5144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[51] VREF PIX_IN[5144] NB2 NB1 CSA_VREF pixel
xPix5145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[51] VREF PIX_IN[5145] NB2 NB1 CSA_VREF pixel
xPix5146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[51] VREF PIX_IN[5146] NB2 NB1 CSA_VREF pixel
xPix5147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[51] VREF PIX_IN[5147] NB2 NB1 CSA_VREF pixel
xPix5148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[51] VREF PIX_IN[5148] NB2 NB1 CSA_VREF pixel
xPix5149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[51] VREF PIX_IN[5149] NB2 NB1 CSA_VREF pixel
xPix5150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[51] VREF PIX_IN[5150] NB2 NB1 CSA_VREF pixel
xPix5151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[51] VREF PIX_IN[5151] NB2 NB1 CSA_VREF pixel
xPix5152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[51] VREF PIX_IN[5152] NB2 NB1 CSA_VREF pixel
xPix5153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[51] VREF PIX_IN[5153] NB2 NB1 CSA_VREF pixel
xPix5154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[51] VREF PIX_IN[5154] NB2 NB1 CSA_VREF pixel
xPix5155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[51] VREF PIX_IN[5155] NB2 NB1 CSA_VREF pixel
xPix5156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[51] VREF PIX_IN[5156] NB2 NB1 CSA_VREF pixel
xPix5157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[51] VREF PIX_IN[5157] NB2 NB1 CSA_VREF pixel
xPix5158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[51] VREF PIX_IN[5158] NB2 NB1 CSA_VREF pixel
xPix5159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[51] VREF PIX_IN[5159] NB2 NB1 CSA_VREF pixel
xPix5160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[51] VREF PIX_IN[5160] NB2 NB1 CSA_VREF pixel
xPix5161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[51] VREF PIX_IN[5161] NB2 NB1 CSA_VREF pixel
xPix5162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[51] VREF PIX_IN[5162] NB2 NB1 CSA_VREF pixel
xPix5163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[51] VREF PIX_IN[5163] NB2 NB1 CSA_VREF pixel
xPix5164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[51] VREF PIX_IN[5164] NB2 NB1 CSA_VREF pixel
xPix5165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[51] VREF PIX_IN[5165] NB2 NB1 CSA_VREF pixel
xPix5166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[51] VREF PIX_IN[5166] NB2 NB1 CSA_VREF pixel
xPix5167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[51] VREF PIX_IN[5167] NB2 NB1 CSA_VREF pixel
xPix5168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[51] VREF PIX_IN[5168] NB2 NB1 CSA_VREF pixel
xPix5169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[51] VREF PIX_IN[5169] NB2 NB1 CSA_VREF pixel
xPix5170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[51] VREF PIX_IN[5170] NB2 NB1 CSA_VREF pixel
xPix5171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[51] VREF PIX_IN[5171] NB2 NB1 CSA_VREF pixel
xPix5172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[51] VREF PIX_IN[5172] NB2 NB1 CSA_VREF pixel
xPix5173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[51] VREF PIX_IN[5173] NB2 NB1 CSA_VREF pixel
xPix5174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[51] VREF PIX_IN[5174] NB2 NB1 CSA_VREF pixel
xPix5175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[51] VREF PIX_IN[5175] NB2 NB1 CSA_VREF pixel
xPix5176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[51] VREF PIX_IN[5176] NB2 NB1 CSA_VREF pixel
xPix5177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[51] VREF PIX_IN[5177] NB2 NB1 CSA_VREF pixel
xPix5178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[51] VREF PIX_IN[5178] NB2 NB1 CSA_VREF pixel
xPix5179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[51] VREF PIX_IN[5179] NB2 NB1 CSA_VREF pixel
xPix5180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[51] VREF PIX_IN[5180] NB2 NB1 CSA_VREF pixel
xPix5181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[51] VREF PIX_IN[5181] NB2 NB1 CSA_VREF pixel
xPix5182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[51] VREF PIX_IN[5182] NB2 NB1 CSA_VREF pixel
xPix5183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[51] VREF PIX_IN[5183] NB2 NB1 CSA_VREF pixel
xPix5184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[51] VREF PIX_IN[5184] NB2 NB1 CSA_VREF pixel
xPix5185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[51] VREF PIX_IN[5185] NB2 NB1 CSA_VREF pixel
xPix5186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[51] VREF PIX_IN[5186] NB2 NB1 CSA_VREF pixel
xPix5187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[51] VREF PIX_IN[5187] NB2 NB1 CSA_VREF pixel
xPix5188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[51] VREF PIX_IN[5188] NB2 NB1 CSA_VREF pixel
xPix5189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[51] VREF PIX_IN[5189] NB2 NB1 CSA_VREF pixel
xPix5190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[51] VREF PIX_IN[5190] NB2 NB1 CSA_VREF pixel
xPix5191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[51] VREF PIX_IN[5191] NB2 NB1 CSA_VREF pixel
xPix5192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[51] VREF PIX_IN[5192] NB2 NB1 CSA_VREF pixel
xPix5193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[51] VREF PIX_IN[5193] NB2 NB1 CSA_VREF pixel
xPix5194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[51] VREF PIX_IN[5194] NB2 NB1 CSA_VREF pixel
xPix5195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[51] VREF PIX_IN[5195] NB2 NB1 CSA_VREF pixel
xPix5196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[51] VREF PIX_IN[5196] NB2 NB1 CSA_VREF pixel
xPix5197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[51] VREF PIX_IN[5197] NB2 NB1 CSA_VREF pixel
xPix5198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[51] VREF PIX_IN[5198] NB2 NB1 CSA_VREF pixel
xPix5199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[51] VREF PIX_IN[5199] NB2 NB1 CSA_VREF pixel
xPix5200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[52] VREF PIX_IN[5200] NB2 NB1 CSA_VREF pixel
xPix5201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[52] VREF PIX_IN[5201] NB2 NB1 CSA_VREF pixel
xPix5202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[52] VREF PIX_IN[5202] NB2 NB1 CSA_VREF pixel
xPix5203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[52] VREF PIX_IN[5203] NB2 NB1 CSA_VREF pixel
xPix5204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[52] VREF PIX_IN[5204] NB2 NB1 CSA_VREF pixel
xPix5205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[52] VREF PIX_IN[5205] NB2 NB1 CSA_VREF pixel
xPix5206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[52] VREF PIX_IN[5206] NB2 NB1 CSA_VREF pixel
xPix5207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[52] VREF PIX_IN[5207] NB2 NB1 CSA_VREF pixel
xPix5208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[52] VREF PIX_IN[5208] NB2 NB1 CSA_VREF pixel
xPix5209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[52] VREF PIX_IN[5209] NB2 NB1 CSA_VREF pixel
xPix5210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[52] VREF PIX_IN[5210] NB2 NB1 CSA_VREF pixel
xPix5211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[52] VREF PIX_IN[5211] NB2 NB1 CSA_VREF pixel
xPix5212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[52] VREF PIX_IN[5212] NB2 NB1 CSA_VREF pixel
xPix5213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[52] VREF PIX_IN[5213] NB2 NB1 CSA_VREF pixel
xPix5214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[52] VREF PIX_IN[5214] NB2 NB1 CSA_VREF pixel
xPix5215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[52] VREF PIX_IN[5215] NB2 NB1 CSA_VREF pixel
xPix5216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[52] VREF PIX_IN[5216] NB2 NB1 CSA_VREF pixel
xPix5217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[52] VREF PIX_IN[5217] NB2 NB1 CSA_VREF pixel
xPix5218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[52] VREF PIX_IN[5218] NB2 NB1 CSA_VREF pixel
xPix5219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[52] VREF PIX_IN[5219] NB2 NB1 CSA_VREF pixel
xPix5220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[52] VREF PIX_IN[5220] NB2 NB1 CSA_VREF pixel
xPix5221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[52] VREF PIX_IN[5221] NB2 NB1 CSA_VREF pixel
xPix5222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[52] VREF PIX_IN[5222] NB2 NB1 CSA_VREF pixel
xPix5223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[52] VREF PIX_IN[5223] NB2 NB1 CSA_VREF pixel
xPix5224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[52] VREF PIX_IN[5224] NB2 NB1 CSA_VREF pixel
xPix5225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[52] VREF PIX_IN[5225] NB2 NB1 CSA_VREF pixel
xPix5226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[52] VREF PIX_IN[5226] NB2 NB1 CSA_VREF pixel
xPix5227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[52] VREF PIX_IN[5227] NB2 NB1 CSA_VREF pixel
xPix5228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[52] VREF PIX_IN[5228] NB2 NB1 CSA_VREF pixel
xPix5229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[52] VREF PIX_IN[5229] NB2 NB1 CSA_VREF pixel
xPix5230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[52] VREF PIX_IN[5230] NB2 NB1 CSA_VREF pixel
xPix5231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[52] VREF PIX_IN[5231] NB2 NB1 CSA_VREF pixel
xPix5232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[52] VREF PIX_IN[5232] NB2 NB1 CSA_VREF pixel
xPix5233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[52] VREF PIX_IN[5233] NB2 NB1 CSA_VREF pixel
xPix5234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[52] VREF PIX_IN[5234] NB2 NB1 CSA_VREF pixel
xPix5235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[52] VREF PIX_IN[5235] NB2 NB1 CSA_VREF pixel
xPix5236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[52] VREF PIX_IN[5236] NB2 NB1 CSA_VREF pixel
xPix5237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[52] VREF PIX_IN[5237] NB2 NB1 CSA_VREF pixel
xPix5238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[52] VREF PIX_IN[5238] NB2 NB1 CSA_VREF pixel
xPix5239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[52] VREF PIX_IN[5239] NB2 NB1 CSA_VREF pixel
xPix5240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[52] VREF PIX_IN[5240] NB2 NB1 CSA_VREF pixel
xPix5241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[52] VREF PIX_IN[5241] NB2 NB1 CSA_VREF pixel
xPix5242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[52] VREF PIX_IN[5242] NB2 NB1 CSA_VREF pixel
xPix5243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[52] VREF PIX_IN[5243] NB2 NB1 CSA_VREF pixel
xPix5244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[52] VREF PIX_IN[5244] NB2 NB1 CSA_VREF pixel
xPix5245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[52] VREF PIX_IN[5245] NB2 NB1 CSA_VREF pixel
xPix5246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[52] VREF PIX_IN[5246] NB2 NB1 CSA_VREF pixel
xPix5247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[52] VREF PIX_IN[5247] NB2 NB1 CSA_VREF pixel
xPix5248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[52] VREF PIX_IN[5248] NB2 NB1 CSA_VREF pixel
xPix5249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[52] VREF PIX_IN[5249] NB2 NB1 CSA_VREF pixel
xPix5250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[52] VREF PIX_IN[5250] NB2 NB1 CSA_VREF pixel
xPix5251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[52] VREF PIX_IN[5251] NB2 NB1 CSA_VREF pixel
xPix5252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[52] VREF PIX_IN[5252] NB2 NB1 CSA_VREF pixel
xPix5253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[52] VREF PIX_IN[5253] NB2 NB1 CSA_VREF pixel
xPix5254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[52] VREF PIX_IN[5254] NB2 NB1 CSA_VREF pixel
xPix5255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[52] VREF PIX_IN[5255] NB2 NB1 CSA_VREF pixel
xPix5256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[52] VREF PIX_IN[5256] NB2 NB1 CSA_VREF pixel
xPix5257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[52] VREF PIX_IN[5257] NB2 NB1 CSA_VREF pixel
xPix5258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[52] VREF PIX_IN[5258] NB2 NB1 CSA_VREF pixel
xPix5259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[52] VREF PIX_IN[5259] NB2 NB1 CSA_VREF pixel
xPix5260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[52] VREF PIX_IN[5260] NB2 NB1 CSA_VREF pixel
xPix5261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[52] VREF PIX_IN[5261] NB2 NB1 CSA_VREF pixel
xPix5262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[52] VREF PIX_IN[5262] NB2 NB1 CSA_VREF pixel
xPix5263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[52] VREF PIX_IN[5263] NB2 NB1 CSA_VREF pixel
xPix5264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[52] VREF PIX_IN[5264] NB2 NB1 CSA_VREF pixel
xPix5265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[52] VREF PIX_IN[5265] NB2 NB1 CSA_VREF pixel
xPix5266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[52] VREF PIX_IN[5266] NB2 NB1 CSA_VREF pixel
xPix5267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[52] VREF PIX_IN[5267] NB2 NB1 CSA_VREF pixel
xPix5268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[52] VREF PIX_IN[5268] NB2 NB1 CSA_VREF pixel
xPix5269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[52] VREF PIX_IN[5269] NB2 NB1 CSA_VREF pixel
xPix5270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[52] VREF PIX_IN[5270] NB2 NB1 CSA_VREF pixel
xPix5271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[52] VREF PIX_IN[5271] NB2 NB1 CSA_VREF pixel
xPix5272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[52] VREF PIX_IN[5272] NB2 NB1 CSA_VREF pixel
xPix5273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[52] VREF PIX_IN[5273] NB2 NB1 CSA_VREF pixel
xPix5274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[52] VREF PIX_IN[5274] NB2 NB1 CSA_VREF pixel
xPix5275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[52] VREF PIX_IN[5275] NB2 NB1 CSA_VREF pixel
xPix5276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[52] VREF PIX_IN[5276] NB2 NB1 CSA_VREF pixel
xPix5277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[52] VREF PIX_IN[5277] NB2 NB1 CSA_VREF pixel
xPix5278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[52] VREF PIX_IN[5278] NB2 NB1 CSA_VREF pixel
xPix5279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[52] VREF PIX_IN[5279] NB2 NB1 CSA_VREF pixel
xPix5280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[52] VREF PIX_IN[5280] NB2 NB1 CSA_VREF pixel
xPix5281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[52] VREF PIX_IN[5281] NB2 NB1 CSA_VREF pixel
xPix5282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[52] VREF PIX_IN[5282] NB2 NB1 CSA_VREF pixel
xPix5283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[52] VREF PIX_IN[5283] NB2 NB1 CSA_VREF pixel
xPix5284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[52] VREF PIX_IN[5284] NB2 NB1 CSA_VREF pixel
xPix5285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[52] VREF PIX_IN[5285] NB2 NB1 CSA_VREF pixel
xPix5286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[52] VREF PIX_IN[5286] NB2 NB1 CSA_VREF pixel
xPix5287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[52] VREF PIX_IN[5287] NB2 NB1 CSA_VREF pixel
xPix5288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[52] VREF PIX_IN[5288] NB2 NB1 CSA_VREF pixel
xPix5289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[52] VREF PIX_IN[5289] NB2 NB1 CSA_VREF pixel
xPix5290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[52] VREF PIX_IN[5290] NB2 NB1 CSA_VREF pixel
xPix5291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[52] VREF PIX_IN[5291] NB2 NB1 CSA_VREF pixel
xPix5292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[52] VREF PIX_IN[5292] NB2 NB1 CSA_VREF pixel
xPix5293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[52] VREF PIX_IN[5293] NB2 NB1 CSA_VREF pixel
xPix5294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[52] VREF PIX_IN[5294] NB2 NB1 CSA_VREF pixel
xPix5295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[52] VREF PIX_IN[5295] NB2 NB1 CSA_VREF pixel
xPix5296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[52] VREF PIX_IN[5296] NB2 NB1 CSA_VREF pixel
xPix5297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[52] VREF PIX_IN[5297] NB2 NB1 CSA_VREF pixel
xPix5298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[52] VREF PIX_IN[5298] NB2 NB1 CSA_VREF pixel
xPix5299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[52] VREF PIX_IN[5299] NB2 NB1 CSA_VREF pixel
xPix5300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[53] VREF PIX_IN[5300] NB2 NB1 CSA_VREF pixel
xPix5301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[53] VREF PIX_IN[5301] NB2 NB1 CSA_VREF pixel
xPix5302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[53] VREF PIX_IN[5302] NB2 NB1 CSA_VREF pixel
xPix5303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[53] VREF PIX_IN[5303] NB2 NB1 CSA_VREF pixel
xPix5304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[53] VREF PIX_IN[5304] NB2 NB1 CSA_VREF pixel
xPix5305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[53] VREF PIX_IN[5305] NB2 NB1 CSA_VREF pixel
xPix5306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[53] VREF PIX_IN[5306] NB2 NB1 CSA_VREF pixel
xPix5307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[53] VREF PIX_IN[5307] NB2 NB1 CSA_VREF pixel
xPix5308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[53] VREF PIX_IN[5308] NB2 NB1 CSA_VREF pixel
xPix5309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[53] VREF PIX_IN[5309] NB2 NB1 CSA_VREF pixel
xPix5310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[53] VREF PIX_IN[5310] NB2 NB1 CSA_VREF pixel
xPix5311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[53] VREF PIX_IN[5311] NB2 NB1 CSA_VREF pixel
xPix5312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[53] VREF PIX_IN[5312] NB2 NB1 CSA_VREF pixel
xPix5313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[53] VREF PIX_IN[5313] NB2 NB1 CSA_VREF pixel
xPix5314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[53] VREF PIX_IN[5314] NB2 NB1 CSA_VREF pixel
xPix5315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[53] VREF PIX_IN[5315] NB2 NB1 CSA_VREF pixel
xPix5316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[53] VREF PIX_IN[5316] NB2 NB1 CSA_VREF pixel
xPix5317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[53] VREF PIX_IN[5317] NB2 NB1 CSA_VREF pixel
xPix5318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[53] VREF PIX_IN[5318] NB2 NB1 CSA_VREF pixel
xPix5319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[53] VREF PIX_IN[5319] NB2 NB1 CSA_VREF pixel
xPix5320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[53] VREF PIX_IN[5320] NB2 NB1 CSA_VREF pixel
xPix5321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[53] VREF PIX_IN[5321] NB2 NB1 CSA_VREF pixel
xPix5322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[53] VREF PIX_IN[5322] NB2 NB1 CSA_VREF pixel
xPix5323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[53] VREF PIX_IN[5323] NB2 NB1 CSA_VREF pixel
xPix5324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[53] VREF PIX_IN[5324] NB2 NB1 CSA_VREF pixel
xPix5325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[53] VREF PIX_IN[5325] NB2 NB1 CSA_VREF pixel
xPix5326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[53] VREF PIX_IN[5326] NB2 NB1 CSA_VREF pixel
xPix5327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[53] VREF PIX_IN[5327] NB2 NB1 CSA_VREF pixel
xPix5328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[53] VREF PIX_IN[5328] NB2 NB1 CSA_VREF pixel
xPix5329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[53] VREF PIX_IN[5329] NB2 NB1 CSA_VREF pixel
xPix5330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[53] VREF PIX_IN[5330] NB2 NB1 CSA_VREF pixel
xPix5331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[53] VREF PIX_IN[5331] NB2 NB1 CSA_VREF pixel
xPix5332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[53] VREF PIX_IN[5332] NB2 NB1 CSA_VREF pixel
xPix5333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[53] VREF PIX_IN[5333] NB2 NB1 CSA_VREF pixel
xPix5334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[53] VREF PIX_IN[5334] NB2 NB1 CSA_VREF pixel
xPix5335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[53] VREF PIX_IN[5335] NB2 NB1 CSA_VREF pixel
xPix5336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[53] VREF PIX_IN[5336] NB2 NB1 CSA_VREF pixel
xPix5337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[53] VREF PIX_IN[5337] NB2 NB1 CSA_VREF pixel
xPix5338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[53] VREF PIX_IN[5338] NB2 NB1 CSA_VREF pixel
xPix5339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[53] VREF PIX_IN[5339] NB2 NB1 CSA_VREF pixel
xPix5340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[53] VREF PIX_IN[5340] NB2 NB1 CSA_VREF pixel
xPix5341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[53] VREF PIX_IN[5341] NB2 NB1 CSA_VREF pixel
xPix5342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[53] VREF PIX_IN[5342] NB2 NB1 CSA_VREF pixel
xPix5343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[53] VREF PIX_IN[5343] NB2 NB1 CSA_VREF pixel
xPix5344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[53] VREF PIX_IN[5344] NB2 NB1 CSA_VREF pixel
xPix5345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[53] VREF PIX_IN[5345] NB2 NB1 CSA_VREF pixel
xPix5346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[53] VREF PIX_IN[5346] NB2 NB1 CSA_VREF pixel
xPix5347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[53] VREF PIX_IN[5347] NB2 NB1 CSA_VREF pixel
xPix5348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[53] VREF PIX_IN[5348] NB2 NB1 CSA_VREF pixel
xPix5349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[53] VREF PIX_IN[5349] NB2 NB1 CSA_VREF pixel
xPix5350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[53] VREF PIX_IN[5350] NB2 NB1 CSA_VREF pixel
xPix5351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[53] VREF PIX_IN[5351] NB2 NB1 CSA_VREF pixel
xPix5352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[53] VREF PIX_IN[5352] NB2 NB1 CSA_VREF pixel
xPix5353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[53] VREF PIX_IN[5353] NB2 NB1 CSA_VREF pixel
xPix5354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[53] VREF PIX_IN[5354] NB2 NB1 CSA_VREF pixel
xPix5355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[53] VREF PIX_IN[5355] NB2 NB1 CSA_VREF pixel
xPix5356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[53] VREF PIX_IN[5356] NB2 NB1 CSA_VREF pixel
xPix5357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[53] VREF PIX_IN[5357] NB2 NB1 CSA_VREF pixel
xPix5358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[53] VREF PIX_IN[5358] NB2 NB1 CSA_VREF pixel
xPix5359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[53] VREF PIX_IN[5359] NB2 NB1 CSA_VREF pixel
xPix5360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[53] VREF PIX_IN[5360] NB2 NB1 CSA_VREF pixel
xPix5361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[53] VREF PIX_IN[5361] NB2 NB1 CSA_VREF pixel
xPix5362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[53] VREF PIX_IN[5362] NB2 NB1 CSA_VREF pixel
xPix5363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[53] VREF PIX_IN[5363] NB2 NB1 CSA_VREF pixel
xPix5364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[53] VREF PIX_IN[5364] NB2 NB1 CSA_VREF pixel
xPix5365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[53] VREF PIX_IN[5365] NB2 NB1 CSA_VREF pixel
xPix5366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[53] VREF PIX_IN[5366] NB2 NB1 CSA_VREF pixel
xPix5367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[53] VREF PIX_IN[5367] NB2 NB1 CSA_VREF pixel
xPix5368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[53] VREF PIX_IN[5368] NB2 NB1 CSA_VREF pixel
xPix5369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[53] VREF PIX_IN[5369] NB2 NB1 CSA_VREF pixel
xPix5370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[53] VREF PIX_IN[5370] NB2 NB1 CSA_VREF pixel
xPix5371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[53] VREF PIX_IN[5371] NB2 NB1 CSA_VREF pixel
xPix5372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[53] VREF PIX_IN[5372] NB2 NB1 CSA_VREF pixel
xPix5373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[53] VREF PIX_IN[5373] NB2 NB1 CSA_VREF pixel
xPix5374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[53] VREF PIX_IN[5374] NB2 NB1 CSA_VREF pixel
xPix5375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[53] VREF PIX_IN[5375] NB2 NB1 CSA_VREF pixel
xPix5376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[53] VREF PIX_IN[5376] NB2 NB1 CSA_VREF pixel
xPix5377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[53] VREF PIX_IN[5377] NB2 NB1 CSA_VREF pixel
xPix5378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[53] VREF PIX_IN[5378] NB2 NB1 CSA_VREF pixel
xPix5379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[53] VREF PIX_IN[5379] NB2 NB1 CSA_VREF pixel
xPix5380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[53] VREF PIX_IN[5380] NB2 NB1 CSA_VREF pixel
xPix5381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[53] VREF PIX_IN[5381] NB2 NB1 CSA_VREF pixel
xPix5382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[53] VREF PIX_IN[5382] NB2 NB1 CSA_VREF pixel
xPix5383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[53] VREF PIX_IN[5383] NB2 NB1 CSA_VREF pixel
xPix5384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[53] VREF PIX_IN[5384] NB2 NB1 CSA_VREF pixel
xPix5385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[53] VREF PIX_IN[5385] NB2 NB1 CSA_VREF pixel
xPix5386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[53] VREF PIX_IN[5386] NB2 NB1 CSA_VREF pixel
xPix5387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[53] VREF PIX_IN[5387] NB2 NB1 CSA_VREF pixel
xPix5388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[53] VREF PIX_IN[5388] NB2 NB1 CSA_VREF pixel
xPix5389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[53] VREF PIX_IN[5389] NB2 NB1 CSA_VREF pixel
xPix5390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[53] VREF PIX_IN[5390] NB2 NB1 CSA_VREF pixel
xPix5391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[53] VREF PIX_IN[5391] NB2 NB1 CSA_VREF pixel
xPix5392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[53] VREF PIX_IN[5392] NB2 NB1 CSA_VREF pixel
xPix5393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[53] VREF PIX_IN[5393] NB2 NB1 CSA_VREF pixel
xPix5394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[53] VREF PIX_IN[5394] NB2 NB1 CSA_VREF pixel
xPix5395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[53] VREF PIX_IN[5395] NB2 NB1 CSA_VREF pixel
xPix5396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[53] VREF PIX_IN[5396] NB2 NB1 CSA_VREF pixel
xPix5397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[53] VREF PIX_IN[5397] NB2 NB1 CSA_VREF pixel
xPix5398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[53] VREF PIX_IN[5398] NB2 NB1 CSA_VREF pixel
xPix5399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[53] VREF PIX_IN[5399] NB2 NB1 CSA_VREF pixel
xPix5400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[54] VREF PIX_IN[5400] NB2 NB1 CSA_VREF pixel
xPix5401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[54] VREF PIX_IN[5401] NB2 NB1 CSA_VREF pixel
xPix5402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[54] VREF PIX_IN[5402] NB2 NB1 CSA_VREF pixel
xPix5403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[54] VREF PIX_IN[5403] NB2 NB1 CSA_VREF pixel
xPix5404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[54] VREF PIX_IN[5404] NB2 NB1 CSA_VREF pixel
xPix5405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[54] VREF PIX_IN[5405] NB2 NB1 CSA_VREF pixel
xPix5406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[54] VREF PIX_IN[5406] NB2 NB1 CSA_VREF pixel
xPix5407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[54] VREF PIX_IN[5407] NB2 NB1 CSA_VREF pixel
xPix5408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[54] VREF PIX_IN[5408] NB2 NB1 CSA_VREF pixel
xPix5409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[54] VREF PIX_IN[5409] NB2 NB1 CSA_VREF pixel
xPix5410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[54] VREF PIX_IN[5410] NB2 NB1 CSA_VREF pixel
xPix5411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[54] VREF PIX_IN[5411] NB2 NB1 CSA_VREF pixel
xPix5412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[54] VREF PIX_IN[5412] NB2 NB1 CSA_VREF pixel
xPix5413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[54] VREF PIX_IN[5413] NB2 NB1 CSA_VREF pixel
xPix5414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[54] VREF PIX_IN[5414] NB2 NB1 CSA_VREF pixel
xPix5415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[54] VREF PIX_IN[5415] NB2 NB1 CSA_VREF pixel
xPix5416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[54] VREF PIX_IN[5416] NB2 NB1 CSA_VREF pixel
xPix5417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[54] VREF PIX_IN[5417] NB2 NB1 CSA_VREF pixel
xPix5418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[54] VREF PIX_IN[5418] NB2 NB1 CSA_VREF pixel
xPix5419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[54] VREF PIX_IN[5419] NB2 NB1 CSA_VREF pixel
xPix5420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[54] VREF PIX_IN[5420] NB2 NB1 CSA_VREF pixel
xPix5421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[54] VREF PIX_IN[5421] NB2 NB1 CSA_VREF pixel
xPix5422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[54] VREF PIX_IN[5422] NB2 NB1 CSA_VREF pixel
xPix5423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[54] VREF PIX_IN[5423] NB2 NB1 CSA_VREF pixel
xPix5424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[54] VREF PIX_IN[5424] NB2 NB1 CSA_VREF pixel
xPix5425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[54] VREF PIX_IN[5425] NB2 NB1 CSA_VREF pixel
xPix5426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[54] VREF PIX_IN[5426] NB2 NB1 CSA_VREF pixel
xPix5427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[54] VREF PIX_IN[5427] NB2 NB1 CSA_VREF pixel
xPix5428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[54] VREF PIX_IN[5428] NB2 NB1 CSA_VREF pixel
xPix5429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[54] VREF PIX_IN[5429] NB2 NB1 CSA_VREF pixel
xPix5430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[54] VREF PIX_IN[5430] NB2 NB1 CSA_VREF pixel
xPix5431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[54] VREF PIX_IN[5431] NB2 NB1 CSA_VREF pixel
xPix5432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[54] VREF PIX_IN[5432] NB2 NB1 CSA_VREF pixel
xPix5433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[54] VREF PIX_IN[5433] NB2 NB1 CSA_VREF pixel
xPix5434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[54] VREF PIX_IN[5434] NB2 NB1 CSA_VREF pixel
xPix5435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[54] VREF PIX_IN[5435] NB2 NB1 CSA_VREF pixel
xPix5436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[54] VREF PIX_IN[5436] NB2 NB1 CSA_VREF pixel
xPix5437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[54] VREF PIX_IN[5437] NB2 NB1 CSA_VREF pixel
xPix5438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[54] VREF PIX_IN[5438] NB2 NB1 CSA_VREF pixel
xPix5439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[54] VREF PIX_IN[5439] NB2 NB1 CSA_VREF pixel
xPix5440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[54] VREF PIX_IN[5440] NB2 NB1 CSA_VREF pixel
xPix5441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[54] VREF PIX_IN[5441] NB2 NB1 CSA_VREF pixel
xPix5442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[54] VREF PIX_IN[5442] NB2 NB1 CSA_VREF pixel
xPix5443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[54] VREF PIX_IN[5443] NB2 NB1 CSA_VREF pixel
xPix5444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[54] VREF PIX_IN[5444] NB2 NB1 CSA_VREF pixel
xPix5445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[54] VREF PIX_IN[5445] NB2 NB1 CSA_VREF pixel
xPix5446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[54] VREF PIX_IN[5446] NB2 NB1 CSA_VREF pixel
xPix5447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[54] VREF PIX_IN[5447] NB2 NB1 CSA_VREF pixel
xPix5448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[54] VREF PIX_IN[5448] NB2 NB1 CSA_VREF pixel
xPix5449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[54] VREF PIX_IN[5449] NB2 NB1 CSA_VREF pixel
xPix5450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[54] VREF PIX_IN[5450] NB2 NB1 CSA_VREF pixel
xPix5451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[54] VREF PIX_IN[5451] NB2 NB1 CSA_VREF pixel
xPix5452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[54] VREF PIX_IN[5452] NB2 NB1 CSA_VREF pixel
xPix5453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[54] VREF PIX_IN[5453] NB2 NB1 CSA_VREF pixel
xPix5454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[54] VREF PIX_IN[5454] NB2 NB1 CSA_VREF pixel
xPix5455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[54] VREF PIX_IN[5455] NB2 NB1 CSA_VREF pixel
xPix5456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[54] VREF PIX_IN[5456] NB2 NB1 CSA_VREF pixel
xPix5457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[54] VREF PIX_IN[5457] NB2 NB1 CSA_VREF pixel
xPix5458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[54] VREF PIX_IN[5458] NB2 NB1 CSA_VREF pixel
xPix5459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[54] VREF PIX_IN[5459] NB2 NB1 CSA_VREF pixel
xPix5460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[54] VREF PIX_IN[5460] NB2 NB1 CSA_VREF pixel
xPix5461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[54] VREF PIX_IN[5461] NB2 NB1 CSA_VREF pixel
xPix5462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[54] VREF PIX_IN[5462] NB2 NB1 CSA_VREF pixel
xPix5463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[54] VREF PIX_IN[5463] NB2 NB1 CSA_VREF pixel
xPix5464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[54] VREF PIX_IN[5464] NB2 NB1 CSA_VREF pixel
xPix5465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[54] VREF PIX_IN[5465] NB2 NB1 CSA_VREF pixel
xPix5466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[54] VREF PIX_IN[5466] NB2 NB1 CSA_VREF pixel
xPix5467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[54] VREF PIX_IN[5467] NB2 NB1 CSA_VREF pixel
xPix5468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[54] VREF PIX_IN[5468] NB2 NB1 CSA_VREF pixel
xPix5469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[54] VREF PIX_IN[5469] NB2 NB1 CSA_VREF pixel
xPix5470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[54] VREF PIX_IN[5470] NB2 NB1 CSA_VREF pixel
xPix5471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[54] VREF PIX_IN[5471] NB2 NB1 CSA_VREF pixel
xPix5472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[54] VREF PIX_IN[5472] NB2 NB1 CSA_VREF pixel
xPix5473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[54] VREF PIX_IN[5473] NB2 NB1 CSA_VREF pixel
xPix5474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[54] VREF PIX_IN[5474] NB2 NB1 CSA_VREF pixel
xPix5475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[54] VREF PIX_IN[5475] NB2 NB1 CSA_VREF pixel
xPix5476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[54] VREF PIX_IN[5476] NB2 NB1 CSA_VREF pixel
xPix5477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[54] VREF PIX_IN[5477] NB2 NB1 CSA_VREF pixel
xPix5478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[54] VREF PIX_IN[5478] NB2 NB1 CSA_VREF pixel
xPix5479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[54] VREF PIX_IN[5479] NB2 NB1 CSA_VREF pixel
xPix5480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[54] VREF PIX_IN[5480] NB2 NB1 CSA_VREF pixel
xPix5481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[54] VREF PIX_IN[5481] NB2 NB1 CSA_VREF pixel
xPix5482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[54] VREF PIX_IN[5482] NB2 NB1 CSA_VREF pixel
xPix5483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[54] VREF PIX_IN[5483] NB2 NB1 CSA_VREF pixel
xPix5484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[54] VREF PIX_IN[5484] NB2 NB1 CSA_VREF pixel
xPix5485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[54] VREF PIX_IN[5485] NB2 NB1 CSA_VREF pixel
xPix5486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[54] VREF PIX_IN[5486] NB2 NB1 CSA_VREF pixel
xPix5487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[54] VREF PIX_IN[5487] NB2 NB1 CSA_VREF pixel
xPix5488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[54] VREF PIX_IN[5488] NB2 NB1 CSA_VREF pixel
xPix5489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[54] VREF PIX_IN[5489] NB2 NB1 CSA_VREF pixel
xPix5490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[54] VREF PIX_IN[5490] NB2 NB1 CSA_VREF pixel
xPix5491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[54] VREF PIX_IN[5491] NB2 NB1 CSA_VREF pixel
xPix5492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[54] VREF PIX_IN[5492] NB2 NB1 CSA_VREF pixel
xPix5493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[54] VREF PIX_IN[5493] NB2 NB1 CSA_VREF pixel
xPix5494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[54] VREF PIX_IN[5494] NB2 NB1 CSA_VREF pixel
xPix5495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[54] VREF PIX_IN[5495] NB2 NB1 CSA_VREF pixel
xPix5496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[54] VREF PIX_IN[5496] NB2 NB1 CSA_VREF pixel
xPix5497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[54] VREF PIX_IN[5497] NB2 NB1 CSA_VREF pixel
xPix5498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[54] VREF PIX_IN[5498] NB2 NB1 CSA_VREF pixel
xPix5499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[54] VREF PIX_IN[5499] NB2 NB1 CSA_VREF pixel
xPix5500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[55] VREF PIX_IN[5500] NB2 NB1 CSA_VREF pixel
xPix5501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[55] VREF PIX_IN[5501] NB2 NB1 CSA_VREF pixel
xPix5502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[55] VREF PIX_IN[5502] NB2 NB1 CSA_VREF pixel
xPix5503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[55] VREF PIX_IN[5503] NB2 NB1 CSA_VREF pixel
xPix5504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[55] VREF PIX_IN[5504] NB2 NB1 CSA_VREF pixel
xPix5505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[55] VREF PIX_IN[5505] NB2 NB1 CSA_VREF pixel
xPix5506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[55] VREF PIX_IN[5506] NB2 NB1 CSA_VREF pixel
xPix5507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[55] VREF PIX_IN[5507] NB2 NB1 CSA_VREF pixel
xPix5508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[55] VREF PIX_IN[5508] NB2 NB1 CSA_VREF pixel
xPix5509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[55] VREF PIX_IN[5509] NB2 NB1 CSA_VREF pixel
xPix5510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[55] VREF PIX_IN[5510] NB2 NB1 CSA_VREF pixel
xPix5511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[55] VREF PIX_IN[5511] NB2 NB1 CSA_VREF pixel
xPix5512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[55] VREF PIX_IN[5512] NB2 NB1 CSA_VREF pixel
xPix5513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[55] VREF PIX_IN[5513] NB2 NB1 CSA_VREF pixel
xPix5514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[55] VREF PIX_IN[5514] NB2 NB1 CSA_VREF pixel
xPix5515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[55] VREF PIX_IN[5515] NB2 NB1 CSA_VREF pixel
xPix5516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[55] VREF PIX_IN[5516] NB2 NB1 CSA_VREF pixel
xPix5517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[55] VREF PIX_IN[5517] NB2 NB1 CSA_VREF pixel
xPix5518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[55] VREF PIX_IN[5518] NB2 NB1 CSA_VREF pixel
xPix5519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[55] VREF PIX_IN[5519] NB2 NB1 CSA_VREF pixel
xPix5520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[55] VREF PIX_IN[5520] NB2 NB1 CSA_VREF pixel
xPix5521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[55] VREF PIX_IN[5521] NB2 NB1 CSA_VREF pixel
xPix5522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[55] VREF PIX_IN[5522] NB2 NB1 CSA_VREF pixel
xPix5523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[55] VREF PIX_IN[5523] NB2 NB1 CSA_VREF pixel
xPix5524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[55] VREF PIX_IN[5524] NB2 NB1 CSA_VREF pixel
xPix5525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[55] VREF PIX_IN[5525] NB2 NB1 CSA_VREF pixel
xPix5526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[55] VREF PIX_IN[5526] NB2 NB1 CSA_VREF pixel
xPix5527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[55] VREF PIX_IN[5527] NB2 NB1 CSA_VREF pixel
xPix5528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[55] VREF PIX_IN[5528] NB2 NB1 CSA_VREF pixel
xPix5529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[55] VREF PIX_IN[5529] NB2 NB1 CSA_VREF pixel
xPix5530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[55] VREF PIX_IN[5530] NB2 NB1 CSA_VREF pixel
xPix5531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[55] VREF PIX_IN[5531] NB2 NB1 CSA_VREF pixel
xPix5532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[55] VREF PIX_IN[5532] NB2 NB1 CSA_VREF pixel
xPix5533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[55] VREF PIX_IN[5533] NB2 NB1 CSA_VREF pixel
xPix5534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[55] VREF PIX_IN[5534] NB2 NB1 CSA_VREF pixel
xPix5535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[55] VREF PIX_IN[5535] NB2 NB1 CSA_VREF pixel
xPix5536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[55] VREF PIX_IN[5536] NB2 NB1 CSA_VREF pixel
xPix5537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[55] VREF PIX_IN[5537] NB2 NB1 CSA_VREF pixel
xPix5538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[55] VREF PIX_IN[5538] NB2 NB1 CSA_VREF pixel
xPix5539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[55] VREF PIX_IN[5539] NB2 NB1 CSA_VREF pixel
xPix5540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[55] VREF PIX_IN[5540] NB2 NB1 CSA_VREF pixel
xPix5541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[55] VREF PIX_IN[5541] NB2 NB1 CSA_VREF pixel
xPix5542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[55] VREF PIX_IN[5542] NB2 NB1 CSA_VREF pixel
xPix5543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[55] VREF PIX_IN[5543] NB2 NB1 CSA_VREF pixel
xPix5544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[55] VREF PIX_IN[5544] NB2 NB1 CSA_VREF pixel
xPix5545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[55] VREF PIX_IN[5545] NB2 NB1 CSA_VREF pixel
xPix5546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[55] VREF PIX_IN[5546] NB2 NB1 CSA_VREF pixel
xPix5547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[55] VREF PIX_IN[5547] NB2 NB1 CSA_VREF pixel
xPix5548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[55] VREF PIX_IN[5548] NB2 NB1 CSA_VREF pixel
xPix5549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[55] VREF PIX_IN[5549] NB2 NB1 CSA_VREF pixel
xPix5550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[55] VREF PIX_IN[5550] NB2 NB1 CSA_VREF pixel
xPix5551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[55] VREF PIX_IN[5551] NB2 NB1 CSA_VREF pixel
xPix5552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[55] VREF PIX_IN[5552] NB2 NB1 CSA_VREF pixel
xPix5553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[55] VREF PIX_IN[5553] NB2 NB1 CSA_VREF pixel
xPix5554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[55] VREF PIX_IN[5554] NB2 NB1 CSA_VREF pixel
xPix5555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[55] VREF PIX_IN[5555] NB2 NB1 CSA_VREF pixel
xPix5556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[55] VREF PIX_IN[5556] NB2 NB1 CSA_VREF pixel
xPix5557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[55] VREF PIX_IN[5557] NB2 NB1 CSA_VREF pixel
xPix5558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[55] VREF PIX_IN[5558] NB2 NB1 CSA_VREF pixel
xPix5559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[55] VREF PIX_IN[5559] NB2 NB1 CSA_VREF pixel
xPix5560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[55] VREF PIX_IN[5560] NB2 NB1 CSA_VREF pixel
xPix5561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[55] VREF PIX_IN[5561] NB2 NB1 CSA_VREF pixel
xPix5562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[55] VREF PIX_IN[5562] NB2 NB1 CSA_VREF pixel
xPix5563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[55] VREF PIX_IN[5563] NB2 NB1 CSA_VREF pixel
xPix5564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[55] VREF PIX_IN[5564] NB2 NB1 CSA_VREF pixel
xPix5565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[55] VREF PIX_IN[5565] NB2 NB1 CSA_VREF pixel
xPix5566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[55] VREF PIX_IN[5566] NB2 NB1 CSA_VREF pixel
xPix5567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[55] VREF PIX_IN[5567] NB2 NB1 CSA_VREF pixel
xPix5568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[55] VREF PIX_IN[5568] NB2 NB1 CSA_VREF pixel
xPix5569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[55] VREF PIX_IN[5569] NB2 NB1 CSA_VREF pixel
xPix5570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[55] VREF PIX_IN[5570] NB2 NB1 CSA_VREF pixel
xPix5571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[55] VREF PIX_IN[5571] NB2 NB1 CSA_VREF pixel
xPix5572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[55] VREF PIX_IN[5572] NB2 NB1 CSA_VREF pixel
xPix5573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[55] VREF PIX_IN[5573] NB2 NB1 CSA_VREF pixel
xPix5574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[55] VREF PIX_IN[5574] NB2 NB1 CSA_VREF pixel
xPix5575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[55] VREF PIX_IN[5575] NB2 NB1 CSA_VREF pixel
xPix5576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[55] VREF PIX_IN[5576] NB2 NB1 CSA_VREF pixel
xPix5577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[55] VREF PIX_IN[5577] NB2 NB1 CSA_VREF pixel
xPix5578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[55] VREF PIX_IN[5578] NB2 NB1 CSA_VREF pixel
xPix5579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[55] VREF PIX_IN[5579] NB2 NB1 CSA_VREF pixel
xPix5580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[55] VREF PIX_IN[5580] NB2 NB1 CSA_VREF pixel
xPix5581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[55] VREF PIX_IN[5581] NB2 NB1 CSA_VREF pixel
xPix5582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[55] VREF PIX_IN[5582] NB2 NB1 CSA_VREF pixel
xPix5583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[55] VREF PIX_IN[5583] NB2 NB1 CSA_VREF pixel
xPix5584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[55] VREF PIX_IN[5584] NB2 NB1 CSA_VREF pixel
xPix5585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[55] VREF PIX_IN[5585] NB2 NB1 CSA_VREF pixel
xPix5586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[55] VREF PIX_IN[5586] NB2 NB1 CSA_VREF pixel
xPix5587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[55] VREF PIX_IN[5587] NB2 NB1 CSA_VREF pixel
xPix5588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[55] VREF PIX_IN[5588] NB2 NB1 CSA_VREF pixel
xPix5589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[55] VREF PIX_IN[5589] NB2 NB1 CSA_VREF pixel
xPix5590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[55] VREF PIX_IN[5590] NB2 NB1 CSA_VREF pixel
xPix5591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[55] VREF PIX_IN[5591] NB2 NB1 CSA_VREF pixel
xPix5592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[55] VREF PIX_IN[5592] NB2 NB1 CSA_VREF pixel
xPix5593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[55] VREF PIX_IN[5593] NB2 NB1 CSA_VREF pixel
xPix5594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[55] VREF PIX_IN[5594] NB2 NB1 CSA_VREF pixel
xPix5595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[55] VREF PIX_IN[5595] NB2 NB1 CSA_VREF pixel
xPix5596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[55] VREF PIX_IN[5596] NB2 NB1 CSA_VREF pixel
xPix5597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[55] VREF PIX_IN[5597] NB2 NB1 CSA_VREF pixel
xPix5598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[55] VREF PIX_IN[5598] NB2 NB1 CSA_VREF pixel
xPix5599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[55] VREF PIX_IN[5599] NB2 NB1 CSA_VREF pixel
xPix5600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[56] VREF PIX_IN[5600] NB2 NB1 CSA_VREF pixel
xPix5601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[56] VREF PIX_IN[5601] NB2 NB1 CSA_VREF pixel
xPix5602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[56] VREF PIX_IN[5602] NB2 NB1 CSA_VREF pixel
xPix5603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[56] VREF PIX_IN[5603] NB2 NB1 CSA_VREF pixel
xPix5604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[56] VREF PIX_IN[5604] NB2 NB1 CSA_VREF pixel
xPix5605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[56] VREF PIX_IN[5605] NB2 NB1 CSA_VREF pixel
xPix5606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[56] VREF PIX_IN[5606] NB2 NB1 CSA_VREF pixel
xPix5607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[56] VREF PIX_IN[5607] NB2 NB1 CSA_VREF pixel
xPix5608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[56] VREF PIX_IN[5608] NB2 NB1 CSA_VREF pixel
xPix5609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[56] VREF PIX_IN[5609] NB2 NB1 CSA_VREF pixel
xPix5610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[56] VREF PIX_IN[5610] NB2 NB1 CSA_VREF pixel
xPix5611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[56] VREF PIX_IN[5611] NB2 NB1 CSA_VREF pixel
xPix5612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[56] VREF PIX_IN[5612] NB2 NB1 CSA_VREF pixel
xPix5613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[56] VREF PIX_IN[5613] NB2 NB1 CSA_VREF pixel
xPix5614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[56] VREF PIX_IN[5614] NB2 NB1 CSA_VREF pixel
xPix5615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[56] VREF PIX_IN[5615] NB2 NB1 CSA_VREF pixel
xPix5616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[56] VREF PIX_IN[5616] NB2 NB1 CSA_VREF pixel
xPix5617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[56] VREF PIX_IN[5617] NB2 NB1 CSA_VREF pixel
xPix5618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[56] VREF PIX_IN[5618] NB2 NB1 CSA_VREF pixel
xPix5619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[56] VREF PIX_IN[5619] NB2 NB1 CSA_VREF pixel
xPix5620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[56] VREF PIX_IN[5620] NB2 NB1 CSA_VREF pixel
xPix5621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[56] VREF PIX_IN[5621] NB2 NB1 CSA_VREF pixel
xPix5622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[56] VREF PIX_IN[5622] NB2 NB1 CSA_VREF pixel
xPix5623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[56] VREF PIX_IN[5623] NB2 NB1 CSA_VREF pixel
xPix5624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[56] VREF PIX_IN[5624] NB2 NB1 CSA_VREF pixel
xPix5625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[56] VREF PIX_IN[5625] NB2 NB1 CSA_VREF pixel
xPix5626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[56] VREF PIX_IN[5626] NB2 NB1 CSA_VREF pixel
xPix5627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[56] VREF PIX_IN[5627] NB2 NB1 CSA_VREF pixel
xPix5628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[56] VREF PIX_IN[5628] NB2 NB1 CSA_VREF pixel
xPix5629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[56] VREF PIX_IN[5629] NB2 NB1 CSA_VREF pixel
xPix5630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[56] VREF PIX_IN[5630] NB2 NB1 CSA_VREF pixel
xPix5631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[56] VREF PIX_IN[5631] NB2 NB1 CSA_VREF pixel
xPix5632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[56] VREF PIX_IN[5632] NB2 NB1 CSA_VREF pixel
xPix5633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[56] VREF PIX_IN[5633] NB2 NB1 CSA_VREF pixel
xPix5634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[56] VREF PIX_IN[5634] NB2 NB1 CSA_VREF pixel
xPix5635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[56] VREF PIX_IN[5635] NB2 NB1 CSA_VREF pixel
xPix5636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[56] VREF PIX_IN[5636] NB2 NB1 CSA_VREF pixel
xPix5637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[56] VREF PIX_IN[5637] NB2 NB1 CSA_VREF pixel
xPix5638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[56] VREF PIX_IN[5638] NB2 NB1 CSA_VREF pixel
xPix5639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[56] VREF PIX_IN[5639] NB2 NB1 CSA_VREF pixel
xPix5640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[56] VREF PIX_IN[5640] NB2 NB1 CSA_VREF pixel
xPix5641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[56] VREF PIX_IN[5641] NB2 NB1 CSA_VREF pixel
xPix5642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[56] VREF PIX_IN[5642] NB2 NB1 CSA_VREF pixel
xPix5643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[56] VREF PIX_IN[5643] NB2 NB1 CSA_VREF pixel
xPix5644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[56] VREF PIX_IN[5644] NB2 NB1 CSA_VREF pixel
xPix5645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[56] VREF PIX_IN[5645] NB2 NB1 CSA_VREF pixel
xPix5646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[56] VREF PIX_IN[5646] NB2 NB1 CSA_VREF pixel
xPix5647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[56] VREF PIX_IN[5647] NB2 NB1 CSA_VREF pixel
xPix5648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[56] VREF PIX_IN[5648] NB2 NB1 CSA_VREF pixel
xPix5649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[56] VREF PIX_IN[5649] NB2 NB1 CSA_VREF pixel
xPix5650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[56] VREF PIX_IN[5650] NB2 NB1 CSA_VREF pixel
xPix5651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[56] VREF PIX_IN[5651] NB2 NB1 CSA_VREF pixel
xPix5652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[56] VREF PIX_IN[5652] NB2 NB1 CSA_VREF pixel
xPix5653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[56] VREF PIX_IN[5653] NB2 NB1 CSA_VREF pixel
xPix5654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[56] VREF PIX_IN[5654] NB2 NB1 CSA_VREF pixel
xPix5655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[56] VREF PIX_IN[5655] NB2 NB1 CSA_VREF pixel
xPix5656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[56] VREF PIX_IN[5656] NB2 NB1 CSA_VREF pixel
xPix5657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[56] VREF PIX_IN[5657] NB2 NB1 CSA_VREF pixel
xPix5658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[56] VREF PIX_IN[5658] NB2 NB1 CSA_VREF pixel
xPix5659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[56] VREF PIX_IN[5659] NB2 NB1 CSA_VREF pixel
xPix5660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[56] VREF PIX_IN[5660] NB2 NB1 CSA_VREF pixel
xPix5661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[56] VREF PIX_IN[5661] NB2 NB1 CSA_VREF pixel
xPix5662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[56] VREF PIX_IN[5662] NB2 NB1 CSA_VREF pixel
xPix5663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[56] VREF PIX_IN[5663] NB2 NB1 CSA_VREF pixel
xPix5664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[56] VREF PIX_IN[5664] NB2 NB1 CSA_VREF pixel
xPix5665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[56] VREF PIX_IN[5665] NB2 NB1 CSA_VREF pixel
xPix5666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[56] VREF PIX_IN[5666] NB2 NB1 CSA_VREF pixel
xPix5667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[56] VREF PIX_IN[5667] NB2 NB1 CSA_VREF pixel
xPix5668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[56] VREF PIX_IN[5668] NB2 NB1 CSA_VREF pixel
xPix5669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[56] VREF PIX_IN[5669] NB2 NB1 CSA_VREF pixel
xPix5670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[56] VREF PIX_IN[5670] NB2 NB1 CSA_VREF pixel
xPix5671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[56] VREF PIX_IN[5671] NB2 NB1 CSA_VREF pixel
xPix5672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[56] VREF PIX_IN[5672] NB2 NB1 CSA_VREF pixel
xPix5673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[56] VREF PIX_IN[5673] NB2 NB1 CSA_VREF pixel
xPix5674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[56] VREF PIX_IN[5674] NB2 NB1 CSA_VREF pixel
xPix5675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[56] VREF PIX_IN[5675] NB2 NB1 CSA_VREF pixel
xPix5676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[56] VREF PIX_IN[5676] NB2 NB1 CSA_VREF pixel
xPix5677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[56] VREF PIX_IN[5677] NB2 NB1 CSA_VREF pixel
xPix5678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[56] VREF PIX_IN[5678] NB2 NB1 CSA_VREF pixel
xPix5679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[56] VREF PIX_IN[5679] NB2 NB1 CSA_VREF pixel
xPix5680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[56] VREF PIX_IN[5680] NB2 NB1 CSA_VREF pixel
xPix5681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[56] VREF PIX_IN[5681] NB2 NB1 CSA_VREF pixel
xPix5682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[56] VREF PIX_IN[5682] NB2 NB1 CSA_VREF pixel
xPix5683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[56] VREF PIX_IN[5683] NB2 NB1 CSA_VREF pixel
xPix5684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[56] VREF PIX_IN[5684] NB2 NB1 CSA_VREF pixel
xPix5685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[56] VREF PIX_IN[5685] NB2 NB1 CSA_VREF pixel
xPix5686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[56] VREF PIX_IN[5686] NB2 NB1 CSA_VREF pixel
xPix5687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[56] VREF PIX_IN[5687] NB2 NB1 CSA_VREF pixel
xPix5688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[56] VREF PIX_IN[5688] NB2 NB1 CSA_VREF pixel
xPix5689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[56] VREF PIX_IN[5689] NB2 NB1 CSA_VREF pixel
xPix5690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[56] VREF PIX_IN[5690] NB2 NB1 CSA_VREF pixel
xPix5691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[56] VREF PIX_IN[5691] NB2 NB1 CSA_VREF pixel
xPix5692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[56] VREF PIX_IN[5692] NB2 NB1 CSA_VREF pixel
xPix5693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[56] VREF PIX_IN[5693] NB2 NB1 CSA_VREF pixel
xPix5694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[56] VREF PIX_IN[5694] NB2 NB1 CSA_VREF pixel
xPix5695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[56] VREF PIX_IN[5695] NB2 NB1 CSA_VREF pixel
xPix5696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[56] VREF PIX_IN[5696] NB2 NB1 CSA_VREF pixel
xPix5697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[56] VREF PIX_IN[5697] NB2 NB1 CSA_VREF pixel
xPix5698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[56] VREF PIX_IN[5698] NB2 NB1 CSA_VREF pixel
xPix5699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[56] VREF PIX_IN[5699] NB2 NB1 CSA_VREF pixel
xPix5700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[57] VREF PIX_IN[5700] NB2 NB1 CSA_VREF pixel
xPix5701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[57] VREF PIX_IN[5701] NB2 NB1 CSA_VREF pixel
xPix5702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[57] VREF PIX_IN[5702] NB2 NB1 CSA_VREF pixel
xPix5703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[57] VREF PIX_IN[5703] NB2 NB1 CSA_VREF pixel
xPix5704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[57] VREF PIX_IN[5704] NB2 NB1 CSA_VREF pixel
xPix5705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[57] VREF PIX_IN[5705] NB2 NB1 CSA_VREF pixel
xPix5706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[57] VREF PIX_IN[5706] NB2 NB1 CSA_VREF pixel
xPix5707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[57] VREF PIX_IN[5707] NB2 NB1 CSA_VREF pixel
xPix5708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[57] VREF PIX_IN[5708] NB2 NB1 CSA_VREF pixel
xPix5709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[57] VREF PIX_IN[5709] NB2 NB1 CSA_VREF pixel
xPix5710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[57] VREF PIX_IN[5710] NB2 NB1 CSA_VREF pixel
xPix5711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[57] VREF PIX_IN[5711] NB2 NB1 CSA_VREF pixel
xPix5712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[57] VREF PIX_IN[5712] NB2 NB1 CSA_VREF pixel
xPix5713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[57] VREF PIX_IN[5713] NB2 NB1 CSA_VREF pixel
xPix5714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[57] VREF PIX_IN[5714] NB2 NB1 CSA_VREF pixel
xPix5715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[57] VREF PIX_IN[5715] NB2 NB1 CSA_VREF pixel
xPix5716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[57] VREF PIX_IN[5716] NB2 NB1 CSA_VREF pixel
xPix5717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[57] VREF PIX_IN[5717] NB2 NB1 CSA_VREF pixel
xPix5718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[57] VREF PIX_IN[5718] NB2 NB1 CSA_VREF pixel
xPix5719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[57] VREF PIX_IN[5719] NB2 NB1 CSA_VREF pixel
xPix5720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[57] VREF PIX_IN[5720] NB2 NB1 CSA_VREF pixel
xPix5721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[57] VREF PIX_IN[5721] NB2 NB1 CSA_VREF pixel
xPix5722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[57] VREF PIX_IN[5722] NB2 NB1 CSA_VREF pixel
xPix5723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[57] VREF PIX_IN[5723] NB2 NB1 CSA_VREF pixel
xPix5724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[57] VREF PIX_IN[5724] NB2 NB1 CSA_VREF pixel
xPix5725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[57] VREF PIX_IN[5725] NB2 NB1 CSA_VREF pixel
xPix5726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[57] VREF PIX_IN[5726] NB2 NB1 CSA_VREF pixel
xPix5727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[57] VREF PIX_IN[5727] NB2 NB1 CSA_VREF pixel
xPix5728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[57] VREF PIX_IN[5728] NB2 NB1 CSA_VREF pixel
xPix5729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[57] VREF PIX_IN[5729] NB2 NB1 CSA_VREF pixel
xPix5730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[57] VREF PIX_IN[5730] NB2 NB1 CSA_VREF pixel
xPix5731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[57] VREF PIX_IN[5731] NB2 NB1 CSA_VREF pixel
xPix5732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[57] VREF PIX_IN[5732] NB2 NB1 CSA_VREF pixel
xPix5733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[57] VREF PIX_IN[5733] NB2 NB1 CSA_VREF pixel
xPix5734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[57] VREF PIX_IN[5734] NB2 NB1 CSA_VREF pixel
xPix5735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[57] VREF PIX_IN[5735] NB2 NB1 CSA_VREF pixel
xPix5736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[57] VREF PIX_IN[5736] NB2 NB1 CSA_VREF pixel
xPix5737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[57] VREF PIX_IN[5737] NB2 NB1 CSA_VREF pixel
xPix5738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[57] VREF PIX_IN[5738] NB2 NB1 CSA_VREF pixel
xPix5739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[57] VREF PIX_IN[5739] NB2 NB1 CSA_VREF pixel
xPix5740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[57] VREF PIX_IN[5740] NB2 NB1 CSA_VREF pixel
xPix5741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[57] VREF PIX_IN[5741] NB2 NB1 CSA_VREF pixel
xPix5742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[57] VREF PIX_IN[5742] NB2 NB1 CSA_VREF pixel
xPix5743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[57] VREF PIX_IN[5743] NB2 NB1 CSA_VREF pixel
xPix5744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[57] VREF PIX_IN[5744] NB2 NB1 CSA_VREF pixel
xPix5745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[57] VREF PIX_IN[5745] NB2 NB1 CSA_VREF pixel
xPix5746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[57] VREF PIX_IN[5746] NB2 NB1 CSA_VREF pixel
xPix5747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[57] VREF PIX_IN[5747] NB2 NB1 CSA_VREF pixel
xPix5748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[57] VREF PIX_IN[5748] NB2 NB1 CSA_VREF pixel
xPix5749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[57] VREF PIX_IN[5749] NB2 NB1 CSA_VREF pixel
xPix5750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[57] VREF PIX_IN[5750] NB2 NB1 CSA_VREF pixel
xPix5751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[57] VREF PIX_IN[5751] NB2 NB1 CSA_VREF pixel
xPix5752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[57] VREF PIX_IN[5752] NB2 NB1 CSA_VREF pixel
xPix5753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[57] VREF PIX_IN[5753] NB2 NB1 CSA_VREF pixel
xPix5754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[57] VREF PIX_IN[5754] NB2 NB1 CSA_VREF pixel
xPix5755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[57] VREF PIX_IN[5755] NB2 NB1 CSA_VREF pixel
xPix5756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[57] VREF PIX_IN[5756] NB2 NB1 CSA_VREF pixel
xPix5757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[57] VREF PIX_IN[5757] NB2 NB1 CSA_VREF pixel
xPix5758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[57] VREF PIX_IN[5758] NB2 NB1 CSA_VREF pixel
xPix5759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[57] VREF PIX_IN[5759] NB2 NB1 CSA_VREF pixel
xPix5760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[57] VREF PIX_IN[5760] NB2 NB1 CSA_VREF pixel
xPix5761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[57] VREF PIX_IN[5761] NB2 NB1 CSA_VREF pixel
xPix5762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[57] VREF PIX_IN[5762] NB2 NB1 CSA_VREF pixel
xPix5763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[57] VREF PIX_IN[5763] NB2 NB1 CSA_VREF pixel
xPix5764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[57] VREF PIX_IN[5764] NB2 NB1 CSA_VREF pixel
xPix5765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[57] VREF PIX_IN[5765] NB2 NB1 CSA_VREF pixel
xPix5766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[57] VREF PIX_IN[5766] NB2 NB1 CSA_VREF pixel
xPix5767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[57] VREF PIX_IN[5767] NB2 NB1 CSA_VREF pixel
xPix5768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[57] VREF PIX_IN[5768] NB2 NB1 CSA_VREF pixel
xPix5769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[57] VREF PIX_IN[5769] NB2 NB1 CSA_VREF pixel
xPix5770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[57] VREF PIX_IN[5770] NB2 NB1 CSA_VREF pixel
xPix5771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[57] VREF PIX_IN[5771] NB2 NB1 CSA_VREF pixel
xPix5772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[57] VREF PIX_IN[5772] NB2 NB1 CSA_VREF pixel
xPix5773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[57] VREF PIX_IN[5773] NB2 NB1 CSA_VREF pixel
xPix5774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[57] VREF PIX_IN[5774] NB2 NB1 CSA_VREF pixel
xPix5775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[57] VREF PIX_IN[5775] NB2 NB1 CSA_VREF pixel
xPix5776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[57] VREF PIX_IN[5776] NB2 NB1 CSA_VREF pixel
xPix5777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[57] VREF PIX_IN[5777] NB2 NB1 CSA_VREF pixel
xPix5778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[57] VREF PIX_IN[5778] NB2 NB1 CSA_VREF pixel
xPix5779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[57] VREF PIX_IN[5779] NB2 NB1 CSA_VREF pixel
xPix5780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[57] VREF PIX_IN[5780] NB2 NB1 CSA_VREF pixel
xPix5781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[57] VREF PIX_IN[5781] NB2 NB1 CSA_VREF pixel
xPix5782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[57] VREF PIX_IN[5782] NB2 NB1 CSA_VREF pixel
xPix5783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[57] VREF PIX_IN[5783] NB2 NB1 CSA_VREF pixel
xPix5784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[57] VREF PIX_IN[5784] NB2 NB1 CSA_VREF pixel
xPix5785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[57] VREF PIX_IN[5785] NB2 NB1 CSA_VREF pixel
xPix5786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[57] VREF PIX_IN[5786] NB2 NB1 CSA_VREF pixel
xPix5787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[57] VREF PIX_IN[5787] NB2 NB1 CSA_VREF pixel
xPix5788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[57] VREF PIX_IN[5788] NB2 NB1 CSA_VREF pixel
xPix5789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[57] VREF PIX_IN[5789] NB2 NB1 CSA_VREF pixel
xPix5790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[57] VREF PIX_IN[5790] NB2 NB1 CSA_VREF pixel
xPix5791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[57] VREF PIX_IN[5791] NB2 NB1 CSA_VREF pixel
xPix5792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[57] VREF PIX_IN[5792] NB2 NB1 CSA_VREF pixel
xPix5793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[57] VREF PIX_IN[5793] NB2 NB1 CSA_VREF pixel
xPix5794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[57] VREF PIX_IN[5794] NB2 NB1 CSA_VREF pixel
xPix5795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[57] VREF PIX_IN[5795] NB2 NB1 CSA_VREF pixel
xPix5796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[57] VREF PIX_IN[5796] NB2 NB1 CSA_VREF pixel
xPix5797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[57] VREF PIX_IN[5797] NB2 NB1 CSA_VREF pixel
xPix5798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[57] VREF PIX_IN[5798] NB2 NB1 CSA_VREF pixel
xPix5799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[57] VREF PIX_IN[5799] NB2 NB1 CSA_VREF pixel
xPix5800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[58] VREF PIX_IN[5800] NB2 NB1 CSA_VREF pixel
xPix5801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[58] VREF PIX_IN[5801] NB2 NB1 CSA_VREF pixel
xPix5802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[58] VREF PIX_IN[5802] NB2 NB1 CSA_VREF pixel
xPix5803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[58] VREF PIX_IN[5803] NB2 NB1 CSA_VREF pixel
xPix5804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[58] VREF PIX_IN[5804] NB2 NB1 CSA_VREF pixel
xPix5805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[58] VREF PIX_IN[5805] NB2 NB1 CSA_VREF pixel
xPix5806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[58] VREF PIX_IN[5806] NB2 NB1 CSA_VREF pixel
xPix5807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[58] VREF PIX_IN[5807] NB2 NB1 CSA_VREF pixel
xPix5808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[58] VREF PIX_IN[5808] NB2 NB1 CSA_VREF pixel
xPix5809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[58] VREF PIX_IN[5809] NB2 NB1 CSA_VREF pixel
xPix5810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[58] VREF PIX_IN[5810] NB2 NB1 CSA_VREF pixel
xPix5811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[58] VREF PIX_IN[5811] NB2 NB1 CSA_VREF pixel
xPix5812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[58] VREF PIX_IN[5812] NB2 NB1 CSA_VREF pixel
xPix5813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[58] VREF PIX_IN[5813] NB2 NB1 CSA_VREF pixel
xPix5814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[58] VREF PIX_IN[5814] NB2 NB1 CSA_VREF pixel
xPix5815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[58] VREF PIX_IN[5815] NB2 NB1 CSA_VREF pixel
xPix5816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[58] VREF PIX_IN[5816] NB2 NB1 CSA_VREF pixel
xPix5817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[58] VREF PIX_IN[5817] NB2 NB1 CSA_VREF pixel
xPix5818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[58] VREF PIX_IN[5818] NB2 NB1 CSA_VREF pixel
xPix5819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[58] VREF PIX_IN[5819] NB2 NB1 CSA_VREF pixel
xPix5820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[58] VREF PIX_IN[5820] NB2 NB1 CSA_VREF pixel
xPix5821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[58] VREF PIX_IN[5821] NB2 NB1 CSA_VREF pixel
xPix5822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[58] VREF PIX_IN[5822] NB2 NB1 CSA_VREF pixel
xPix5823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[58] VREF PIX_IN[5823] NB2 NB1 CSA_VREF pixel
xPix5824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[58] VREF PIX_IN[5824] NB2 NB1 CSA_VREF pixel
xPix5825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[58] VREF PIX_IN[5825] NB2 NB1 CSA_VREF pixel
xPix5826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[58] VREF PIX_IN[5826] NB2 NB1 CSA_VREF pixel
xPix5827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[58] VREF PIX_IN[5827] NB2 NB1 CSA_VREF pixel
xPix5828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[58] VREF PIX_IN[5828] NB2 NB1 CSA_VREF pixel
xPix5829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[58] VREF PIX_IN[5829] NB2 NB1 CSA_VREF pixel
xPix5830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[58] VREF PIX_IN[5830] NB2 NB1 CSA_VREF pixel
xPix5831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[58] VREF PIX_IN[5831] NB2 NB1 CSA_VREF pixel
xPix5832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[58] VREF PIX_IN[5832] NB2 NB1 CSA_VREF pixel
xPix5833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[58] VREF PIX_IN[5833] NB2 NB1 CSA_VREF pixel
xPix5834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[58] VREF PIX_IN[5834] NB2 NB1 CSA_VREF pixel
xPix5835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[58] VREF PIX_IN[5835] NB2 NB1 CSA_VREF pixel
xPix5836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[58] VREF PIX_IN[5836] NB2 NB1 CSA_VREF pixel
xPix5837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[58] VREF PIX_IN[5837] NB2 NB1 CSA_VREF pixel
xPix5838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[58] VREF PIX_IN[5838] NB2 NB1 CSA_VREF pixel
xPix5839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[58] VREF PIX_IN[5839] NB2 NB1 CSA_VREF pixel
xPix5840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[58] VREF PIX_IN[5840] NB2 NB1 CSA_VREF pixel
xPix5841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[58] VREF PIX_IN[5841] NB2 NB1 CSA_VREF pixel
xPix5842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[58] VREF PIX_IN[5842] NB2 NB1 CSA_VREF pixel
xPix5843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[58] VREF PIX_IN[5843] NB2 NB1 CSA_VREF pixel
xPix5844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[58] VREF PIX_IN[5844] NB2 NB1 CSA_VREF pixel
xPix5845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[58] VREF PIX_IN[5845] NB2 NB1 CSA_VREF pixel
xPix5846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[58] VREF PIX_IN[5846] NB2 NB1 CSA_VREF pixel
xPix5847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[58] VREF PIX_IN[5847] NB2 NB1 CSA_VREF pixel
xPix5848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[58] VREF PIX_IN[5848] NB2 NB1 CSA_VREF pixel
xPix5849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[58] VREF PIX_IN[5849] NB2 NB1 CSA_VREF pixel
xPix5850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[58] VREF PIX_IN[5850] NB2 NB1 CSA_VREF pixel
xPix5851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[58] VREF PIX_IN[5851] NB2 NB1 CSA_VREF pixel
xPix5852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[58] VREF PIX_IN[5852] NB2 NB1 CSA_VREF pixel
xPix5853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[58] VREF PIX_IN[5853] NB2 NB1 CSA_VREF pixel
xPix5854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[58] VREF PIX_IN[5854] NB2 NB1 CSA_VREF pixel
xPix5855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[58] VREF PIX_IN[5855] NB2 NB1 CSA_VREF pixel
xPix5856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[58] VREF PIX_IN[5856] NB2 NB1 CSA_VREF pixel
xPix5857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[58] VREF PIX_IN[5857] NB2 NB1 CSA_VREF pixel
xPix5858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[58] VREF PIX_IN[5858] NB2 NB1 CSA_VREF pixel
xPix5859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[58] VREF PIX_IN[5859] NB2 NB1 CSA_VREF pixel
xPix5860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[58] VREF PIX_IN[5860] NB2 NB1 CSA_VREF pixel
xPix5861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[58] VREF PIX_IN[5861] NB2 NB1 CSA_VREF pixel
xPix5862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[58] VREF PIX_IN[5862] NB2 NB1 CSA_VREF pixel
xPix5863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[58] VREF PIX_IN[5863] NB2 NB1 CSA_VREF pixel
xPix5864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[58] VREF PIX_IN[5864] NB2 NB1 CSA_VREF pixel
xPix5865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[58] VREF PIX_IN[5865] NB2 NB1 CSA_VREF pixel
xPix5866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[58] VREF PIX_IN[5866] NB2 NB1 CSA_VREF pixel
xPix5867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[58] VREF PIX_IN[5867] NB2 NB1 CSA_VREF pixel
xPix5868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[58] VREF PIX_IN[5868] NB2 NB1 CSA_VREF pixel
xPix5869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[58] VREF PIX_IN[5869] NB2 NB1 CSA_VREF pixel
xPix5870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[58] VREF PIX_IN[5870] NB2 NB1 CSA_VREF pixel
xPix5871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[58] VREF PIX_IN[5871] NB2 NB1 CSA_VREF pixel
xPix5872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[58] VREF PIX_IN[5872] NB2 NB1 CSA_VREF pixel
xPix5873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[58] VREF PIX_IN[5873] NB2 NB1 CSA_VREF pixel
xPix5874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[58] VREF PIX_IN[5874] NB2 NB1 CSA_VREF pixel
xPix5875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[58] VREF PIX_IN[5875] NB2 NB1 CSA_VREF pixel
xPix5876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[58] VREF PIX_IN[5876] NB2 NB1 CSA_VREF pixel
xPix5877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[58] VREF PIX_IN[5877] NB2 NB1 CSA_VREF pixel
xPix5878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[58] VREF PIX_IN[5878] NB2 NB1 CSA_VREF pixel
xPix5879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[58] VREF PIX_IN[5879] NB2 NB1 CSA_VREF pixel
xPix5880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[58] VREF PIX_IN[5880] NB2 NB1 CSA_VREF pixel
xPix5881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[58] VREF PIX_IN[5881] NB2 NB1 CSA_VREF pixel
xPix5882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[58] VREF PIX_IN[5882] NB2 NB1 CSA_VREF pixel
xPix5883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[58] VREF PIX_IN[5883] NB2 NB1 CSA_VREF pixel
xPix5884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[58] VREF PIX_IN[5884] NB2 NB1 CSA_VREF pixel
xPix5885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[58] VREF PIX_IN[5885] NB2 NB1 CSA_VREF pixel
xPix5886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[58] VREF PIX_IN[5886] NB2 NB1 CSA_VREF pixel
xPix5887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[58] VREF PIX_IN[5887] NB2 NB1 CSA_VREF pixel
xPix5888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[58] VREF PIX_IN[5888] NB2 NB1 CSA_VREF pixel
xPix5889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[58] VREF PIX_IN[5889] NB2 NB1 CSA_VREF pixel
xPix5890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[58] VREF PIX_IN[5890] NB2 NB1 CSA_VREF pixel
xPix5891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[58] VREF PIX_IN[5891] NB2 NB1 CSA_VREF pixel
xPix5892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[58] VREF PIX_IN[5892] NB2 NB1 CSA_VREF pixel
xPix5893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[58] VREF PIX_IN[5893] NB2 NB1 CSA_VREF pixel
xPix5894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[58] VREF PIX_IN[5894] NB2 NB1 CSA_VREF pixel
xPix5895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[58] VREF PIX_IN[5895] NB2 NB1 CSA_VREF pixel
xPix5896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[58] VREF PIX_IN[5896] NB2 NB1 CSA_VREF pixel
xPix5897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[58] VREF PIX_IN[5897] NB2 NB1 CSA_VREF pixel
xPix5898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[58] VREF PIX_IN[5898] NB2 NB1 CSA_VREF pixel
xPix5899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[58] VREF PIX_IN[5899] NB2 NB1 CSA_VREF pixel
xPix5900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[59] VREF PIX_IN[5900] NB2 NB1 CSA_VREF pixel
xPix5901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[59] VREF PIX_IN[5901] NB2 NB1 CSA_VREF pixel
xPix5902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[59] VREF PIX_IN[5902] NB2 NB1 CSA_VREF pixel
xPix5903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[59] VREF PIX_IN[5903] NB2 NB1 CSA_VREF pixel
xPix5904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[59] VREF PIX_IN[5904] NB2 NB1 CSA_VREF pixel
xPix5905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[59] VREF PIX_IN[5905] NB2 NB1 CSA_VREF pixel
xPix5906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[59] VREF PIX_IN[5906] NB2 NB1 CSA_VREF pixel
xPix5907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[59] VREF PIX_IN[5907] NB2 NB1 CSA_VREF pixel
xPix5908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[59] VREF PIX_IN[5908] NB2 NB1 CSA_VREF pixel
xPix5909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[59] VREF PIX_IN[5909] NB2 NB1 CSA_VREF pixel
xPix5910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[59] VREF PIX_IN[5910] NB2 NB1 CSA_VREF pixel
xPix5911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[59] VREF PIX_IN[5911] NB2 NB1 CSA_VREF pixel
xPix5912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[59] VREF PIX_IN[5912] NB2 NB1 CSA_VREF pixel
xPix5913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[59] VREF PIX_IN[5913] NB2 NB1 CSA_VREF pixel
xPix5914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[59] VREF PIX_IN[5914] NB2 NB1 CSA_VREF pixel
xPix5915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[59] VREF PIX_IN[5915] NB2 NB1 CSA_VREF pixel
xPix5916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[59] VREF PIX_IN[5916] NB2 NB1 CSA_VREF pixel
xPix5917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[59] VREF PIX_IN[5917] NB2 NB1 CSA_VREF pixel
xPix5918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[59] VREF PIX_IN[5918] NB2 NB1 CSA_VREF pixel
xPix5919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[59] VREF PIX_IN[5919] NB2 NB1 CSA_VREF pixel
xPix5920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[59] VREF PIX_IN[5920] NB2 NB1 CSA_VREF pixel
xPix5921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[59] VREF PIX_IN[5921] NB2 NB1 CSA_VREF pixel
xPix5922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[59] VREF PIX_IN[5922] NB2 NB1 CSA_VREF pixel
xPix5923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[59] VREF PIX_IN[5923] NB2 NB1 CSA_VREF pixel
xPix5924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[59] VREF PIX_IN[5924] NB2 NB1 CSA_VREF pixel
xPix5925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[59] VREF PIX_IN[5925] NB2 NB1 CSA_VREF pixel
xPix5926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[59] VREF PIX_IN[5926] NB2 NB1 CSA_VREF pixel
xPix5927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[59] VREF PIX_IN[5927] NB2 NB1 CSA_VREF pixel
xPix5928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[59] VREF PIX_IN[5928] NB2 NB1 CSA_VREF pixel
xPix5929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[59] VREF PIX_IN[5929] NB2 NB1 CSA_VREF pixel
xPix5930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[59] VREF PIX_IN[5930] NB2 NB1 CSA_VREF pixel
xPix5931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[59] VREF PIX_IN[5931] NB2 NB1 CSA_VREF pixel
xPix5932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[59] VREF PIX_IN[5932] NB2 NB1 CSA_VREF pixel
xPix5933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[59] VREF PIX_IN[5933] NB2 NB1 CSA_VREF pixel
xPix5934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[59] VREF PIX_IN[5934] NB2 NB1 CSA_VREF pixel
xPix5935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[59] VREF PIX_IN[5935] NB2 NB1 CSA_VREF pixel
xPix5936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[59] VREF PIX_IN[5936] NB2 NB1 CSA_VREF pixel
xPix5937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[59] VREF PIX_IN[5937] NB2 NB1 CSA_VREF pixel
xPix5938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[59] VREF PIX_IN[5938] NB2 NB1 CSA_VREF pixel
xPix5939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[59] VREF PIX_IN[5939] NB2 NB1 CSA_VREF pixel
xPix5940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[59] VREF PIX_IN[5940] NB2 NB1 CSA_VREF pixel
xPix5941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[59] VREF PIX_IN[5941] NB2 NB1 CSA_VREF pixel
xPix5942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[59] VREF PIX_IN[5942] NB2 NB1 CSA_VREF pixel
xPix5943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[59] VREF PIX_IN[5943] NB2 NB1 CSA_VREF pixel
xPix5944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[59] VREF PIX_IN[5944] NB2 NB1 CSA_VREF pixel
xPix5945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[59] VREF PIX_IN[5945] NB2 NB1 CSA_VREF pixel
xPix5946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[59] VREF PIX_IN[5946] NB2 NB1 CSA_VREF pixel
xPix5947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[59] VREF PIX_IN[5947] NB2 NB1 CSA_VREF pixel
xPix5948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[59] VREF PIX_IN[5948] NB2 NB1 CSA_VREF pixel
xPix5949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[59] VREF PIX_IN[5949] NB2 NB1 CSA_VREF pixel
xPix5950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[59] VREF PIX_IN[5950] NB2 NB1 CSA_VREF pixel
xPix5951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[59] VREF PIX_IN[5951] NB2 NB1 CSA_VREF pixel
xPix5952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[59] VREF PIX_IN[5952] NB2 NB1 CSA_VREF pixel
xPix5953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[59] VREF PIX_IN[5953] NB2 NB1 CSA_VREF pixel
xPix5954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[59] VREF PIX_IN[5954] NB2 NB1 CSA_VREF pixel
xPix5955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[59] VREF PIX_IN[5955] NB2 NB1 CSA_VREF pixel
xPix5956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[59] VREF PIX_IN[5956] NB2 NB1 CSA_VREF pixel
xPix5957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[59] VREF PIX_IN[5957] NB2 NB1 CSA_VREF pixel
xPix5958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[59] VREF PIX_IN[5958] NB2 NB1 CSA_VREF pixel
xPix5959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[59] VREF PIX_IN[5959] NB2 NB1 CSA_VREF pixel
xPix5960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[59] VREF PIX_IN[5960] NB2 NB1 CSA_VREF pixel
xPix5961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[59] VREF PIX_IN[5961] NB2 NB1 CSA_VREF pixel
xPix5962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[59] VREF PIX_IN[5962] NB2 NB1 CSA_VREF pixel
xPix5963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[59] VREF PIX_IN[5963] NB2 NB1 CSA_VREF pixel
xPix5964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[59] VREF PIX_IN[5964] NB2 NB1 CSA_VREF pixel
xPix5965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[59] VREF PIX_IN[5965] NB2 NB1 CSA_VREF pixel
xPix5966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[59] VREF PIX_IN[5966] NB2 NB1 CSA_VREF pixel
xPix5967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[59] VREF PIX_IN[5967] NB2 NB1 CSA_VREF pixel
xPix5968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[59] VREF PIX_IN[5968] NB2 NB1 CSA_VREF pixel
xPix5969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[59] VREF PIX_IN[5969] NB2 NB1 CSA_VREF pixel
xPix5970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[59] VREF PIX_IN[5970] NB2 NB1 CSA_VREF pixel
xPix5971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[59] VREF PIX_IN[5971] NB2 NB1 CSA_VREF pixel
xPix5972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[59] VREF PIX_IN[5972] NB2 NB1 CSA_VREF pixel
xPix5973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[59] VREF PIX_IN[5973] NB2 NB1 CSA_VREF pixel
xPix5974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[59] VREF PIX_IN[5974] NB2 NB1 CSA_VREF pixel
xPix5975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[59] VREF PIX_IN[5975] NB2 NB1 CSA_VREF pixel
xPix5976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[59] VREF PIX_IN[5976] NB2 NB1 CSA_VREF pixel
xPix5977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[59] VREF PIX_IN[5977] NB2 NB1 CSA_VREF pixel
xPix5978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[59] VREF PIX_IN[5978] NB2 NB1 CSA_VREF pixel
xPix5979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[59] VREF PIX_IN[5979] NB2 NB1 CSA_VREF pixel
xPix5980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[59] VREF PIX_IN[5980] NB2 NB1 CSA_VREF pixel
xPix5981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[59] VREF PIX_IN[5981] NB2 NB1 CSA_VREF pixel
xPix5982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[59] VREF PIX_IN[5982] NB2 NB1 CSA_VREF pixel
xPix5983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[59] VREF PIX_IN[5983] NB2 NB1 CSA_VREF pixel
xPix5984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[59] VREF PIX_IN[5984] NB2 NB1 CSA_VREF pixel
xPix5985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[59] VREF PIX_IN[5985] NB2 NB1 CSA_VREF pixel
xPix5986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[59] VREF PIX_IN[5986] NB2 NB1 CSA_VREF pixel
xPix5987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[59] VREF PIX_IN[5987] NB2 NB1 CSA_VREF pixel
xPix5988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[59] VREF PIX_IN[5988] NB2 NB1 CSA_VREF pixel
xPix5989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[59] VREF PIX_IN[5989] NB2 NB1 CSA_VREF pixel
xPix5990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[59] VREF PIX_IN[5990] NB2 NB1 CSA_VREF pixel
xPix5991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[59] VREF PIX_IN[5991] NB2 NB1 CSA_VREF pixel
xPix5992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[59] VREF PIX_IN[5992] NB2 NB1 CSA_VREF pixel
xPix5993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[59] VREF PIX_IN[5993] NB2 NB1 CSA_VREF pixel
xPix5994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[59] VREF PIX_IN[5994] NB2 NB1 CSA_VREF pixel
xPix5995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[59] VREF PIX_IN[5995] NB2 NB1 CSA_VREF pixel
xPix5996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[59] VREF PIX_IN[5996] NB2 NB1 CSA_VREF pixel
xPix5997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[59] VREF PIX_IN[5997] NB2 NB1 CSA_VREF pixel
xPix5998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[59] VREF PIX_IN[5998] NB2 NB1 CSA_VREF pixel
xPix5999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[59] VREF PIX_IN[5999] NB2 NB1 CSA_VREF pixel
xPix6000 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[60] VREF PIX_IN[6000] NB2 NB1 CSA_VREF pixel
xPix6001 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[60] VREF PIX_IN[6001] NB2 NB1 CSA_VREF pixel
xPix6002 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[60] VREF PIX_IN[6002] NB2 NB1 CSA_VREF pixel
xPix6003 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[60] VREF PIX_IN[6003] NB2 NB1 CSA_VREF pixel
xPix6004 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[60] VREF PIX_IN[6004] NB2 NB1 CSA_VREF pixel
xPix6005 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[60] VREF PIX_IN[6005] NB2 NB1 CSA_VREF pixel
xPix6006 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[60] VREF PIX_IN[6006] NB2 NB1 CSA_VREF pixel
xPix6007 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[60] VREF PIX_IN[6007] NB2 NB1 CSA_VREF pixel
xPix6008 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[60] VREF PIX_IN[6008] NB2 NB1 CSA_VREF pixel
xPix6009 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[60] VREF PIX_IN[6009] NB2 NB1 CSA_VREF pixel
xPix6010 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[60] VREF PIX_IN[6010] NB2 NB1 CSA_VREF pixel
xPix6011 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[60] VREF PIX_IN[6011] NB2 NB1 CSA_VREF pixel
xPix6012 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[60] VREF PIX_IN[6012] NB2 NB1 CSA_VREF pixel
xPix6013 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[60] VREF PIX_IN[6013] NB2 NB1 CSA_VREF pixel
xPix6014 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[60] VREF PIX_IN[6014] NB2 NB1 CSA_VREF pixel
xPix6015 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[60] VREF PIX_IN[6015] NB2 NB1 CSA_VREF pixel
xPix6016 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[60] VREF PIX_IN[6016] NB2 NB1 CSA_VREF pixel
xPix6017 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[60] VREF PIX_IN[6017] NB2 NB1 CSA_VREF pixel
xPix6018 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[60] VREF PIX_IN[6018] NB2 NB1 CSA_VREF pixel
xPix6019 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[60] VREF PIX_IN[6019] NB2 NB1 CSA_VREF pixel
xPix6020 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[60] VREF PIX_IN[6020] NB2 NB1 CSA_VREF pixel
xPix6021 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[60] VREF PIX_IN[6021] NB2 NB1 CSA_VREF pixel
xPix6022 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[60] VREF PIX_IN[6022] NB2 NB1 CSA_VREF pixel
xPix6023 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[60] VREF PIX_IN[6023] NB2 NB1 CSA_VREF pixel
xPix6024 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[60] VREF PIX_IN[6024] NB2 NB1 CSA_VREF pixel
xPix6025 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[60] VREF PIX_IN[6025] NB2 NB1 CSA_VREF pixel
xPix6026 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[60] VREF PIX_IN[6026] NB2 NB1 CSA_VREF pixel
xPix6027 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[60] VREF PIX_IN[6027] NB2 NB1 CSA_VREF pixel
xPix6028 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[60] VREF PIX_IN[6028] NB2 NB1 CSA_VREF pixel
xPix6029 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[60] VREF PIX_IN[6029] NB2 NB1 CSA_VREF pixel
xPix6030 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[60] VREF PIX_IN[6030] NB2 NB1 CSA_VREF pixel
xPix6031 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[60] VREF PIX_IN[6031] NB2 NB1 CSA_VREF pixel
xPix6032 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[60] VREF PIX_IN[6032] NB2 NB1 CSA_VREF pixel
xPix6033 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[60] VREF PIX_IN[6033] NB2 NB1 CSA_VREF pixel
xPix6034 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[60] VREF PIX_IN[6034] NB2 NB1 CSA_VREF pixel
xPix6035 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[60] VREF PIX_IN[6035] NB2 NB1 CSA_VREF pixel
xPix6036 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[60] VREF PIX_IN[6036] NB2 NB1 CSA_VREF pixel
xPix6037 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[60] VREF PIX_IN[6037] NB2 NB1 CSA_VREF pixel
xPix6038 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[60] VREF PIX_IN[6038] NB2 NB1 CSA_VREF pixel
xPix6039 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[60] VREF PIX_IN[6039] NB2 NB1 CSA_VREF pixel
xPix6040 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[60] VREF PIX_IN[6040] NB2 NB1 CSA_VREF pixel
xPix6041 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[60] VREF PIX_IN[6041] NB2 NB1 CSA_VREF pixel
xPix6042 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[60] VREF PIX_IN[6042] NB2 NB1 CSA_VREF pixel
xPix6043 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[60] VREF PIX_IN[6043] NB2 NB1 CSA_VREF pixel
xPix6044 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[60] VREF PIX_IN[6044] NB2 NB1 CSA_VREF pixel
xPix6045 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[60] VREF PIX_IN[6045] NB2 NB1 CSA_VREF pixel
xPix6046 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[60] VREF PIX_IN[6046] NB2 NB1 CSA_VREF pixel
xPix6047 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[60] VREF PIX_IN[6047] NB2 NB1 CSA_VREF pixel
xPix6048 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[60] VREF PIX_IN[6048] NB2 NB1 CSA_VREF pixel
xPix6049 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[60] VREF PIX_IN[6049] NB2 NB1 CSA_VREF pixel
xPix6050 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[60] VREF PIX_IN[6050] NB2 NB1 CSA_VREF pixel
xPix6051 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[60] VREF PIX_IN[6051] NB2 NB1 CSA_VREF pixel
xPix6052 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[60] VREF PIX_IN[6052] NB2 NB1 CSA_VREF pixel
xPix6053 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[60] VREF PIX_IN[6053] NB2 NB1 CSA_VREF pixel
xPix6054 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[60] VREF PIX_IN[6054] NB2 NB1 CSA_VREF pixel
xPix6055 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[60] VREF PIX_IN[6055] NB2 NB1 CSA_VREF pixel
xPix6056 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[60] VREF PIX_IN[6056] NB2 NB1 CSA_VREF pixel
xPix6057 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[60] VREF PIX_IN[6057] NB2 NB1 CSA_VREF pixel
xPix6058 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[60] VREF PIX_IN[6058] NB2 NB1 CSA_VREF pixel
xPix6059 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[60] VREF PIX_IN[6059] NB2 NB1 CSA_VREF pixel
xPix6060 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[60] VREF PIX_IN[6060] NB2 NB1 CSA_VREF pixel
xPix6061 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[60] VREF PIX_IN[6061] NB2 NB1 CSA_VREF pixel
xPix6062 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[60] VREF PIX_IN[6062] NB2 NB1 CSA_VREF pixel
xPix6063 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[60] VREF PIX_IN[6063] NB2 NB1 CSA_VREF pixel
xPix6064 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[60] VREF PIX_IN[6064] NB2 NB1 CSA_VREF pixel
xPix6065 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[60] VREF PIX_IN[6065] NB2 NB1 CSA_VREF pixel
xPix6066 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[60] VREF PIX_IN[6066] NB2 NB1 CSA_VREF pixel
xPix6067 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[60] VREF PIX_IN[6067] NB2 NB1 CSA_VREF pixel
xPix6068 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[60] VREF PIX_IN[6068] NB2 NB1 CSA_VREF pixel
xPix6069 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[60] VREF PIX_IN[6069] NB2 NB1 CSA_VREF pixel
xPix6070 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[60] VREF PIX_IN[6070] NB2 NB1 CSA_VREF pixel
xPix6071 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[60] VREF PIX_IN[6071] NB2 NB1 CSA_VREF pixel
xPix6072 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[60] VREF PIX_IN[6072] NB2 NB1 CSA_VREF pixel
xPix6073 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[60] VREF PIX_IN[6073] NB2 NB1 CSA_VREF pixel
xPix6074 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[60] VREF PIX_IN[6074] NB2 NB1 CSA_VREF pixel
xPix6075 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[60] VREF PIX_IN[6075] NB2 NB1 CSA_VREF pixel
xPix6076 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[60] VREF PIX_IN[6076] NB2 NB1 CSA_VREF pixel
xPix6077 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[60] VREF PIX_IN[6077] NB2 NB1 CSA_VREF pixel
xPix6078 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[60] VREF PIX_IN[6078] NB2 NB1 CSA_VREF pixel
xPix6079 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[60] VREF PIX_IN[6079] NB2 NB1 CSA_VREF pixel
xPix6080 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[60] VREF PIX_IN[6080] NB2 NB1 CSA_VREF pixel
xPix6081 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[60] VREF PIX_IN[6081] NB2 NB1 CSA_VREF pixel
xPix6082 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[60] VREF PIX_IN[6082] NB2 NB1 CSA_VREF pixel
xPix6083 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[60] VREF PIX_IN[6083] NB2 NB1 CSA_VREF pixel
xPix6084 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[60] VREF PIX_IN[6084] NB2 NB1 CSA_VREF pixel
xPix6085 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[60] VREF PIX_IN[6085] NB2 NB1 CSA_VREF pixel
xPix6086 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[60] VREF PIX_IN[6086] NB2 NB1 CSA_VREF pixel
xPix6087 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[60] VREF PIX_IN[6087] NB2 NB1 CSA_VREF pixel
xPix6088 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[60] VREF PIX_IN[6088] NB2 NB1 CSA_VREF pixel
xPix6089 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[60] VREF PIX_IN[6089] NB2 NB1 CSA_VREF pixel
xPix6090 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[60] VREF PIX_IN[6090] NB2 NB1 CSA_VREF pixel
xPix6091 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[60] VREF PIX_IN[6091] NB2 NB1 CSA_VREF pixel
xPix6092 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[60] VREF PIX_IN[6092] NB2 NB1 CSA_VREF pixel
xPix6093 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[60] VREF PIX_IN[6093] NB2 NB1 CSA_VREF pixel
xPix6094 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[60] VREF PIX_IN[6094] NB2 NB1 CSA_VREF pixel
xPix6095 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[60] VREF PIX_IN[6095] NB2 NB1 CSA_VREF pixel
xPix6096 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[60] VREF PIX_IN[6096] NB2 NB1 CSA_VREF pixel
xPix6097 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[60] VREF PIX_IN[6097] NB2 NB1 CSA_VREF pixel
xPix6098 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[60] VREF PIX_IN[6098] NB2 NB1 CSA_VREF pixel
xPix6099 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[60] VREF PIX_IN[6099] NB2 NB1 CSA_VREF pixel
xPix6100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[61] VREF PIX_IN[6100] NB2 NB1 CSA_VREF pixel
xPix6101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[61] VREF PIX_IN[6101] NB2 NB1 CSA_VREF pixel
xPix6102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[61] VREF PIX_IN[6102] NB2 NB1 CSA_VREF pixel
xPix6103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[61] VREF PIX_IN[6103] NB2 NB1 CSA_VREF pixel
xPix6104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[61] VREF PIX_IN[6104] NB2 NB1 CSA_VREF pixel
xPix6105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[61] VREF PIX_IN[6105] NB2 NB1 CSA_VREF pixel
xPix6106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[61] VREF PIX_IN[6106] NB2 NB1 CSA_VREF pixel
xPix6107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[61] VREF PIX_IN[6107] NB2 NB1 CSA_VREF pixel
xPix6108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[61] VREF PIX_IN[6108] NB2 NB1 CSA_VREF pixel
xPix6109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[61] VREF PIX_IN[6109] NB2 NB1 CSA_VREF pixel
xPix6110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[61] VREF PIX_IN[6110] NB2 NB1 CSA_VREF pixel
xPix6111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[61] VREF PIX_IN[6111] NB2 NB1 CSA_VREF pixel
xPix6112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[61] VREF PIX_IN[6112] NB2 NB1 CSA_VREF pixel
xPix6113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[61] VREF PIX_IN[6113] NB2 NB1 CSA_VREF pixel
xPix6114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[61] VREF PIX_IN[6114] NB2 NB1 CSA_VREF pixel
xPix6115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[61] VREF PIX_IN[6115] NB2 NB1 CSA_VREF pixel
xPix6116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[61] VREF PIX_IN[6116] NB2 NB1 CSA_VREF pixel
xPix6117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[61] VREF PIX_IN[6117] NB2 NB1 CSA_VREF pixel
xPix6118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[61] VREF PIX_IN[6118] NB2 NB1 CSA_VREF pixel
xPix6119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[61] VREF PIX_IN[6119] NB2 NB1 CSA_VREF pixel
xPix6120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[61] VREF PIX_IN[6120] NB2 NB1 CSA_VREF pixel
xPix6121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[61] VREF PIX_IN[6121] NB2 NB1 CSA_VREF pixel
xPix6122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[61] VREF PIX_IN[6122] NB2 NB1 CSA_VREF pixel
xPix6123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[61] VREF PIX_IN[6123] NB2 NB1 CSA_VREF pixel
xPix6124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[61] VREF PIX_IN[6124] NB2 NB1 CSA_VREF pixel
xPix6125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[61] VREF PIX_IN[6125] NB2 NB1 CSA_VREF pixel
xPix6126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[61] VREF PIX_IN[6126] NB2 NB1 CSA_VREF pixel
xPix6127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[61] VREF PIX_IN[6127] NB2 NB1 CSA_VREF pixel
xPix6128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[61] VREF PIX_IN[6128] NB2 NB1 CSA_VREF pixel
xPix6129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[61] VREF PIX_IN[6129] NB2 NB1 CSA_VREF pixel
xPix6130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[61] VREF PIX_IN[6130] NB2 NB1 CSA_VREF pixel
xPix6131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[61] VREF PIX_IN[6131] NB2 NB1 CSA_VREF pixel
xPix6132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[61] VREF PIX_IN[6132] NB2 NB1 CSA_VREF pixel
xPix6133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[61] VREF PIX_IN[6133] NB2 NB1 CSA_VREF pixel
xPix6134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[61] VREF PIX_IN[6134] NB2 NB1 CSA_VREF pixel
xPix6135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[61] VREF PIX_IN[6135] NB2 NB1 CSA_VREF pixel
xPix6136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[61] VREF PIX_IN[6136] NB2 NB1 CSA_VREF pixel
xPix6137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[61] VREF PIX_IN[6137] NB2 NB1 CSA_VREF pixel
xPix6138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[61] VREF PIX_IN[6138] NB2 NB1 CSA_VREF pixel
xPix6139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[61] VREF PIX_IN[6139] NB2 NB1 CSA_VREF pixel
xPix6140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[61] VREF PIX_IN[6140] NB2 NB1 CSA_VREF pixel
xPix6141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[61] VREF PIX_IN[6141] NB2 NB1 CSA_VREF pixel
xPix6142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[61] VREF PIX_IN[6142] NB2 NB1 CSA_VREF pixel
xPix6143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[61] VREF PIX_IN[6143] NB2 NB1 CSA_VREF pixel
xPix6144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[61] VREF PIX_IN[6144] NB2 NB1 CSA_VREF pixel
xPix6145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[61] VREF PIX_IN[6145] NB2 NB1 CSA_VREF pixel
xPix6146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[61] VREF PIX_IN[6146] NB2 NB1 CSA_VREF pixel
xPix6147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[61] VREF PIX_IN[6147] NB2 NB1 CSA_VREF pixel
xPix6148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[61] VREF PIX_IN[6148] NB2 NB1 CSA_VREF pixel
xPix6149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[61] VREF PIX_IN[6149] NB2 NB1 CSA_VREF pixel
xPix6150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[61] VREF PIX_IN[6150] NB2 NB1 CSA_VREF pixel
xPix6151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[61] VREF PIX_IN[6151] NB2 NB1 CSA_VREF pixel
xPix6152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[61] VREF PIX_IN[6152] NB2 NB1 CSA_VREF pixel
xPix6153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[61] VREF PIX_IN[6153] NB2 NB1 CSA_VREF pixel
xPix6154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[61] VREF PIX_IN[6154] NB2 NB1 CSA_VREF pixel
xPix6155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[61] VREF PIX_IN[6155] NB2 NB1 CSA_VREF pixel
xPix6156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[61] VREF PIX_IN[6156] NB2 NB1 CSA_VREF pixel
xPix6157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[61] VREF PIX_IN[6157] NB2 NB1 CSA_VREF pixel
xPix6158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[61] VREF PIX_IN[6158] NB2 NB1 CSA_VREF pixel
xPix6159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[61] VREF PIX_IN[6159] NB2 NB1 CSA_VREF pixel
xPix6160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[61] VREF PIX_IN[6160] NB2 NB1 CSA_VREF pixel
xPix6161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[61] VREF PIX_IN[6161] NB2 NB1 CSA_VREF pixel
xPix6162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[61] VREF PIX_IN[6162] NB2 NB1 CSA_VREF pixel
xPix6163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[61] VREF PIX_IN[6163] NB2 NB1 CSA_VREF pixel
xPix6164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[61] VREF PIX_IN[6164] NB2 NB1 CSA_VREF pixel
xPix6165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[61] VREF PIX_IN[6165] NB2 NB1 CSA_VREF pixel
xPix6166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[61] VREF PIX_IN[6166] NB2 NB1 CSA_VREF pixel
xPix6167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[61] VREF PIX_IN[6167] NB2 NB1 CSA_VREF pixel
xPix6168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[61] VREF PIX_IN[6168] NB2 NB1 CSA_VREF pixel
xPix6169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[61] VREF PIX_IN[6169] NB2 NB1 CSA_VREF pixel
xPix6170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[61] VREF PIX_IN[6170] NB2 NB1 CSA_VREF pixel
xPix6171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[61] VREF PIX_IN[6171] NB2 NB1 CSA_VREF pixel
xPix6172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[61] VREF PIX_IN[6172] NB2 NB1 CSA_VREF pixel
xPix6173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[61] VREF PIX_IN[6173] NB2 NB1 CSA_VREF pixel
xPix6174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[61] VREF PIX_IN[6174] NB2 NB1 CSA_VREF pixel
xPix6175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[61] VREF PIX_IN[6175] NB2 NB1 CSA_VREF pixel
xPix6176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[61] VREF PIX_IN[6176] NB2 NB1 CSA_VREF pixel
xPix6177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[61] VREF PIX_IN[6177] NB2 NB1 CSA_VREF pixel
xPix6178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[61] VREF PIX_IN[6178] NB2 NB1 CSA_VREF pixel
xPix6179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[61] VREF PIX_IN[6179] NB2 NB1 CSA_VREF pixel
xPix6180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[61] VREF PIX_IN[6180] NB2 NB1 CSA_VREF pixel
xPix6181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[61] VREF PIX_IN[6181] NB2 NB1 CSA_VREF pixel
xPix6182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[61] VREF PIX_IN[6182] NB2 NB1 CSA_VREF pixel
xPix6183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[61] VREF PIX_IN[6183] NB2 NB1 CSA_VREF pixel
xPix6184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[61] VREF PIX_IN[6184] NB2 NB1 CSA_VREF pixel
xPix6185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[61] VREF PIX_IN[6185] NB2 NB1 CSA_VREF pixel
xPix6186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[61] VREF PIX_IN[6186] NB2 NB1 CSA_VREF pixel
xPix6187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[61] VREF PIX_IN[6187] NB2 NB1 CSA_VREF pixel
xPix6188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[61] VREF PIX_IN[6188] NB2 NB1 CSA_VREF pixel
xPix6189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[61] VREF PIX_IN[6189] NB2 NB1 CSA_VREF pixel
xPix6190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[61] VREF PIX_IN[6190] NB2 NB1 CSA_VREF pixel
xPix6191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[61] VREF PIX_IN[6191] NB2 NB1 CSA_VREF pixel
xPix6192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[61] VREF PIX_IN[6192] NB2 NB1 CSA_VREF pixel
xPix6193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[61] VREF PIX_IN[6193] NB2 NB1 CSA_VREF pixel
xPix6194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[61] VREF PIX_IN[6194] NB2 NB1 CSA_VREF pixel
xPix6195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[61] VREF PIX_IN[6195] NB2 NB1 CSA_VREF pixel
xPix6196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[61] VREF PIX_IN[6196] NB2 NB1 CSA_VREF pixel
xPix6197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[61] VREF PIX_IN[6197] NB2 NB1 CSA_VREF pixel
xPix6198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[61] VREF PIX_IN[6198] NB2 NB1 CSA_VREF pixel
xPix6199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[61] VREF PIX_IN[6199] NB2 NB1 CSA_VREF pixel
xPix6200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[62] VREF PIX_IN[6200] NB2 NB1 CSA_VREF pixel
xPix6201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[62] VREF PIX_IN[6201] NB2 NB1 CSA_VREF pixel
xPix6202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[62] VREF PIX_IN[6202] NB2 NB1 CSA_VREF pixel
xPix6203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[62] VREF PIX_IN[6203] NB2 NB1 CSA_VREF pixel
xPix6204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[62] VREF PIX_IN[6204] NB2 NB1 CSA_VREF pixel
xPix6205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[62] VREF PIX_IN[6205] NB2 NB1 CSA_VREF pixel
xPix6206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[62] VREF PIX_IN[6206] NB2 NB1 CSA_VREF pixel
xPix6207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[62] VREF PIX_IN[6207] NB2 NB1 CSA_VREF pixel
xPix6208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[62] VREF PIX_IN[6208] NB2 NB1 CSA_VREF pixel
xPix6209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[62] VREF PIX_IN[6209] NB2 NB1 CSA_VREF pixel
xPix6210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[62] VREF PIX_IN[6210] NB2 NB1 CSA_VREF pixel
xPix6211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[62] VREF PIX_IN[6211] NB2 NB1 CSA_VREF pixel
xPix6212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[62] VREF PIX_IN[6212] NB2 NB1 CSA_VREF pixel
xPix6213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[62] VREF PIX_IN[6213] NB2 NB1 CSA_VREF pixel
xPix6214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[62] VREF PIX_IN[6214] NB2 NB1 CSA_VREF pixel
xPix6215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[62] VREF PIX_IN[6215] NB2 NB1 CSA_VREF pixel
xPix6216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[62] VREF PIX_IN[6216] NB2 NB1 CSA_VREF pixel
xPix6217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[62] VREF PIX_IN[6217] NB2 NB1 CSA_VREF pixel
xPix6218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[62] VREF PIX_IN[6218] NB2 NB1 CSA_VREF pixel
xPix6219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[62] VREF PIX_IN[6219] NB2 NB1 CSA_VREF pixel
xPix6220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[62] VREF PIX_IN[6220] NB2 NB1 CSA_VREF pixel
xPix6221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[62] VREF PIX_IN[6221] NB2 NB1 CSA_VREF pixel
xPix6222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[62] VREF PIX_IN[6222] NB2 NB1 CSA_VREF pixel
xPix6223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[62] VREF PIX_IN[6223] NB2 NB1 CSA_VREF pixel
xPix6224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[62] VREF PIX_IN[6224] NB2 NB1 CSA_VREF pixel
xPix6225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[62] VREF PIX_IN[6225] NB2 NB1 CSA_VREF pixel
xPix6226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[62] VREF PIX_IN[6226] NB2 NB1 CSA_VREF pixel
xPix6227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[62] VREF PIX_IN[6227] NB2 NB1 CSA_VREF pixel
xPix6228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[62] VREF PIX_IN[6228] NB2 NB1 CSA_VREF pixel
xPix6229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[62] VREF PIX_IN[6229] NB2 NB1 CSA_VREF pixel
xPix6230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[62] VREF PIX_IN[6230] NB2 NB1 CSA_VREF pixel
xPix6231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[62] VREF PIX_IN[6231] NB2 NB1 CSA_VREF pixel
xPix6232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[62] VREF PIX_IN[6232] NB2 NB1 CSA_VREF pixel
xPix6233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[62] VREF PIX_IN[6233] NB2 NB1 CSA_VREF pixel
xPix6234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[62] VREF PIX_IN[6234] NB2 NB1 CSA_VREF pixel
xPix6235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[62] VREF PIX_IN[6235] NB2 NB1 CSA_VREF pixel
xPix6236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[62] VREF PIX_IN[6236] NB2 NB1 CSA_VREF pixel
xPix6237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[62] VREF PIX_IN[6237] NB2 NB1 CSA_VREF pixel
xPix6238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[62] VREF PIX_IN[6238] NB2 NB1 CSA_VREF pixel
xPix6239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[62] VREF PIX_IN[6239] NB2 NB1 CSA_VREF pixel
xPix6240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[62] VREF PIX_IN[6240] NB2 NB1 CSA_VREF pixel
xPix6241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[62] VREF PIX_IN[6241] NB2 NB1 CSA_VREF pixel
xPix6242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[62] VREF PIX_IN[6242] NB2 NB1 CSA_VREF pixel
xPix6243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[62] VREF PIX_IN[6243] NB2 NB1 CSA_VREF pixel
xPix6244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[62] VREF PIX_IN[6244] NB2 NB1 CSA_VREF pixel
xPix6245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[62] VREF PIX_IN[6245] NB2 NB1 CSA_VREF pixel
xPix6246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[62] VREF PIX_IN[6246] NB2 NB1 CSA_VREF pixel
xPix6247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[62] VREF PIX_IN[6247] NB2 NB1 CSA_VREF pixel
xPix6248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[62] VREF PIX_IN[6248] NB2 NB1 CSA_VREF pixel
xPix6249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[62] VREF PIX_IN[6249] NB2 NB1 CSA_VREF pixel
xPix6250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[62] VREF PIX_IN[6250] NB2 NB1 CSA_VREF pixel
xPix6251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[62] VREF PIX_IN[6251] NB2 NB1 CSA_VREF pixel
xPix6252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[62] VREF PIX_IN[6252] NB2 NB1 CSA_VREF pixel
xPix6253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[62] VREF PIX_IN[6253] NB2 NB1 CSA_VREF pixel
xPix6254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[62] VREF PIX_IN[6254] NB2 NB1 CSA_VREF pixel
xPix6255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[62] VREF PIX_IN[6255] NB2 NB1 CSA_VREF pixel
xPix6256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[62] VREF PIX_IN[6256] NB2 NB1 CSA_VREF pixel
xPix6257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[62] VREF PIX_IN[6257] NB2 NB1 CSA_VREF pixel
xPix6258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[62] VREF PIX_IN[6258] NB2 NB1 CSA_VREF pixel
xPix6259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[62] VREF PIX_IN[6259] NB2 NB1 CSA_VREF pixel
xPix6260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[62] VREF PIX_IN[6260] NB2 NB1 CSA_VREF pixel
xPix6261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[62] VREF PIX_IN[6261] NB2 NB1 CSA_VREF pixel
xPix6262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[62] VREF PIX_IN[6262] NB2 NB1 CSA_VREF pixel
xPix6263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[62] VREF PIX_IN[6263] NB2 NB1 CSA_VREF pixel
xPix6264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[62] VREF PIX_IN[6264] NB2 NB1 CSA_VREF pixel
xPix6265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[62] VREF PIX_IN[6265] NB2 NB1 CSA_VREF pixel
xPix6266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[62] VREF PIX_IN[6266] NB2 NB1 CSA_VREF pixel
xPix6267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[62] VREF PIX_IN[6267] NB2 NB1 CSA_VREF pixel
xPix6268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[62] VREF PIX_IN[6268] NB2 NB1 CSA_VREF pixel
xPix6269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[62] VREF PIX_IN[6269] NB2 NB1 CSA_VREF pixel
xPix6270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[62] VREF PIX_IN[6270] NB2 NB1 CSA_VREF pixel
xPix6271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[62] VREF PIX_IN[6271] NB2 NB1 CSA_VREF pixel
xPix6272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[62] VREF PIX_IN[6272] NB2 NB1 CSA_VREF pixel
xPix6273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[62] VREF PIX_IN[6273] NB2 NB1 CSA_VREF pixel
xPix6274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[62] VREF PIX_IN[6274] NB2 NB1 CSA_VREF pixel
xPix6275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[62] VREF PIX_IN[6275] NB2 NB1 CSA_VREF pixel
xPix6276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[62] VREF PIX_IN[6276] NB2 NB1 CSA_VREF pixel
xPix6277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[62] VREF PIX_IN[6277] NB2 NB1 CSA_VREF pixel
xPix6278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[62] VREF PIX_IN[6278] NB2 NB1 CSA_VREF pixel
xPix6279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[62] VREF PIX_IN[6279] NB2 NB1 CSA_VREF pixel
xPix6280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[62] VREF PIX_IN[6280] NB2 NB1 CSA_VREF pixel
xPix6281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[62] VREF PIX_IN[6281] NB2 NB1 CSA_VREF pixel
xPix6282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[62] VREF PIX_IN[6282] NB2 NB1 CSA_VREF pixel
xPix6283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[62] VREF PIX_IN[6283] NB2 NB1 CSA_VREF pixel
xPix6284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[62] VREF PIX_IN[6284] NB2 NB1 CSA_VREF pixel
xPix6285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[62] VREF PIX_IN[6285] NB2 NB1 CSA_VREF pixel
xPix6286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[62] VREF PIX_IN[6286] NB2 NB1 CSA_VREF pixel
xPix6287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[62] VREF PIX_IN[6287] NB2 NB1 CSA_VREF pixel
xPix6288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[62] VREF PIX_IN[6288] NB2 NB1 CSA_VREF pixel
xPix6289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[62] VREF PIX_IN[6289] NB2 NB1 CSA_VREF pixel
xPix6290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[62] VREF PIX_IN[6290] NB2 NB1 CSA_VREF pixel
xPix6291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[62] VREF PIX_IN[6291] NB2 NB1 CSA_VREF pixel
xPix6292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[62] VREF PIX_IN[6292] NB2 NB1 CSA_VREF pixel
xPix6293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[62] VREF PIX_IN[6293] NB2 NB1 CSA_VREF pixel
xPix6294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[62] VREF PIX_IN[6294] NB2 NB1 CSA_VREF pixel
xPix6295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[62] VREF PIX_IN[6295] NB2 NB1 CSA_VREF pixel
xPix6296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[62] VREF PIX_IN[6296] NB2 NB1 CSA_VREF pixel
xPix6297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[62] VREF PIX_IN[6297] NB2 NB1 CSA_VREF pixel
xPix6298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[62] VREF PIX_IN[6298] NB2 NB1 CSA_VREF pixel
xPix6299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[62] VREF PIX_IN[6299] NB2 NB1 CSA_VREF pixel
xPix6300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[63] VREF PIX_IN[6300] NB2 NB1 CSA_VREF pixel
xPix6301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[63] VREF PIX_IN[6301] NB2 NB1 CSA_VREF pixel
xPix6302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[63] VREF PIX_IN[6302] NB2 NB1 CSA_VREF pixel
xPix6303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[63] VREF PIX_IN[6303] NB2 NB1 CSA_VREF pixel
xPix6304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[63] VREF PIX_IN[6304] NB2 NB1 CSA_VREF pixel
xPix6305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[63] VREF PIX_IN[6305] NB2 NB1 CSA_VREF pixel
xPix6306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[63] VREF PIX_IN[6306] NB2 NB1 CSA_VREF pixel
xPix6307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[63] VREF PIX_IN[6307] NB2 NB1 CSA_VREF pixel
xPix6308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[63] VREF PIX_IN[6308] NB2 NB1 CSA_VREF pixel
xPix6309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[63] VREF PIX_IN[6309] NB2 NB1 CSA_VREF pixel
xPix6310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[63] VREF PIX_IN[6310] NB2 NB1 CSA_VREF pixel
xPix6311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[63] VREF PIX_IN[6311] NB2 NB1 CSA_VREF pixel
xPix6312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[63] VREF PIX_IN[6312] NB2 NB1 CSA_VREF pixel
xPix6313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[63] VREF PIX_IN[6313] NB2 NB1 CSA_VREF pixel
xPix6314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[63] VREF PIX_IN[6314] NB2 NB1 CSA_VREF pixel
xPix6315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[63] VREF PIX_IN[6315] NB2 NB1 CSA_VREF pixel
xPix6316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[63] VREF PIX_IN[6316] NB2 NB1 CSA_VREF pixel
xPix6317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[63] VREF PIX_IN[6317] NB2 NB1 CSA_VREF pixel
xPix6318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[63] VREF PIX_IN[6318] NB2 NB1 CSA_VREF pixel
xPix6319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[63] VREF PIX_IN[6319] NB2 NB1 CSA_VREF pixel
xPix6320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[63] VREF PIX_IN[6320] NB2 NB1 CSA_VREF pixel
xPix6321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[63] VREF PIX_IN[6321] NB2 NB1 CSA_VREF pixel
xPix6322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[63] VREF PIX_IN[6322] NB2 NB1 CSA_VREF pixel
xPix6323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[63] VREF PIX_IN[6323] NB2 NB1 CSA_VREF pixel
xPix6324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[63] VREF PIX_IN[6324] NB2 NB1 CSA_VREF pixel
xPix6325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[63] VREF PIX_IN[6325] NB2 NB1 CSA_VREF pixel
xPix6326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[63] VREF PIX_IN[6326] NB2 NB1 CSA_VREF pixel
xPix6327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[63] VREF PIX_IN[6327] NB2 NB1 CSA_VREF pixel
xPix6328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[63] VREF PIX_IN[6328] NB2 NB1 CSA_VREF pixel
xPix6329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[63] VREF PIX_IN[6329] NB2 NB1 CSA_VREF pixel
xPix6330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[63] VREF PIX_IN[6330] NB2 NB1 CSA_VREF pixel
xPix6331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[63] VREF PIX_IN[6331] NB2 NB1 CSA_VREF pixel
xPix6332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[63] VREF PIX_IN[6332] NB2 NB1 CSA_VREF pixel
xPix6333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[63] VREF PIX_IN[6333] NB2 NB1 CSA_VREF pixel
xPix6334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[63] VREF PIX_IN[6334] NB2 NB1 CSA_VREF pixel
xPix6335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[63] VREF PIX_IN[6335] NB2 NB1 CSA_VREF pixel
xPix6336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[63] VREF PIX_IN[6336] NB2 NB1 CSA_VREF pixel
xPix6337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[63] VREF PIX_IN[6337] NB2 NB1 CSA_VREF pixel
xPix6338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[63] VREF PIX_IN[6338] NB2 NB1 CSA_VREF pixel
xPix6339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[63] VREF PIX_IN[6339] NB2 NB1 CSA_VREF pixel
xPix6340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[63] VREF PIX_IN[6340] NB2 NB1 CSA_VREF pixel
xPix6341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[63] VREF PIX_IN[6341] NB2 NB1 CSA_VREF pixel
xPix6342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[63] VREF PIX_IN[6342] NB2 NB1 CSA_VREF pixel
xPix6343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[63] VREF PIX_IN[6343] NB2 NB1 CSA_VREF pixel
xPix6344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[63] VREF PIX_IN[6344] NB2 NB1 CSA_VREF pixel
xPix6345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[63] VREF PIX_IN[6345] NB2 NB1 CSA_VREF pixel
xPix6346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[63] VREF PIX_IN[6346] NB2 NB1 CSA_VREF pixel
xPix6347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[63] VREF PIX_IN[6347] NB2 NB1 CSA_VREF pixel
xPix6348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[63] VREF PIX_IN[6348] NB2 NB1 CSA_VREF pixel
xPix6349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[63] VREF PIX_IN[6349] NB2 NB1 CSA_VREF pixel
xPix6350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[63] VREF PIX_IN[6350] NB2 NB1 CSA_VREF pixel
xPix6351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[63] VREF PIX_IN[6351] NB2 NB1 CSA_VREF pixel
xPix6352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[63] VREF PIX_IN[6352] NB2 NB1 CSA_VREF pixel
xPix6353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[63] VREF PIX_IN[6353] NB2 NB1 CSA_VREF pixel
xPix6354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[63] VREF PIX_IN[6354] NB2 NB1 CSA_VREF pixel
xPix6355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[63] VREF PIX_IN[6355] NB2 NB1 CSA_VREF pixel
xPix6356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[63] VREF PIX_IN[6356] NB2 NB1 CSA_VREF pixel
xPix6357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[63] VREF PIX_IN[6357] NB2 NB1 CSA_VREF pixel
xPix6358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[63] VREF PIX_IN[6358] NB2 NB1 CSA_VREF pixel
xPix6359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[63] VREF PIX_IN[6359] NB2 NB1 CSA_VREF pixel
xPix6360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[63] VREF PIX_IN[6360] NB2 NB1 CSA_VREF pixel
xPix6361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[63] VREF PIX_IN[6361] NB2 NB1 CSA_VREF pixel
xPix6362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[63] VREF PIX_IN[6362] NB2 NB1 CSA_VREF pixel
xPix6363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[63] VREF PIX_IN[6363] NB2 NB1 CSA_VREF pixel
xPix6364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[63] VREF PIX_IN[6364] NB2 NB1 CSA_VREF pixel
xPix6365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[63] VREF PIX_IN[6365] NB2 NB1 CSA_VREF pixel
xPix6366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[63] VREF PIX_IN[6366] NB2 NB1 CSA_VREF pixel
xPix6367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[63] VREF PIX_IN[6367] NB2 NB1 CSA_VREF pixel
xPix6368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[63] VREF PIX_IN[6368] NB2 NB1 CSA_VREF pixel
xPix6369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[63] VREF PIX_IN[6369] NB2 NB1 CSA_VREF pixel
xPix6370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[63] VREF PIX_IN[6370] NB2 NB1 CSA_VREF pixel
xPix6371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[63] VREF PIX_IN[6371] NB2 NB1 CSA_VREF pixel
xPix6372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[63] VREF PIX_IN[6372] NB2 NB1 CSA_VREF pixel
xPix6373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[63] VREF PIX_IN[6373] NB2 NB1 CSA_VREF pixel
xPix6374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[63] VREF PIX_IN[6374] NB2 NB1 CSA_VREF pixel
xPix6375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[63] VREF PIX_IN[6375] NB2 NB1 CSA_VREF pixel
xPix6376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[63] VREF PIX_IN[6376] NB2 NB1 CSA_VREF pixel
xPix6377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[63] VREF PIX_IN[6377] NB2 NB1 CSA_VREF pixel
xPix6378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[63] VREF PIX_IN[6378] NB2 NB1 CSA_VREF pixel
xPix6379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[63] VREF PIX_IN[6379] NB2 NB1 CSA_VREF pixel
xPix6380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[63] VREF PIX_IN[6380] NB2 NB1 CSA_VREF pixel
xPix6381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[63] VREF PIX_IN[6381] NB2 NB1 CSA_VREF pixel
xPix6382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[63] VREF PIX_IN[6382] NB2 NB1 CSA_VREF pixel
xPix6383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[63] VREF PIX_IN[6383] NB2 NB1 CSA_VREF pixel
xPix6384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[63] VREF PIX_IN[6384] NB2 NB1 CSA_VREF pixel
xPix6385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[63] VREF PIX_IN[6385] NB2 NB1 CSA_VREF pixel
xPix6386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[63] VREF PIX_IN[6386] NB2 NB1 CSA_VREF pixel
xPix6387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[63] VREF PIX_IN[6387] NB2 NB1 CSA_VREF pixel
xPix6388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[63] VREF PIX_IN[6388] NB2 NB1 CSA_VREF pixel
xPix6389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[63] VREF PIX_IN[6389] NB2 NB1 CSA_VREF pixel
xPix6390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[63] VREF PIX_IN[6390] NB2 NB1 CSA_VREF pixel
xPix6391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[63] VREF PIX_IN[6391] NB2 NB1 CSA_VREF pixel
xPix6392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[63] VREF PIX_IN[6392] NB2 NB1 CSA_VREF pixel
xPix6393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[63] VREF PIX_IN[6393] NB2 NB1 CSA_VREF pixel
xPix6394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[63] VREF PIX_IN[6394] NB2 NB1 CSA_VREF pixel
xPix6395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[63] VREF PIX_IN[6395] NB2 NB1 CSA_VREF pixel
xPix6396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[63] VREF PIX_IN[6396] NB2 NB1 CSA_VREF pixel
xPix6397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[63] VREF PIX_IN[6397] NB2 NB1 CSA_VREF pixel
xPix6398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[63] VREF PIX_IN[6398] NB2 NB1 CSA_VREF pixel
xPix6399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[63] VREF PIX_IN[6399] NB2 NB1 CSA_VREF pixel
xPix6400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[64] VREF PIX_IN[6400] NB2 NB1 CSA_VREF pixel
xPix6401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[64] VREF PIX_IN[6401] NB2 NB1 CSA_VREF pixel
xPix6402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[64] VREF PIX_IN[6402] NB2 NB1 CSA_VREF pixel
xPix6403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[64] VREF PIX_IN[6403] NB2 NB1 CSA_VREF pixel
xPix6404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[64] VREF PIX_IN[6404] NB2 NB1 CSA_VREF pixel
xPix6405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[64] VREF PIX_IN[6405] NB2 NB1 CSA_VREF pixel
xPix6406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[64] VREF PIX_IN[6406] NB2 NB1 CSA_VREF pixel
xPix6407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[64] VREF PIX_IN[6407] NB2 NB1 CSA_VREF pixel
xPix6408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[64] VREF PIX_IN[6408] NB2 NB1 CSA_VREF pixel
xPix6409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[64] VREF PIX_IN[6409] NB2 NB1 CSA_VREF pixel
xPix6410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[64] VREF PIX_IN[6410] NB2 NB1 CSA_VREF pixel
xPix6411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[64] VREF PIX_IN[6411] NB2 NB1 CSA_VREF pixel
xPix6412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[64] VREF PIX_IN[6412] NB2 NB1 CSA_VREF pixel
xPix6413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[64] VREF PIX_IN[6413] NB2 NB1 CSA_VREF pixel
xPix6414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[64] VREF PIX_IN[6414] NB2 NB1 CSA_VREF pixel
xPix6415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[64] VREF PIX_IN[6415] NB2 NB1 CSA_VREF pixel
xPix6416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[64] VREF PIX_IN[6416] NB2 NB1 CSA_VREF pixel
xPix6417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[64] VREF PIX_IN[6417] NB2 NB1 CSA_VREF pixel
xPix6418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[64] VREF PIX_IN[6418] NB2 NB1 CSA_VREF pixel
xPix6419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[64] VREF PIX_IN[6419] NB2 NB1 CSA_VREF pixel
xPix6420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[64] VREF PIX_IN[6420] NB2 NB1 CSA_VREF pixel
xPix6421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[64] VREF PIX_IN[6421] NB2 NB1 CSA_VREF pixel
xPix6422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[64] VREF PIX_IN[6422] NB2 NB1 CSA_VREF pixel
xPix6423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[64] VREF PIX_IN[6423] NB2 NB1 CSA_VREF pixel
xPix6424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[64] VREF PIX_IN[6424] NB2 NB1 CSA_VREF pixel
xPix6425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[64] VREF PIX_IN[6425] NB2 NB1 CSA_VREF pixel
xPix6426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[64] VREF PIX_IN[6426] NB2 NB1 CSA_VREF pixel
xPix6427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[64] VREF PIX_IN[6427] NB2 NB1 CSA_VREF pixel
xPix6428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[64] VREF PIX_IN[6428] NB2 NB1 CSA_VREF pixel
xPix6429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[64] VREF PIX_IN[6429] NB2 NB1 CSA_VREF pixel
xPix6430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[64] VREF PIX_IN[6430] NB2 NB1 CSA_VREF pixel
xPix6431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[64] VREF PIX_IN[6431] NB2 NB1 CSA_VREF pixel
xPix6432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[64] VREF PIX_IN[6432] NB2 NB1 CSA_VREF pixel
xPix6433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[64] VREF PIX_IN[6433] NB2 NB1 CSA_VREF pixel
xPix6434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[64] VREF PIX_IN[6434] NB2 NB1 CSA_VREF pixel
xPix6435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[64] VREF PIX_IN[6435] NB2 NB1 CSA_VREF pixel
xPix6436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[64] VREF PIX_IN[6436] NB2 NB1 CSA_VREF pixel
xPix6437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[64] VREF PIX_IN[6437] NB2 NB1 CSA_VREF pixel
xPix6438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[64] VREF PIX_IN[6438] NB2 NB1 CSA_VREF pixel
xPix6439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[64] VREF PIX_IN[6439] NB2 NB1 CSA_VREF pixel
xPix6440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[64] VREF PIX_IN[6440] NB2 NB1 CSA_VREF pixel
xPix6441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[64] VREF PIX_IN[6441] NB2 NB1 CSA_VREF pixel
xPix6442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[64] VREF PIX_IN[6442] NB2 NB1 CSA_VREF pixel
xPix6443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[64] VREF PIX_IN[6443] NB2 NB1 CSA_VREF pixel
xPix6444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[64] VREF PIX_IN[6444] NB2 NB1 CSA_VREF pixel
xPix6445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[64] VREF PIX_IN[6445] NB2 NB1 CSA_VREF pixel
xPix6446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[64] VREF PIX_IN[6446] NB2 NB1 CSA_VREF pixel
xPix6447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[64] VREF PIX_IN[6447] NB2 NB1 CSA_VREF pixel
xPix6448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[64] VREF PIX_IN[6448] NB2 NB1 CSA_VREF pixel
xPix6449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[64] VREF PIX_IN[6449] NB2 NB1 CSA_VREF pixel
xPix6450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[64] VREF PIX_IN[6450] NB2 NB1 CSA_VREF pixel
xPix6451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[64] VREF PIX_IN[6451] NB2 NB1 CSA_VREF pixel
xPix6452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[64] VREF PIX_IN[6452] NB2 NB1 CSA_VREF pixel
xPix6453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[64] VREF PIX_IN[6453] NB2 NB1 CSA_VREF pixel
xPix6454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[64] VREF PIX_IN[6454] NB2 NB1 CSA_VREF pixel
xPix6455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[64] VREF PIX_IN[6455] NB2 NB1 CSA_VREF pixel
xPix6456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[64] VREF PIX_IN[6456] NB2 NB1 CSA_VREF pixel
xPix6457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[64] VREF PIX_IN[6457] NB2 NB1 CSA_VREF pixel
xPix6458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[64] VREF PIX_IN[6458] NB2 NB1 CSA_VREF pixel
xPix6459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[64] VREF PIX_IN[6459] NB2 NB1 CSA_VREF pixel
xPix6460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[64] VREF PIX_IN[6460] NB2 NB1 CSA_VREF pixel
xPix6461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[64] VREF PIX_IN[6461] NB2 NB1 CSA_VREF pixel
xPix6462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[64] VREF PIX_IN[6462] NB2 NB1 CSA_VREF pixel
xPix6463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[64] VREF PIX_IN[6463] NB2 NB1 CSA_VREF pixel
xPix6464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[64] VREF PIX_IN[6464] NB2 NB1 CSA_VREF pixel
xPix6465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[64] VREF PIX_IN[6465] NB2 NB1 CSA_VREF pixel
xPix6466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[64] VREF PIX_IN[6466] NB2 NB1 CSA_VREF pixel
xPix6467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[64] VREF PIX_IN[6467] NB2 NB1 CSA_VREF pixel
xPix6468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[64] VREF PIX_IN[6468] NB2 NB1 CSA_VREF pixel
xPix6469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[64] VREF PIX_IN[6469] NB2 NB1 CSA_VREF pixel
xPix6470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[64] VREF PIX_IN[6470] NB2 NB1 CSA_VREF pixel
xPix6471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[64] VREF PIX_IN[6471] NB2 NB1 CSA_VREF pixel
xPix6472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[64] VREF PIX_IN[6472] NB2 NB1 CSA_VREF pixel
xPix6473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[64] VREF PIX_IN[6473] NB2 NB1 CSA_VREF pixel
xPix6474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[64] VREF PIX_IN[6474] NB2 NB1 CSA_VREF pixel
xPix6475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[64] VREF PIX_IN[6475] NB2 NB1 CSA_VREF pixel
xPix6476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[64] VREF PIX_IN[6476] NB2 NB1 CSA_VREF pixel
xPix6477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[64] VREF PIX_IN[6477] NB2 NB1 CSA_VREF pixel
xPix6478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[64] VREF PIX_IN[6478] NB2 NB1 CSA_VREF pixel
xPix6479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[64] VREF PIX_IN[6479] NB2 NB1 CSA_VREF pixel
xPix6480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[64] VREF PIX_IN[6480] NB2 NB1 CSA_VREF pixel
xPix6481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[64] VREF PIX_IN[6481] NB2 NB1 CSA_VREF pixel
xPix6482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[64] VREF PIX_IN[6482] NB2 NB1 CSA_VREF pixel
xPix6483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[64] VREF PIX_IN[6483] NB2 NB1 CSA_VREF pixel
xPix6484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[64] VREF PIX_IN[6484] NB2 NB1 CSA_VREF pixel
xPix6485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[64] VREF PIX_IN[6485] NB2 NB1 CSA_VREF pixel
xPix6486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[64] VREF PIX_IN[6486] NB2 NB1 CSA_VREF pixel
xPix6487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[64] VREF PIX_IN[6487] NB2 NB1 CSA_VREF pixel
xPix6488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[64] VREF PIX_IN[6488] NB2 NB1 CSA_VREF pixel
xPix6489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[64] VREF PIX_IN[6489] NB2 NB1 CSA_VREF pixel
xPix6490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[64] VREF PIX_IN[6490] NB2 NB1 CSA_VREF pixel
xPix6491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[64] VREF PIX_IN[6491] NB2 NB1 CSA_VREF pixel
xPix6492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[64] VREF PIX_IN[6492] NB2 NB1 CSA_VREF pixel
xPix6493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[64] VREF PIX_IN[6493] NB2 NB1 CSA_VREF pixel
xPix6494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[64] VREF PIX_IN[6494] NB2 NB1 CSA_VREF pixel
xPix6495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[64] VREF PIX_IN[6495] NB2 NB1 CSA_VREF pixel
xPix6496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[64] VREF PIX_IN[6496] NB2 NB1 CSA_VREF pixel
xPix6497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[64] VREF PIX_IN[6497] NB2 NB1 CSA_VREF pixel
xPix6498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[64] VREF PIX_IN[6498] NB2 NB1 CSA_VREF pixel
xPix6499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[64] VREF PIX_IN[6499] NB2 NB1 CSA_VREF pixel
xPix6500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[65] VREF PIX_IN[6500] NB2 NB1 CSA_VREF pixel
xPix6501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[65] VREF PIX_IN[6501] NB2 NB1 CSA_VREF pixel
xPix6502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[65] VREF PIX_IN[6502] NB2 NB1 CSA_VREF pixel
xPix6503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[65] VREF PIX_IN[6503] NB2 NB1 CSA_VREF pixel
xPix6504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[65] VREF PIX_IN[6504] NB2 NB1 CSA_VREF pixel
xPix6505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[65] VREF PIX_IN[6505] NB2 NB1 CSA_VREF pixel
xPix6506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[65] VREF PIX_IN[6506] NB2 NB1 CSA_VREF pixel
xPix6507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[65] VREF PIX_IN[6507] NB2 NB1 CSA_VREF pixel
xPix6508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[65] VREF PIX_IN[6508] NB2 NB1 CSA_VREF pixel
xPix6509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[65] VREF PIX_IN[6509] NB2 NB1 CSA_VREF pixel
xPix6510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[65] VREF PIX_IN[6510] NB2 NB1 CSA_VREF pixel
xPix6511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[65] VREF PIX_IN[6511] NB2 NB1 CSA_VREF pixel
xPix6512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[65] VREF PIX_IN[6512] NB2 NB1 CSA_VREF pixel
xPix6513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[65] VREF PIX_IN[6513] NB2 NB1 CSA_VREF pixel
xPix6514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[65] VREF PIX_IN[6514] NB2 NB1 CSA_VREF pixel
xPix6515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[65] VREF PIX_IN[6515] NB2 NB1 CSA_VREF pixel
xPix6516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[65] VREF PIX_IN[6516] NB2 NB1 CSA_VREF pixel
xPix6517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[65] VREF PIX_IN[6517] NB2 NB1 CSA_VREF pixel
xPix6518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[65] VREF PIX_IN[6518] NB2 NB1 CSA_VREF pixel
xPix6519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[65] VREF PIX_IN[6519] NB2 NB1 CSA_VREF pixel
xPix6520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[65] VREF PIX_IN[6520] NB2 NB1 CSA_VREF pixel
xPix6521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[65] VREF PIX_IN[6521] NB2 NB1 CSA_VREF pixel
xPix6522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[65] VREF PIX_IN[6522] NB2 NB1 CSA_VREF pixel
xPix6523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[65] VREF PIX_IN[6523] NB2 NB1 CSA_VREF pixel
xPix6524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[65] VREF PIX_IN[6524] NB2 NB1 CSA_VREF pixel
xPix6525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[65] VREF PIX_IN[6525] NB2 NB1 CSA_VREF pixel
xPix6526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[65] VREF PIX_IN[6526] NB2 NB1 CSA_VREF pixel
xPix6527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[65] VREF PIX_IN[6527] NB2 NB1 CSA_VREF pixel
xPix6528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[65] VREF PIX_IN[6528] NB2 NB1 CSA_VREF pixel
xPix6529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[65] VREF PIX_IN[6529] NB2 NB1 CSA_VREF pixel
xPix6530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[65] VREF PIX_IN[6530] NB2 NB1 CSA_VREF pixel
xPix6531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[65] VREF PIX_IN[6531] NB2 NB1 CSA_VREF pixel
xPix6532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[65] VREF PIX_IN[6532] NB2 NB1 CSA_VREF pixel
xPix6533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[65] VREF PIX_IN[6533] NB2 NB1 CSA_VREF pixel
xPix6534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[65] VREF PIX_IN[6534] NB2 NB1 CSA_VREF pixel
xPix6535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[65] VREF PIX_IN[6535] NB2 NB1 CSA_VREF pixel
xPix6536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[65] VREF PIX_IN[6536] NB2 NB1 CSA_VREF pixel
xPix6537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[65] VREF PIX_IN[6537] NB2 NB1 CSA_VREF pixel
xPix6538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[65] VREF PIX_IN[6538] NB2 NB1 CSA_VREF pixel
xPix6539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[65] VREF PIX_IN[6539] NB2 NB1 CSA_VREF pixel
xPix6540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[65] VREF PIX_IN[6540] NB2 NB1 CSA_VREF pixel
xPix6541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[65] VREF PIX_IN[6541] NB2 NB1 CSA_VREF pixel
xPix6542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[65] VREF PIX_IN[6542] NB2 NB1 CSA_VREF pixel
xPix6543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[65] VREF PIX_IN[6543] NB2 NB1 CSA_VREF pixel
xPix6544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[65] VREF PIX_IN[6544] NB2 NB1 CSA_VREF pixel
xPix6545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[65] VREF PIX_IN[6545] NB2 NB1 CSA_VREF pixel
xPix6546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[65] VREF PIX_IN[6546] NB2 NB1 CSA_VREF pixel
xPix6547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[65] VREF PIX_IN[6547] NB2 NB1 CSA_VREF pixel
xPix6548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[65] VREF PIX_IN[6548] NB2 NB1 CSA_VREF pixel
xPix6549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[65] VREF PIX_IN[6549] NB2 NB1 CSA_VREF pixel
xPix6550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[65] VREF PIX_IN[6550] NB2 NB1 CSA_VREF pixel
xPix6551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[65] VREF PIX_IN[6551] NB2 NB1 CSA_VREF pixel
xPix6552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[65] VREF PIX_IN[6552] NB2 NB1 CSA_VREF pixel
xPix6553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[65] VREF PIX_IN[6553] NB2 NB1 CSA_VREF pixel
xPix6554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[65] VREF PIX_IN[6554] NB2 NB1 CSA_VREF pixel
xPix6555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[65] VREF PIX_IN[6555] NB2 NB1 CSA_VREF pixel
xPix6556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[65] VREF PIX_IN[6556] NB2 NB1 CSA_VREF pixel
xPix6557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[65] VREF PIX_IN[6557] NB2 NB1 CSA_VREF pixel
xPix6558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[65] VREF PIX_IN[6558] NB2 NB1 CSA_VREF pixel
xPix6559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[65] VREF PIX_IN[6559] NB2 NB1 CSA_VREF pixel
xPix6560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[65] VREF PIX_IN[6560] NB2 NB1 CSA_VREF pixel
xPix6561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[65] VREF PIX_IN[6561] NB2 NB1 CSA_VREF pixel
xPix6562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[65] VREF PIX_IN[6562] NB2 NB1 CSA_VREF pixel
xPix6563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[65] VREF PIX_IN[6563] NB2 NB1 CSA_VREF pixel
xPix6564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[65] VREF PIX_IN[6564] NB2 NB1 CSA_VREF pixel
xPix6565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[65] VREF PIX_IN[6565] NB2 NB1 CSA_VREF pixel
xPix6566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[65] VREF PIX_IN[6566] NB2 NB1 CSA_VREF pixel
xPix6567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[65] VREF PIX_IN[6567] NB2 NB1 CSA_VREF pixel
xPix6568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[65] VREF PIX_IN[6568] NB2 NB1 CSA_VREF pixel
xPix6569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[65] VREF PIX_IN[6569] NB2 NB1 CSA_VREF pixel
xPix6570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[65] VREF PIX_IN[6570] NB2 NB1 CSA_VREF pixel
xPix6571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[65] VREF PIX_IN[6571] NB2 NB1 CSA_VREF pixel
xPix6572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[65] VREF PIX_IN[6572] NB2 NB1 CSA_VREF pixel
xPix6573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[65] VREF PIX_IN[6573] NB2 NB1 CSA_VREF pixel
xPix6574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[65] VREF PIX_IN[6574] NB2 NB1 CSA_VREF pixel
xPix6575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[65] VREF PIX_IN[6575] NB2 NB1 CSA_VREF pixel
xPix6576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[65] VREF PIX_IN[6576] NB2 NB1 CSA_VREF pixel
xPix6577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[65] VREF PIX_IN[6577] NB2 NB1 CSA_VREF pixel
xPix6578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[65] VREF PIX_IN[6578] NB2 NB1 CSA_VREF pixel
xPix6579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[65] VREF PIX_IN[6579] NB2 NB1 CSA_VREF pixel
xPix6580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[65] VREF PIX_IN[6580] NB2 NB1 CSA_VREF pixel
xPix6581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[65] VREF PIX_IN[6581] NB2 NB1 CSA_VREF pixel
xPix6582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[65] VREF PIX_IN[6582] NB2 NB1 CSA_VREF pixel
xPix6583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[65] VREF PIX_IN[6583] NB2 NB1 CSA_VREF pixel
xPix6584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[65] VREF PIX_IN[6584] NB2 NB1 CSA_VREF pixel
xPix6585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[65] VREF PIX_IN[6585] NB2 NB1 CSA_VREF pixel
xPix6586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[65] VREF PIX_IN[6586] NB2 NB1 CSA_VREF pixel
xPix6587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[65] VREF PIX_IN[6587] NB2 NB1 CSA_VREF pixel
xPix6588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[65] VREF PIX_IN[6588] NB2 NB1 CSA_VREF pixel
xPix6589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[65] VREF PIX_IN[6589] NB2 NB1 CSA_VREF pixel
xPix6590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[65] VREF PIX_IN[6590] NB2 NB1 CSA_VREF pixel
xPix6591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[65] VREF PIX_IN[6591] NB2 NB1 CSA_VREF pixel
xPix6592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[65] VREF PIX_IN[6592] NB2 NB1 CSA_VREF pixel
xPix6593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[65] VREF PIX_IN[6593] NB2 NB1 CSA_VREF pixel
xPix6594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[65] VREF PIX_IN[6594] NB2 NB1 CSA_VREF pixel
xPix6595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[65] VREF PIX_IN[6595] NB2 NB1 CSA_VREF pixel
xPix6596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[65] VREF PIX_IN[6596] NB2 NB1 CSA_VREF pixel
xPix6597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[65] VREF PIX_IN[6597] NB2 NB1 CSA_VREF pixel
xPix6598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[65] VREF PIX_IN[6598] NB2 NB1 CSA_VREF pixel
xPix6599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[65] VREF PIX_IN[6599] NB2 NB1 CSA_VREF pixel
xPix6600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[66] VREF PIX_IN[6600] NB2 NB1 CSA_VREF pixel
xPix6601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[66] VREF PIX_IN[6601] NB2 NB1 CSA_VREF pixel
xPix6602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[66] VREF PIX_IN[6602] NB2 NB1 CSA_VREF pixel
xPix6603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[66] VREF PIX_IN[6603] NB2 NB1 CSA_VREF pixel
xPix6604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[66] VREF PIX_IN[6604] NB2 NB1 CSA_VREF pixel
xPix6605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[66] VREF PIX_IN[6605] NB2 NB1 CSA_VREF pixel
xPix6606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[66] VREF PIX_IN[6606] NB2 NB1 CSA_VREF pixel
xPix6607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[66] VREF PIX_IN[6607] NB2 NB1 CSA_VREF pixel
xPix6608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[66] VREF PIX_IN[6608] NB2 NB1 CSA_VREF pixel
xPix6609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[66] VREF PIX_IN[6609] NB2 NB1 CSA_VREF pixel
xPix6610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[66] VREF PIX_IN[6610] NB2 NB1 CSA_VREF pixel
xPix6611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[66] VREF PIX_IN[6611] NB2 NB1 CSA_VREF pixel
xPix6612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[66] VREF PIX_IN[6612] NB2 NB1 CSA_VREF pixel
xPix6613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[66] VREF PIX_IN[6613] NB2 NB1 CSA_VREF pixel
xPix6614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[66] VREF PIX_IN[6614] NB2 NB1 CSA_VREF pixel
xPix6615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[66] VREF PIX_IN[6615] NB2 NB1 CSA_VREF pixel
xPix6616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[66] VREF PIX_IN[6616] NB2 NB1 CSA_VREF pixel
xPix6617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[66] VREF PIX_IN[6617] NB2 NB1 CSA_VREF pixel
xPix6618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[66] VREF PIX_IN[6618] NB2 NB1 CSA_VREF pixel
xPix6619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[66] VREF PIX_IN[6619] NB2 NB1 CSA_VREF pixel
xPix6620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[66] VREF PIX_IN[6620] NB2 NB1 CSA_VREF pixel
xPix6621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[66] VREF PIX_IN[6621] NB2 NB1 CSA_VREF pixel
xPix6622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[66] VREF PIX_IN[6622] NB2 NB1 CSA_VREF pixel
xPix6623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[66] VREF PIX_IN[6623] NB2 NB1 CSA_VREF pixel
xPix6624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[66] VREF PIX_IN[6624] NB2 NB1 CSA_VREF pixel
xPix6625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[66] VREF PIX_IN[6625] NB2 NB1 CSA_VREF pixel
xPix6626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[66] VREF PIX_IN[6626] NB2 NB1 CSA_VREF pixel
xPix6627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[66] VREF PIX_IN[6627] NB2 NB1 CSA_VREF pixel
xPix6628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[66] VREF PIX_IN[6628] NB2 NB1 CSA_VREF pixel
xPix6629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[66] VREF PIX_IN[6629] NB2 NB1 CSA_VREF pixel
xPix6630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[66] VREF PIX_IN[6630] NB2 NB1 CSA_VREF pixel
xPix6631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[66] VREF PIX_IN[6631] NB2 NB1 CSA_VREF pixel
xPix6632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[66] VREF PIX_IN[6632] NB2 NB1 CSA_VREF pixel
xPix6633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[66] VREF PIX_IN[6633] NB2 NB1 CSA_VREF pixel
xPix6634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[66] VREF PIX_IN[6634] NB2 NB1 CSA_VREF pixel
xPix6635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[66] VREF PIX_IN[6635] NB2 NB1 CSA_VREF pixel
xPix6636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[66] VREF PIX_IN[6636] NB2 NB1 CSA_VREF pixel
xPix6637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[66] VREF PIX_IN[6637] NB2 NB1 CSA_VREF pixel
xPix6638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[66] VREF PIX_IN[6638] NB2 NB1 CSA_VREF pixel
xPix6639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[66] VREF PIX_IN[6639] NB2 NB1 CSA_VREF pixel
xPix6640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[66] VREF PIX_IN[6640] NB2 NB1 CSA_VREF pixel
xPix6641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[66] VREF PIX_IN[6641] NB2 NB1 CSA_VREF pixel
xPix6642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[66] VREF PIX_IN[6642] NB2 NB1 CSA_VREF pixel
xPix6643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[66] VREF PIX_IN[6643] NB2 NB1 CSA_VREF pixel
xPix6644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[66] VREF PIX_IN[6644] NB2 NB1 CSA_VREF pixel
xPix6645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[66] VREF PIX_IN[6645] NB2 NB1 CSA_VREF pixel
xPix6646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[66] VREF PIX_IN[6646] NB2 NB1 CSA_VREF pixel
xPix6647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[66] VREF PIX_IN[6647] NB2 NB1 CSA_VREF pixel
xPix6648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[66] VREF PIX_IN[6648] NB2 NB1 CSA_VREF pixel
xPix6649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[66] VREF PIX_IN[6649] NB2 NB1 CSA_VREF pixel
xPix6650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[66] VREF PIX_IN[6650] NB2 NB1 CSA_VREF pixel
xPix6651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[66] VREF PIX_IN[6651] NB2 NB1 CSA_VREF pixel
xPix6652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[66] VREF PIX_IN[6652] NB2 NB1 CSA_VREF pixel
xPix6653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[66] VREF PIX_IN[6653] NB2 NB1 CSA_VREF pixel
xPix6654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[66] VREF PIX_IN[6654] NB2 NB1 CSA_VREF pixel
xPix6655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[66] VREF PIX_IN[6655] NB2 NB1 CSA_VREF pixel
xPix6656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[66] VREF PIX_IN[6656] NB2 NB1 CSA_VREF pixel
xPix6657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[66] VREF PIX_IN[6657] NB2 NB1 CSA_VREF pixel
xPix6658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[66] VREF PIX_IN[6658] NB2 NB1 CSA_VREF pixel
xPix6659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[66] VREF PIX_IN[6659] NB2 NB1 CSA_VREF pixel
xPix6660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[66] VREF PIX_IN[6660] NB2 NB1 CSA_VREF pixel
xPix6661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[66] VREF PIX_IN[6661] NB2 NB1 CSA_VREF pixel
xPix6662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[66] VREF PIX_IN[6662] NB2 NB1 CSA_VREF pixel
xPix6663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[66] VREF PIX_IN[6663] NB2 NB1 CSA_VREF pixel
xPix6664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[66] VREF PIX_IN[6664] NB2 NB1 CSA_VREF pixel
xPix6665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[66] VREF PIX_IN[6665] NB2 NB1 CSA_VREF pixel
xPix6666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[66] VREF PIX_IN[6666] NB2 NB1 CSA_VREF pixel
xPix6667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[66] VREF PIX_IN[6667] NB2 NB1 CSA_VREF pixel
xPix6668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[66] VREF PIX_IN[6668] NB2 NB1 CSA_VREF pixel
xPix6669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[66] VREF PIX_IN[6669] NB2 NB1 CSA_VREF pixel
xPix6670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[66] VREF PIX_IN[6670] NB2 NB1 CSA_VREF pixel
xPix6671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[66] VREF PIX_IN[6671] NB2 NB1 CSA_VREF pixel
xPix6672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[66] VREF PIX_IN[6672] NB2 NB1 CSA_VREF pixel
xPix6673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[66] VREF PIX_IN[6673] NB2 NB1 CSA_VREF pixel
xPix6674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[66] VREF PIX_IN[6674] NB2 NB1 CSA_VREF pixel
xPix6675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[66] VREF PIX_IN[6675] NB2 NB1 CSA_VREF pixel
xPix6676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[66] VREF PIX_IN[6676] NB2 NB1 CSA_VREF pixel
xPix6677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[66] VREF PIX_IN[6677] NB2 NB1 CSA_VREF pixel
xPix6678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[66] VREF PIX_IN[6678] NB2 NB1 CSA_VREF pixel
xPix6679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[66] VREF PIX_IN[6679] NB2 NB1 CSA_VREF pixel
xPix6680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[66] VREF PIX_IN[6680] NB2 NB1 CSA_VREF pixel
xPix6681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[66] VREF PIX_IN[6681] NB2 NB1 CSA_VREF pixel
xPix6682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[66] VREF PIX_IN[6682] NB2 NB1 CSA_VREF pixel
xPix6683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[66] VREF PIX_IN[6683] NB2 NB1 CSA_VREF pixel
xPix6684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[66] VREF PIX_IN[6684] NB2 NB1 CSA_VREF pixel
xPix6685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[66] VREF PIX_IN[6685] NB2 NB1 CSA_VREF pixel
xPix6686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[66] VREF PIX_IN[6686] NB2 NB1 CSA_VREF pixel
xPix6687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[66] VREF PIX_IN[6687] NB2 NB1 CSA_VREF pixel
xPix6688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[66] VREF PIX_IN[6688] NB2 NB1 CSA_VREF pixel
xPix6689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[66] VREF PIX_IN[6689] NB2 NB1 CSA_VREF pixel
xPix6690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[66] VREF PIX_IN[6690] NB2 NB1 CSA_VREF pixel
xPix6691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[66] VREF PIX_IN[6691] NB2 NB1 CSA_VREF pixel
xPix6692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[66] VREF PIX_IN[6692] NB2 NB1 CSA_VREF pixel
xPix6693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[66] VREF PIX_IN[6693] NB2 NB1 CSA_VREF pixel
xPix6694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[66] VREF PIX_IN[6694] NB2 NB1 CSA_VREF pixel
xPix6695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[66] VREF PIX_IN[6695] NB2 NB1 CSA_VREF pixel
xPix6696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[66] VREF PIX_IN[6696] NB2 NB1 CSA_VREF pixel
xPix6697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[66] VREF PIX_IN[6697] NB2 NB1 CSA_VREF pixel
xPix6698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[66] VREF PIX_IN[6698] NB2 NB1 CSA_VREF pixel
xPix6699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[66] VREF PIX_IN[6699] NB2 NB1 CSA_VREF pixel
xPix6700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[67] VREF PIX_IN[6700] NB2 NB1 CSA_VREF pixel
xPix6701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[67] VREF PIX_IN[6701] NB2 NB1 CSA_VREF pixel
xPix6702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[67] VREF PIX_IN[6702] NB2 NB1 CSA_VREF pixel
xPix6703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[67] VREF PIX_IN[6703] NB2 NB1 CSA_VREF pixel
xPix6704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[67] VREF PIX_IN[6704] NB2 NB1 CSA_VREF pixel
xPix6705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[67] VREF PIX_IN[6705] NB2 NB1 CSA_VREF pixel
xPix6706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[67] VREF PIX_IN[6706] NB2 NB1 CSA_VREF pixel
xPix6707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[67] VREF PIX_IN[6707] NB2 NB1 CSA_VREF pixel
xPix6708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[67] VREF PIX_IN[6708] NB2 NB1 CSA_VREF pixel
xPix6709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[67] VREF PIX_IN[6709] NB2 NB1 CSA_VREF pixel
xPix6710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[67] VREF PIX_IN[6710] NB2 NB1 CSA_VREF pixel
xPix6711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[67] VREF PIX_IN[6711] NB2 NB1 CSA_VREF pixel
xPix6712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[67] VREF PIX_IN[6712] NB2 NB1 CSA_VREF pixel
xPix6713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[67] VREF PIX_IN[6713] NB2 NB1 CSA_VREF pixel
xPix6714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[67] VREF PIX_IN[6714] NB2 NB1 CSA_VREF pixel
xPix6715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[67] VREF PIX_IN[6715] NB2 NB1 CSA_VREF pixel
xPix6716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[67] VREF PIX_IN[6716] NB2 NB1 CSA_VREF pixel
xPix6717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[67] VREF PIX_IN[6717] NB2 NB1 CSA_VREF pixel
xPix6718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[67] VREF PIX_IN[6718] NB2 NB1 CSA_VREF pixel
xPix6719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[67] VREF PIX_IN[6719] NB2 NB1 CSA_VREF pixel
xPix6720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[67] VREF PIX_IN[6720] NB2 NB1 CSA_VREF pixel
xPix6721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[67] VREF PIX_IN[6721] NB2 NB1 CSA_VREF pixel
xPix6722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[67] VREF PIX_IN[6722] NB2 NB1 CSA_VREF pixel
xPix6723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[67] VREF PIX_IN[6723] NB2 NB1 CSA_VREF pixel
xPix6724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[67] VREF PIX_IN[6724] NB2 NB1 CSA_VREF pixel
xPix6725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[67] VREF PIX_IN[6725] NB2 NB1 CSA_VREF pixel
xPix6726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[67] VREF PIX_IN[6726] NB2 NB1 CSA_VREF pixel
xPix6727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[67] VREF PIX_IN[6727] NB2 NB1 CSA_VREF pixel
xPix6728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[67] VREF PIX_IN[6728] NB2 NB1 CSA_VREF pixel
xPix6729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[67] VREF PIX_IN[6729] NB2 NB1 CSA_VREF pixel
xPix6730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[67] VREF PIX_IN[6730] NB2 NB1 CSA_VREF pixel
xPix6731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[67] VREF PIX_IN[6731] NB2 NB1 CSA_VREF pixel
xPix6732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[67] VREF PIX_IN[6732] NB2 NB1 CSA_VREF pixel
xPix6733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[67] VREF PIX_IN[6733] NB2 NB1 CSA_VREF pixel
xPix6734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[67] VREF PIX_IN[6734] NB2 NB1 CSA_VREF pixel
xPix6735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[67] VREF PIX_IN[6735] NB2 NB1 CSA_VREF pixel
xPix6736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[67] VREF PIX_IN[6736] NB2 NB1 CSA_VREF pixel
xPix6737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[67] VREF PIX_IN[6737] NB2 NB1 CSA_VREF pixel
xPix6738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[67] VREF PIX_IN[6738] NB2 NB1 CSA_VREF pixel
xPix6739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[67] VREF PIX_IN[6739] NB2 NB1 CSA_VREF pixel
xPix6740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[67] VREF PIX_IN[6740] NB2 NB1 CSA_VREF pixel
xPix6741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[67] VREF PIX_IN[6741] NB2 NB1 CSA_VREF pixel
xPix6742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[67] VREF PIX_IN[6742] NB2 NB1 CSA_VREF pixel
xPix6743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[67] VREF PIX_IN[6743] NB2 NB1 CSA_VREF pixel
xPix6744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[67] VREF PIX_IN[6744] NB2 NB1 CSA_VREF pixel
xPix6745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[67] VREF PIX_IN[6745] NB2 NB1 CSA_VREF pixel
xPix6746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[67] VREF PIX_IN[6746] NB2 NB1 CSA_VREF pixel
xPix6747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[67] VREF PIX_IN[6747] NB2 NB1 CSA_VREF pixel
xPix6748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[67] VREF PIX_IN[6748] NB2 NB1 CSA_VREF pixel
xPix6749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[67] VREF PIX_IN[6749] NB2 NB1 CSA_VREF pixel
xPix6750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[67] VREF PIX_IN[6750] NB2 NB1 CSA_VREF pixel
xPix6751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[67] VREF PIX_IN[6751] NB2 NB1 CSA_VREF pixel
xPix6752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[67] VREF PIX_IN[6752] NB2 NB1 CSA_VREF pixel
xPix6753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[67] VREF PIX_IN[6753] NB2 NB1 CSA_VREF pixel
xPix6754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[67] VREF PIX_IN[6754] NB2 NB1 CSA_VREF pixel
xPix6755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[67] VREF PIX_IN[6755] NB2 NB1 CSA_VREF pixel
xPix6756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[67] VREF PIX_IN[6756] NB2 NB1 CSA_VREF pixel
xPix6757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[67] VREF PIX_IN[6757] NB2 NB1 CSA_VREF pixel
xPix6758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[67] VREF PIX_IN[6758] NB2 NB1 CSA_VREF pixel
xPix6759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[67] VREF PIX_IN[6759] NB2 NB1 CSA_VREF pixel
xPix6760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[67] VREF PIX_IN[6760] NB2 NB1 CSA_VREF pixel
xPix6761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[67] VREF PIX_IN[6761] NB2 NB1 CSA_VREF pixel
xPix6762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[67] VREF PIX_IN[6762] NB2 NB1 CSA_VREF pixel
xPix6763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[67] VREF PIX_IN[6763] NB2 NB1 CSA_VREF pixel
xPix6764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[67] VREF PIX_IN[6764] NB2 NB1 CSA_VREF pixel
xPix6765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[67] VREF PIX_IN[6765] NB2 NB1 CSA_VREF pixel
xPix6766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[67] VREF PIX_IN[6766] NB2 NB1 CSA_VREF pixel
xPix6767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[67] VREF PIX_IN[6767] NB2 NB1 CSA_VREF pixel
xPix6768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[67] VREF PIX_IN[6768] NB2 NB1 CSA_VREF pixel
xPix6769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[67] VREF PIX_IN[6769] NB2 NB1 CSA_VREF pixel
xPix6770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[67] VREF PIX_IN[6770] NB2 NB1 CSA_VREF pixel
xPix6771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[67] VREF PIX_IN[6771] NB2 NB1 CSA_VREF pixel
xPix6772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[67] VREF PIX_IN[6772] NB2 NB1 CSA_VREF pixel
xPix6773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[67] VREF PIX_IN[6773] NB2 NB1 CSA_VREF pixel
xPix6774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[67] VREF PIX_IN[6774] NB2 NB1 CSA_VREF pixel
xPix6775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[67] VREF PIX_IN[6775] NB2 NB1 CSA_VREF pixel
xPix6776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[67] VREF PIX_IN[6776] NB2 NB1 CSA_VREF pixel
xPix6777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[67] VREF PIX_IN[6777] NB2 NB1 CSA_VREF pixel
xPix6778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[67] VREF PIX_IN[6778] NB2 NB1 CSA_VREF pixel
xPix6779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[67] VREF PIX_IN[6779] NB2 NB1 CSA_VREF pixel
xPix6780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[67] VREF PIX_IN[6780] NB2 NB1 CSA_VREF pixel
xPix6781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[67] VREF PIX_IN[6781] NB2 NB1 CSA_VREF pixel
xPix6782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[67] VREF PIX_IN[6782] NB2 NB1 CSA_VREF pixel
xPix6783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[67] VREF PIX_IN[6783] NB2 NB1 CSA_VREF pixel
xPix6784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[67] VREF PIX_IN[6784] NB2 NB1 CSA_VREF pixel
xPix6785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[67] VREF PIX_IN[6785] NB2 NB1 CSA_VREF pixel
xPix6786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[67] VREF PIX_IN[6786] NB2 NB1 CSA_VREF pixel
xPix6787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[67] VREF PIX_IN[6787] NB2 NB1 CSA_VREF pixel
xPix6788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[67] VREF PIX_IN[6788] NB2 NB1 CSA_VREF pixel
xPix6789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[67] VREF PIX_IN[6789] NB2 NB1 CSA_VREF pixel
xPix6790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[67] VREF PIX_IN[6790] NB2 NB1 CSA_VREF pixel
xPix6791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[67] VREF PIX_IN[6791] NB2 NB1 CSA_VREF pixel
xPix6792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[67] VREF PIX_IN[6792] NB2 NB1 CSA_VREF pixel
xPix6793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[67] VREF PIX_IN[6793] NB2 NB1 CSA_VREF pixel
xPix6794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[67] VREF PIX_IN[6794] NB2 NB1 CSA_VREF pixel
xPix6795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[67] VREF PIX_IN[6795] NB2 NB1 CSA_VREF pixel
xPix6796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[67] VREF PIX_IN[6796] NB2 NB1 CSA_VREF pixel
xPix6797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[67] VREF PIX_IN[6797] NB2 NB1 CSA_VREF pixel
xPix6798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[67] VREF PIX_IN[6798] NB2 NB1 CSA_VREF pixel
xPix6799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[67] VREF PIX_IN[6799] NB2 NB1 CSA_VREF pixel
xPix6800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[68] VREF PIX_IN[6800] NB2 NB1 CSA_VREF pixel
xPix6801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[68] VREF PIX_IN[6801] NB2 NB1 CSA_VREF pixel
xPix6802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[68] VREF PIX_IN[6802] NB2 NB1 CSA_VREF pixel
xPix6803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[68] VREF PIX_IN[6803] NB2 NB1 CSA_VREF pixel
xPix6804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[68] VREF PIX_IN[6804] NB2 NB1 CSA_VREF pixel
xPix6805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[68] VREF PIX_IN[6805] NB2 NB1 CSA_VREF pixel
xPix6806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[68] VREF PIX_IN[6806] NB2 NB1 CSA_VREF pixel
xPix6807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[68] VREF PIX_IN[6807] NB2 NB1 CSA_VREF pixel
xPix6808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[68] VREF PIX_IN[6808] NB2 NB1 CSA_VREF pixel
xPix6809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[68] VREF PIX_IN[6809] NB2 NB1 CSA_VREF pixel
xPix6810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[68] VREF PIX_IN[6810] NB2 NB1 CSA_VREF pixel
xPix6811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[68] VREF PIX_IN[6811] NB2 NB1 CSA_VREF pixel
xPix6812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[68] VREF PIX_IN[6812] NB2 NB1 CSA_VREF pixel
xPix6813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[68] VREF PIX_IN[6813] NB2 NB1 CSA_VREF pixel
xPix6814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[68] VREF PIX_IN[6814] NB2 NB1 CSA_VREF pixel
xPix6815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[68] VREF PIX_IN[6815] NB2 NB1 CSA_VREF pixel
xPix6816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[68] VREF PIX_IN[6816] NB2 NB1 CSA_VREF pixel
xPix6817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[68] VREF PIX_IN[6817] NB2 NB1 CSA_VREF pixel
xPix6818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[68] VREF PIX_IN[6818] NB2 NB1 CSA_VREF pixel
xPix6819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[68] VREF PIX_IN[6819] NB2 NB1 CSA_VREF pixel
xPix6820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[68] VREF PIX_IN[6820] NB2 NB1 CSA_VREF pixel
xPix6821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[68] VREF PIX_IN[6821] NB2 NB1 CSA_VREF pixel
xPix6822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[68] VREF PIX_IN[6822] NB2 NB1 CSA_VREF pixel
xPix6823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[68] VREF PIX_IN[6823] NB2 NB1 CSA_VREF pixel
xPix6824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[68] VREF PIX_IN[6824] NB2 NB1 CSA_VREF pixel
xPix6825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[68] VREF PIX_IN[6825] NB2 NB1 CSA_VREF pixel
xPix6826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[68] VREF PIX_IN[6826] NB2 NB1 CSA_VREF pixel
xPix6827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[68] VREF PIX_IN[6827] NB2 NB1 CSA_VREF pixel
xPix6828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[68] VREF PIX_IN[6828] NB2 NB1 CSA_VREF pixel
xPix6829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[68] VREF PIX_IN[6829] NB2 NB1 CSA_VREF pixel
xPix6830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[68] VREF PIX_IN[6830] NB2 NB1 CSA_VREF pixel
xPix6831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[68] VREF PIX_IN[6831] NB2 NB1 CSA_VREF pixel
xPix6832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[68] VREF PIX_IN[6832] NB2 NB1 CSA_VREF pixel
xPix6833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[68] VREF PIX_IN[6833] NB2 NB1 CSA_VREF pixel
xPix6834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[68] VREF PIX_IN[6834] NB2 NB1 CSA_VREF pixel
xPix6835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[68] VREF PIX_IN[6835] NB2 NB1 CSA_VREF pixel
xPix6836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[68] VREF PIX_IN[6836] NB2 NB1 CSA_VREF pixel
xPix6837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[68] VREF PIX_IN[6837] NB2 NB1 CSA_VREF pixel
xPix6838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[68] VREF PIX_IN[6838] NB2 NB1 CSA_VREF pixel
xPix6839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[68] VREF PIX_IN[6839] NB2 NB1 CSA_VREF pixel
xPix6840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[68] VREF PIX_IN[6840] NB2 NB1 CSA_VREF pixel
xPix6841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[68] VREF PIX_IN[6841] NB2 NB1 CSA_VREF pixel
xPix6842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[68] VREF PIX_IN[6842] NB2 NB1 CSA_VREF pixel
xPix6843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[68] VREF PIX_IN[6843] NB2 NB1 CSA_VREF pixel
xPix6844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[68] VREF PIX_IN[6844] NB2 NB1 CSA_VREF pixel
xPix6845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[68] VREF PIX_IN[6845] NB2 NB1 CSA_VREF pixel
xPix6846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[68] VREF PIX_IN[6846] NB2 NB1 CSA_VREF pixel
xPix6847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[68] VREF PIX_IN[6847] NB2 NB1 CSA_VREF pixel
xPix6848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[68] VREF PIX_IN[6848] NB2 NB1 CSA_VREF pixel
xPix6849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[68] VREF PIX_IN[6849] NB2 NB1 CSA_VREF pixel
xPix6850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[68] VREF PIX_IN[6850] NB2 NB1 CSA_VREF pixel
xPix6851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[68] VREF PIX_IN[6851] NB2 NB1 CSA_VREF pixel
xPix6852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[68] VREF PIX_IN[6852] NB2 NB1 CSA_VREF pixel
xPix6853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[68] VREF PIX_IN[6853] NB2 NB1 CSA_VREF pixel
xPix6854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[68] VREF PIX_IN[6854] NB2 NB1 CSA_VREF pixel
xPix6855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[68] VREF PIX_IN[6855] NB2 NB1 CSA_VREF pixel
xPix6856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[68] VREF PIX_IN[6856] NB2 NB1 CSA_VREF pixel
xPix6857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[68] VREF PIX_IN[6857] NB2 NB1 CSA_VREF pixel
xPix6858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[68] VREF PIX_IN[6858] NB2 NB1 CSA_VREF pixel
xPix6859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[68] VREF PIX_IN[6859] NB2 NB1 CSA_VREF pixel
xPix6860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[68] VREF PIX_IN[6860] NB2 NB1 CSA_VREF pixel
xPix6861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[68] VREF PIX_IN[6861] NB2 NB1 CSA_VREF pixel
xPix6862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[68] VREF PIX_IN[6862] NB2 NB1 CSA_VREF pixel
xPix6863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[68] VREF PIX_IN[6863] NB2 NB1 CSA_VREF pixel
xPix6864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[68] VREF PIX_IN[6864] NB2 NB1 CSA_VREF pixel
xPix6865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[68] VREF PIX_IN[6865] NB2 NB1 CSA_VREF pixel
xPix6866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[68] VREF PIX_IN[6866] NB2 NB1 CSA_VREF pixel
xPix6867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[68] VREF PIX_IN[6867] NB2 NB1 CSA_VREF pixel
xPix6868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[68] VREF PIX_IN[6868] NB2 NB1 CSA_VREF pixel
xPix6869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[68] VREF PIX_IN[6869] NB2 NB1 CSA_VREF pixel
xPix6870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[68] VREF PIX_IN[6870] NB2 NB1 CSA_VREF pixel
xPix6871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[68] VREF PIX_IN[6871] NB2 NB1 CSA_VREF pixel
xPix6872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[68] VREF PIX_IN[6872] NB2 NB1 CSA_VREF pixel
xPix6873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[68] VREF PIX_IN[6873] NB2 NB1 CSA_VREF pixel
xPix6874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[68] VREF PIX_IN[6874] NB2 NB1 CSA_VREF pixel
xPix6875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[68] VREF PIX_IN[6875] NB2 NB1 CSA_VREF pixel
xPix6876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[68] VREF PIX_IN[6876] NB2 NB1 CSA_VREF pixel
xPix6877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[68] VREF PIX_IN[6877] NB2 NB1 CSA_VREF pixel
xPix6878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[68] VREF PIX_IN[6878] NB2 NB1 CSA_VREF pixel
xPix6879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[68] VREF PIX_IN[6879] NB2 NB1 CSA_VREF pixel
xPix6880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[68] VREF PIX_IN[6880] NB2 NB1 CSA_VREF pixel
xPix6881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[68] VREF PIX_IN[6881] NB2 NB1 CSA_VREF pixel
xPix6882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[68] VREF PIX_IN[6882] NB2 NB1 CSA_VREF pixel
xPix6883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[68] VREF PIX_IN[6883] NB2 NB1 CSA_VREF pixel
xPix6884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[68] VREF PIX_IN[6884] NB2 NB1 CSA_VREF pixel
xPix6885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[68] VREF PIX_IN[6885] NB2 NB1 CSA_VREF pixel
xPix6886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[68] VREF PIX_IN[6886] NB2 NB1 CSA_VREF pixel
xPix6887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[68] VREF PIX_IN[6887] NB2 NB1 CSA_VREF pixel
xPix6888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[68] VREF PIX_IN[6888] NB2 NB1 CSA_VREF pixel
xPix6889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[68] VREF PIX_IN[6889] NB2 NB1 CSA_VREF pixel
xPix6890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[68] VREF PIX_IN[6890] NB2 NB1 CSA_VREF pixel
xPix6891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[68] VREF PIX_IN[6891] NB2 NB1 CSA_VREF pixel
xPix6892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[68] VREF PIX_IN[6892] NB2 NB1 CSA_VREF pixel
xPix6893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[68] VREF PIX_IN[6893] NB2 NB1 CSA_VREF pixel
xPix6894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[68] VREF PIX_IN[6894] NB2 NB1 CSA_VREF pixel
xPix6895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[68] VREF PIX_IN[6895] NB2 NB1 CSA_VREF pixel
xPix6896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[68] VREF PIX_IN[6896] NB2 NB1 CSA_VREF pixel
xPix6897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[68] VREF PIX_IN[6897] NB2 NB1 CSA_VREF pixel
xPix6898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[68] VREF PIX_IN[6898] NB2 NB1 CSA_VREF pixel
xPix6899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[68] VREF PIX_IN[6899] NB2 NB1 CSA_VREF pixel
xPix6900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[69] VREF PIX_IN[6900] NB2 NB1 CSA_VREF pixel
xPix6901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[69] VREF PIX_IN[6901] NB2 NB1 CSA_VREF pixel
xPix6902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[69] VREF PIX_IN[6902] NB2 NB1 CSA_VREF pixel
xPix6903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[69] VREF PIX_IN[6903] NB2 NB1 CSA_VREF pixel
xPix6904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[69] VREF PIX_IN[6904] NB2 NB1 CSA_VREF pixel
xPix6905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[69] VREF PIX_IN[6905] NB2 NB1 CSA_VREF pixel
xPix6906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[69] VREF PIX_IN[6906] NB2 NB1 CSA_VREF pixel
xPix6907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[69] VREF PIX_IN[6907] NB2 NB1 CSA_VREF pixel
xPix6908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[69] VREF PIX_IN[6908] NB2 NB1 CSA_VREF pixel
xPix6909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[69] VREF PIX_IN[6909] NB2 NB1 CSA_VREF pixel
xPix6910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[69] VREF PIX_IN[6910] NB2 NB1 CSA_VREF pixel
xPix6911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[69] VREF PIX_IN[6911] NB2 NB1 CSA_VREF pixel
xPix6912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[69] VREF PIX_IN[6912] NB2 NB1 CSA_VREF pixel
xPix6913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[69] VREF PIX_IN[6913] NB2 NB1 CSA_VREF pixel
xPix6914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[69] VREF PIX_IN[6914] NB2 NB1 CSA_VREF pixel
xPix6915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[69] VREF PIX_IN[6915] NB2 NB1 CSA_VREF pixel
xPix6916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[69] VREF PIX_IN[6916] NB2 NB1 CSA_VREF pixel
xPix6917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[69] VREF PIX_IN[6917] NB2 NB1 CSA_VREF pixel
xPix6918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[69] VREF PIX_IN[6918] NB2 NB1 CSA_VREF pixel
xPix6919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[69] VREF PIX_IN[6919] NB2 NB1 CSA_VREF pixel
xPix6920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[69] VREF PIX_IN[6920] NB2 NB1 CSA_VREF pixel
xPix6921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[69] VREF PIX_IN[6921] NB2 NB1 CSA_VREF pixel
xPix6922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[69] VREF PIX_IN[6922] NB2 NB1 CSA_VREF pixel
xPix6923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[69] VREF PIX_IN[6923] NB2 NB1 CSA_VREF pixel
xPix6924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[69] VREF PIX_IN[6924] NB2 NB1 CSA_VREF pixel
xPix6925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[69] VREF PIX_IN[6925] NB2 NB1 CSA_VREF pixel
xPix6926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[69] VREF PIX_IN[6926] NB2 NB1 CSA_VREF pixel
xPix6927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[69] VREF PIX_IN[6927] NB2 NB1 CSA_VREF pixel
xPix6928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[69] VREF PIX_IN[6928] NB2 NB1 CSA_VREF pixel
xPix6929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[69] VREF PIX_IN[6929] NB2 NB1 CSA_VREF pixel
xPix6930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[69] VREF PIX_IN[6930] NB2 NB1 CSA_VREF pixel
xPix6931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[69] VREF PIX_IN[6931] NB2 NB1 CSA_VREF pixel
xPix6932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[69] VREF PIX_IN[6932] NB2 NB1 CSA_VREF pixel
xPix6933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[69] VREF PIX_IN[6933] NB2 NB1 CSA_VREF pixel
xPix6934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[69] VREF PIX_IN[6934] NB2 NB1 CSA_VREF pixel
xPix6935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[69] VREF PIX_IN[6935] NB2 NB1 CSA_VREF pixel
xPix6936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[69] VREF PIX_IN[6936] NB2 NB1 CSA_VREF pixel
xPix6937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[69] VREF PIX_IN[6937] NB2 NB1 CSA_VREF pixel
xPix6938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[69] VREF PIX_IN[6938] NB2 NB1 CSA_VREF pixel
xPix6939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[69] VREF PIX_IN[6939] NB2 NB1 CSA_VREF pixel
xPix6940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[69] VREF PIX_IN[6940] NB2 NB1 CSA_VREF pixel
xPix6941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[69] VREF PIX_IN[6941] NB2 NB1 CSA_VREF pixel
xPix6942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[69] VREF PIX_IN[6942] NB2 NB1 CSA_VREF pixel
xPix6943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[69] VREF PIX_IN[6943] NB2 NB1 CSA_VREF pixel
xPix6944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[69] VREF PIX_IN[6944] NB2 NB1 CSA_VREF pixel
xPix6945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[69] VREF PIX_IN[6945] NB2 NB1 CSA_VREF pixel
xPix6946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[69] VREF PIX_IN[6946] NB2 NB1 CSA_VREF pixel
xPix6947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[69] VREF PIX_IN[6947] NB2 NB1 CSA_VREF pixel
xPix6948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[69] VREF PIX_IN[6948] NB2 NB1 CSA_VREF pixel
xPix6949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[69] VREF PIX_IN[6949] NB2 NB1 CSA_VREF pixel
xPix6950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[69] VREF PIX_IN[6950] NB2 NB1 CSA_VREF pixel
xPix6951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[69] VREF PIX_IN[6951] NB2 NB1 CSA_VREF pixel
xPix6952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[69] VREF PIX_IN[6952] NB2 NB1 CSA_VREF pixel
xPix6953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[69] VREF PIX_IN[6953] NB2 NB1 CSA_VREF pixel
xPix6954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[69] VREF PIX_IN[6954] NB2 NB1 CSA_VREF pixel
xPix6955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[69] VREF PIX_IN[6955] NB2 NB1 CSA_VREF pixel
xPix6956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[69] VREF PIX_IN[6956] NB2 NB1 CSA_VREF pixel
xPix6957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[69] VREF PIX_IN[6957] NB2 NB1 CSA_VREF pixel
xPix6958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[69] VREF PIX_IN[6958] NB2 NB1 CSA_VREF pixel
xPix6959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[69] VREF PIX_IN[6959] NB2 NB1 CSA_VREF pixel
xPix6960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[69] VREF PIX_IN[6960] NB2 NB1 CSA_VREF pixel
xPix6961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[69] VREF PIX_IN[6961] NB2 NB1 CSA_VREF pixel
xPix6962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[69] VREF PIX_IN[6962] NB2 NB1 CSA_VREF pixel
xPix6963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[69] VREF PIX_IN[6963] NB2 NB1 CSA_VREF pixel
xPix6964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[69] VREF PIX_IN[6964] NB2 NB1 CSA_VREF pixel
xPix6965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[69] VREF PIX_IN[6965] NB2 NB1 CSA_VREF pixel
xPix6966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[69] VREF PIX_IN[6966] NB2 NB1 CSA_VREF pixel
xPix6967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[69] VREF PIX_IN[6967] NB2 NB1 CSA_VREF pixel
xPix6968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[69] VREF PIX_IN[6968] NB2 NB1 CSA_VREF pixel
xPix6969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[69] VREF PIX_IN[6969] NB2 NB1 CSA_VREF pixel
xPix6970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[69] VREF PIX_IN[6970] NB2 NB1 CSA_VREF pixel
xPix6971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[69] VREF PIX_IN[6971] NB2 NB1 CSA_VREF pixel
xPix6972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[69] VREF PIX_IN[6972] NB2 NB1 CSA_VREF pixel
xPix6973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[69] VREF PIX_IN[6973] NB2 NB1 CSA_VREF pixel
xPix6974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[69] VREF PIX_IN[6974] NB2 NB1 CSA_VREF pixel
xPix6975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[69] VREF PIX_IN[6975] NB2 NB1 CSA_VREF pixel
xPix6976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[69] VREF PIX_IN[6976] NB2 NB1 CSA_VREF pixel
xPix6977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[69] VREF PIX_IN[6977] NB2 NB1 CSA_VREF pixel
xPix6978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[69] VREF PIX_IN[6978] NB2 NB1 CSA_VREF pixel
xPix6979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[69] VREF PIX_IN[6979] NB2 NB1 CSA_VREF pixel
xPix6980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[69] VREF PIX_IN[6980] NB2 NB1 CSA_VREF pixel
xPix6981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[69] VREF PIX_IN[6981] NB2 NB1 CSA_VREF pixel
xPix6982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[69] VREF PIX_IN[6982] NB2 NB1 CSA_VREF pixel
xPix6983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[69] VREF PIX_IN[6983] NB2 NB1 CSA_VREF pixel
xPix6984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[69] VREF PIX_IN[6984] NB2 NB1 CSA_VREF pixel
xPix6985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[69] VREF PIX_IN[6985] NB2 NB1 CSA_VREF pixel
xPix6986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[69] VREF PIX_IN[6986] NB2 NB1 CSA_VREF pixel
xPix6987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[69] VREF PIX_IN[6987] NB2 NB1 CSA_VREF pixel
xPix6988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[69] VREF PIX_IN[6988] NB2 NB1 CSA_VREF pixel
xPix6989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[69] VREF PIX_IN[6989] NB2 NB1 CSA_VREF pixel
xPix6990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[69] VREF PIX_IN[6990] NB2 NB1 CSA_VREF pixel
xPix6991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[69] VREF PIX_IN[6991] NB2 NB1 CSA_VREF pixel
xPix6992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[69] VREF PIX_IN[6992] NB2 NB1 CSA_VREF pixel
xPix6993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[69] VREF PIX_IN[6993] NB2 NB1 CSA_VREF pixel
xPix6994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[69] VREF PIX_IN[6994] NB2 NB1 CSA_VREF pixel
xPix6995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[69] VREF PIX_IN[6995] NB2 NB1 CSA_VREF pixel
xPix6996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[69] VREF PIX_IN[6996] NB2 NB1 CSA_VREF pixel
xPix6997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[69] VREF PIX_IN[6997] NB2 NB1 CSA_VREF pixel
xPix6998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[69] VREF PIX_IN[6998] NB2 NB1 CSA_VREF pixel
xPix6999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[69] VREF PIX_IN[6999] NB2 NB1 CSA_VREF pixel
xPix7000 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[70] VREF PIX_IN[7000] NB2 NB1 CSA_VREF pixel
xPix7001 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[70] VREF PIX_IN[7001] NB2 NB1 CSA_VREF pixel
xPix7002 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[70] VREF PIX_IN[7002] NB2 NB1 CSA_VREF pixel
xPix7003 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[70] VREF PIX_IN[7003] NB2 NB1 CSA_VREF pixel
xPix7004 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[70] VREF PIX_IN[7004] NB2 NB1 CSA_VREF pixel
xPix7005 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[70] VREF PIX_IN[7005] NB2 NB1 CSA_VREF pixel
xPix7006 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[70] VREF PIX_IN[7006] NB2 NB1 CSA_VREF pixel
xPix7007 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[70] VREF PIX_IN[7007] NB2 NB1 CSA_VREF pixel
xPix7008 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[70] VREF PIX_IN[7008] NB2 NB1 CSA_VREF pixel
xPix7009 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[70] VREF PIX_IN[7009] NB2 NB1 CSA_VREF pixel
xPix7010 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[70] VREF PIX_IN[7010] NB2 NB1 CSA_VREF pixel
xPix7011 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[70] VREF PIX_IN[7011] NB2 NB1 CSA_VREF pixel
xPix7012 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[70] VREF PIX_IN[7012] NB2 NB1 CSA_VREF pixel
xPix7013 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[70] VREF PIX_IN[7013] NB2 NB1 CSA_VREF pixel
xPix7014 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[70] VREF PIX_IN[7014] NB2 NB1 CSA_VREF pixel
xPix7015 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[70] VREF PIX_IN[7015] NB2 NB1 CSA_VREF pixel
xPix7016 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[70] VREF PIX_IN[7016] NB2 NB1 CSA_VREF pixel
xPix7017 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[70] VREF PIX_IN[7017] NB2 NB1 CSA_VREF pixel
xPix7018 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[70] VREF PIX_IN[7018] NB2 NB1 CSA_VREF pixel
xPix7019 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[70] VREF PIX_IN[7019] NB2 NB1 CSA_VREF pixel
xPix7020 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[70] VREF PIX_IN[7020] NB2 NB1 CSA_VREF pixel
xPix7021 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[70] VREF PIX_IN[7021] NB2 NB1 CSA_VREF pixel
xPix7022 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[70] VREF PIX_IN[7022] NB2 NB1 CSA_VREF pixel
xPix7023 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[70] VREF PIX_IN[7023] NB2 NB1 CSA_VREF pixel
xPix7024 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[70] VREF PIX_IN[7024] NB2 NB1 CSA_VREF pixel
xPix7025 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[70] VREF PIX_IN[7025] NB2 NB1 CSA_VREF pixel
xPix7026 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[70] VREF PIX_IN[7026] NB2 NB1 CSA_VREF pixel
xPix7027 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[70] VREF PIX_IN[7027] NB2 NB1 CSA_VREF pixel
xPix7028 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[70] VREF PIX_IN[7028] NB2 NB1 CSA_VREF pixel
xPix7029 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[70] VREF PIX_IN[7029] NB2 NB1 CSA_VREF pixel
xPix7030 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[70] VREF PIX_IN[7030] NB2 NB1 CSA_VREF pixel
xPix7031 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[70] VREF PIX_IN[7031] NB2 NB1 CSA_VREF pixel
xPix7032 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[70] VREF PIX_IN[7032] NB2 NB1 CSA_VREF pixel
xPix7033 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[70] VREF PIX_IN[7033] NB2 NB1 CSA_VREF pixel
xPix7034 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[70] VREF PIX_IN[7034] NB2 NB1 CSA_VREF pixel
xPix7035 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[70] VREF PIX_IN[7035] NB2 NB1 CSA_VREF pixel
xPix7036 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[70] VREF PIX_IN[7036] NB2 NB1 CSA_VREF pixel
xPix7037 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[70] VREF PIX_IN[7037] NB2 NB1 CSA_VREF pixel
xPix7038 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[70] VREF PIX_IN[7038] NB2 NB1 CSA_VREF pixel
xPix7039 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[70] VREF PIX_IN[7039] NB2 NB1 CSA_VREF pixel
xPix7040 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[70] VREF PIX_IN[7040] NB2 NB1 CSA_VREF pixel
xPix7041 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[70] VREF PIX_IN[7041] NB2 NB1 CSA_VREF pixel
xPix7042 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[70] VREF PIX_IN[7042] NB2 NB1 CSA_VREF pixel
xPix7043 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[70] VREF PIX_IN[7043] NB2 NB1 CSA_VREF pixel
xPix7044 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[70] VREF PIX_IN[7044] NB2 NB1 CSA_VREF pixel
xPix7045 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[70] VREF PIX_IN[7045] NB2 NB1 CSA_VREF pixel
xPix7046 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[70] VREF PIX_IN[7046] NB2 NB1 CSA_VREF pixel
xPix7047 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[70] VREF PIX_IN[7047] NB2 NB1 CSA_VREF pixel
xPix7048 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[70] VREF PIX_IN[7048] NB2 NB1 CSA_VREF pixel
xPix7049 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[70] VREF PIX_IN[7049] NB2 NB1 CSA_VREF pixel
xPix7050 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[70] VREF PIX_IN[7050] NB2 NB1 CSA_VREF pixel
xPix7051 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[70] VREF PIX_IN[7051] NB2 NB1 CSA_VREF pixel
xPix7052 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[70] VREF PIX_IN[7052] NB2 NB1 CSA_VREF pixel
xPix7053 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[70] VREF PIX_IN[7053] NB2 NB1 CSA_VREF pixel
xPix7054 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[70] VREF PIX_IN[7054] NB2 NB1 CSA_VREF pixel
xPix7055 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[70] VREF PIX_IN[7055] NB2 NB1 CSA_VREF pixel
xPix7056 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[70] VREF PIX_IN[7056] NB2 NB1 CSA_VREF pixel
xPix7057 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[70] VREF PIX_IN[7057] NB2 NB1 CSA_VREF pixel
xPix7058 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[70] VREF PIX_IN[7058] NB2 NB1 CSA_VREF pixel
xPix7059 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[70] VREF PIX_IN[7059] NB2 NB1 CSA_VREF pixel
xPix7060 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[70] VREF PIX_IN[7060] NB2 NB1 CSA_VREF pixel
xPix7061 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[70] VREF PIX_IN[7061] NB2 NB1 CSA_VREF pixel
xPix7062 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[70] VREF PIX_IN[7062] NB2 NB1 CSA_VREF pixel
xPix7063 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[70] VREF PIX_IN[7063] NB2 NB1 CSA_VREF pixel
xPix7064 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[70] VREF PIX_IN[7064] NB2 NB1 CSA_VREF pixel
xPix7065 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[70] VREF PIX_IN[7065] NB2 NB1 CSA_VREF pixel
xPix7066 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[70] VREF PIX_IN[7066] NB2 NB1 CSA_VREF pixel
xPix7067 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[70] VREF PIX_IN[7067] NB2 NB1 CSA_VREF pixel
xPix7068 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[70] VREF PIX_IN[7068] NB2 NB1 CSA_VREF pixel
xPix7069 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[70] VREF PIX_IN[7069] NB2 NB1 CSA_VREF pixel
xPix7070 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[70] VREF PIX_IN[7070] NB2 NB1 CSA_VREF pixel
xPix7071 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[70] VREF PIX_IN[7071] NB2 NB1 CSA_VREF pixel
xPix7072 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[70] VREF PIX_IN[7072] NB2 NB1 CSA_VREF pixel
xPix7073 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[70] VREF PIX_IN[7073] NB2 NB1 CSA_VREF pixel
xPix7074 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[70] VREF PIX_IN[7074] NB2 NB1 CSA_VREF pixel
xPix7075 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[70] VREF PIX_IN[7075] NB2 NB1 CSA_VREF pixel
xPix7076 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[70] VREF PIX_IN[7076] NB2 NB1 CSA_VREF pixel
xPix7077 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[70] VREF PIX_IN[7077] NB2 NB1 CSA_VREF pixel
xPix7078 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[70] VREF PIX_IN[7078] NB2 NB1 CSA_VREF pixel
xPix7079 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[70] VREF PIX_IN[7079] NB2 NB1 CSA_VREF pixel
xPix7080 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[70] VREF PIX_IN[7080] NB2 NB1 CSA_VREF pixel
xPix7081 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[70] VREF PIX_IN[7081] NB2 NB1 CSA_VREF pixel
xPix7082 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[70] VREF PIX_IN[7082] NB2 NB1 CSA_VREF pixel
xPix7083 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[70] VREF PIX_IN[7083] NB2 NB1 CSA_VREF pixel
xPix7084 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[70] VREF PIX_IN[7084] NB2 NB1 CSA_VREF pixel
xPix7085 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[70] VREF PIX_IN[7085] NB2 NB1 CSA_VREF pixel
xPix7086 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[70] VREF PIX_IN[7086] NB2 NB1 CSA_VREF pixel
xPix7087 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[70] VREF PIX_IN[7087] NB2 NB1 CSA_VREF pixel
xPix7088 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[70] VREF PIX_IN[7088] NB2 NB1 CSA_VREF pixel
xPix7089 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[70] VREF PIX_IN[7089] NB2 NB1 CSA_VREF pixel
xPix7090 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[70] VREF PIX_IN[7090] NB2 NB1 CSA_VREF pixel
xPix7091 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[70] VREF PIX_IN[7091] NB2 NB1 CSA_VREF pixel
xPix7092 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[70] VREF PIX_IN[7092] NB2 NB1 CSA_VREF pixel
xPix7093 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[70] VREF PIX_IN[7093] NB2 NB1 CSA_VREF pixel
xPix7094 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[70] VREF PIX_IN[7094] NB2 NB1 CSA_VREF pixel
xPix7095 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[70] VREF PIX_IN[7095] NB2 NB1 CSA_VREF pixel
xPix7096 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[70] VREF PIX_IN[7096] NB2 NB1 CSA_VREF pixel
xPix7097 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[70] VREF PIX_IN[7097] NB2 NB1 CSA_VREF pixel
xPix7098 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[70] VREF PIX_IN[7098] NB2 NB1 CSA_VREF pixel
xPix7099 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[70] VREF PIX_IN[7099] NB2 NB1 CSA_VREF pixel
xPix7100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[71] VREF PIX_IN[7100] NB2 NB1 CSA_VREF pixel
xPix7101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[71] VREF PIX_IN[7101] NB2 NB1 CSA_VREF pixel
xPix7102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[71] VREF PIX_IN[7102] NB2 NB1 CSA_VREF pixel
xPix7103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[71] VREF PIX_IN[7103] NB2 NB1 CSA_VREF pixel
xPix7104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[71] VREF PIX_IN[7104] NB2 NB1 CSA_VREF pixel
xPix7105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[71] VREF PIX_IN[7105] NB2 NB1 CSA_VREF pixel
xPix7106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[71] VREF PIX_IN[7106] NB2 NB1 CSA_VREF pixel
xPix7107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[71] VREF PIX_IN[7107] NB2 NB1 CSA_VREF pixel
xPix7108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[71] VREF PIX_IN[7108] NB2 NB1 CSA_VREF pixel
xPix7109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[71] VREF PIX_IN[7109] NB2 NB1 CSA_VREF pixel
xPix7110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[71] VREF PIX_IN[7110] NB2 NB1 CSA_VREF pixel
xPix7111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[71] VREF PIX_IN[7111] NB2 NB1 CSA_VREF pixel
xPix7112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[71] VREF PIX_IN[7112] NB2 NB1 CSA_VREF pixel
xPix7113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[71] VREF PIX_IN[7113] NB2 NB1 CSA_VREF pixel
xPix7114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[71] VREF PIX_IN[7114] NB2 NB1 CSA_VREF pixel
xPix7115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[71] VREF PIX_IN[7115] NB2 NB1 CSA_VREF pixel
xPix7116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[71] VREF PIX_IN[7116] NB2 NB1 CSA_VREF pixel
xPix7117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[71] VREF PIX_IN[7117] NB2 NB1 CSA_VREF pixel
xPix7118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[71] VREF PIX_IN[7118] NB2 NB1 CSA_VREF pixel
xPix7119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[71] VREF PIX_IN[7119] NB2 NB1 CSA_VREF pixel
xPix7120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[71] VREF PIX_IN[7120] NB2 NB1 CSA_VREF pixel
xPix7121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[71] VREF PIX_IN[7121] NB2 NB1 CSA_VREF pixel
xPix7122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[71] VREF PIX_IN[7122] NB2 NB1 CSA_VREF pixel
xPix7123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[71] VREF PIX_IN[7123] NB2 NB1 CSA_VREF pixel
xPix7124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[71] VREF PIX_IN[7124] NB2 NB1 CSA_VREF pixel
xPix7125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[71] VREF PIX_IN[7125] NB2 NB1 CSA_VREF pixel
xPix7126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[71] VREF PIX_IN[7126] NB2 NB1 CSA_VREF pixel
xPix7127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[71] VREF PIX_IN[7127] NB2 NB1 CSA_VREF pixel
xPix7128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[71] VREF PIX_IN[7128] NB2 NB1 CSA_VREF pixel
xPix7129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[71] VREF PIX_IN[7129] NB2 NB1 CSA_VREF pixel
xPix7130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[71] VREF PIX_IN[7130] NB2 NB1 CSA_VREF pixel
xPix7131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[71] VREF PIX_IN[7131] NB2 NB1 CSA_VREF pixel
xPix7132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[71] VREF PIX_IN[7132] NB2 NB1 CSA_VREF pixel
xPix7133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[71] VREF PIX_IN[7133] NB2 NB1 CSA_VREF pixel
xPix7134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[71] VREF PIX_IN[7134] NB2 NB1 CSA_VREF pixel
xPix7135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[71] VREF PIX_IN[7135] NB2 NB1 CSA_VREF pixel
xPix7136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[71] VREF PIX_IN[7136] NB2 NB1 CSA_VREF pixel
xPix7137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[71] VREF PIX_IN[7137] NB2 NB1 CSA_VREF pixel
xPix7138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[71] VREF PIX_IN[7138] NB2 NB1 CSA_VREF pixel
xPix7139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[71] VREF PIX_IN[7139] NB2 NB1 CSA_VREF pixel
xPix7140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[71] VREF PIX_IN[7140] NB2 NB1 CSA_VREF pixel
xPix7141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[71] VREF PIX_IN[7141] NB2 NB1 CSA_VREF pixel
xPix7142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[71] VREF PIX_IN[7142] NB2 NB1 CSA_VREF pixel
xPix7143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[71] VREF PIX_IN[7143] NB2 NB1 CSA_VREF pixel
xPix7144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[71] VREF PIX_IN[7144] NB2 NB1 CSA_VREF pixel
xPix7145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[71] VREF PIX_IN[7145] NB2 NB1 CSA_VREF pixel
xPix7146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[71] VREF PIX_IN[7146] NB2 NB1 CSA_VREF pixel
xPix7147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[71] VREF PIX_IN[7147] NB2 NB1 CSA_VREF pixel
xPix7148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[71] VREF PIX_IN[7148] NB2 NB1 CSA_VREF pixel
xPix7149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[71] VREF PIX_IN[7149] NB2 NB1 CSA_VREF pixel
xPix7150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[71] VREF PIX_IN[7150] NB2 NB1 CSA_VREF pixel
xPix7151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[71] VREF PIX_IN[7151] NB2 NB1 CSA_VREF pixel
xPix7152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[71] VREF PIX_IN[7152] NB2 NB1 CSA_VREF pixel
xPix7153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[71] VREF PIX_IN[7153] NB2 NB1 CSA_VREF pixel
xPix7154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[71] VREF PIX_IN[7154] NB2 NB1 CSA_VREF pixel
xPix7155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[71] VREF PIX_IN[7155] NB2 NB1 CSA_VREF pixel
xPix7156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[71] VREF PIX_IN[7156] NB2 NB1 CSA_VREF pixel
xPix7157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[71] VREF PIX_IN[7157] NB2 NB1 CSA_VREF pixel
xPix7158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[71] VREF PIX_IN[7158] NB2 NB1 CSA_VREF pixel
xPix7159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[71] VREF PIX_IN[7159] NB2 NB1 CSA_VREF pixel
xPix7160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[71] VREF PIX_IN[7160] NB2 NB1 CSA_VREF pixel
xPix7161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[71] VREF PIX_IN[7161] NB2 NB1 CSA_VREF pixel
xPix7162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[71] VREF PIX_IN[7162] NB2 NB1 CSA_VREF pixel
xPix7163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[71] VREF PIX_IN[7163] NB2 NB1 CSA_VREF pixel
xPix7164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[71] VREF PIX_IN[7164] NB2 NB1 CSA_VREF pixel
xPix7165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[71] VREF PIX_IN[7165] NB2 NB1 CSA_VREF pixel
xPix7166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[71] VREF PIX_IN[7166] NB2 NB1 CSA_VREF pixel
xPix7167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[71] VREF PIX_IN[7167] NB2 NB1 CSA_VREF pixel
xPix7168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[71] VREF PIX_IN[7168] NB2 NB1 CSA_VREF pixel
xPix7169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[71] VREF PIX_IN[7169] NB2 NB1 CSA_VREF pixel
xPix7170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[71] VREF PIX_IN[7170] NB2 NB1 CSA_VREF pixel
xPix7171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[71] VREF PIX_IN[7171] NB2 NB1 CSA_VREF pixel
xPix7172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[71] VREF PIX_IN[7172] NB2 NB1 CSA_VREF pixel
xPix7173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[71] VREF PIX_IN[7173] NB2 NB1 CSA_VREF pixel
xPix7174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[71] VREF PIX_IN[7174] NB2 NB1 CSA_VREF pixel
xPix7175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[71] VREF PIX_IN[7175] NB2 NB1 CSA_VREF pixel
xPix7176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[71] VREF PIX_IN[7176] NB2 NB1 CSA_VREF pixel
xPix7177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[71] VREF PIX_IN[7177] NB2 NB1 CSA_VREF pixel
xPix7178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[71] VREF PIX_IN[7178] NB2 NB1 CSA_VREF pixel
xPix7179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[71] VREF PIX_IN[7179] NB2 NB1 CSA_VREF pixel
xPix7180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[71] VREF PIX_IN[7180] NB2 NB1 CSA_VREF pixel
xPix7181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[71] VREF PIX_IN[7181] NB2 NB1 CSA_VREF pixel
xPix7182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[71] VREF PIX_IN[7182] NB2 NB1 CSA_VREF pixel
xPix7183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[71] VREF PIX_IN[7183] NB2 NB1 CSA_VREF pixel
xPix7184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[71] VREF PIX_IN[7184] NB2 NB1 CSA_VREF pixel
xPix7185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[71] VREF PIX_IN[7185] NB2 NB1 CSA_VREF pixel
xPix7186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[71] VREF PIX_IN[7186] NB2 NB1 CSA_VREF pixel
xPix7187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[71] VREF PIX_IN[7187] NB2 NB1 CSA_VREF pixel
xPix7188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[71] VREF PIX_IN[7188] NB2 NB1 CSA_VREF pixel
xPix7189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[71] VREF PIX_IN[7189] NB2 NB1 CSA_VREF pixel
xPix7190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[71] VREF PIX_IN[7190] NB2 NB1 CSA_VREF pixel
xPix7191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[71] VREF PIX_IN[7191] NB2 NB1 CSA_VREF pixel
xPix7192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[71] VREF PIX_IN[7192] NB2 NB1 CSA_VREF pixel
xPix7193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[71] VREF PIX_IN[7193] NB2 NB1 CSA_VREF pixel
xPix7194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[71] VREF PIX_IN[7194] NB2 NB1 CSA_VREF pixel
xPix7195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[71] VREF PIX_IN[7195] NB2 NB1 CSA_VREF pixel
xPix7196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[71] VREF PIX_IN[7196] NB2 NB1 CSA_VREF pixel
xPix7197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[71] VREF PIX_IN[7197] NB2 NB1 CSA_VREF pixel
xPix7198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[71] VREF PIX_IN[7198] NB2 NB1 CSA_VREF pixel
xPix7199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[71] VREF PIX_IN[7199] NB2 NB1 CSA_VREF pixel
xPix7200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[72] VREF PIX_IN[7200] NB2 NB1 CSA_VREF pixel
xPix7201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[72] VREF PIX_IN[7201] NB2 NB1 CSA_VREF pixel
xPix7202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[72] VREF PIX_IN[7202] NB2 NB1 CSA_VREF pixel
xPix7203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[72] VREF PIX_IN[7203] NB2 NB1 CSA_VREF pixel
xPix7204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[72] VREF PIX_IN[7204] NB2 NB1 CSA_VREF pixel
xPix7205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[72] VREF PIX_IN[7205] NB2 NB1 CSA_VREF pixel
xPix7206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[72] VREF PIX_IN[7206] NB2 NB1 CSA_VREF pixel
xPix7207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[72] VREF PIX_IN[7207] NB2 NB1 CSA_VREF pixel
xPix7208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[72] VREF PIX_IN[7208] NB2 NB1 CSA_VREF pixel
xPix7209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[72] VREF PIX_IN[7209] NB2 NB1 CSA_VREF pixel
xPix7210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[72] VREF PIX_IN[7210] NB2 NB1 CSA_VREF pixel
xPix7211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[72] VREF PIX_IN[7211] NB2 NB1 CSA_VREF pixel
xPix7212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[72] VREF PIX_IN[7212] NB2 NB1 CSA_VREF pixel
xPix7213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[72] VREF PIX_IN[7213] NB2 NB1 CSA_VREF pixel
xPix7214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[72] VREF PIX_IN[7214] NB2 NB1 CSA_VREF pixel
xPix7215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[72] VREF PIX_IN[7215] NB2 NB1 CSA_VREF pixel
xPix7216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[72] VREF PIX_IN[7216] NB2 NB1 CSA_VREF pixel
xPix7217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[72] VREF PIX_IN[7217] NB2 NB1 CSA_VREF pixel
xPix7218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[72] VREF PIX_IN[7218] NB2 NB1 CSA_VREF pixel
xPix7219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[72] VREF PIX_IN[7219] NB2 NB1 CSA_VREF pixel
xPix7220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[72] VREF PIX_IN[7220] NB2 NB1 CSA_VREF pixel
xPix7221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[72] VREF PIX_IN[7221] NB2 NB1 CSA_VREF pixel
xPix7222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[72] VREF PIX_IN[7222] NB2 NB1 CSA_VREF pixel
xPix7223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[72] VREF PIX_IN[7223] NB2 NB1 CSA_VREF pixel
xPix7224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[72] VREF PIX_IN[7224] NB2 NB1 CSA_VREF pixel
xPix7225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[72] VREF PIX_IN[7225] NB2 NB1 CSA_VREF pixel
xPix7226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[72] VREF PIX_IN[7226] NB2 NB1 CSA_VREF pixel
xPix7227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[72] VREF PIX_IN[7227] NB2 NB1 CSA_VREF pixel
xPix7228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[72] VREF PIX_IN[7228] NB2 NB1 CSA_VREF pixel
xPix7229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[72] VREF PIX_IN[7229] NB2 NB1 CSA_VREF pixel
xPix7230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[72] VREF PIX_IN[7230] NB2 NB1 CSA_VREF pixel
xPix7231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[72] VREF PIX_IN[7231] NB2 NB1 CSA_VREF pixel
xPix7232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[72] VREF PIX_IN[7232] NB2 NB1 CSA_VREF pixel
xPix7233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[72] VREF PIX_IN[7233] NB2 NB1 CSA_VREF pixel
xPix7234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[72] VREF PIX_IN[7234] NB2 NB1 CSA_VREF pixel
xPix7235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[72] VREF PIX_IN[7235] NB2 NB1 CSA_VREF pixel
xPix7236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[72] VREF PIX_IN[7236] NB2 NB1 CSA_VREF pixel
xPix7237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[72] VREF PIX_IN[7237] NB2 NB1 CSA_VREF pixel
xPix7238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[72] VREF PIX_IN[7238] NB2 NB1 CSA_VREF pixel
xPix7239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[72] VREF PIX_IN[7239] NB2 NB1 CSA_VREF pixel
xPix7240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[72] VREF PIX_IN[7240] NB2 NB1 CSA_VREF pixel
xPix7241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[72] VREF PIX_IN[7241] NB2 NB1 CSA_VREF pixel
xPix7242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[72] VREF PIX_IN[7242] NB2 NB1 CSA_VREF pixel
xPix7243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[72] VREF PIX_IN[7243] NB2 NB1 CSA_VREF pixel
xPix7244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[72] VREF PIX_IN[7244] NB2 NB1 CSA_VREF pixel
xPix7245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[72] VREF PIX_IN[7245] NB2 NB1 CSA_VREF pixel
xPix7246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[72] VREF PIX_IN[7246] NB2 NB1 CSA_VREF pixel
xPix7247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[72] VREF PIX_IN[7247] NB2 NB1 CSA_VREF pixel
xPix7248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[72] VREF PIX_IN[7248] NB2 NB1 CSA_VREF pixel
xPix7249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[72] VREF PIX_IN[7249] NB2 NB1 CSA_VREF pixel
xPix7250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[72] VREF PIX_IN[7250] NB2 NB1 CSA_VREF pixel
xPix7251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[72] VREF PIX_IN[7251] NB2 NB1 CSA_VREF pixel
xPix7252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[72] VREF PIX_IN[7252] NB2 NB1 CSA_VREF pixel
xPix7253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[72] VREF PIX_IN[7253] NB2 NB1 CSA_VREF pixel
xPix7254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[72] VREF PIX_IN[7254] NB2 NB1 CSA_VREF pixel
xPix7255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[72] VREF PIX_IN[7255] NB2 NB1 CSA_VREF pixel
xPix7256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[72] VREF PIX_IN[7256] NB2 NB1 CSA_VREF pixel
xPix7257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[72] VREF PIX_IN[7257] NB2 NB1 CSA_VREF pixel
xPix7258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[72] VREF PIX_IN[7258] NB2 NB1 CSA_VREF pixel
xPix7259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[72] VREF PIX_IN[7259] NB2 NB1 CSA_VREF pixel
xPix7260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[72] VREF PIX_IN[7260] NB2 NB1 CSA_VREF pixel
xPix7261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[72] VREF PIX_IN[7261] NB2 NB1 CSA_VREF pixel
xPix7262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[72] VREF PIX_IN[7262] NB2 NB1 CSA_VREF pixel
xPix7263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[72] VREF PIX_IN[7263] NB2 NB1 CSA_VREF pixel
xPix7264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[72] VREF PIX_IN[7264] NB2 NB1 CSA_VREF pixel
xPix7265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[72] VREF PIX_IN[7265] NB2 NB1 CSA_VREF pixel
xPix7266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[72] VREF PIX_IN[7266] NB2 NB1 CSA_VREF pixel
xPix7267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[72] VREF PIX_IN[7267] NB2 NB1 CSA_VREF pixel
xPix7268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[72] VREF PIX_IN[7268] NB2 NB1 CSA_VREF pixel
xPix7269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[72] VREF PIX_IN[7269] NB2 NB1 CSA_VREF pixel
xPix7270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[72] VREF PIX_IN[7270] NB2 NB1 CSA_VREF pixel
xPix7271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[72] VREF PIX_IN[7271] NB2 NB1 CSA_VREF pixel
xPix7272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[72] VREF PIX_IN[7272] NB2 NB1 CSA_VREF pixel
xPix7273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[72] VREF PIX_IN[7273] NB2 NB1 CSA_VREF pixel
xPix7274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[72] VREF PIX_IN[7274] NB2 NB1 CSA_VREF pixel
xPix7275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[72] VREF PIX_IN[7275] NB2 NB1 CSA_VREF pixel
xPix7276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[72] VREF PIX_IN[7276] NB2 NB1 CSA_VREF pixel
xPix7277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[72] VREF PIX_IN[7277] NB2 NB1 CSA_VREF pixel
xPix7278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[72] VREF PIX_IN[7278] NB2 NB1 CSA_VREF pixel
xPix7279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[72] VREF PIX_IN[7279] NB2 NB1 CSA_VREF pixel
xPix7280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[72] VREF PIX_IN[7280] NB2 NB1 CSA_VREF pixel
xPix7281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[72] VREF PIX_IN[7281] NB2 NB1 CSA_VREF pixel
xPix7282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[72] VREF PIX_IN[7282] NB2 NB1 CSA_VREF pixel
xPix7283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[72] VREF PIX_IN[7283] NB2 NB1 CSA_VREF pixel
xPix7284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[72] VREF PIX_IN[7284] NB2 NB1 CSA_VREF pixel
xPix7285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[72] VREF PIX_IN[7285] NB2 NB1 CSA_VREF pixel
xPix7286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[72] VREF PIX_IN[7286] NB2 NB1 CSA_VREF pixel
xPix7287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[72] VREF PIX_IN[7287] NB2 NB1 CSA_VREF pixel
xPix7288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[72] VREF PIX_IN[7288] NB2 NB1 CSA_VREF pixel
xPix7289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[72] VREF PIX_IN[7289] NB2 NB1 CSA_VREF pixel
xPix7290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[72] VREF PIX_IN[7290] NB2 NB1 CSA_VREF pixel
xPix7291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[72] VREF PIX_IN[7291] NB2 NB1 CSA_VREF pixel
xPix7292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[72] VREF PIX_IN[7292] NB2 NB1 CSA_VREF pixel
xPix7293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[72] VREF PIX_IN[7293] NB2 NB1 CSA_VREF pixel
xPix7294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[72] VREF PIX_IN[7294] NB2 NB1 CSA_VREF pixel
xPix7295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[72] VREF PIX_IN[7295] NB2 NB1 CSA_VREF pixel
xPix7296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[72] VREF PIX_IN[7296] NB2 NB1 CSA_VREF pixel
xPix7297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[72] VREF PIX_IN[7297] NB2 NB1 CSA_VREF pixel
xPix7298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[72] VREF PIX_IN[7298] NB2 NB1 CSA_VREF pixel
xPix7299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[72] VREF PIX_IN[7299] NB2 NB1 CSA_VREF pixel
xPix7300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[73] VREF PIX_IN[7300] NB2 NB1 CSA_VREF pixel
xPix7301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[73] VREF PIX_IN[7301] NB2 NB1 CSA_VREF pixel
xPix7302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[73] VREF PIX_IN[7302] NB2 NB1 CSA_VREF pixel
xPix7303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[73] VREF PIX_IN[7303] NB2 NB1 CSA_VREF pixel
xPix7304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[73] VREF PIX_IN[7304] NB2 NB1 CSA_VREF pixel
xPix7305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[73] VREF PIX_IN[7305] NB2 NB1 CSA_VREF pixel
xPix7306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[73] VREF PIX_IN[7306] NB2 NB1 CSA_VREF pixel
xPix7307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[73] VREF PIX_IN[7307] NB2 NB1 CSA_VREF pixel
xPix7308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[73] VREF PIX_IN[7308] NB2 NB1 CSA_VREF pixel
xPix7309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[73] VREF PIX_IN[7309] NB2 NB1 CSA_VREF pixel
xPix7310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[73] VREF PIX_IN[7310] NB2 NB1 CSA_VREF pixel
xPix7311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[73] VREF PIX_IN[7311] NB2 NB1 CSA_VREF pixel
xPix7312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[73] VREF PIX_IN[7312] NB2 NB1 CSA_VREF pixel
xPix7313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[73] VREF PIX_IN[7313] NB2 NB1 CSA_VREF pixel
xPix7314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[73] VREF PIX_IN[7314] NB2 NB1 CSA_VREF pixel
xPix7315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[73] VREF PIX_IN[7315] NB2 NB1 CSA_VREF pixel
xPix7316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[73] VREF PIX_IN[7316] NB2 NB1 CSA_VREF pixel
xPix7317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[73] VREF PIX_IN[7317] NB2 NB1 CSA_VREF pixel
xPix7318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[73] VREF PIX_IN[7318] NB2 NB1 CSA_VREF pixel
xPix7319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[73] VREF PIX_IN[7319] NB2 NB1 CSA_VREF pixel
xPix7320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[73] VREF PIX_IN[7320] NB2 NB1 CSA_VREF pixel
xPix7321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[73] VREF PIX_IN[7321] NB2 NB1 CSA_VREF pixel
xPix7322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[73] VREF PIX_IN[7322] NB2 NB1 CSA_VREF pixel
xPix7323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[73] VREF PIX_IN[7323] NB2 NB1 CSA_VREF pixel
xPix7324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[73] VREF PIX_IN[7324] NB2 NB1 CSA_VREF pixel
xPix7325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[73] VREF PIX_IN[7325] NB2 NB1 CSA_VREF pixel
xPix7326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[73] VREF PIX_IN[7326] NB2 NB1 CSA_VREF pixel
xPix7327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[73] VREF PIX_IN[7327] NB2 NB1 CSA_VREF pixel
xPix7328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[73] VREF PIX_IN[7328] NB2 NB1 CSA_VREF pixel
xPix7329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[73] VREF PIX_IN[7329] NB2 NB1 CSA_VREF pixel
xPix7330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[73] VREF PIX_IN[7330] NB2 NB1 CSA_VREF pixel
xPix7331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[73] VREF PIX_IN[7331] NB2 NB1 CSA_VREF pixel
xPix7332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[73] VREF PIX_IN[7332] NB2 NB1 CSA_VREF pixel
xPix7333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[73] VREF PIX_IN[7333] NB2 NB1 CSA_VREF pixel
xPix7334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[73] VREF PIX_IN[7334] NB2 NB1 CSA_VREF pixel
xPix7335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[73] VREF PIX_IN[7335] NB2 NB1 CSA_VREF pixel
xPix7336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[73] VREF PIX_IN[7336] NB2 NB1 CSA_VREF pixel
xPix7337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[73] VREF PIX_IN[7337] NB2 NB1 CSA_VREF pixel
xPix7338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[73] VREF PIX_IN[7338] NB2 NB1 CSA_VREF pixel
xPix7339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[73] VREF PIX_IN[7339] NB2 NB1 CSA_VREF pixel
xPix7340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[73] VREF PIX_IN[7340] NB2 NB1 CSA_VREF pixel
xPix7341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[73] VREF PIX_IN[7341] NB2 NB1 CSA_VREF pixel
xPix7342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[73] VREF PIX_IN[7342] NB2 NB1 CSA_VREF pixel
xPix7343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[73] VREF PIX_IN[7343] NB2 NB1 CSA_VREF pixel
xPix7344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[73] VREF PIX_IN[7344] NB2 NB1 CSA_VREF pixel
xPix7345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[73] VREF PIX_IN[7345] NB2 NB1 CSA_VREF pixel
xPix7346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[73] VREF PIX_IN[7346] NB2 NB1 CSA_VREF pixel
xPix7347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[73] VREF PIX_IN[7347] NB2 NB1 CSA_VREF pixel
xPix7348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[73] VREF PIX_IN[7348] NB2 NB1 CSA_VREF pixel
xPix7349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[73] VREF PIX_IN[7349] NB2 NB1 CSA_VREF pixel
xPix7350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[73] VREF PIX_IN[7350] NB2 NB1 CSA_VREF pixel
xPix7351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[73] VREF PIX_IN[7351] NB2 NB1 CSA_VREF pixel
xPix7352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[73] VREF PIX_IN[7352] NB2 NB1 CSA_VREF pixel
xPix7353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[73] VREF PIX_IN[7353] NB2 NB1 CSA_VREF pixel
xPix7354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[73] VREF PIX_IN[7354] NB2 NB1 CSA_VREF pixel
xPix7355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[73] VREF PIX_IN[7355] NB2 NB1 CSA_VREF pixel
xPix7356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[73] VREF PIX_IN[7356] NB2 NB1 CSA_VREF pixel
xPix7357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[73] VREF PIX_IN[7357] NB2 NB1 CSA_VREF pixel
xPix7358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[73] VREF PIX_IN[7358] NB2 NB1 CSA_VREF pixel
xPix7359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[73] VREF PIX_IN[7359] NB2 NB1 CSA_VREF pixel
xPix7360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[73] VREF PIX_IN[7360] NB2 NB1 CSA_VREF pixel
xPix7361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[73] VREF PIX_IN[7361] NB2 NB1 CSA_VREF pixel
xPix7362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[73] VREF PIX_IN[7362] NB2 NB1 CSA_VREF pixel
xPix7363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[73] VREF PIX_IN[7363] NB2 NB1 CSA_VREF pixel
xPix7364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[73] VREF PIX_IN[7364] NB2 NB1 CSA_VREF pixel
xPix7365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[73] VREF PIX_IN[7365] NB2 NB1 CSA_VREF pixel
xPix7366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[73] VREF PIX_IN[7366] NB2 NB1 CSA_VREF pixel
xPix7367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[73] VREF PIX_IN[7367] NB2 NB1 CSA_VREF pixel
xPix7368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[73] VREF PIX_IN[7368] NB2 NB1 CSA_VREF pixel
xPix7369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[73] VREF PIX_IN[7369] NB2 NB1 CSA_VREF pixel
xPix7370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[73] VREF PIX_IN[7370] NB2 NB1 CSA_VREF pixel
xPix7371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[73] VREF PIX_IN[7371] NB2 NB1 CSA_VREF pixel
xPix7372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[73] VREF PIX_IN[7372] NB2 NB1 CSA_VREF pixel
xPix7373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[73] VREF PIX_IN[7373] NB2 NB1 CSA_VREF pixel
xPix7374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[73] VREF PIX_IN[7374] NB2 NB1 CSA_VREF pixel
xPix7375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[73] VREF PIX_IN[7375] NB2 NB1 CSA_VREF pixel
xPix7376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[73] VREF PIX_IN[7376] NB2 NB1 CSA_VREF pixel
xPix7377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[73] VREF PIX_IN[7377] NB2 NB1 CSA_VREF pixel
xPix7378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[73] VREF PIX_IN[7378] NB2 NB1 CSA_VREF pixel
xPix7379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[73] VREF PIX_IN[7379] NB2 NB1 CSA_VREF pixel
xPix7380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[73] VREF PIX_IN[7380] NB2 NB1 CSA_VREF pixel
xPix7381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[73] VREF PIX_IN[7381] NB2 NB1 CSA_VREF pixel
xPix7382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[73] VREF PIX_IN[7382] NB2 NB1 CSA_VREF pixel
xPix7383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[73] VREF PIX_IN[7383] NB2 NB1 CSA_VREF pixel
xPix7384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[73] VREF PIX_IN[7384] NB2 NB1 CSA_VREF pixel
xPix7385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[73] VREF PIX_IN[7385] NB2 NB1 CSA_VREF pixel
xPix7386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[73] VREF PIX_IN[7386] NB2 NB1 CSA_VREF pixel
xPix7387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[73] VREF PIX_IN[7387] NB2 NB1 CSA_VREF pixel
xPix7388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[73] VREF PIX_IN[7388] NB2 NB1 CSA_VREF pixel
xPix7389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[73] VREF PIX_IN[7389] NB2 NB1 CSA_VREF pixel
xPix7390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[73] VREF PIX_IN[7390] NB2 NB1 CSA_VREF pixel
xPix7391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[73] VREF PIX_IN[7391] NB2 NB1 CSA_VREF pixel
xPix7392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[73] VREF PIX_IN[7392] NB2 NB1 CSA_VREF pixel
xPix7393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[73] VREF PIX_IN[7393] NB2 NB1 CSA_VREF pixel
xPix7394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[73] VREF PIX_IN[7394] NB2 NB1 CSA_VREF pixel
xPix7395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[73] VREF PIX_IN[7395] NB2 NB1 CSA_VREF pixel
xPix7396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[73] VREF PIX_IN[7396] NB2 NB1 CSA_VREF pixel
xPix7397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[73] VREF PIX_IN[7397] NB2 NB1 CSA_VREF pixel
xPix7398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[73] VREF PIX_IN[7398] NB2 NB1 CSA_VREF pixel
xPix7399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[73] VREF PIX_IN[7399] NB2 NB1 CSA_VREF pixel
xPix7400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[74] VREF PIX_IN[7400] NB2 NB1 CSA_VREF pixel
xPix7401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[74] VREF PIX_IN[7401] NB2 NB1 CSA_VREF pixel
xPix7402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[74] VREF PIX_IN[7402] NB2 NB1 CSA_VREF pixel
xPix7403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[74] VREF PIX_IN[7403] NB2 NB1 CSA_VREF pixel
xPix7404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[74] VREF PIX_IN[7404] NB2 NB1 CSA_VREF pixel
xPix7405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[74] VREF PIX_IN[7405] NB2 NB1 CSA_VREF pixel
xPix7406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[74] VREF PIX_IN[7406] NB2 NB1 CSA_VREF pixel
xPix7407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[74] VREF PIX_IN[7407] NB2 NB1 CSA_VREF pixel
xPix7408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[74] VREF PIX_IN[7408] NB2 NB1 CSA_VREF pixel
xPix7409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[74] VREF PIX_IN[7409] NB2 NB1 CSA_VREF pixel
xPix7410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[74] VREF PIX_IN[7410] NB2 NB1 CSA_VREF pixel
xPix7411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[74] VREF PIX_IN[7411] NB2 NB1 CSA_VREF pixel
xPix7412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[74] VREF PIX_IN[7412] NB2 NB1 CSA_VREF pixel
xPix7413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[74] VREF PIX_IN[7413] NB2 NB1 CSA_VREF pixel
xPix7414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[74] VREF PIX_IN[7414] NB2 NB1 CSA_VREF pixel
xPix7415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[74] VREF PIX_IN[7415] NB2 NB1 CSA_VREF pixel
xPix7416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[74] VREF PIX_IN[7416] NB2 NB1 CSA_VREF pixel
xPix7417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[74] VREF PIX_IN[7417] NB2 NB1 CSA_VREF pixel
xPix7418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[74] VREF PIX_IN[7418] NB2 NB1 CSA_VREF pixel
xPix7419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[74] VREF PIX_IN[7419] NB2 NB1 CSA_VREF pixel
xPix7420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[74] VREF PIX_IN[7420] NB2 NB1 CSA_VREF pixel
xPix7421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[74] VREF PIX_IN[7421] NB2 NB1 CSA_VREF pixel
xPix7422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[74] VREF PIX_IN[7422] NB2 NB1 CSA_VREF pixel
xPix7423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[74] VREF PIX_IN[7423] NB2 NB1 CSA_VREF pixel
xPix7424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[74] VREF PIX_IN[7424] NB2 NB1 CSA_VREF pixel
xPix7425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[74] VREF PIX_IN[7425] NB2 NB1 CSA_VREF pixel
xPix7426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[74] VREF PIX_IN[7426] NB2 NB1 CSA_VREF pixel
xPix7427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[74] VREF PIX_IN[7427] NB2 NB1 CSA_VREF pixel
xPix7428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[74] VREF PIX_IN[7428] NB2 NB1 CSA_VREF pixel
xPix7429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[74] VREF PIX_IN[7429] NB2 NB1 CSA_VREF pixel
xPix7430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[74] VREF PIX_IN[7430] NB2 NB1 CSA_VREF pixel
xPix7431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[74] VREF PIX_IN[7431] NB2 NB1 CSA_VREF pixel
xPix7432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[74] VREF PIX_IN[7432] NB2 NB1 CSA_VREF pixel
xPix7433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[74] VREF PIX_IN[7433] NB2 NB1 CSA_VREF pixel
xPix7434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[74] VREF PIX_IN[7434] NB2 NB1 CSA_VREF pixel
xPix7435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[74] VREF PIX_IN[7435] NB2 NB1 CSA_VREF pixel
xPix7436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[74] VREF PIX_IN[7436] NB2 NB1 CSA_VREF pixel
xPix7437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[74] VREF PIX_IN[7437] NB2 NB1 CSA_VREF pixel
xPix7438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[74] VREF PIX_IN[7438] NB2 NB1 CSA_VREF pixel
xPix7439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[74] VREF PIX_IN[7439] NB2 NB1 CSA_VREF pixel
xPix7440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[74] VREF PIX_IN[7440] NB2 NB1 CSA_VREF pixel
xPix7441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[74] VREF PIX_IN[7441] NB2 NB1 CSA_VREF pixel
xPix7442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[74] VREF PIX_IN[7442] NB2 NB1 CSA_VREF pixel
xPix7443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[74] VREF PIX_IN[7443] NB2 NB1 CSA_VREF pixel
xPix7444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[74] VREF PIX_IN[7444] NB2 NB1 CSA_VREF pixel
xPix7445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[74] VREF PIX_IN[7445] NB2 NB1 CSA_VREF pixel
xPix7446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[74] VREF PIX_IN[7446] NB2 NB1 CSA_VREF pixel
xPix7447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[74] VREF PIX_IN[7447] NB2 NB1 CSA_VREF pixel
xPix7448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[74] VREF PIX_IN[7448] NB2 NB1 CSA_VREF pixel
xPix7449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[74] VREF PIX_IN[7449] NB2 NB1 CSA_VREF pixel
xPix7450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[74] VREF PIX_IN[7450] NB2 NB1 CSA_VREF pixel
xPix7451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[74] VREF PIX_IN[7451] NB2 NB1 CSA_VREF pixel
xPix7452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[74] VREF PIX_IN[7452] NB2 NB1 CSA_VREF pixel
xPix7453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[74] VREF PIX_IN[7453] NB2 NB1 CSA_VREF pixel
xPix7454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[74] VREF PIX_IN[7454] NB2 NB1 CSA_VREF pixel
xPix7455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[74] VREF PIX_IN[7455] NB2 NB1 CSA_VREF pixel
xPix7456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[74] VREF PIX_IN[7456] NB2 NB1 CSA_VREF pixel
xPix7457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[74] VREF PIX_IN[7457] NB2 NB1 CSA_VREF pixel
xPix7458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[74] VREF PIX_IN[7458] NB2 NB1 CSA_VREF pixel
xPix7459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[74] VREF PIX_IN[7459] NB2 NB1 CSA_VREF pixel
xPix7460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[74] VREF PIX_IN[7460] NB2 NB1 CSA_VREF pixel
xPix7461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[74] VREF PIX_IN[7461] NB2 NB1 CSA_VREF pixel
xPix7462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[74] VREF PIX_IN[7462] NB2 NB1 CSA_VREF pixel
xPix7463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[74] VREF PIX_IN[7463] NB2 NB1 CSA_VREF pixel
xPix7464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[74] VREF PIX_IN[7464] NB2 NB1 CSA_VREF pixel
xPix7465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[74] VREF PIX_IN[7465] NB2 NB1 CSA_VREF pixel
xPix7466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[74] VREF PIX_IN[7466] NB2 NB1 CSA_VREF pixel
xPix7467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[74] VREF PIX_IN[7467] NB2 NB1 CSA_VREF pixel
xPix7468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[74] VREF PIX_IN[7468] NB2 NB1 CSA_VREF pixel
xPix7469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[74] VREF PIX_IN[7469] NB2 NB1 CSA_VREF pixel
xPix7470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[74] VREF PIX_IN[7470] NB2 NB1 CSA_VREF pixel
xPix7471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[74] VREF PIX_IN[7471] NB2 NB1 CSA_VREF pixel
xPix7472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[74] VREF PIX_IN[7472] NB2 NB1 CSA_VREF pixel
xPix7473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[74] VREF PIX_IN[7473] NB2 NB1 CSA_VREF pixel
xPix7474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[74] VREF PIX_IN[7474] NB2 NB1 CSA_VREF pixel
xPix7475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[74] VREF PIX_IN[7475] NB2 NB1 CSA_VREF pixel
xPix7476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[74] VREF PIX_IN[7476] NB2 NB1 CSA_VREF pixel
xPix7477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[74] VREF PIX_IN[7477] NB2 NB1 CSA_VREF pixel
xPix7478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[74] VREF PIX_IN[7478] NB2 NB1 CSA_VREF pixel
xPix7479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[74] VREF PIX_IN[7479] NB2 NB1 CSA_VREF pixel
xPix7480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[74] VREF PIX_IN[7480] NB2 NB1 CSA_VREF pixel
xPix7481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[74] VREF PIX_IN[7481] NB2 NB1 CSA_VREF pixel
xPix7482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[74] VREF PIX_IN[7482] NB2 NB1 CSA_VREF pixel
xPix7483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[74] VREF PIX_IN[7483] NB2 NB1 CSA_VREF pixel
xPix7484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[74] VREF PIX_IN[7484] NB2 NB1 CSA_VREF pixel
xPix7485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[74] VREF PIX_IN[7485] NB2 NB1 CSA_VREF pixel
xPix7486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[74] VREF PIX_IN[7486] NB2 NB1 CSA_VREF pixel
xPix7487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[74] VREF PIX_IN[7487] NB2 NB1 CSA_VREF pixel
xPix7488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[74] VREF PIX_IN[7488] NB2 NB1 CSA_VREF pixel
xPix7489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[74] VREF PIX_IN[7489] NB2 NB1 CSA_VREF pixel
xPix7490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[74] VREF PIX_IN[7490] NB2 NB1 CSA_VREF pixel
xPix7491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[74] VREF PIX_IN[7491] NB2 NB1 CSA_VREF pixel
xPix7492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[74] VREF PIX_IN[7492] NB2 NB1 CSA_VREF pixel
xPix7493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[74] VREF PIX_IN[7493] NB2 NB1 CSA_VREF pixel
xPix7494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[74] VREF PIX_IN[7494] NB2 NB1 CSA_VREF pixel
xPix7495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[74] VREF PIX_IN[7495] NB2 NB1 CSA_VREF pixel
xPix7496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[74] VREF PIX_IN[7496] NB2 NB1 CSA_VREF pixel
xPix7497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[74] VREF PIX_IN[7497] NB2 NB1 CSA_VREF pixel
xPix7498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[74] VREF PIX_IN[7498] NB2 NB1 CSA_VREF pixel
xPix7499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[74] VREF PIX_IN[7499] NB2 NB1 CSA_VREF pixel
xPix7500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[75] VREF PIX_IN[7500] NB2 NB1 CSA_VREF pixel
xPix7501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[75] VREF PIX_IN[7501] NB2 NB1 CSA_VREF pixel
xPix7502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[75] VREF PIX_IN[7502] NB2 NB1 CSA_VREF pixel
xPix7503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[75] VREF PIX_IN[7503] NB2 NB1 CSA_VREF pixel
xPix7504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[75] VREF PIX_IN[7504] NB2 NB1 CSA_VREF pixel
xPix7505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[75] VREF PIX_IN[7505] NB2 NB1 CSA_VREF pixel
xPix7506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[75] VREF PIX_IN[7506] NB2 NB1 CSA_VREF pixel
xPix7507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[75] VREF PIX_IN[7507] NB2 NB1 CSA_VREF pixel
xPix7508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[75] VREF PIX_IN[7508] NB2 NB1 CSA_VREF pixel
xPix7509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[75] VREF PIX_IN[7509] NB2 NB1 CSA_VREF pixel
xPix7510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[75] VREF PIX_IN[7510] NB2 NB1 CSA_VREF pixel
xPix7511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[75] VREF PIX_IN[7511] NB2 NB1 CSA_VREF pixel
xPix7512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[75] VREF PIX_IN[7512] NB2 NB1 CSA_VREF pixel
xPix7513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[75] VREF PIX_IN[7513] NB2 NB1 CSA_VREF pixel
xPix7514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[75] VREF PIX_IN[7514] NB2 NB1 CSA_VREF pixel
xPix7515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[75] VREF PIX_IN[7515] NB2 NB1 CSA_VREF pixel
xPix7516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[75] VREF PIX_IN[7516] NB2 NB1 CSA_VREF pixel
xPix7517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[75] VREF PIX_IN[7517] NB2 NB1 CSA_VREF pixel
xPix7518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[75] VREF PIX_IN[7518] NB2 NB1 CSA_VREF pixel
xPix7519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[75] VREF PIX_IN[7519] NB2 NB1 CSA_VREF pixel
xPix7520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[75] VREF PIX_IN[7520] NB2 NB1 CSA_VREF pixel
xPix7521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[75] VREF PIX_IN[7521] NB2 NB1 CSA_VREF pixel
xPix7522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[75] VREF PIX_IN[7522] NB2 NB1 CSA_VREF pixel
xPix7523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[75] VREF PIX_IN[7523] NB2 NB1 CSA_VREF pixel
xPix7524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[75] VREF PIX_IN[7524] NB2 NB1 CSA_VREF pixel
xPix7525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[75] VREF PIX_IN[7525] NB2 NB1 CSA_VREF pixel
xPix7526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[75] VREF PIX_IN[7526] NB2 NB1 CSA_VREF pixel
xPix7527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[75] VREF PIX_IN[7527] NB2 NB1 CSA_VREF pixel
xPix7528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[75] VREF PIX_IN[7528] NB2 NB1 CSA_VREF pixel
xPix7529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[75] VREF PIX_IN[7529] NB2 NB1 CSA_VREF pixel
xPix7530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[75] VREF PIX_IN[7530] NB2 NB1 CSA_VREF pixel
xPix7531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[75] VREF PIX_IN[7531] NB2 NB1 CSA_VREF pixel
xPix7532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[75] VREF PIX_IN[7532] NB2 NB1 CSA_VREF pixel
xPix7533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[75] VREF PIX_IN[7533] NB2 NB1 CSA_VREF pixel
xPix7534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[75] VREF PIX_IN[7534] NB2 NB1 CSA_VREF pixel
xPix7535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[75] VREF PIX_IN[7535] NB2 NB1 CSA_VREF pixel
xPix7536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[75] VREF PIX_IN[7536] NB2 NB1 CSA_VREF pixel
xPix7537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[75] VREF PIX_IN[7537] NB2 NB1 CSA_VREF pixel
xPix7538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[75] VREF PIX_IN[7538] NB2 NB1 CSA_VREF pixel
xPix7539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[75] VREF PIX_IN[7539] NB2 NB1 CSA_VREF pixel
xPix7540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[75] VREF PIX_IN[7540] NB2 NB1 CSA_VREF pixel
xPix7541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[75] VREF PIX_IN[7541] NB2 NB1 CSA_VREF pixel
xPix7542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[75] VREF PIX_IN[7542] NB2 NB1 CSA_VREF pixel
xPix7543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[75] VREF PIX_IN[7543] NB2 NB1 CSA_VREF pixel
xPix7544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[75] VREF PIX_IN[7544] NB2 NB1 CSA_VREF pixel
xPix7545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[75] VREF PIX_IN[7545] NB2 NB1 CSA_VREF pixel
xPix7546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[75] VREF PIX_IN[7546] NB2 NB1 CSA_VREF pixel
xPix7547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[75] VREF PIX_IN[7547] NB2 NB1 CSA_VREF pixel
xPix7548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[75] VREF PIX_IN[7548] NB2 NB1 CSA_VREF pixel
xPix7549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[75] VREF PIX_IN[7549] NB2 NB1 CSA_VREF pixel
xPix7550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[75] VREF PIX_IN[7550] NB2 NB1 CSA_VREF pixel
xPix7551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[75] VREF PIX_IN[7551] NB2 NB1 CSA_VREF pixel
xPix7552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[75] VREF PIX_IN[7552] NB2 NB1 CSA_VREF pixel
xPix7553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[75] VREF PIX_IN[7553] NB2 NB1 CSA_VREF pixel
xPix7554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[75] VREF PIX_IN[7554] NB2 NB1 CSA_VREF pixel
xPix7555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[75] VREF PIX_IN[7555] NB2 NB1 CSA_VREF pixel
xPix7556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[75] VREF PIX_IN[7556] NB2 NB1 CSA_VREF pixel
xPix7557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[75] VREF PIX_IN[7557] NB2 NB1 CSA_VREF pixel
xPix7558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[75] VREF PIX_IN[7558] NB2 NB1 CSA_VREF pixel
xPix7559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[75] VREF PIX_IN[7559] NB2 NB1 CSA_VREF pixel
xPix7560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[75] VREF PIX_IN[7560] NB2 NB1 CSA_VREF pixel
xPix7561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[75] VREF PIX_IN[7561] NB2 NB1 CSA_VREF pixel
xPix7562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[75] VREF PIX_IN[7562] NB2 NB1 CSA_VREF pixel
xPix7563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[75] VREF PIX_IN[7563] NB2 NB1 CSA_VREF pixel
xPix7564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[75] VREF PIX_IN[7564] NB2 NB1 CSA_VREF pixel
xPix7565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[75] VREF PIX_IN[7565] NB2 NB1 CSA_VREF pixel
xPix7566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[75] VREF PIX_IN[7566] NB2 NB1 CSA_VREF pixel
xPix7567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[75] VREF PIX_IN[7567] NB2 NB1 CSA_VREF pixel
xPix7568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[75] VREF PIX_IN[7568] NB2 NB1 CSA_VREF pixel
xPix7569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[75] VREF PIX_IN[7569] NB2 NB1 CSA_VREF pixel
xPix7570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[75] VREF PIX_IN[7570] NB2 NB1 CSA_VREF pixel
xPix7571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[75] VREF PIX_IN[7571] NB2 NB1 CSA_VREF pixel
xPix7572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[75] VREF PIX_IN[7572] NB2 NB1 CSA_VREF pixel
xPix7573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[75] VREF PIX_IN[7573] NB2 NB1 CSA_VREF pixel
xPix7574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[75] VREF PIX_IN[7574] NB2 NB1 CSA_VREF pixel
xPix7575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[75] VREF PIX_IN[7575] NB2 NB1 CSA_VREF pixel
xPix7576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[75] VREF PIX_IN[7576] NB2 NB1 CSA_VREF pixel
xPix7577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[75] VREF PIX_IN[7577] NB2 NB1 CSA_VREF pixel
xPix7578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[75] VREF PIX_IN[7578] NB2 NB1 CSA_VREF pixel
xPix7579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[75] VREF PIX_IN[7579] NB2 NB1 CSA_VREF pixel
xPix7580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[75] VREF PIX_IN[7580] NB2 NB1 CSA_VREF pixel
xPix7581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[75] VREF PIX_IN[7581] NB2 NB1 CSA_VREF pixel
xPix7582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[75] VREF PIX_IN[7582] NB2 NB1 CSA_VREF pixel
xPix7583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[75] VREF PIX_IN[7583] NB2 NB1 CSA_VREF pixel
xPix7584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[75] VREF PIX_IN[7584] NB2 NB1 CSA_VREF pixel
xPix7585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[75] VREF PIX_IN[7585] NB2 NB1 CSA_VREF pixel
xPix7586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[75] VREF PIX_IN[7586] NB2 NB1 CSA_VREF pixel
xPix7587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[75] VREF PIX_IN[7587] NB2 NB1 CSA_VREF pixel
xPix7588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[75] VREF PIX_IN[7588] NB2 NB1 CSA_VREF pixel
xPix7589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[75] VREF PIX_IN[7589] NB2 NB1 CSA_VREF pixel
xPix7590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[75] VREF PIX_IN[7590] NB2 NB1 CSA_VREF pixel
xPix7591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[75] VREF PIX_IN[7591] NB2 NB1 CSA_VREF pixel
xPix7592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[75] VREF PIX_IN[7592] NB2 NB1 CSA_VREF pixel
xPix7593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[75] VREF PIX_IN[7593] NB2 NB1 CSA_VREF pixel
xPix7594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[75] VREF PIX_IN[7594] NB2 NB1 CSA_VREF pixel
xPix7595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[75] VREF PIX_IN[7595] NB2 NB1 CSA_VREF pixel
xPix7596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[75] VREF PIX_IN[7596] NB2 NB1 CSA_VREF pixel
xPix7597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[75] VREF PIX_IN[7597] NB2 NB1 CSA_VREF pixel
xPix7598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[75] VREF PIX_IN[7598] NB2 NB1 CSA_VREF pixel
xPix7599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[75] VREF PIX_IN[7599] NB2 NB1 CSA_VREF pixel
xPix7600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[76] VREF PIX_IN[7600] NB2 NB1 CSA_VREF pixel
xPix7601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[76] VREF PIX_IN[7601] NB2 NB1 CSA_VREF pixel
xPix7602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[76] VREF PIX_IN[7602] NB2 NB1 CSA_VREF pixel
xPix7603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[76] VREF PIX_IN[7603] NB2 NB1 CSA_VREF pixel
xPix7604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[76] VREF PIX_IN[7604] NB2 NB1 CSA_VREF pixel
xPix7605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[76] VREF PIX_IN[7605] NB2 NB1 CSA_VREF pixel
xPix7606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[76] VREF PIX_IN[7606] NB2 NB1 CSA_VREF pixel
xPix7607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[76] VREF PIX_IN[7607] NB2 NB1 CSA_VREF pixel
xPix7608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[76] VREF PIX_IN[7608] NB2 NB1 CSA_VREF pixel
xPix7609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[76] VREF PIX_IN[7609] NB2 NB1 CSA_VREF pixel
xPix7610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[76] VREF PIX_IN[7610] NB2 NB1 CSA_VREF pixel
xPix7611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[76] VREF PIX_IN[7611] NB2 NB1 CSA_VREF pixel
xPix7612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[76] VREF PIX_IN[7612] NB2 NB1 CSA_VREF pixel
xPix7613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[76] VREF PIX_IN[7613] NB2 NB1 CSA_VREF pixel
xPix7614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[76] VREF PIX_IN[7614] NB2 NB1 CSA_VREF pixel
xPix7615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[76] VREF PIX_IN[7615] NB2 NB1 CSA_VREF pixel
xPix7616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[76] VREF PIX_IN[7616] NB2 NB1 CSA_VREF pixel
xPix7617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[76] VREF PIX_IN[7617] NB2 NB1 CSA_VREF pixel
xPix7618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[76] VREF PIX_IN[7618] NB2 NB1 CSA_VREF pixel
xPix7619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[76] VREF PIX_IN[7619] NB2 NB1 CSA_VREF pixel
xPix7620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[76] VREF PIX_IN[7620] NB2 NB1 CSA_VREF pixel
xPix7621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[76] VREF PIX_IN[7621] NB2 NB1 CSA_VREF pixel
xPix7622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[76] VREF PIX_IN[7622] NB2 NB1 CSA_VREF pixel
xPix7623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[76] VREF PIX_IN[7623] NB2 NB1 CSA_VREF pixel
xPix7624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[76] VREF PIX_IN[7624] NB2 NB1 CSA_VREF pixel
xPix7625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[76] VREF PIX_IN[7625] NB2 NB1 CSA_VREF pixel
xPix7626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[76] VREF PIX_IN[7626] NB2 NB1 CSA_VREF pixel
xPix7627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[76] VREF PIX_IN[7627] NB2 NB1 CSA_VREF pixel
xPix7628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[76] VREF PIX_IN[7628] NB2 NB1 CSA_VREF pixel
xPix7629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[76] VREF PIX_IN[7629] NB2 NB1 CSA_VREF pixel
xPix7630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[76] VREF PIX_IN[7630] NB2 NB1 CSA_VREF pixel
xPix7631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[76] VREF PIX_IN[7631] NB2 NB1 CSA_VREF pixel
xPix7632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[76] VREF PIX_IN[7632] NB2 NB1 CSA_VREF pixel
xPix7633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[76] VREF PIX_IN[7633] NB2 NB1 CSA_VREF pixel
xPix7634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[76] VREF PIX_IN[7634] NB2 NB1 CSA_VREF pixel
xPix7635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[76] VREF PIX_IN[7635] NB2 NB1 CSA_VREF pixel
xPix7636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[76] VREF PIX_IN[7636] NB2 NB1 CSA_VREF pixel
xPix7637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[76] VREF PIX_IN[7637] NB2 NB1 CSA_VREF pixel
xPix7638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[76] VREF PIX_IN[7638] NB2 NB1 CSA_VREF pixel
xPix7639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[76] VREF PIX_IN[7639] NB2 NB1 CSA_VREF pixel
xPix7640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[76] VREF PIX_IN[7640] NB2 NB1 CSA_VREF pixel
xPix7641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[76] VREF PIX_IN[7641] NB2 NB1 CSA_VREF pixel
xPix7642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[76] VREF PIX_IN[7642] NB2 NB1 CSA_VREF pixel
xPix7643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[76] VREF PIX_IN[7643] NB2 NB1 CSA_VREF pixel
xPix7644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[76] VREF PIX_IN[7644] NB2 NB1 CSA_VREF pixel
xPix7645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[76] VREF PIX_IN[7645] NB2 NB1 CSA_VREF pixel
xPix7646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[76] VREF PIX_IN[7646] NB2 NB1 CSA_VREF pixel
xPix7647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[76] VREF PIX_IN[7647] NB2 NB1 CSA_VREF pixel
xPix7648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[76] VREF PIX_IN[7648] NB2 NB1 CSA_VREF pixel
xPix7649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[76] VREF PIX_IN[7649] NB2 NB1 CSA_VREF pixel
xPix7650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[76] VREF PIX_IN[7650] NB2 NB1 CSA_VREF pixel
xPix7651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[76] VREF PIX_IN[7651] NB2 NB1 CSA_VREF pixel
xPix7652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[76] VREF PIX_IN[7652] NB2 NB1 CSA_VREF pixel
xPix7653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[76] VREF PIX_IN[7653] NB2 NB1 CSA_VREF pixel
xPix7654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[76] VREF PIX_IN[7654] NB2 NB1 CSA_VREF pixel
xPix7655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[76] VREF PIX_IN[7655] NB2 NB1 CSA_VREF pixel
xPix7656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[76] VREF PIX_IN[7656] NB2 NB1 CSA_VREF pixel
xPix7657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[76] VREF PIX_IN[7657] NB2 NB1 CSA_VREF pixel
xPix7658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[76] VREF PIX_IN[7658] NB2 NB1 CSA_VREF pixel
xPix7659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[76] VREF PIX_IN[7659] NB2 NB1 CSA_VREF pixel
xPix7660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[76] VREF PIX_IN[7660] NB2 NB1 CSA_VREF pixel
xPix7661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[76] VREF PIX_IN[7661] NB2 NB1 CSA_VREF pixel
xPix7662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[76] VREF PIX_IN[7662] NB2 NB1 CSA_VREF pixel
xPix7663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[76] VREF PIX_IN[7663] NB2 NB1 CSA_VREF pixel
xPix7664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[76] VREF PIX_IN[7664] NB2 NB1 CSA_VREF pixel
xPix7665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[76] VREF PIX_IN[7665] NB2 NB1 CSA_VREF pixel
xPix7666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[76] VREF PIX_IN[7666] NB2 NB1 CSA_VREF pixel
xPix7667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[76] VREF PIX_IN[7667] NB2 NB1 CSA_VREF pixel
xPix7668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[76] VREF PIX_IN[7668] NB2 NB1 CSA_VREF pixel
xPix7669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[76] VREF PIX_IN[7669] NB2 NB1 CSA_VREF pixel
xPix7670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[76] VREF PIX_IN[7670] NB2 NB1 CSA_VREF pixel
xPix7671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[76] VREF PIX_IN[7671] NB2 NB1 CSA_VREF pixel
xPix7672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[76] VREF PIX_IN[7672] NB2 NB1 CSA_VREF pixel
xPix7673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[76] VREF PIX_IN[7673] NB2 NB1 CSA_VREF pixel
xPix7674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[76] VREF PIX_IN[7674] NB2 NB1 CSA_VREF pixel
xPix7675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[76] VREF PIX_IN[7675] NB2 NB1 CSA_VREF pixel
xPix7676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[76] VREF PIX_IN[7676] NB2 NB1 CSA_VREF pixel
xPix7677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[76] VREF PIX_IN[7677] NB2 NB1 CSA_VREF pixel
xPix7678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[76] VREF PIX_IN[7678] NB2 NB1 CSA_VREF pixel
xPix7679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[76] VREF PIX_IN[7679] NB2 NB1 CSA_VREF pixel
xPix7680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[76] VREF PIX_IN[7680] NB2 NB1 CSA_VREF pixel
xPix7681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[76] VREF PIX_IN[7681] NB2 NB1 CSA_VREF pixel
xPix7682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[76] VREF PIX_IN[7682] NB2 NB1 CSA_VREF pixel
xPix7683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[76] VREF PIX_IN[7683] NB2 NB1 CSA_VREF pixel
xPix7684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[76] VREF PIX_IN[7684] NB2 NB1 CSA_VREF pixel
xPix7685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[76] VREF PIX_IN[7685] NB2 NB1 CSA_VREF pixel
xPix7686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[76] VREF PIX_IN[7686] NB2 NB1 CSA_VREF pixel
xPix7687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[76] VREF PIX_IN[7687] NB2 NB1 CSA_VREF pixel
xPix7688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[76] VREF PIX_IN[7688] NB2 NB1 CSA_VREF pixel
xPix7689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[76] VREF PIX_IN[7689] NB2 NB1 CSA_VREF pixel
xPix7690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[76] VREF PIX_IN[7690] NB2 NB1 CSA_VREF pixel
xPix7691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[76] VREF PIX_IN[7691] NB2 NB1 CSA_VREF pixel
xPix7692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[76] VREF PIX_IN[7692] NB2 NB1 CSA_VREF pixel
xPix7693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[76] VREF PIX_IN[7693] NB2 NB1 CSA_VREF pixel
xPix7694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[76] VREF PIX_IN[7694] NB2 NB1 CSA_VREF pixel
xPix7695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[76] VREF PIX_IN[7695] NB2 NB1 CSA_VREF pixel
xPix7696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[76] VREF PIX_IN[7696] NB2 NB1 CSA_VREF pixel
xPix7697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[76] VREF PIX_IN[7697] NB2 NB1 CSA_VREF pixel
xPix7698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[76] VREF PIX_IN[7698] NB2 NB1 CSA_VREF pixel
xPix7699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[76] VREF PIX_IN[7699] NB2 NB1 CSA_VREF pixel
xPix7700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[77] VREF PIX_IN[7700] NB2 NB1 CSA_VREF pixel
xPix7701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[77] VREF PIX_IN[7701] NB2 NB1 CSA_VREF pixel
xPix7702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[77] VREF PIX_IN[7702] NB2 NB1 CSA_VREF pixel
xPix7703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[77] VREF PIX_IN[7703] NB2 NB1 CSA_VREF pixel
xPix7704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[77] VREF PIX_IN[7704] NB2 NB1 CSA_VREF pixel
xPix7705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[77] VREF PIX_IN[7705] NB2 NB1 CSA_VREF pixel
xPix7706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[77] VREF PIX_IN[7706] NB2 NB1 CSA_VREF pixel
xPix7707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[77] VREF PIX_IN[7707] NB2 NB1 CSA_VREF pixel
xPix7708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[77] VREF PIX_IN[7708] NB2 NB1 CSA_VREF pixel
xPix7709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[77] VREF PIX_IN[7709] NB2 NB1 CSA_VREF pixel
xPix7710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[77] VREF PIX_IN[7710] NB2 NB1 CSA_VREF pixel
xPix7711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[77] VREF PIX_IN[7711] NB2 NB1 CSA_VREF pixel
xPix7712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[77] VREF PIX_IN[7712] NB2 NB1 CSA_VREF pixel
xPix7713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[77] VREF PIX_IN[7713] NB2 NB1 CSA_VREF pixel
xPix7714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[77] VREF PIX_IN[7714] NB2 NB1 CSA_VREF pixel
xPix7715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[77] VREF PIX_IN[7715] NB2 NB1 CSA_VREF pixel
xPix7716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[77] VREF PIX_IN[7716] NB2 NB1 CSA_VREF pixel
xPix7717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[77] VREF PIX_IN[7717] NB2 NB1 CSA_VREF pixel
xPix7718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[77] VREF PIX_IN[7718] NB2 NB1 CSA_VREF pixel
xPix7719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[77] VREF PIX_IN[7719] NB2 NB1 CSA_VREF pixel
xPix7720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[77] VREF PIX_IN[7720] NB2 NB1 CSA_VREF pixel
xPix7721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[77] VREF PIX_IN[7721] NB2 NB1 CSA_VREF pixel
xPix7722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[77] VREF PIX_IN[7722] NB2 NB1 CSA_VREF pixel
xPix7723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[77] VREF PIX_IN[7723] NB2 NB1 CSA_VREF pixel
xPix7724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[77] VREF PIX_IN[7724] NB2 NB1 CSA_VREF pixel
xPix7725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[77] VREF PIX_IN[7725] NB2 NB1 CSA_VREF pixel
xPix7726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[77] VREF PIX_IN[7726] NB2 NB1 CSA_VREF pixel
xPix7727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[77] VREF PIX_IN[7727] NB2 NB1 CSA_VREF pixel
xPix7728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[77] VREF PIX_IN[7728] NB2 NB1 CSA_VREF pixel
xPix7729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[77] VREF PIX_IN[7729] NB2 NB1 CSA_VREF pixel
xPix7730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[77] VREF PIX_IN[7730] NB2 NB1 CSA_VREF pixel
xPix7731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[77] VREF PIX_IN[7731] NB2 NB1 CSA_VREF pixel
xPix7732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[77] VREF PIX_IN[7732] NB2 NB1 CSA_VREF pixel
xPix7733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[77] VREF PIX_IN[7733] NB2 NB1 CSA_VREF pixel
xPix7734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[77] VREF PIX_IN[7734] NB2 NB1 CSA_VREF pixel
xPix7735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[77] VREF PIX_IN[7735] NB2 NB1 CSA_VREF pixel
xPix7736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[77] VREF PIX_IN[7736] NB2 NB1 CSA_VREF pixel
xPix7737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[77] VREF PIX_IN[7737] NB2 NB1 CSA_VREF pixel
xPix7738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[77] VREF PIX_IN[7738] NB2 NB1 CSA_VREF pixel
xPix7739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[77] VREF PIX_IN[7739] NB2 NB1 CSA_VREF pixel
xPix7740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[77] VREF PIX_IN[7740] NB2 NB1 CSA_VREF pixel
xPix7741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[77] VREF PIX_IN[7741] NB2 NB1 CSA_VREF pixel
xPix7742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[77] VREF PIX_IN[7742] NB2 NB1 CSA_VREF pixel
xPix7743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[77] VREF PIX_IN[7743] NB2 NB1 CSA_VREF pixel
xPix7744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[77] VREF PIX_IN[7744] NB2 NB1 CSA_VREF pixel
xPix7745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[77] VREF PIX_IN[7745] NB2 NB1 CSA_VREF pixel
xPix7746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[77] VREF PIX_IN[7746] NB2 NB1 CSA_VREF pixel
xPix7747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[77] VREF PIX_IN[7747] NB2 NB1 CSA_VREF pixel
xPix7748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[77] VREF PIX_IN[7748] NB2 NB1 CSA_VREF pixel
xPix7749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[77] VREF PIX_IN[7749] NB2 NB1 CSA_VREF pixel
xPix7750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[77] VREF PIX_IN[7750] NB2 NB1 CSA_VREF pixel
xPix7751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[77] VREF PIX_IN[7751] NB2 NB1 CSA_VREF pixel
xPix7752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[77] VREF PIX_IN[7752] NB2 NB1 CSA_VREF pixel
xPix7753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[77] VREF PIX_IN[7753] NB2 NB1 CSA_VREF pixel
xPix7754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[77] VREF PIX_IN[7754] NB2 NB1 CSA_VREF pixel
xPix7755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[77] VREF PIX_IN[7755] NB2 NB1 CSA_VREF pixel
xPix7756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[77] VREF PIX_IN[7756] NB2 NB1 CSA_VREF pixel
xPix7757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[77] VREF PIX_IN[7757] NB2 NB1 CSA_VREF pixel
xPix7758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[77] VREF PIX_IN[7758] NB2 NB1 CSA_VREF pixel
xPix7759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[77] VREF PIX_IN[7759] NB2 NB1 CSA_VREF pixel
xPix7760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[77] VREF PIX_IN[7760] NB2 NB1 CSA_VREF pixel
xPix7761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[77] VREF PIX_IN[7761] NB2 NB1 CSA_VREF pixel
xPix7762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[77] VREF PIX_IN[7762] NB2 NB1 CSA_VREF pixel
xPix7763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[77] VREF PIX_IN[7763] NB2 NB1 CSA_VREF pixel
xPix7764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[77] VREF PIX_IN[7764] NB2 NB1 CSA_VREF pixel
xPix7765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[77] VREF PIX_IN[7765] NB2 NB1 CSA_VREF pixel
xPix7766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[77] VREF PIX_IN[7766] NB2 NB1 CSA_VREF pixel
xPix7767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[77] VREF PIX_IN[7767] NB2 NB1 CSA_VREF pixel
xPix7768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[77] VREF PIX_IN[7768] NB2 NB1 CSA_VREF pixel
xPix7769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[77] VREF PIX_IN[7769] NB2 NB1 CSA_VREF pixel
xPix7770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[77] VREF PIX_IN[7770] NB2 NB1 CSA_VREF pixel
xPix7771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[77] VREF PIX_IN[7771] NB2 NB1 CSA_VREF pixel
xPix7772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[77] VREF PIX_IN[7772] NB2 NB1 CSA_VREF pixel
xPix7773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[77] VREF PIX_IN[7773] NB2 NB1 CSA_VREF pixel
xPix7774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[77] VREF PIX_IN[7774] NB2 NB1 CSA_VREF pixel
xPix7775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[77] VREF PIX_IN[7775] NB2 NB1 CSA_VREF pixel
xPix7776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[77] VREF PIX_IN[7776] NB2 NB1 CSA_VREF pixel
xPix7777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[77] VREF PIX_IN[7777] NB2 NB1 CSA_VREF pixel
xPix7778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[77] VREF PIX_IN[7778] NB2 NB1 CSA_VREF pixel
xPix7779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[77] VREF PIX_IN[7779] NB2 NB1 CSA_VREF pixel
xPix7780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[77] VREF PIX_IN[7780] NB2 NB1 CSA_VREF pixel
xPix7781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[77] VREF PIX_IN[7781] NB2 NB1 CSA_VREF pixel
xPix7782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[77] VREF PIX_IN[7782] NB2 NB1 CSA_VREF pixel
xPix7783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[77] VREF PIX_IN[7783] NB2 NB1 CSA_VREF pixel
xPix7784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[77] VREF PIX_IN[7784] NB2 NB1 CSA_VREF pixel
xPix7785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[77] VREF PIX_IN[7785] NB2 NB1 CSA_VREF pixel
xPix7786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[77] VREF PIX_IN[7786] NB2 NB1 CSA_VREF pixel
xPix7787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[77] VREF PIX_IN[7787] NB2 NB1 CSA_VREF pixel
xPix7788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[77] VREF PIX_IN[7788] NB2 NB1 CSA_VREF pixel
xPix7789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[77] VREF PIX_IN[7789] NB2 NB1 CSA_VREF pixel
xPix7790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[77] VREF PIX_IN[7790] NB2 NB1 CSA_VREF pixel
xPix7791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[77] VREF PIX_IN[7791] NB2 NB1 CSA_VREF pixel
xPix7792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[77] VREF PIX_IN[7792] NB2 NB1 CSA_VREF pixel
xPix7793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[77] VREF PIX_IN[7793] NB2 NB1 CSA_VREF pixel
xPix7794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[77] VREF PIX_IN[7794] NB2 NB1 CSA_VREF pixel
xPix7795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[77] VREF PIX_IN[7795] NB2 NB1 CSA_VREF pixel
xPix7796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[77] VREF PIX_IN[7796] NB2 NB1 CSA_VREF pixel
xPix7797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[77] VREF PIX_IN[7797] NB2 NB1 CSA_VREF pixel
xPix7798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[77] VREF PIX_IN[7798] NB2 NB1 CSA_VREF pixel
xPix7799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[77] VREF PIX_IN[7799] NB2 NB1 CSA_VREF pixel
xPix7800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[78] VREF PIX_IN[7800] NB2 NB1 CSA_VREF pixel
xPix7801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[78] VREF PIX_IN[7801] NB2 NB1 CSA_VREF pixel
xPix7802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[78] VREF PIX_IN[7802] NB2 NB1 CSA_VREF pixel
xPix7803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[78] VREF PIX_IN[7803] NB2 NB1 CSA_VREF pixel
xPix7804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[78] VREF PIX_IN[7804] NB2 NB1 CSA_VREF pixel
xPix7805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[78] VREF PIX_IN[7805] NB2 NB1 CSA_VREF pixel
xPix7806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[78] VREF PIX_IN[7806] NB2 NB1 CSA_VREF pixel
xPix7807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[78] VREF PIX_IN[7807] NB2 NB1 CSA_VREF pixel
xPix7808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[78] VREF PIX_IN[7808] NB2 NB1 CSA_VREF pixel
xPix7809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[78] VREF PIX_IN[7809] NB2 NB1 CSA_VREF pixel
xPix7810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[78] VREF PIX_IN[7810] NB2 NB1 CSA_VREF pixel
xPix7811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[78] VREF PIX_IN[7811] NB2 NB1 CSA_VREF pixel
xPix7812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[78] VREF PIX_IN[7812] NB2 NB1 CSA_VREF pixel
xPix7813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[78] VREF PIX_IN[7813] NB2 NB1 CSA_VREF pixel
xPix7814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[78] VREF PIX_IN[7814] NB2 NB1 CSA_VREF pixel
xPix7815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[78] VREF PIX_IN[7815] NB2 NB1 CSA_VREF pixel
xPix7816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[78] VREF PIX_IN[7816] NB2 NB1 CSA_VREF pixel
xPix7817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[78] VREF PIX_IN[7817] NB2 NB1 CSA_VREF pixel
xPix7818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[78] VREF PIX_IN[7818] NB2 NB1 CSA_VREF pixel
xPix7819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[78] VREF PIX_IN[7819] NB2 NB1 CSA_VREF pixel
xPix7820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[78] VREF PIX_IN[7820] NB2 NB1 CSA_VREF pixel
xPix7821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[78] VREF PIX_IN[7821] NB2 NB1 CSA_VREF pixel
xPix7822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[78] VREF PIX_IN[7822] NB2 NB1 CSA_VREF pixel
xPix7823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[78] VREF PIX_IN[7823] NB2 NB1 CSA_VREF pixel
xPix7824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[78] VREF PIX_IN[7824] NB2 NB1 CSA_VREF pixel
xPix7825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[78] VREF PIX_IN[7825] NB2 NB1 CSA_VREF pixel
xPix7826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[78] VREF PIX_IN[7826] NB2 NB1 CSA_VREF pixel
xPix7827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[78] VREF PIX_IN[7827] NB2 NB1 CSA_VREF pixel
xPix7828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[78] VREF PIX_IN[7828] NB2 NB1 CSA_VREF pixel
xPix7829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[78] VREF PIX_IN[7829] NB2 NB1 CSA_VREF pixel
xPix7830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[78] VREF PIX_IN[7830] NB2 NB1 CSA_VREF pixel
xPix7831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[78] VREF PIX_IN[7831] NB2 NB1 CSA_VREF pixel
xPix7832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[78] VREF PIX_IN[7832] NB2 NB1 CSA_VREF pixel
xPix7833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[78] VREF PIX_IN[7833] NB2 NB1 CSA_VREF pixel
xPix7834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[78] VREF PIX_IN[7834] NB2 NB1 CSA_VREF pixel
xPix7835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[78] VREF PIX_IN[7835] NB2 NB1 CSA_VREF pixel
xPix7836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[78] VREF PIX_IN[7836] NB2 NB1 CSA_VREF pixel
xPix7837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[78] VREF PIX_IN[7837] NB2 NB1 CSA_VREF pixel
xPix7838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[78] VREF PIX_IN[7838] NB2 NB1 CSA_VREF pixel
xPix7839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[78] VREF PIX_IN[7839] NB2 NB1 CSA_VREF pixel
xPix7840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[78] VREF PIX_IN[7840] NB2 NB1 CSA_VREF pixel
xPix7841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[78] VREF PIX_IN[7841] NB2 NB1 CSA_VREF pixel
xPix7842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[78] VREF PIX_IN[7842] NB2 NB1 CSA_VREF pixel
xPix7843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[78] VREF PIX_IN[7843] NB2 NB1 CSA_VREF pixel
xPix7844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[78] VREF PIX_IN[7844] NB2 NB1 CSA_VREF pixel
xPix7845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[78] VREF PIX_IN[7845] NB2 NB1 CSA_VREF pixel
xPix7846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[78] VREF PIX_IN[7846] NB2 NB1 CSA_VREF pixel
xPix7847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[78] VREF PIX_IN[7847] NB2 NB1 CSA_VREF pixel
xPix7848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[78] VREF PIX_IN[7848] NB2 NB1 CSA_VREF pixel
xPix7849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[78] VREF PIX_IN[7849] NB2 NB1 CSA_VREF pixel
xPix7850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[78] VREF PIX_IN[7850] NB2 NB1 CSA_VREF pixel
xPix7851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[78] VREF PIX_IN[7851] NB2 NB1 CSA_VREF pixel
xPix7852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[78] VREF PIX_IN[7852] NB2 NB1 CSA_VREF pixel
xPix7853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[78] VREF PIX_IN[7853] NB2 NB1 CSA_VREF pixel
xPix7854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[78] VREF PIX_IN[7854] NB2 NB1 CSA_VREF pixel
xPix7855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[78] VREF PIX_IN[7855] NB2 NB1 CSA_VREF pixel
xPix7856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[78] VREF PIX_IN[7856] NB2 NB1 CSA_VREF pixel
xPix7857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[78] VREF PIX_IN[7857] NB2 NB1 CSA_VREF pixel
xPix7858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[78] VREF PIX_IN[7858] NB2 NB1 CSA_VREF pixel
xPix7859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[78] VREF PIX_IN[7859] NB2 NB1 CSA_VREF pixel
xPix7860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[78] VREF PIX_IN[7860] NB2 NB1 CSA_VREF pixel
xPix7861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[78] VREF PIX_IN[7861] NB2 NB1 CSA_VREF pixel
xPix7862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[78] VREF PIX_IN[7862] NB2 NB1 CSA_VREF pixel
xPix7863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[78] VREF PIX_IN[7863] NB2 NB1 CSA_VREF pixel
xPix7864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[78] VREF PIX_IN[7864] NB2 NB1 CSA_VREF pixel
xPix7865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[78] VREF PIX_IN[7865] NB2 NB1 CSA_VREF pixel
xPix7866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[78] VREF PIX_IN[7866] NB2 NB1 CSA_VREF pixel
xPix7867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[78] VREF PIX_IN[7867] NB2 NB1 CSA_VREF pixel
xPix7868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[78] VREF PIX_IN[7868] NB2 NB1 CSA_VREF pixel
xPix7869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[78] VREF PIX_IN[7869] NB2 NB1 CSA_VREF pixel
xPix7870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[78] VREF PIX_IN[7870] NB2 NB1 CSA_VREF pixel
xPix7871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[78] VREF PIX_IN[7871] NB2 NB1 CSA_VREF pixel
xPix7872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[78] VREF PIX_IN[7872] NB2 NB1 CSA_VREF pixel
xPix7873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[78] VREF PIX_IN[7873] NB2 NB1 CSA_VREF pixel
xPix7874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[78] VREF PIX_IN[7874] NB2 NB1 CSA_VREF pixel
xPix7875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[78] VREF PIX_IN[7875] NB2 NB1 CSA_VREF pixel
xPix7876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[78] VREF PIX_IN[7876] NB2 NB1 CSA_VREF pixel
xPix7877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[78] VREF PIX_IN[7877] NB2 NB1 CSA_VREF pixel
xPix7878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[78] VREF PIX_IN[7878] NB2 NB1 CSA_VREF pixel
xPix7879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[78] VREF PIX_IN[7879] NB2 NB1 CSA_VREF pixel
xPix7880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[78] VREF PIX_IN[7880] NB2 NB1 CSA_VREF pixel
xPix7881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[78] VREF PIX_IN[7881] NB2 NB1 CSA_VREF pixel
xPix7882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[78] VREF PIX_IN[7882] NB2 NB1 CSA_VREF pixel
xPix7883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[78] VREF PIX_IN[7883] NB2 NB1 CSA_VREF pixel
xPix7884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[78] VREF PIX_IN[7884] NB2 NB1 CSA_VREF pixel
xPix7885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[78] VREF PIX_IN[7885] NB2 NB1 CSA_VREF pixel
xPix7886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[78] VREF PIX_IN[7886] NB2 NB1 CSA_VREF pixel
xPix7887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[78] VREF PIX_IN[7887] NB2 NB1 CSA_VREF pixel
xPix7888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[78] VREF PIX_IN[7888] NB2 NB1 CSA_VREF pixel
xPix7889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[78] VREF PIX_IN[7889] NB2 NB1 CSA_VREF pixel
xPix7890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[78] VREF PIX_IN[7890] NB2 NB1 CSA_VREF pixel
xPix7891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[78] VREF PIX_IN[7891] NB2 NB1 CSA_VREF pixel
xPix7892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[78] VREF PIX_IN[7892] NB2 NB1 CSA_VREF pixel
xPix7893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[78] VREF PIX_IN[7893] NB2 NB1 CSA_VREF pixel
xPix7894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[78] VREF PIX_IN[7894] NB2 NB1 CSA_VREF pixel
xPix7895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[78] VREF PIX_IN[7895] NB2 NB1 CSA_VREF pixel
xPix7896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[78] VREF PIX_IN[7896] NB2 NB1 CSA_VREF pixel
xPix7897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[78] VREF PIX_IN[7897] NB2 NB1 CSA_VREF pixel
xPix7898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[78] VREF PIX_IN[7898] NB2 NB1 CSA_VREF pixel
xPix7899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[78] VREF PIX_IN[7899] NB2 NB1 CSA_VREF pixel
xPix7900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[79] VREF PIX_IN[7900] NB2 NB1 CSA_VREF pixel
xPix7901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[79] VREF PIX_IN[7901] NB2 NB1 CSA_VREF pixel
xPix7902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[79] VREF PIX_IN[7902] NB2 NB1 CSA_VREF pixel
xPix7903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[79] VREF PIX_IN[7903] NB2 NB1 CSA_VREF pixel
xPix7904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[79] VREF PIX_IN[7904] NB2 NB1 CSA_VREF pixel
xPix7905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[79] VREF PIX_IN[7905] NB2 NB1 CSA_VREF pixel
xPix7906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[79] VREF PIX_IN[7906] NB2 NB1 CSA_VREF pixel
xPix7907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[79] VREF PIX_IN[7907] NB2 NB1 CSA_VREF pixel
xPix7908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[79] VREF PIX_IN[7908] NB2 NB1 CSA_VREF pixel
xPix7909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[79] VREF PIX_IN[7909] NB2 NB1 CSA_VREF pixel
xPix7910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[79] VREF PIX_IN[7910] NB2 NB1 CSA_VREF pixel
xPix7911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[79] VREF PIX_IN[7911] NB2 NB1 CSA_VREF pixel
xPix7912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[79] VREF PIX_IN[7912] NB2 NB1 CSA_VREF pixel
xPix7913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[79] VREF PIX_IN[7913] NB2 NB1 CSA_VREF pixel
xPix7914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[79] VREF PIX_IN[7914] NB2 NB1 CSA_VREF pixel
xPix7915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[79] VREF PIX_IN[7915] NB2 NB1 CSA_VREF pixel
xPix7916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[79] VREF PIX_IN[7916] NB2 NB1 CSA_VREF pixel
xPix7917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[79] VREF PIX_IN[7917] NB2 NB1 CSA_VREF pixel
xPix7918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[79] VREF PIX_IN[7918] NB2 NB1 CSA_VREF pixel
xPix7919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[79] VREF PIX_IN[7919] NB2 NB1 CSA_VREF pixel
xPix7920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[79] VREF PIX_IN[7920] NB2 NB1 CSA_VREF pixel
xPix7921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[79] VREF PIX_IN[7921] NB2 NB1 CSA_VREF pixel
xPix7922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[79] VREF PIX_IN[7922] NB2 NB1 CSA_VREF pixel
xPix7923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[79] VREF PIX_IN[7923] NB2 NB1 CSA_VREF pixel
xPix7924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[79] VREF PIX_IN[7924] NB2 NB1 CSA_VREF pixel
xPix7925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[79] VREF PIX_IN[7925] NB2 NB1 CSA_VREF pixel
xPix7926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[79] VREF PIX_IN[7926] NB2 NB1 CSA_VREF pixel
xPix7927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[79] VREF PIX_IN[7927] NB2 NB1 CSA_VREF pixel
xPix7928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[79] VREF PIX_IN[7928] NB2 NB1 CSA_VREF pixel
xPix7929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[79] VREF PIX_IN[7929] NB2 NB1 CSA_VREF pixel
xPix7930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[79] VREF PIX_IN[7930] NB2 NB1 CSA_VREF pixel
xPix7931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[79] VREF PIX_IN[7931] NB2 NB1 CSA_VREF pixel
xPix7932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[79] VREF PIX_IN[7932] NB2 NB1 CSA_VREF pixel
xPix7933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[79] VREF PIX_IN[7933] NB2 NB1 CSA_VREF pixel
xPix7934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[79] VREF PIX_IN[7934] NB2 NB1 CSA_VREF pixel
xPix7935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[79] VREF PIX_IN[7935] NB2 NB1 CSA_VREF pixel
xPix7936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[79] VREF PIX_IN[7936] NB2 NB1 CSA_VREF pixel
xPix7937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[79] VREF PIX_IN[7937] NB2 NB1 CSA_VREF pixel
xPix7938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[79] VREF PIX_IN[7938] NB2 NB1 CSA_VREF pixel
xPix7939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[79] VREF PIX_IN[7939] NB2 NB1 CSA_VREF pixel
xPix7940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[79] VREF PIX_IN[7940] NB2 NB1 CSA_VREF pixel
xPix7941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[79] VREF PIX_IN[7941] NB2 NB1 CSA_VREF pixel
xPix7942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[79] VREF PIX_IN[7942] NB2 NB1 CSA_VREF pixel
xPix7943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[79] VREF PIX_IN[7943] NB2 NB1 CSA_VREF pixel
xPix7944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[79] VREF PIX_IN[7944] NB2 NB1 CSA_VREF pixel
xPix7945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[79] VREF PIX_IN[7945] NB2 NB1 CSA_VREF pixel
xPix7946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[79] VREF PIX_IN[7946] NB2 NB1 CSA_VREF pixel
xPix7947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[79] VREF PIX_IN[7947] NB2 NB1 CSA_VREF pixel
xPix7948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[79] VREF PIX_IN[7948] NB2 NB1 CSA_VREF pixel
xPix7949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[79] VREF PIX_IN[7949] NB2 NB1 CSA_VREF pixel
xPix7950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[79] VREF PIX_IN[7950] NB2 NB1 CSA_VREF pixel
xPix7951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[79] VREF PIX_IN[7951] NB2 NB1 CSA_VREF pixel
xPix7952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[79] VREF PIX_IN[7952] NB2 NB1 CSA_VREF pixel
xPix7953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[79] VREF PIX_IN[7953] NB2 NB1 CSA_VREF pixel
xPix7954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[79] VREF PIX_IN[7954] NB2 NB1 CSA_VREF pixel
xPix7955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[79] VREF PIX_IN[7955] NB2 NB1 CSA_VREF pixel
xPix7956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[79] VREF PIX_IN[7956] NB2 NB1 CSA_VREF pixel
xPix7957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[79] VREF PIX_IN[7957] NB2 NB1 CSA_VREF pixel
xPix7958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[79] VREF PIX_IN[7958] NB2 NB1 CSA_VREF pixel
xPix7959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[79] VREF PIX_IN[7959] NB2 NB1 CSA_VREF pixel
xPix7960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[79] VREF PIX_IN[7960] NB2 NB1 CSA_VREF pixel
xPix7961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[79] VREF PIX_IN[7961] NB2 NB1 CSA_VREF pixel
xPix7962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[79] VREF PIX_IN[7962] NB2 NB1 CSA_VREF pixel
xPix7963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[79] VREF PIX_IN[7963] NB2 NB1 CSA_VREF pixel
xPix7964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[79] VREF PIX_IN[7964] NB2 NB1 CSA_VREF pixel
xPix7965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[79] VREF PIX_IN[7965] NB2 NB1 CSA_VREF pixel
xPix7966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[79] VREF PIX_IN[7966] NB2 NB1 CSA_VREF pixel
xPix7967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[79] VREF PIX_IN[7967] NB2 NB1 CSA_VREF pixel
xPix7968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[79] VREF PIX_IN[7968] NB2 NB1 CSA_VREF pixel
xPix7969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[79] VREF PIX_IN[7969] NB2 NB1 CSA_VREF pixel
xPix7970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[79] VREF PIX_IN[7970] NB2 NB1 CSA_VREF pixel
xPix7971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[79] VREF PIX_IN[7971] NB2 NB1 CSA_VREF pixel
xPix7972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[79] VREF PIX_IN[7972] NB2 NB1 CSA_VREF pixel
xPix7973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[79] VREF PIX_IN[7973] NB2 NB1 CSA_VREF pixel
xPix7974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[79] VREF PIX_IN[7974] NB2 NB1 CSA_VREF pixel
xPix7975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[79] VREF PIX_IN[7975] NB2 NB1 CSA_VREF pixel
xPix7976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[79] VREF PIX_IN[7976] NB2 NB1 CSA_VREF pixel
xPix7977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[79] VREF PIX_IN[7977] NB2 NB1 CSA_VREF pixel
xPix7978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[79] VREF PIX_IN[7978] NB2 NB1 CSA_VREF pixel
xPix7979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[79] VREF PIX_IN[7979] NB2 NB1 CSA_VREF pixel
xPix7980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[79] VREF PIX_IN[7980] NB2 NB1 CSA_VREF pixel
xPix7981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[79] VREF PIX_IN[7981] NB2 NB1 CSA_VREF pixel
xPix7982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[79] VREF PIX_IN[7982] NB2 NB1 CSA_VREF pixel
xPix7983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[79] VREF PIX_IN[7983] NB2 NB1 CSA_VREF pixel
xPix7984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[79] VREF PIX_IN[7984] NB2 NB1 CSA_VREF pixel
xPix7985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[79] VREF PIX_IN[7985] NB2 NB1 CSA_VREF pixel
xPix7986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[79] VREF PIX_IN[7986] NB2 NB1 CSA_VREF pixel
xPix7987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[79] VREF PIX_IN[7987] NB2 NB1 CSA_VREF pixel
xPix7988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[79] VREF PIX_IN[7988] NB2 NB1 CSA_VREF pixel
xPix7989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[79] VREF PIX_IN[7989] NB2 NB1 CSA_VREF pixel
xPix7990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[79] VREF PIX_IN[7990] NB2 NB1 CSA_VREF pixel
xPix7991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[79] VREF PIX_IN[7991] NB2 NB1 CSA_VREF pixel
xPix7992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[79] VREF PIX_IN[7992] NB2 NB1 CSA_VREF pixel
xPix7993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[79] VREF PIX_IN[7993] NB2 NB1 CSA_VREF pixel
xPix7994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[79] VREF PIX_IN[7994] NB2 NB1 CSA_VREF pixel
xPix7995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[79] VREF PIX_IN[7995] NB2 NB1 CSA_VREF pixel
xPix7996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[79] VREF PIX_IN[7996] NB2 NB1 CSA_VREF pixel
xPix7997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[79] VREF PIX_IN[7997] NB2 NB1 CSA_VREF pixel
xPix7998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[79] VREF PIX_IN[7998] NB2 NB1 CSA_VREF pixel
xPix7999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[79] VREF PIX_IN[7999] NB2 NB1 CSA_VREF pixel
xPix8000 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[80] VREF PIX_IN[8000] NB2 NB1 CSA_VREF pixel
xPix8001 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[80] VREF PIX_IN[8001] NB2 NB1 CSA_VREF pixel
xPix8002 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[80] VREF PIX_IN[8002] NB2 NB1 CSA_VREF pixel
xPix8003 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[80] VREF PIX_IN[8003] NB2 NB1 CSA_VREF pixel
xPix8004 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[80] VREF PIX_IN[8004] NB2 NB1 CSA_VREF pixel
xPix8005 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[80] VREF PIX_IN[8005] NB2 NB1 CSA_VREF pixel
xPix8006 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[80] VREF PIX_IN[8006] NB2 NB1 CSA_VREF pixel
xPix8007 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[80] VREF PIX_IN[8007] NB2 NB1 CSA_VREF pixel
xPix8008 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[80] VREF PIX_IN[8008] NB2 NB1 CSA_VREF pixel
xPix8009 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[80] VREF PIX_IN[8009] NB2 NB1 CSA_VREF pixel
xPix8010 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[80] VREF PIX_IN[8010] NB2 NB1 CSA_VREF pixel
xPix8011 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[80] VREF PIX_IN[8011] NB2 NB1 CSA_VREF pixel
xPix8012 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[80] VREF PIX_IN[8012] NB2 NB1 CSA_VREF pixel
xPix8013 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[80] VREF PIX_IN[8013] NB2 NB1 CSA_VREF pixel
xPix8014 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[80] VREF PIX_IN[8014] NB2 NB1 CSA_VREF pixel
xPix8015 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[80] VREF PIX_IN[8015] NB2 NB1 CSA_VREF pixel
xPix8016 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[80] VREF PIX_IN[8016] NB2 NB1 CSA_VREF pixel
xPix8017 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[80] VREF PIX_IN[8017] NB2 NB1 CSA_VREF pixel
xPix8018 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[80] VREF PIX_IN[8018] NB2 NB1 CSA_VREF pixel
xPix8019 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[80] VREF PIX_IN[8019] NB2 NB1 CSA_VREF pixel
xPix8020 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[80] VREF PIX_IN[8020] NB2 NB1 CSA_VREF pixel
xPix8021 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[80] VREF PIX_IN[8021] NB2 NB1 CSA_VREF pixel
xPix8022 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[80] VREF PIX_IN[8022] NB2 NB1 CSA_VREF pixel
xPix8023 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[80] VREF PIX_IN[8023] NB2 NB1 CSA_VREF pixel
xPix8024 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[80] VREF PIX_IN[8024] NB2 NB1 CSA_VREF pixel
xPix8025 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[80] VREF PIX_IN[8025] NB2 NB1 CSA_VREF pixel
xPix8026 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[80] VREF PIX_IN[8026] NB2 NB1 CSA_VREF pixel
xPix8027 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[80] VREF PIX_IN[8027] NB2 NB1 CSA_VREF pixel
xPix8028 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[80] VREF PIX_IN[8028] NB2 NB1 CSA_VREF pixel
xPix8029 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[80] VREF PIX_IN[8029] NB2 NB1 CSA_VREF pixel
xPix8030 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[80] VREF PIX_IN[8030] NB2 NB1 CSA_VREF pixel
xPix8031 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[80] VREF PIX_IN[8031] NB2 NB1 CSA_VREF pixel
xPix8032 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[80] VREF PIX_IN[8032] NB2 NB1 CSA_VREF pixel
xPix8033 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[80] VREF PIX_IN[8033] NB2 NB1 CSA_VREF pixel
xPix8034 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[80] VREF PIX_IN[8034] NB2 NB1 CSA_VREF pixel
xPix8035 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[80] VREF PIX_IN[8035] NB2 NB1 CSA_VREF pixel
xPix8036 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[80] VREF PIX_IN[8036] NB2 NB1 CSA_VREF pixel
xPix8037 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[80] VREF PIX_IN[8037] NB2 NB1 CSA_VREF pixel
xPix8038 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[80] VREF PIX_IN[8038] NB2 NB1 CSA_VREF pixel
xPix8039 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[80] VREF PIX_IN[8039] NB2 NB1 CSA_VREF pixel
xPix8040 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[80] VREF PIX_IN[8040] NB2 NB1 CSA_VREF pixel
xPix8041 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[80] VREF PIX_IN[8041] NB2 NB1 CSA_VREF pixel
xPix8042 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[80] VREF PIX_IN[8042] NB2 NB1 CSA_VREF pixel
xPix8043 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[80] VREF PIX_IN[8043] NB2 NB1 CSA_VREF pixel
xPix8044 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[80] VREF PIX_IN[8044] NB2 NB1 CSA_VREF pixel
xPix8045 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[80] VREF PIX_IN[8045] NB2 NB1 CSA_VREF pixel
xPix8046 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[80] VREF PIX_IN[8046] NB2 NB1 CSA_VREF pixel
xPix8047 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[80] VREF PIX_IN[8047] NB2 NB1 CSA_VREF pixel
xPix8048 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[80] VREF PIX_IN[8048] NB2 NB1 CSA_VREF pixel
xPix8049 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[80] VREF PIX_IN[8049] NB2 NB1 CSA_VREF pixel
xPix8050 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[80] VREF PIX_IN[8050] NB2 NB1 CSA_VREF pixel
xPix8051 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[80] VREF PIX_IN[8051] NB2 NB1 CSA_VREF pixel
xPix8052 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[80] VREF PIX_IN[8052] NB2 NB1 CSA_VREF pixel
xPix8053 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[80] VREF PIX_IN[8053] NB2 NB1 CSA_VREF pixel
xPix8054 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[80] VREF PIX_IN[8054] NB2 NB1 CSA_VREF pixel
xPix8055 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[80] VREF PIX_IN[8055] NB2 NB1 CSA_VREF pixel
xPix8056 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[80] VREF PIX_IN[8056] NB2 NB1 CSA_VREF pixel
xPix8057 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[80] VREF PIX_IN[8057] NB2 NB1 CSA_VREF pixel
xPix8058 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[80] VREF PIX_IN[8058] NB2 NB1 CSA_VREF pixel
xPix8059 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[80] VREF PIX_IN[8059] NB2 NB1 CSA_VREF pixel
xPix8060 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[80] VREF PIX_IN[8060] NB2 NB1 CSA_VREF pixel
xPix8061 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[80] VREF PIX_IN[8061] NB2 NB1 CSA_VREF pixel
xPix8062 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[80] VREF PIX_IN[8062] NB2 NB1 CSA_VREF pixel
xPix8063 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[80] VREF PIX_IN[8063] NB2 NB1 CSA_VREF pixel
xPix8064 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[80] VREF PIX_IN[8064] NB2 NB1 CSA_VREF pixel
xPix8065 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[80] VREF PIX_IN[8065] NB2 NB1 CSA_VREF pixel
xPix8066 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[80] VREF PIX_IN[8066] NB2 NB1 CSA_VREF pixel
xPix8067 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[80] VREF PIX_IN[8067] NB2 NB1 CSA_VREF pixel
xPix8068 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[80] VREF PIX_IN[8068] NB2 NB1 CSA_VREF pixel
xPix8069 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[80] VREF PIX_IN[8069] NB2 NB1 CSA_VREF pixel
xPix8070 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[80] VREF PIX_IN[8070] NB2 NB1 CSA_VREF pixel
xPix8071 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[80] VREF PIX_IN[8071] NB2 NB1 CSA_VREF pixel
xPix8072 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[80] VREF PIX_IN[8072] NB2 NB1 CSA_VREF pixel
xPix8073 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[80] VREF PIX_IN[8073] NB2 NB1 CSA_VREF pixel
xPix8074 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[80] VREF PIX_IN[8074] NB2 NB1 CSA_VREF pixel
xPix8075 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[80] VREF PIX_IN[8075] NB2 NB1 CSA_VREF pixel
xPix8076 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[80] VREF PIX_IN[8076] NB2 NB1 CSA_VREF pixel
xPix8077 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[80] VREF PIX_IN[8077] NB2 NB1 CSA_VREF pixel
xPix8078 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[80] VREF PIX_IN[8078] NB2 NB1 CSA_VREF pixel
xPix8079 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[80] VREF PIX_IN[8079] NB2 NB1 CSA_VREF pixel
xPix8080 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[80] VREF PIX_IN[8080] NB2 NB1 CSA_VREF pixel
xPix8081 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[80] VREF PIX_IN[8081] NB2 NB1 CSA_VREF pixel
xPix8082 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[80] VREF PIX_IN[8082] NB2 NB1 CSA_VREF pixel
xPix8083 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[80] VREF PIX_IN[8083] NB2 NB1 CSA_VREF pixel
xPix8084 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[80] VREF PIX_IN[8084] NB2 NB1 CSA_VREF pixel
xPix8085 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[80] VREF PIX_IN[8085] NB2 NB1 CSA_VREF pixel
xPix8086 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[80] VREF PIX_IN[8086] NB2 NB1 CSA_VREF pixel
xPix8087 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[80] VREF PIX_IN[8087] NB2 NB1 CSA_VREF pixel
xPix8088 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[80] VREF PIX_IN[8088] NB2 NB1 CSA_VREF pixel
xPix8089 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[80] VREF PIX_IN[8089] NB2 NB1 CSA_VREF pixel
xPix8090 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[80] VREF PIX_IN[8090] NB2 NB1 CSA_VREF pixel
xPix8091 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[80] VREF PIX_IN[8091] NB2 NB1 CSA_VREF pixel
xPix8092 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[80] VREF PIX_IN[8092] NB2 NB1 CSA_VREF pixel
xPix8093 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[80] VREF PIX_IN[8093] NB2 NB1 CSA_VREF pixel
xPix8094 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[80] VREF PIX_IN[8094] NB2 NB1 CSA_VREF pixel
xPix8095 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[80] VREF PIX_IN[8095] NB2 NB1 CSA_VREF pixel
xPix8096 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[80] VREF PIX_IN[8096] NB2 NB1 CSA_VREF pixel
xPix8097 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[80] VREF PIX_IN[8097] NB2 NB1 CSA_VREF pixel
xPix8098 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[80] VREF PIX_IN[8098] NB2 NB1 CSA_VREF pixel
xPix8099 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[80] VREF PIX_IN[8099] NB2 NB1 CSA_VREF pixel
xPix8100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[81] VREF PIX_IN[8100] NB2 NB1 CSA_VREF pixel
xPix8101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[81] VREF PIX_IN[8101] NB2 NB1 CSA_VREF pixel
xPix8102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[81] VREF PIX_IN[8102] NB2 NB1 CSA_VREF pixel
xPix8103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[81] VREF PIX_IN[8103] NB2 NB1 CSA_VREF pixel
xPix8104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[81] VREF PIX_IN[8104] NB2 NB1 CSA_VREF pixel
xPix8105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[81] VREF PIX_IN[8105] NB2 NB1 CSA_VREF pixel
xPix8106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[81] VREF PIX_IN[8106] NB2 NB1 CSA_VREF pixel
xPix8107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[81] VREF PIX_IN[8107] NB2 NB1 CSA_VREF pixel
xPix8108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[81] VREF PIX_IN[8108] NB2 NB1 CSA_VREF pixel
xPix8109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[81] VREF PIX_IN[8109] NB2 NB1 CSA_VREF pixel
xPix8110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[81] VREF PIX_IN[8110] NB2 NB1 CSA_VREF pixel
xPix8111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[81] VREF PIX_IN[8111] NB2 NB1 CSA_VREF pixel
xPix8112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[81] VREF PIX_IN[8112] NB2 NB1 CSA_VREF pixel
xPix8113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[81] VREF PIX_IN[8113] NB2 NB1 CSA_VREF pixel
xPix8114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[81] VREF PIX_IN[8114] NB2 NB1 CSA_VREF pixel
xPix8115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[81] VREF PIX_IN[8115] NB2 NB1 CSA_VREF pixel
xPix8116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[81] VREF PIX_IN[8116] NB2 NB1 CSA_VREF pixel
xPix8117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[81] VREF PIX_IN[8117] NB2 NB1 CSA_VREF pixel
xPix8118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[81] VREF PIX_IN[8118] NB2 NB1 CSA_VREF pixel
xPix8119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[81] VREF PIX_IN[8119] NB2 NB1 CSA_VREF pixel
xPix8120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[81] VREF PIX_IN[8120] NB2 NB1 CSA_VREF pixel
xPix8121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[81] VREF PIX_IN[8121] NB2 NB1 CSA_VREF pixel
xPix8122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[81] VREF PIX_IN[8122] NB2 NB1 CSA_VREF pixel
xPix8123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[81] VREF PIX_IN[8123] NB2 NB1 CSA_VREF pixel
xPix8124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[81] VREF PIX_IN[8124] NB2 NB1 CSA_VREF pixel
xPix8125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[81] VREF PIX_IN[8125] NB2 NB1 CSA_VREF pixel
xPix8126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[81] VREF PIX_IN[8126] NB2 NB1 CSA_VREF pixel
xPix8127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[81] VREF PIX_IN[8127] NB2 NB1 CSA_VREF pixel
xPix8128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[81] VREF PIX_IN[8128] NB2 NB1 CSA_VREF pixel
xPix8129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[81] VREF PIX_IN[8129] NB2 NB1 CSA_VREF pixel
xPix8130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[81] VREF PIX_IN[8130] NB2 NB1 CSA_VREF pixel
xPix8131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[81] VREF PIX_IN[8131] NB2 NB1 CSA_VREF pixel
xPix8132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[81] VREF PIX_IN[8132] NB2 NB1 CSA_VREF pixel
xPix8133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[81] VREF PIX_IN[8133] NB2 NB1 CSA_VREF pixel
xPix8134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[81] VREF PIX_IN[8134] NB2 NB1 CSA_VREF pixel
xPix8135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[81] VREF PIX_IN[8135] NB2 NB1 CSA_VREF pixel
xPix8136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[81] VREF PIX_IN[8136] NB2 NB1 CSA_VREF pixel
xPix8137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[81] VREF PIX_IN[8137] NB2 NB1 CSA_VREF pixel
xPix8138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[81] VREF PIX_IN[8138] NB2 NB1 CSA_VREF pixel
xPix8139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[81] VREF PIX_IN[8139] NB2 NB1 CSA_VREF pixel
xPix8140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[81] VREF PIX_IN[8140] NB2 NB1 CSA_VREF pixel
xPix8141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[81] VREF PIX_IN[8141] NB2 NB1 CSA_VREF pixel
xPix8142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[81] VREF PIX_IN[8142] NB2 NB1 CSA_VREF pixel
xPix8143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[81] VREF PIX_IN[8143] NB2 NB1 CSA_VREF pixel
xPix8144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[81] VREF PIX_IN[8144] NB2 NB1 CSA_VREF pixel
xPix8145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[81] VREF PIX_IN[8145] NB2 NB1 CSA_VREF pixel
xPix8146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[81] VREF PIX_IN[8146] NB2 NB1 CSA_VREF pixel
xPix8147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[81] VREF PIX_IN[8147] NB2 NB1 CSA_VREF pixel
xPix8148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[81] VREF PIX_IN[8148] NB2 NB1 CSA_VREF pixel
xPix8149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[81] VREF PIX_IN[8149] NB2 NB1 CSA_VREF pixel
xPix8150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[81] VREF PIX_IN[8150] NB2 NB1 CSA_VREF pixel
xPix8151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[81] VREF PIX_IN[8151] NB2 NB1 CSA_VREF pixel
xPix8152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[81] VREF PIX_IN[8152] NB2 NB1 CSA_VREF pixel
xPix8153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[81] VREF PIX_IN[8153] NB2 NB1 CSA_VREF pixel
xPix8154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[81] VREF PIX_IN[8154] NB2 NB1 CSA_VREF pixel
xPix8155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[81] VREF PIX_IN[8155] NB2 NB1 CSA_VREF pixel
xPix8156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[81] VREF PIX_IN[8156] NB2 NB1 CSA_VREF pixel
xPix8157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[81] VREF PIX_IN[8157] NB2 NB1 CSA_VREF pixel
xPix8158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[81] VREF PIX_IN[8158] NB2 NB1 CSA_VREF pixel
xPix8159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[81] VREF PIX_IN[8159] NB2 NB1 CSA_VREF pixel
xPix8160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[81] VREF PIX_IN[8160] NB2 NB1 CSA_VREF pixel
xPix8161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[81] VREF PIX_IN[8161] NB2 NB1 CSA_VREF pixel
xPix8162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[81] VREF PIX_IN[8162] NB2 NB1 CSA_VREF pixel
xPix8163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[81] VREF PIX_IN[8163] NB2 NB1 CSA_VREF pixel
xPix8164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[81] VREF PIX_IN[8164] NB2 NB1 CSA_VREF pixel
xPix8165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[81] VREF PIX_IN[8165] NB2 NB1 CSA_VREF pixel
xPix8166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[81] VREF PIX_IN[8166] NB2 NB1 CSA_VREF pixel
xPix8167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[81] VREF PIX_IN[8167] NB2 NB1 CSA_VREF pixel
xPix8168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[81] VREF PIX_IN[8168] NB2 NB1 CSA_VREF pixel
xPix8169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[81] VREF PIX_IN[8169] NB2 NB1 CSA_VREF pixel
xPix8170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[81] VREF PIX_IN[8170] NB2 NB1 CSA_VREF pixel
xPix8171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[81] VREF PIX_IN[8171] NB2 NB1 CSA_VREF pixel
xPix8172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[81] VREF PIX_IN[8172] NB2 NB1 CSA_VREF pixel
xPix8173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[81] VREF PIX_IN[8173] NB2 NB1 CSA_VREF pixel
xPix8174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[81] VREF PIX_IN[8174] NB2 NB1 CSA_VREF pixel
xPix8175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[81] VREF PIX_IN[8175] NB2 NB1 CSA_VREF pixel
xPix8176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[81] VREF PIX_IN[8176] NB2 NB1 CSA_VREF pixel
xPix8177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[81] VREF PIX_IN[8177] NB2 NB1 CSA_VREF pixel
xPix8178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[81] VREF PIX_IN[8178] NB2 NB1 CSA_VREF pixel
xPix8179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[81] VREF PIX_IN[8179] NB2 NB1 CSA_VREF pixel
xPix8180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[81] VREF PIX_IN[8180] NB2 NB1 CSA_VREF pixel
xPix8181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[81] VREF PIX_IN[8181] NB2 NB1 CSA_VREF pixel
xPix8182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[81] VREF PIX_IN[8182] NB2 NB1 CSA_VREF pixel
xPix8183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[81] VREF PIX_IN[8183] NB2 NB1 CSA_VREF pixel
xPix8184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[81] VREF PIX_IN[8184] NB2 NB1 CSA_VREF pixel
xPix8185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[81] VREF PIX_IN[8185] NB2 NB1 CSA_VREF pixel
xPix8186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[81] VREF PIX_IN[8186] NB2 NB1 CSA_VREF pixel
xPix8187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[81] VREF PIX_IN[8187] NB2 NB1 CSA_VREF pixel
xPix8188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[81] VREF PIX_IN[8188] NB2 NB1 CSA_VREF pixel
xPix8189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[81] VREF PIX_IN[8189] NB2 NB1 CSA_VREF pixel
xPix8190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[81] VREF PIX_IN[8190] NB2 NB1 CSA_VREF pixel
xPix8191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[81] VREF PIX_IN[8191] NB2 NB1 CSA_VREF pixel
xPix8192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[81] VREF PIX_IN[8192] NB2 NB1 CSA_VREF pixel
xPix8193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[81] VREF PIX_IN[8193] NB2 NB1 CSA_VREF pixel
xPix8194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[81] VREF PIX_IN[8194] NB2 NB1 CSA_VREF pixel
xPix8195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[81] VREF PIX_IN[8195] NB2 NB1 CSA_VREF pixel
xPix8196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[81] VREF PIX_IN[8196] NB2 NB1 CSA_VREF pixel
xPix8197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[81] VREF PIX_IN[8197] NB2 NB1 CSA_VREF pixel
xPix8198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[81] VREF PIX_IN[8198] NB2 NB1 CSA_VREF pixel
xPix8199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[81] VREF PIX_IN[8199] NB2 NB1 CSA_VREF pixel
xPix8200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[82] VREF PIX_IN[8200] NB2 NB1 CSA_VREF pixel
xPix8201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[82] VREF PIX_IN[8201] NB2 NB1 CSA_VREF pixel
xPix8202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[82] VREF PIX_IN[8202] NB2 NB1 CSA_VREF pixel
xPix8203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[82] VREF PIX_IN[8203] NB2 NB1 CSA_VREF pixel
xPix8204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[82] VREF PIX_IN[8204] NB2 NB1 CSA_VREF pixel
xPix8205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[82] VREF PIX_IN[8205] NB2 NB1 CSA_VREF pixel
xPix8206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[82] VREF PIX_IN[8206] NB2 NB1 CSA_VREF pixel
xPix8207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[82] VREF PIX_IN[8207] NB2 NB1 CSA_VREF pixel
xPix8208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[82] VREF PIX_IN[8208] NB2 NB1 CSA_VREF pixel
xPix8209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[82] VREF PIX_IN[8209] NB2 NB1 CSA_VREF pixel
xPix8210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[82] VREF PIX_IN[8210] NB2 NB1 CSA_VREF pixel
xPix8211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[82] VREF PIX_IN[8211] NB2 NB1 CSA_VREF pixel
xPix8212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[82] VREF PIX_IN[8212] NB2 NB1 CSA_VREF pixel
xPix8213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[82] VREF PIX_IN[8213] NB2 NB1 CSA_VREF pixel
xPix8214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[82] VREF PIX_IN[8214] NB2 NB1 CSA_VREF pixel
xPix8215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[82] VREF PIX_IN[8215] NB2 NB1 CSA_VREF pixel
xPix8216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[82] VREF PIX_IN[8216] NB2 NB1 CSA_VREF pixel
xPix8217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[82] VREF PIX_IN[8217] NB2 NB1 CSA_VREF pixel
xPix8218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[82] VREF PIX_IN[8218] NB2 NB1 CSA_VREF pixel
xPix8219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[82] VREF PIX_IN[8219] NB2 NB1 CSA_VREF pixel
xPix8220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[82] VREF PIX_IN[8220] NB2 NB1 CSA_VREF pixel
xPix8221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[82] VREF PIX_IN[8221] NB2 NB1 CSA_VREF pixel
xPix8222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[82] VREF PIX_IN[8222] NB2 NB1 CSA_VREF pixel
xPix8223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[82] VREF PIX_IN[8223] NB2 NB1 CSA_VREF pixel
xPix8224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[82] VREF PIX_IN[8224] NB2 NB1 CSA_VREF pixel
xPix8225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[82] VREF PIX_IN[8225] NB2 NB1 CSA_VREF pixel
xPix8226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[82] VREF PIX_IN[8226] NB2 NB1 CSA_VREF pixel
xPix8227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[82] VREF PIX_IN[8227] NB2 NB1 CSA_VREF pixel
xPix8228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[82] VREF PIX_IN[8228] NB2 NB1 CSA_VREF pixel
xPix8229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[82] VREF PIX_IN[8229] NB2 NB1 CSA_VREF pixel
xPix8230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[82] VREF PIX_IN[8230] NB2 NB1 CSA_VREF pixel
xPix8231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[82] VREF PIX_IN[8231] NB2 NB1 CSA_VREF pixel
xPix8232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[82] VREF PIX_IN[8232] NB2 NB1 CSA_VREF pixel
xPix8233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[82] VREF PIX_IN[8233] NB2 NB1 CSA_VREF pixel
xPix8234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[82] VREF PIX_IN[8234] NB2 NB1 CSA_VREF pixel
xPix8235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[82] VREF PIX_IN[8235] NB2 NB1 CSA_VREF pixel
xPix8236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[82] VREF PIX_IN[8236] NB2 NB1 CSA_VREF pixel
xPix8237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[82] VREF PIX_IN[8237] NB2 NB1 CSA_VREF pixel
xPix8238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[82] VREF PIX_IN[8238] NB2 NB1 CSA_VREF pixel
xPix8239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[82] VREF PIX_IN[8239] NB2 NB1 CSA_VREF pixel
xPix8240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[82] VREF PIX_IN[8240] NB2 NB1 CSA_VREF pixel
xPix8241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[82] VREF PIX_IN[8241] NB2 NB1 CSA_VREF pixel
xPix8242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[82] VREF PIX_IN[8242] NB2 NB1 CSA_VREF pixel
xPix8243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[82] VREF PIX_IN[8243] NB2 NB1 CSA_VREF pixel
xPix8244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[82] VREF PIX_IN[8244] NB2 NB1 CSA_VREF pixel
xPix8245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[82] VREF PIX_IN[8245] NB2 NB1 CSA_VREF pixel
xPix8246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[82] VREF PIX_IN[8246] NB2 NB1 CSA_VREF pixel
xPix8247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[82] VREF PIX_IN[8247] NB2 NB1 CSA_VREF pixel
xPix8248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[82] VREF PIX_IN[8248] NB2 NB1 CSA_VREF pixel
xPix8249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[82] VREF PIX_IN[8249] NB2 NB1 CSA_VREF pixel
xPix8250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[82] VREF PIX_IN[8250] NB2 NB1 CSA_VREF pixel
xPix8251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[82] VREF PIX_IN[8251] NB2 NB1 CSA_VREF pixel
xPix8252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[82] VREF PIX_IN[8252] NB2 NB1 CSA_VREF pixel
xPix8253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[82] VREF PIX_IN[8253] NB2 NB1 CSA_VREF pixel
xPix8254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[82] VREF PIX_IN[8254] NB2 NB1 CSA_VREF pixel
xPix8255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[82] VREF PIX_IN[8255] NB2 NB1 CSA_VREF pixel
xPix8256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[82] VREF PIX_IN[8256] NB2 NB1 CSA_VREF pixel
xPix8257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[82] VREF PIX_IN[8257] NB2 NB1 CSA_VREF pixel
xPix8258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[82] VREF PIX_IN[8258] NB2 NB1 CSA_VREF pixel
xPix8259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[82] VREF PIX_IN[8259] NB2 NB1 CSA_VREF pixel
xPix8260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[82] VREF PIX_IN[8260] NB2 NB1 CSA_VREF pixel
xPix8261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[82] VREF PIX_IN[8261] NB2 NB1 CSA_VREF pixel
xPix8262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[82] VREF PIX_IN[8262] NB2 NB1 CSA_VREF pixel
xPix8263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[82] VREF PIX_IN[8263] NB2 NB1 CSA_VREF pixel
xPix8264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[82] VREF PIX_IN[8264] NB2 NB1 CSA_VREF pixel
xPix8265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[82] VREF PIX_IN[8265] NB2 NB1 CSA_VREF pixel
xPix8266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[82] VREF PIX_IN[8266] NB2 NB1 CSA_VREF pixel
xPix8267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[82] VREF PIX_IN[8267] NB2 NB1 CSA_VREF pixel
xPix8268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[82] VREF PIX_IN[8268] NB2 NB1 CSA_VREF pixel
xPix8269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[82] VREF PIX_IN[8269] NB2 NB1 CSA_VREF pixel
xPix8270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[82] VREF PIX_IN[8270] NB2 NB1 CSA_VREF pixel
xPix8271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[82] VREF PIX_IN[8271] NB2 NB1 CSA_VREF pixel
xPix8272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[82] VREF PIX_IN[8272] NB2 NB1 CSA_VREF pixel
xPix8273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[82] VREF PIX_IN[8273] NB2 NB1 CSA_VREF pixel
xPix8274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[82] VREF PIX_IN[8274] NB2 NB1 CSA_VREF pixel
xPix8275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[82] VREF PIX_IN[8275] NB2 NB1 CSA_VREF pixel
xPix8276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[82] VREF PIX_IN[8276] NB2 NB1 CSA_VREF pixel
xPix8277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[82] VREF PIX_IN[8277] NB2 NB1 CSA_VREF pixel
xPix8278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[82] VREF PIX_IN[8278] NB2 NB1 CSA_VREF pixel
xPix8279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[82] VREF PIX_IN[8279] NB2 NB1 CSA_VREF pixel
xPix8280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[82] VREF PIX_IN[8280] NB2 NB1 CSA_VREF pixel
xPix8281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[82] VREF PIX_IN[8281] NB2 NB1 CSA_VREF pixel
xPix8282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[82] VREF PIX_IN[8282] NB2 NB1 CSA_VREF pixel
xPix8283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[82] VREF PIX_IN[8283] NB2 NB1 CSA_VREF pixel
xPix8284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[82] VREF PIX_IN[8284] NB2 NB1 CSA_VREF pixel
xPix8285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[82] VREF PIX_IN[8285] NB2 NB1 CSA_VREF pixel
xPix8286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[82] VREF PIX_IN[8286] NB2 NB1 CSA_VREF pixel
xPix8287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[82] VREF PIX_IN[8287] NB2 NB1 CSA_VREF pixel
xPix8288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[82] VREF PIX_IN[8288] NB2 NB1 CSA_VREF pixel
xPix8289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[82] VREF PIX_IN[8289] NB2 NB1 CSA_VREF pixel
xPix8290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[82] VREF PIX_IN[8290] NB2 NB1 CSA_VREF pixel
xPix8291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[82] VREF PIX_IN[8291] NB2 NB1 CSA_VREF pixel
xPix8292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[82] VREF PIX_IN[8292] NB2 NB1 CSA_VREF pixel
xPix8293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[82] VREF PIX_IN[8293] NB2 NB1 CSA_VREF pixel
xPix8294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[82] VREF PIX_IN[8294] NB2 NB1 CSA_VREF pixel
xPix8295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[82] VREF PIX_IN[8295] NB2 NB1 CSA_VREF pixel
xPix8296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[82] VREF PIX_IN[8296] NB2 NB1 CSA_VREF pixel
xPix8297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[82] VREF PIX_IN[8297] NB2 NB1 CSA_VREF pixel
xPix8298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[82] VREF PIX_IN[8298] NB2 NB1 CSA_VREF pixel
xPix8299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[82] VREF PIX_IN[8299] NB2 NB1 CSA_VREF pixel
xPix8300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[83] VREF PIX_IN[8300] NB2 NB1 CSA_VREF pixel
xPix8301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[83] VREF PIX_IN[8301] NB2 NB1 CSA_VREF pixel
xPix8302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[83] VREF PIX_IN[8302] NB2 NB1 CSA_VREF pixel
xPix8303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[83] VREF PIX_IN[8303] NB2 NB1 CSA_VREF pixel
xPix8304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[83] VREF PIX_IN[8304] NB2 NB1 CSA_VREF pixel
xPix8305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[83] VREF PIX_IN[8305] NB2 NB1 CSA_VREF pixel
xPix8306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[83] VREF PIX_IN[8306] NB2 NB1 CSA_VREF pixel
xPix8307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[83] VREF PIX_IN[8307] NB2 NB1 CSA_VREF pixel
xPix8308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[83] VREF PIX_IN[8308] NB2 NB1 CSA_VREF pixel
xPix8309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[83] VREF PIX_IN[8309] NB2 NB1 CSA_VREF pixel
xPix8310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[83] VREF PIX_IN[8310] NB2 NB1 CSA_VREF pixel
xPix8311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[83] VREF PIX_IN[8311] NB2 NB1 CSA_VREF pixel
xPix8312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[83] VREF PIX_IN[8312] NB2 NB1 CSA_VREF pixel
xPix8313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[83] VREF PIX_IN[8313] NB2 NB1 CSA_VREF pixel
xPix8314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[83] VREF PIX_IN[8314] NB2 NB1 CSA_VREF pixel
xPix8315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[83] VREF PIX_IN[8315] NB2 NB1 CSA_VREF pixel
xPix8316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[83] VREF PIX_IN[8316] NB2 NB1 CSA_VREF pixel
xPix8317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[83] VREF PIX_IN[8317] NB2 NB1 CSA_VREF pixel
xPix8318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[83] VREF PIX_IN[8318] NB2 NB1 CSA_VREF pixel
xPix8319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[83] VREF PIX_IN[8319] NB2 NB1 CSA_VREF pixel
xPix8320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[83] VREF PIX_IN[8320] NB2 NB1 CSA_VREF pixel
xPix8321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[83] VREF PIX_IN[8321] NB2 NB1 CSA_VREF pixel
xPix8322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[83] VREF PIX_IN[8322] NB2 NB1 CSA_VREF pixel
xPix8323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[83] VREF PIX_IN[8323] NB2 NB1 CSA_VREF pixel
xPix8324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[83] VREF PIX_IN[8324] NB2 NB1 CSA_VREF pixel
xPix8325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[83] VREF PIX_IN[8325] NB2 NB1 CSA_VREF pixel
xPix8326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[83] VREF PIX_IN[8326] NB2 NB1 CSA_VREF pixel
xPix8327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[83] VREF PIX_IN[8327] NB2 NB1 CSA_VREF pixel
xPix8328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[83] VREF PIX_IN[8328] NB2 NB1 CSA_VREF pixel
xPix8329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[83] VREF PIX_IN[8329] NB2 NB1 CSA_VREF pixel
xPix8330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[83] VREF PIX_IN[8330] NB2 NB1 CSA_VREF pixel
xPix8331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[83] VREF PIX_IN[8331] NB2 NB1 CSA_VREF pixel
xPix8332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[83] VREF PIX_IN[8332] NB2 NB1 CSA_VREF pixel
xPix8333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[83] VREF PIX_IN[8333] NB2 NB1 CSA_VREF pixel
xPix8334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[83] VREF PIX_IN[8334] NB2 NB1 CSA_VREF pixel
xPix8335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[83] VREF PIX_IN[8335] NB2 NB1 CSA_VREF pixel
xPix8336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[83] VREF PIX_IN[8336] NB2 NB1 CSA_VREF pixel
xPix8337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[83] VREF PIX_IN[8337] NB2 NB1 CSA_VREF pixel
xPix8338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[83] VREF PIX_IN[8338] NB2 NB1 CSA_VREF pixel
xPix8339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[83] VREF PIX_IN[8339] NB2 NB1 CSA_VREF pixel
xPix8340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[83] VREF PIX_IN[8340] NB2 NB1 CSA_VREF pixel
xPix8341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[83] VREF PIX_IN[8341] NB2 NB1 CSA_VREF pixel
xPix8342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[83] VREF PIX_IN[8342] NB2 NB1 CSA_VREF pixel
xPix8343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[83] VREF PIX_IN[8343] NB2 NB1 CSA_VREF pixel
xPix8344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[83] VREF PIX_IN[8344] NB2 NB1 CSA_VREF pixel
xPix8345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[83] VREF PIX_IN[8345] NB2 NB1 CSA_VREF pixel
xPix8346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[83] VREF PIX_IN[8346] NB2 NB1 CSA_VREF pixel
xPix8347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[83] VREF PIX_IN[8347] NB2 NB1 CSA_VREF pixel
xPix8348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[83] VREF PIX_IN[8348] NB2 NB1 CSA_VREF pixel
xPix8349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[83] VREF PIX_IN[8349] NB2 NB1 CSA_VREF pixel
xPix8350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[83] VREF PIX_IN[8350] NB2 NB1 CSA_VREF pixel
xPix8351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[83] VREF PIX_IN[8351] NB2 NB1 CSA_VREF pixel
xPix8352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[83] VREF PIX_IN[8352] NB2 NB1 CSA_VREF pixel
xPix8353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[83] VREF PIX_IN[8353] NB2 NB1 CSA_VREF pixel
xPix8354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[83] VREF PIX_IN[8354] NB2 NB1 CSA_VREF pixel
xPix8355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[83] VREF PIX_IN[8355] NB2 NB1 CSA_VREF pixel
xPix8356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[83] VREF PIX_IN[8356] NB2 NB1 CSA_VREF pixel
xPix8357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[83] VREF PIX_IN[8357] NB2 NB1 CSA_VREF pixel
xPix8358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[83] VREF PIX_IN[8358] NB2 NB1 CSA_VREF pixel
xPix8359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[83] VREF PIX_IN[8359] NB2 NB1 CSA_VREF pixel
xPix8360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[83] VREF PIX_IN[8360] NB2 NB1 CSA_VREF pixel
xPix8361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[83] VREF PIX_IN[8361] NB2 NB1 CSA_VREF pixel
xPix8362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[83] VREF PIX_IN[8362] NB2 NB1 CSA_VREF pixel
xPix8363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[83] VREF PIX_IN[8363] NB2 NB1 CSA_VREF pixel
xPix8364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[83] VREF PIX_IN[8364] NB2 NB1 CSA_VREF pixel
xPix8365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[83] VREF PIX_IN[8365] NB2 NB1 CSA_VREF pixel
xPix8366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[83] VREF PIX_IN[8366] NB2 NB1 CSA_VREF pixel
xPix8367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[83] VREF PIX_IN[8367] NB2 NB1 CSA_VREF pixel
xPix8368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[83] VREF PIX_IN[8368] NB2 NB1 CSA_VREF pixel
xPix8369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[83] VREF PIX_IN[8369] NB2 NB1 CSA_VREF pixel
xPix8370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[83] VREF PIX_IN[8370] NB2 NB1 CSA_VREF pixel
xPix8371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[83] VREF PIX_IN[8371] NB2 NB1 CSA_VREF pixel
xPix8372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[83] VREF PIX_IN[8372] NB2 NB1 CSA_VREF pixel
xPix8373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[83] VREF PIX_IN[8373] NB2 NB1 CSA_VREF pixel
xPix8374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[83] VREF PIX_IN[8374] NB2 NB1 CSA_VREF pixel
xPix8375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[83] VREF PIX_IN[8375] NB2 NB1 CSA_VREF pixel
xPix8376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[83] VREF PIX_IN[8376] NB2 NB1 CSA_VREF pixel
xPix8377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[83] VREF PIX_IN[8377] NB2 NB1 CSA_VREF pixel
xPix8378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[83] VREF PIX_IN[8378] NB2 NB1 CSA_VREF pixel
xPix8379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[83] VREF PIX_IN[8379] NB2 NB1 CSA_VREF pixel
xPix8380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[83] VREF PIX_IN[8380] NB2 NB1 CSA_VREF pixel
xPix8381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[83] VREF PIX_IN[8381] NB2 NB1 CSA_VREF pixel
xPix8382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[83] VREF PIX_IN[8382] NB2 NB1 CSA_VREF pixel
xPix8383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[83] VREF PIX_IN[8383] NB2 NB1 CSA_VREF pixel
xPix8384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[83] VREF PIX_IN[8384] NB2 NB1 CSA_VREF pixel
xPix8385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[83] VREF PIX_IN[8385] NB2 NB1 CSA_VREF pixel
xPix8386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[83] VREF PIX_IN[8386] NB2 NB1 CSA_VREF pixel
xPix8387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[83] VREF PIX_IN[8387] NB2 NB1 CSA_VREF pixel
xPix8388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[83] VREF PIX_IN[8388] NB2 NB1 CSA_VREF pixel
xPix8389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[83] VREF PIX_IN[8389] NB2 NB1 CSA_VREF pixel
xPix8390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[83] VREF PIX_IN[8390] NB2 NB1 CSA_VREF pixel
xPix8391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[83] VREF PIX_IN[8391] NB2 NB1 CSA_VREF pixel
xPix8392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[83] VREF PIX_IN[8392] NB2 NB1 CSA_VREF pixel
xPix8393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[83] VREF PIX_IN[8393] NB2 NB1 CSA_VREF pixel
xPix8394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[83] VREF PIX_IN[8394] NB2 NB1 CSA_VREF pixel
xPix8395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[83] VREF PIX_IN[8395] NB2 NB1 CSA_VREF pixel
xPix8396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[83] VREF PIX_IN[8396] NB2 NB1 CSA_VREF pixel
xPix8397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[83] VREF PIX_IN[8397] NB2 NB1 CSA_VREF pixel
xPix8398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[83] VREF PIX_IN[8398] NB2 NB1 CSA_VREF pixel
xPix8399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[83] VREF PIX_IN[8399] NB2 NB1 CSA_VREF pixel
xPix8400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[84] VREF PIX_IN[8400] NB2 NB1 CSA_VREF pixel
xPix8401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[84] VREF PIX_IN[8401] NB2 NB1 CSA_VREF pixel
xPix8402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[84] VREF PIX_IN[8402] NB2 NB1 CSA_VREF pixel
xPix8403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[84] VREF PIX_IN[8403] NB2 NB1 CSA_VREF pixel
xPix8404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[84] VREF PIX_IN[8404] NB2 NB1 CSA_VREF pixel
xPix8405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[84] VREF PIX_IN[8405] NB2 NB1 CSA_VREF pixel
xPix8406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[84] VREF PIX_IN[8406] NB2 NB1 CSA_VREF pixel
xPix8407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[84] VREF PIX_IN[8407] NB2 NB1 CSA_VREF pixel
xPix8408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[84] VREF PIX_IN[8408] NB2 NB1 CSA_VREF pixel
xPix8409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[84] VREF PIX_IN[8409] NB2 NB1 CSA_VREF pixel
xPix8410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[84] VREF PIX_IN[8410] NB2 NB1 CSA_VREF pixel
xPix8411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[84] VREF PIX_IN[8411] NB2 NB1 CSA_VREF pixel
xPix8412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[84] VREF PIX_IN[8412] NB2 NB1 CSA_VREF pixel
xPix8413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[84] VREF PIX_IN[8413] NB2 NB1 CSA_VREF pixel
xPix8414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[84] VREF PIX_IN[8414] NB2 NB1 CSA_VREF pixel
xPix8415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[84] VREF PIX_IN[8415] NB2 NB1 CSA_VREF pixel
xPix8416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[84] VREF PIX_IN[8416] NB2 NB1 CSA_VREF pixel
xPix8417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[84] VREF PIX_IN[8417] NB2 NB1 CSA_VREF pixel
xPix8418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[84] VREF PIX_IN[8418] NB2 NB1 CSA_VREF pixel
xPix8419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[84] VREF PIX_IN[8419] NB2 NB1 CSA_VREF pixel
xPix8420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[84] VREF PIX_IN[8420] NB2 NB1 CSA_VREF pixel
xPix8421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[84] VREF PIX_IN[8421] NB2 NB1 CSA_VREF pixel
xPix8422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[84] VREF PIX_IN[8422] NB2 NB1 CSA_VREF pixel
xPix8423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[84] VREF PIX_IN[8423] NB2 NB1 CSA_VREF pixel
xPix8424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[84] VREF PIX_IN[8424] NB2 NB1 CSA_VREF pixel
xPix8425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[84] VREF PIX_IN[8425] NB2 NB1 CSA_VREF pixel
xPix8426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[84] VREF PIX_IN[8426] NB2 NB1 CSA_VREF pixel
xPix8427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[84] VREF PIX_IN[8427] NB2 NB1 CSA_VREF pixel
xPix8428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[84] VREF PIX_IN[8428] NB2 NB1 CSA_VREF pixel
xPix8429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[84] VREF PIX_IN[8429] NB2 NB1 CSA_VREF pixel
xPix8430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[84] VREF PIX_IN[8430] NB2 NB1 CSA_VREF pixel
xPix8431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[84] VREF PIX_IN[8431] NB2 NB1 CSA_VREF pixel
xPix8432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[84] VREF PIX_IN[8432] NB2 NB1 CSA_VREF pixel
xPix8433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[84] VREF PIX_IN[8433] NB2 NB1 CSA_VREF pixel
xPix8434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[84] VREF PIX_IN[8434] NB2 NB1 CSA_VREF pixel
xPix8435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[84] VREF PIX_IN[8435] NB2 NB1 CSA_VREF pixel
xPix8436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[84] VREF PIX_IN[8436] NB2 NB1 CSA_VREF pixel
xPix8437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[84] VREF PIX_IN[8437] NB2 NB1 CSA_VREF pixel
xPix8438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[84] VREF PIX_IN[8438] NB2 NB1 CSA_VREF pixel
xPix8439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[84] VREF PIX_IN[8439] NB2 NB1 CSA_VREF pixel
xPix8440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[84] VREF PIX_IN[8440] NB2 NB1 CSA_VREF pixel
xPix8441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[84] VREF PIX_IN[8441] NB2 NB1 CSA_VREF pixel
xPix8442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[84] VREF PIX_IN[8442] NB2 NB1 CSA_VREF pixel
xPix8443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[84] VREF PIX_IN[8443] NB2 NB1 CSA_VREF pixel
xPix8444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[84] VREF PIX_IN[8444] NB2 NB1 CSA_VREF pixel
xPix8445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[84] VREF PIX_IN[8445] NB2 NB1 CSA_VREF pixel
xPix8446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[84] VREF PIX_IN[8446] NB2 NB1 CSA_VREF pixel
xPix8447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[84] VREF PIX_IN[8447] NB2 NB1 CSA_VREF pixel
xPix8448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[84] VREF PIX_IN[8448] NB2 NB1 CSA_VREF pixel
xPix8449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[84] VREF PIX_IN[8449] NB2 NB1 CSA_VREF pixel
xPix8450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[84] VREF PIX_IN[8450] NB2 NB1 CSA_VREF pixel
xPix8451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[84] VREF PIX_IN[8451] NB2 NB1 CSA_VREF pixel
xPix8452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[84] VREF PIX_IN[8452] NB2 NB1 CSA_VREF pixel
xPix8453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[84] VREF PIX_IN[8453] NB2 NB1 CSA_VREF pixel
xPix8454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[84] VREF PIX_IN[8454] NB2 NB1 CSA_VREF pixel
xPix8455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[84] VREF PIX_IN[8455] NB2 NB1 CSA_VREF pixel
xPix8456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[84] VREF PIX_IN[8456] NB2 NB1 CSA_VREF pixel
xPix8457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[84] VREF PIX_IN[8457] NB2 NB1 CSA_VREF pixel
xPix8458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[84] VREF PIX_IN[8458] NB2 NB1 CSA_VREF pixel
xPix8459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[84] VREF PIX_IN[8459] NB2 NB1 CSA_VREF pixel
xPix8460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[84] VREF PIX_IN[8460] NB2 NB1 CSA_VREF pixel
xPix8461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[84] VREF PIX_IN[8461] NB2 NB1 CSA_VREF pixel
xPix8462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[84] VREF PIX_IN[8462] NB2 NB1 CSA_VREF pixel
xPix8463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[84] VREF PIX_IN[8463] NB2 NB1 CSA_VREF pixel
xPix8464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[84] VREF PIX_IN[8464] NB2 NB1 CSA_VREF pixel
xPix8465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[84] VREF PIX_IN[8465] NB2 NB1 CSA_VREF pixel
xPix8466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[84] VREF PIX_IN[8466] NB2 NB1 CSA_VREF pixel
xPix8467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[84] VREF PIX_IN[8467] NB2 NB1 CSA_VREF pixel
xPix8468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[84] VREF PIX_IN[8468] NB2 NB1 CSA_VREF pixel
xPix8469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[84] VREF PIX_IN[8469] NB2 NB1 CSA_VREF pixel
xPix8470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[84] VREF PIX_IN[8470] NB2 NB1 CSA_VREF pixel
xPix8471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[84] VREF PIX_IN[8471] NB2 NB1 CSA_VREF pixel
xPix8472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[84] VREF PIX_IN[8472] NB2 NB1 CSA_VREF pixel
xPix8473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[84] VREF PIX_IN[8473] NB2 NB1 CSA_VREF pixel
xPix8474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[84] VREF PIX_IN[8474] NB2 NB1 CSA_VREF pixel
xPix8475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[84] VREF PIX_IN[8475] NB2 NB1 CSA_VREF pixel
xPix8476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[84] VREF PIX_IN[8476] NB2 NB1 CSA_VREF pixel
xPix8477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[84] VREF PIX_IN[8477] NB2 NB1 CSA_VREF pixel
xPix8478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[84] VREF PIX_IN[8478] NB2 NB1 CSA_VREF pixel
xPix8479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[84] VREF PIX_IN[8479] NB2 NB1 CSA_VREF pixel
xPix8480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[84] VREF PIX_IN[8480] NB2 NB1 CSA_VREF pixel
xPix8481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[84] VREF PIX_IN[8481] NB2 NB1 CSA_VREF pixel
xPix8482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[84] VREF PIX_IN[8482] NB2 NB1 CSA_VREF pixel
xPix8483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[84] VREF PIX_IN[8483] NB2 NB1 CSA_VREF pixel
xPix8484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[84] VREF PIX_IN[8484] NB2 NB1 CSA_VREF pixel
xPix8485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[84] VREF PIX_IN[8485] NB2 NB1 CSA_VREF pixel
xPix8486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[84] VREF PIX_IN[8486] NB2 NB1 CSA_VREF pixel
xPix8487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[84] VREF PIX_IN[8487] NB2 NB1 CSA_VREF pixel
xPix8488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[84] VREF PIX_IN[8488] NB2 NB1 CSA_VREF pixel
xPix8489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[84] VREF PIX_IN[8489] NB2 NB1 CSA_VREF pixel
xPix8490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[84] VREF PIX_IN[8490] NB2 NB1 CSA_VREF pixel
xPix8491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[84] VREF PIX_IN[8491] NB2 NB1 CSA_VREF pixel
xPix8492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[84] VREF PIX_IN[8492] NB2 NB1 CSA_VREF pixel
xPix8493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[84] VREF PIX_IN[8493] NB2 NB1 CSA_VREF pixel
xPix8494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[84] VREF PIX_IN[8494] NB2 NB1 CSA_VREF pixel
xPix8495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[84] VREF PIX_IN[8495] NB2 NB1 CSA_VREF pixel
xPix8496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[84] VREF PIX_IN[8496] NB2 NB1 CSA_VREF pixel
xPix8497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[84] VREF PIX_IN[8497] NB2 NB1 CSA_VREF pixel
xPix8498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[84] VREF PIX_IN[8498] NB2 NB1 CSA_VREF pixel
xPix8499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[84] VREF PIX_IN[8499] NB2 NB1 CSA_VREF pixel
xPix8500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[85] VREF PIX_IN[8500] NB2 NB1 CSA_VREF pixel
xPix8501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[85] VREF PIX_IN[8501] NB2 NB1 CSA_VREF pixel
xPix8502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[85] VREF PIX_IN[8502] NB2 NB1 CSA_VREF pixel
xPix8503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[85] VREF PIX_IN[8503] NB2 NB1 CSA_VREF pixel
xPix8504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[85] VREF PIX_IN[8504] NB2 NB1 CSA_VREF pixel
xPix8505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[85] VREF PIX_IN[8505] NB2 NB1 CSA_VREF pixel
xPix8506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[85] VREF PIX_IN[8506] NB2 NB1 CSA_VREF pixel
xPix8507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[85] VREF PIX_IN[8507] NB2 NB1 CSA_VREF pixel
xPix8508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[85] VREF PIX_IN[8508] NB2 NB1 CSA_VREF pixel
xPix8509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[85] VREF PIX_IN[8509] NB2 NB1 CSA_VREF pixel
xPix8510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[85] VREF PIX_IN[8510] NB2 NB1 CSA_VREF pixel
xPix8511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[85] VREF PIX_IN[8511] NB2 NB1 CSA_VREF pixel
xPix8512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[85] VREF PIX_IN[8512] NB2 NB1 CSA_VREF pixel
xPix8513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[85] VREF PIX_IN[8513] NB2 NB1 CSA_VREF pixel
xPix8514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[85] VREF PIX_IN[8514] NB2 NB1 CSA_VREF pixel
xPix8515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[85] VREF PIX_IN[8515] NB2 NB1 CSA_VREF pixel
xPix8516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[85] VREF PIX_IN[8516] NB2 NB1 CSA_VREF pixel
xPix8517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[85] VREF PIX_IN[8517] NB2 NB1 CSA_VREF pixel
xPix8518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[85] VREF PIX_IN[8518] NB2 NB1 CSA_VREF pixel
xPix8519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[85] VREF PIX_IN[8519] NB2 NB1 CSA_VREF pixel
xPix8520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[85] VREF PIX_IN[8520] NB2 NB1 CSA_VREF pixel
xPix8521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[85] VREF PIX_IN[8521] NB2 NB1 CSA_VREF pixel
xPix8522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[85] VREF PIX_IN[8522] NB2 NB1 CSA_VREF pixel
xPix8523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[85] VREF PIX_IN[8523] NB2 NB1 CSA_VREF pixel
xPix8524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[85] VREF PIX_IN[8524] NB2 NB1 CSA_VREF pixel
xPix8525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[85] VREF PIX_IN[8525] NB2 NB1 CSA_VREF pixel
xPix8526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[85] VREF PIX_IN[8526] NB2 NB1 CSA_VREF pixel
xPix8527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[85] VREF PIX_IN[8527] NB2 NB1 CSA_VREF pixel
xPix8528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[85] VREF PIX_IN[8528] NB2 NB1 CSA_VREF pixel
xPix8529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[85] VREF PIX_IN[8529] NB2 NB1 CSA_VREF pixel
xPix8530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[85] VREF PIX_IN[8530] NB2 NB1 CSA_VREF pixel
xPix8531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[85] VREF PIX_IN[8531] NB2 NB1 CSA_VREF pixel
xPix8532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[85] VREF PIX_IN[8532] NB2 NB1 CSA_VREF pixel
xPix8533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[85] VREF PIX_IN[8533] NB2 NB1 CSA_VREF pixel
xPix8534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[85] VREF PIX_IN[8534] NB2 NB1 CSA_VREF pixel
xPix8535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[85] VREF PIX_IN[8535] NB2 NB1 CSA_VREF pixel
xPix8536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[85] VREF PIX_IN[8536] NB2 NB1 CSA_VREF pixel
xPix8537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[85] VREF PIX_IN[8537] NB2 NB1 CSA_VREF pixel
xPix8538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[85] VREF PIX_IN[8538] NB2 NB1 CSA_VREF pixel
xPix8539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[85] VREF PIX_IN[8539] NB2 NB1 CSA_VREF pixel
xPix8540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[85] VREF PIX_IN[8540] NB2 NB1 CSA_VREF pixel
xPix8541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[85] VREF PIX_IN[8541] NB2 NB1 CSA_VREF pixel
xPix8542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[85] VREF PIX_IN[8542] NB2 NB1 CSA_VREF pixel
xPix8543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[85] VREF PIX_IN[8543] NB2 NB1 CSA_VREF pixel
xPix8544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[85] VREF PIX_IN[8544] NB2 NB1 CSA_VREF pixel
xPix8545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[85] VREF PIX_IN[8545] NB2 NB1 CSA_VREF pixel
xPix8546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[85] VREF PIX_IN[8546] NB2 NB1 CSA_VREF pixel
xPix8547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[85] VREF PIX_IN[8547] NB2 NB1 CSA_VREF pixel
xPix8548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[85] VREF PIX_IN[8548] NB2 NB1 CSA_VREF pixel
xPix8549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[85] VREF PIX_IN[8549] NB2 NB1 CSA_VREF pixel
xPix8550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[85] VREF PIX_IN[8550] NB2 NB1 CSA_VREF pixel
xPix8551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[85] VREF PIX_IN[8551] NB2 NB1 CSA_VREF pixel
xPix8552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[85] VREF PIX_IN[8552] NB2 NB1 CSA_VREF pixel
xPix8553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[85] VREF PIX_IN[8553] NB2 NB1 CSA_VREF pixel
xPix8554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[85] VREF PIX_IN[8554] NB2 NB1 CSA_VREF pixel
xPix8555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[85] VREF PIX_IN[8555] NB2 NB1 CSA_VREF pixel
xPix8556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[85] VREF PIX_IN[8556] NB2 NB1 CSA_VREF pixel
xPix8557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[85] VREF PIX_IN[8557] NB2 NB1 CSA_VREF pixel
xPix8558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[85] VREF PIX_IN[8558] NB2 NB1 CSA_VREF pixel
xPix8559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[85] VREF PIX_IN[8559] NB2 NB1 CSA_VREF pixel
xPix8560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[85] VREF PIX_IN[8560] NB2 NB1 CSA_VREF pixel
xPix8561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[85] VREF PIX_IN[8561] NB2 NB1 CSA_VREF pixel
xPix8562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[85] VREF PIX_IN[8562] NB2 NB1 CSA_VREF pixel
xPix8563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[85] VREF PIX_IN[8563] NB2 NB1 CSA_VREF pixel
xPix8564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[85] VREF PIX_IN[8564] NB2 NB1 CSA_VREF pixel
xPix8565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[85] VREF PIX_IN[8565] NB2 NB1 CSA_VREF pixel
xPix8566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[85] VREF PIX_IN[8566] NB2 NB1 CSA_VREF pixel
xPix8567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[85] VREF PIX_IN[8567] NB2 NB1 CSA_VREF pixel
xPix8568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[85] VREF PIX_IN[8568] NB2 NB1 CSA_VREF pixel
xPix8569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[85] VREF PIX_IN[8569] NB2 NB1 CSA_VREF pixel
xPix8570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[85] VREF PIX_IN[8570] NB2 NB1 CSA_VREF pixel
xPix8571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[85] VREF PIX_IN[8571] NB2 NB1 CSA_VREF pixel
xPix8572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[85] VREF PIX_IN[8572] NB2 NB1 CSA_VREF pixel
xPix8573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[85] VREF PIX_IN[8573] NB2 NB1 CSA_VREF pixel
xPix8574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[85] VREF PIX_IN[8574] NB2 NB1 CSA_VREF pixel
xPix8575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[85] VREF PIX_IN[8575] NB2 NB1 CSA_VREF pixel
xPix8576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[85] VREF PIX_IN[8576] NB2 NB1 CSA_VREF pixel
xPix8577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[85] VREF PIX_IN[8577] NB2 NB1 CSA_VREF pixel
xPix8578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[85] VREF PIX_IN[8578] NB2 NB1 CSA_VREF pixel
xPix8579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[85] VREF PIX_IN[8579] NB2 NB1 CSA_VREF pixel
xPix8580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[85] VREF PIX_IN[8580] NB2 NB1 CSA_VREF pixel
xPix8581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[85] VREF PIX_IN[8581] NB2 NB1 CSA_VREF pixel
xPix8582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[85] VREF PIX_IN[8582] NB2 NB1 CSA_VREF pixel
xPix8583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[85] VREF PIX_IN[8583] NB2 NB1 CSA_VREF pixel
xPix8584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[85] VREF PIX_IN[8584] NB2 NB1 CSA_VREF pixel
xPix8585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[85] VREF PIX_IN[8585] NB2 NB1 CSA_VREF pixel
xPix8586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[85] VREF PIX_IN[8586] NB2 NB1 CSA_VREF pixel
xPix8587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[85] VREF PIX_IN[8587] NB2 NB1 CSA_VREF pixel
xPix8588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[85] VREF PIX_IN[8588] NB2 NB1 CSA_VREF pixel
xPix8589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[85] VREF PIX_IN[8589] NB2 NB1 CSA_VREF pixel
xPix8590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[85] VREF PIX_IN[8590] NB2 NB1 CSA_VREF pixel
xPix8591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[85] VREF PIX_IN[8591] NB2 NB1 CSA_VREF pixel
xPix8592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[85] VREF PIX_IN[8592] NB2 NB1 CSA_VREF pixel
xPix8593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[85] VREF PIX_IN[8593] NB2 NB1 CSA_VREF pixel
xPix8594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[85] VREF PIX_IN[8594] NB2 NB1 CSA_VREF pixel
xPix8595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[85] VREF PIX_IN[8595] NB2 NB1 CSA_VREF pixel
xPix8596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[85] VREF PIX_IN[8596] NB2 NB1 CSA_VREF pixel
xPix8597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[85] VREF PIX_IN[8597] NB2 NB1 CSA_VREF pixel
xPix8598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[85] VREF PIX_IN[8598] NB2 NB1 CSA_VREF pixel
xPix8599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[85] VREF PIX_IN[8599] NB2 NB1 CSA_VREF pixel
xPix8600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[86] VREF PIX_IN[8600] NB2 NB1 CSA_VREF pixel
xPix8601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[86] VREF PIX_IN[8601] NB2 NB1 CSA_VREF pixel
xPix8602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[86] VREF PIX_IN[8602] NB2 NB1 CSA_VREF pixel
xPix8603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[86] VREF PIX_IN[8603] NB2 NB1 CSA_VREF pixel
xPix8604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[86] VREF PIX_IN[8604] NB2 NB1 CSA_VREF pixel
xPix8605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[86] VREF PIX_IN[8605] NB2 NB1 CSA_VREF pixel
xPix8606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[86] VREF PIX_IN[8606] NB2 NB1 CSA_VREF pixel
xPix8607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[86] VREF PIX_IN[8607] NB2 NB1 CSA_VREF pixel
xPix8608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[86] VREF PIX_IN[8608] NB2 NB1 CSA_VREF pixel
xPix8609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[86] VREF PIX_IN[8609] NB2 NB1 CSA_VREF pixel
xPix8610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[86] VREF PIX_IN[8610] NB2 NB1 CSA_VREF pixel
xPix8611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[86] VREF PIX_IN[8611] NB2 NB1 CSA_VREF pixel
xPix8612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[86] VREF PIX_IN[8612] NB2 NB1 CSA_VREF pixel
xPix8613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[86] VREF PIX_IN[8613] NB2 NB1 CSA_VREF pixel
xPix8614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[86] VREF PIX_IN[8614] NB2 NB1 CSA_VREF pixel
xPix8615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[86] VREF PIX_IN[8615] NB2 NB1 CSA_VREF pixel
xPix8616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[86] VREF PIX_IN[8616] NB2 NB1 CSA_VREF pixel
xPix8617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[86] VREF PIX_IN[8617] NB2 NB1 CSA_VREF pixel
xPix8618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[86] VREF PIX_IN[8618] NB2 NB1 CSA_VREF pixel
xPix8619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[86] VREF PIX_IN[8619] NB2 NB1 CSA_VREF pixel
xPix8620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[86] VREF PIX_IN[8620] NB2 NB1 CSA_VREF pixel
xPix8621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[86] VREF PIX_IN[8621] NB2 NB1 CSA_VREF pixel
xPix8622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[86] VREF PIX_IN[8622] NB2 NB1 CSA_VREF pixel
xPix8623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[86] VREF PIX_IN[8623] NB2 NB1 CSA_VREF pixel
xPix8624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[86] VREF PIX_IN[8624] NB2 NB1 CSA_VREF pixel
xPix8625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[86] VREF PIX_IN[8625] NB2 NB1 CSA_VREF pixel
xPix8626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[86] VREF PIX_IN[8626] NB2 NB1 CSA_VREF pixel
xPix8627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[86] VREF PIX_IN[8627] NB2 NB1 CSA_VREF pixel
xPix8628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[86] VREF PIX_IN[8628] NB2 NB1 CSA_VREF pixel
xPix8629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[86] VREF PIX_IN[8629] NB2 NB1 CSA_VREF pixel
xPix8630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[86] VREF PIX_IN[8630] NB2 NB1 CSA_VREF pixel
xPix8631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[86] VREF PIX_IN[8631] NB2 NB1 CSA_VREF pixel
xPix8632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[86] VREF PIX_IN[8632] NB2 NB1 CSA_VREF pixel
xPix8633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[86] VREF PIX_IN[8633] NB2 NB1 CSA_VREF pixel
xPix8634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[86] VREF PIX_IN[8634] NB2 NB1 CSA_VREF pixel
xPix8635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[86] VREF PIX_IN[8635] NB2 NB1 CSA_VREF pixel
xPix8636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[86] VREF PIX_IN[8636] NB2 NB1 CSA_VREF pixel
xPix8637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[86] VREF PIX_IN[8637] NB2 NB1 CSA_VREF pixel
xPix8638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[86] VREF PIX_IN[8638] NB2 NB1 CSA_VREF pixel
xPix8639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[86] VREF PIX_IN[8639] NB2 NB1 CSA_VREF pixel
xPix8640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[86] VREF PIX_IN[8640] NB2 NB1 CSA_VREF pixel
xPix8641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[86] VREF PIX_IN[8641] NB2 NB1 CSA_VREF pixel
xPix8642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[86] VREF PIX_IN[8642] NB2 NB1 CSA_VREF pixel
xPix8643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[86] VREF PIX_IN[8643] NB2 NB1 CSA_VREF pixel
xPix8644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[86] VREF PIX_IN[8644] NB2 NB1 CSA_VREF pixel
xPix8645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[86] VREF PIX_IN[8645] NB2 NB1 CSA_VREF pixel
xPix8646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[86] VREF PIX_IN[8646] NB2 NB1 CSA_VREF pixel
xPix8647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[86] VREF PIX_IN[8647] NB2 NB1 CSA_VREF pixel
xPix8648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[86] VREF PIX_IN[8648] NB2 NB1 CSA_VREF pixel
xPix8649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[86] VREF PIX_IN[8649] NB2 NB1 CSA_VREF pixel
xPix8650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[86] VREF PIX_IN[8650] NB2 NB1 CSA_VREF pixel
xPix8651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[86] VREF PIX_IN[8651] NB2 NB1 CSA_VREF pixel
xPix8652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[86] VREF PIX_IN[8652] NB2 NB1 CSA_VREF pixel
xPix8653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[86] VREF PIX_IN[8653] NB2 NB1 CSA_VREF pixel
xPix8654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[86] VREF PIX_IN[8654] NB2 NB1 CSA_VREF pixel
xPix8655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[86] VREF PIX_IN[8655] NB2 NB1 CSA_VREF pixel
xPix8656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[86] VREF PIX_IN[8656] NB2 NB1 CSA_VREF pixel
xPix8657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[86] VREF PIX_IN[8657] NB2 NB1 CSA_VREF pixel
xPix8658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[86] VREF PIX_IN[8658] NB2 NB1 CSA_VREF pixel
xPix8659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[86] VREF PIX_IN[8659] NB2 NB1 CSA_VREF pixel
xPix8660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[86] VREF PIX_IN[8660] NB2 NB1 CSA_VREF pixel
xPix8661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[86] VREF PIX_IN[8661] NB2 NB1 CSA_VREF pixel
xPix8662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[86] VREF PIX_IN[8662] NB2 NB1 CSA_VREF pixel
xPix8663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[86] VREF PIX_IN[8663] NB2 NB1 CSA_VREF pixel
xPix8664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[86] VREF PIX_IN[8664] NB2 NB1 CSA_VREF pixel
xPix8665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[86] VREF PIX_IN[8665] NB2 NB1 CSA_VREF pixel
xPix8666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[86] VREF PIX_IN[8666] NB2 NB1 CSA_VREF pixel
xPix8667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[86] VREF PIX_IN[8667] NB2 NB1 CSA_VREF pixel
xPix8668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[86] VREF PIX_IN[8668] NB2 NB1 CSA_VREF pixel
xPix8669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[86] VREF PIX_IN[8669] NB2 NB1 CSA_VREF pixel
xPix8670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[86] VREF PIX_IN[8670] NB2 NB1 CSA_VREF pixel
xPix8671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[86] VREF PIX_IN[8671] NB2 NB1 CSA_VREF pixel
xPix8672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[86] VREF PIX_IN[8672] NB2 NB1 CSA_VREF pixel
xPix8673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[86] VREF PIX_IN[8673] NB2 NB1 CSA_VREF pixel
xPix8674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[86] VREF PIX_IN[8674] NB2 NB1 CSA_VREF pixel
xPix8675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[86] VREF PIX_IN[8675] NB2 NB1 CSA_VREF pixel
xPix8676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[86] VREF PIX_IN[8676] NB2 NB1 CSA_VREF pixel
xPix8677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[86] VREF PIX_IN[8677] NB2 NB1 CSA_VREF pixel
xPix8678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[86] VREF PIX_IN[8678] NB2 NB1 CSA_VREF pixel
xPix8679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[86] VREF PIX_IN[8679] NB2 NB1 CSA_VREF pixel
xPix8680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[86] VREF PIX_IN[8680] NB2 NB1 CSA_VREF pixel
xPix8681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[86] VREF PIX_IN[8681] NB2 NB1 CSA_VREF pixel
xPix8682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[86] VREF PIX_IN[8682] NB2 NB1 CSA_VREF pixel
xPix8683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[86] VREF PIX_IN[8683] NB2 NB1 CSA_VREF pixel
xPix8684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[86] VREF PIX_IN[8684] NB2 NB1 CSA_VREF pixel
xPix8685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[86] VREF PIX_IN[8685] NB2 NB1 CSA_VREF pixel
xPix8686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[86] VREF PIX_IN[8686] NB2 NB1 CSA_VREF pixel
xPix8687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[86] VREF PIX_IN[8687] NB2 NB1 CSA_VREF pixel
xPix8688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[86] VREF PIX_IN[8688] NB2 NB1 CSA_VREF pixel
xPix8689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[86] VREF PIX_IN[8689] NB2 NB1 CSA_VREF pixel
xPix8690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[86] VREF PIX_IN[8690] NB2 NB1 CSA_VREF pixel
xPix8691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[86] VREF PIX_IN[8691] NB2 NB1 CSA_VREF pixel
xPix8692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[86] VREF PIX_IN[8692] NB2 NB1 CSA_VREF pixel
xPix8693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[86] VREF PIX_IN[8693] NB2 NB1 CSA_VREF pixel
xPix8694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[86] VREF PIX_IN[8694] NB2 NB1 CSA_VREF pixel
xPix8695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[86] VREF PIX_IN[8695] NB2 NB1 CSA_VREF pixel
xPix8696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[86] VREF PIX_IN[8696] NB2 NB1 CSA_VREF pixel
xPix8697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[86] VREF PIX_IN[8697] NB2 NB1 CSA_VREF pixel
xPix8698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[86] VREF PIX_IN[8698] NB2 NB1 CSA_VREF pixel
xPix8699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[86] VREF PIX_IN[8699] NB2 NB1 CSA_VREF pixel
xPix8700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[87] VREF PIX_IN[8700] NB2 NB1 CSA_VREF pixel
xPix8701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[87] VREF PIX_IN[8701] NB2 NB1 CSA_VREF pixel
xPix8702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[87] VREF PIX_IN[8702] NB2 NB1 CSA_VREF pixel
xPix8703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[87] VREF PIX_IN[8703] NB2 NB1 CSA_VREF pixel
xPix8704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[87] VREF PIX_IN[8704] NB2 NB1 CSA_VREF pixel
xPix8705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[87] VREF PIX_IN[8705] NB2 NB1 CSA_VREF pixel
xPix8706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[87] VREF PIX_IN[8706] NB2 NB1 CSA_VREF pixel
xPix8707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[87] VREF PIX_IN[8707] NB2 NB1 CSA_VREF pixel
xPix8708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[87] VREF PIX_IN[8708] NB2 NB1 CSA_VREF pixel
xPix8709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[87] VREF PIX_IN[8709] NB2 NB1 CSA_VREF pixel
xPix8710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[87] VREF PIX_IN[8710] NB2 NB1 CSA_VREF pixel
xPix8711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[87] VREF PIX_IN[8711] NB2 NB1 CSA_VREF pixel
xPix8712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[87] VREF PIX_IN[8712] NB2 NB1 CSA_VREF pixel
xPix8713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[87] VREF PIX_IN[8713] NB2 NB1 CSA_VREF pixel
xPix8714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[87] VREF PIX_IN[8714] NB2 NB1 CSA_VREF pixel
xPix8715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[87] VREF PIX_IN[8715] NB2 NB1 CSA_VREF pixel
xPix8716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[87] VREF PIX_IN[8716] NB2 NB1 CSA_VREF pixel
xPix8717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[87] VREF PIX_IN[8717] NB2 NB1 CSA_VREF pixel
xPix8718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[87] VREF PIX_IN[8718] NB2 NB1 CSA_VREF pixel
xPix8719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[87] VREF PIX_IN[8719] NB2 NB1 CSA_VREF pixel
xPix8720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[87] VREF PIX_IN[8720] NB2 NB1 CSA_VREF pixel
xPix8721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[87] VREF PIX_IN[8721] NB2 NB1 CSA_VREF pixel
xPix8722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[87] VREF PIX_IN[8722] NB2 NB1 CSA_VREF pixel
xPix8723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[87] VREF PIX_IN[8723] NB2 NB1 CSA_VREF pixel
xPix8724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[87] VREF PIX_IN[8724] NB2 NB1 CSA_VREF pixel
xPix8725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[87] VREF PIX_IN[8725] NB2 NB1 CSA_VREF pixel
xPix8726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[87] VREF PIX_IN[8726] NB2 NB1 CSA_VREF pixel
xPix8727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[87] VREF PIX_IN[8727] NB2 NB1 CSA_VREF pixel
xPix8728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[87] VREF PIX_IN[8728] NB2 NB1 CSA_VREF pixel
xPix8729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[87] VREF PIX_IN[8729] NB2 NB1 CSA_VREF pixel
xPix8730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[87] VREF PIX_IN[8730] NB2 NB1 CSA_VREF pixel
xPix8731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[87] VREF PIX_IN[8731] NB2 NB1 CSA_VREF pixel
xPix8732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[87] VREF PIX_IN[8732] NB2 NB1 CSA_VREF pixel
xPix8733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[87] VREF PIX_IN[8733] NB2 NB1 CSA_VREF pixel
xPix8734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[87] VREF PIX_IN[8734] NB2 NB1 CSA_VREF pixel
xPix8735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[87] VREF PIX_IN[8735] NB2 NB1 CSA_VREF pixel
xPix8736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[87] VREF PIX_IN[8736] NB2 NB1 CSA_VREF pixel
xPix8737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[87] VREF PIX_IN[8737] NB2 NB1 CSA_VREF pixel
xPix8738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[87] VREF PIX_IN[8738] NB2 NB1 CSA_VREF pixel
xPix8739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[87] VREF PIX_IN[8739] NB2 NB1 CSA_VREF pixel
xPix8740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[87] VREF PIX_IN[8740] NB2 NB1 CSA_VREF pixel
xPix8741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[87] VREF PIX_IN[8741] NB2 NB1 CSA_VREF pixel
xPix8742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[87] VREF PIX_IN[8742] NB2 NB1 CSA_VREF pixel
xPix8743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[87] VREF PIX_IN[8743] NB2 NB1 CSA_VREF pixel
xPix8744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[87] VREF PIX_IN[8744] NB2 NB1 CSA_VREF pixel
xPix8745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[87] VREF PIX_IN[8745] NB2 NB1 CSA_VREF pixel
xPix8746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[87] VREF PIX_IN[8746] NB2 NB1 CSA_VREF pixel
xPix8747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[87] VREF PIX_IN[8747] NB2 NB1 CSA_VREF pixel
xPix8748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[87] VREF PIX_IN[8748] NB2 NB1 CSA_VREF pixel
xPix8749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[87] VREF PIX_IN[8749] NB2 NB1 CSA_VREF pixel
xPix8750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[87] VREF PIX_IN[8750] NB2 NB1 CSA_VREF pixel
xPix8751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[87] VREF PIX_IN[8751] NB2 NB1 CSA_VREF pixel
xPix8752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[87] VREF PIX_IN[8752] NB2 NB1 CSA_VREF pixel
xPix8753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[87] VREF PIX_IN[8753] NB2 NB1 CSA_VREF pixel
xPix8754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[87] VREF PIX_IN[8754] NB2 NB1 CSA_VREF pixel
xPix8755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[87] VREF PIX_IN[8755] NB2 NB1 CSA_VREF pixel
xPix8756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[87] VREF PIX_IN[8756] NB2 NB1 CSA_VREF pixel
xPix8757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[87] VREF PIX_IN[8757] NB2 NB1 CSA_VREF pixel
xPix8758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[87] VREF PIX_IN[8758] NB2 NB1 CSA_VREF pixel
xPix8759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[87] VREF PIX_IN[8759] NB2 NB1 CSA_VREF pixel
xPix8760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[87] VREF PIX_IN[8760] NB2 NB1 CSA_VREF pixel
xPix8761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[87] VREF PIX_IN[8761] NB2 NB1 CSA_VREF pixel
xPix8762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[87] VREF PIX_IN[8762] NB2 NB1 CSA_VREF pixel
xPix8763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[87] VREF PIX_IN[8763] NB2 NB1 CSA_VREF pixel
xPix8764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[87] VREF PIX_IN[8764] NB2 NB1 CSA_VREF pixel
xPix8765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[87] VREF PIX_IN[8765] NB2 NB1 CSA_VREF pixel
xPix8766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[87] VREF PIX_IN[8766] NB2 NB1 CSA_VREF pixel
xPix8767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[87] VREF PIX_IN[8767] NB2 NB1 CSA_VREF pixel
xPix8768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[87] VREF PIX_IN[8768] NB2 NB1 CSA_VREF pixel
xPix8769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[87] VREF PIX_IN[8769] NB2 NB1 CSA_VREF pixel
xPix8770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[87] VREF PIX_IN[8770] NB2 NB1 CSA_VREF pixel
xPix8771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[87] VREF PIX_IN[8771] NB2 NB1 CSA_VREF pixel
xPix8772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[87] VREF PIX_IN[8772] NB2 NB1 CSA_VREF pixel
xPix8773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[87] VREF PIX_IN[8773] NB2 NB1 CSA_VREF pixel
xPix8774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[87] VREF PIX_IN[8774] NB2 NB1 CSA_VREF pixel
xPix8775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[87] VREF PIX_IN[8775] NB2 NB1 CSA_VREF pixel
xPix8776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[87] VREF PIX_IN[8776] NB2 NB1 CSA_VREF pixel
xPix8777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[87] VREF PIX_IN[8777] NB2 NB1 CSA_VREF pixel
xPix8778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[87] VREF PIX_IN[8778] NB2 NB1 CSA_VREF pixel
xPix8779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[87] VREF PIX_IN[8779] NB2 NB1 CSA_VREF pixel
xPix8780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[87] VREF PIX_IN[8780] NB2 NB1 CSA_VREF pixel
xPix8781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[87] VREF PIX_IN[8781] NB2 NB1 CSA_VREF pixel
xPix8782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[87] VREF PIX_IN[8782] NB2 NB1 CSA_VREF pixel
xPix8783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[87] VREF PIX_IN[8783] NB2 NB1 CSA_VREF pixel
xPix8784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[87] VREF PIX_IN[8784] NB2 NB1 CSA_VREF pixel
xPix8785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[87] VREF PIX_IN[8785] NB2 NB1 CSA_VREF pixel
xPix8786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[87] VREF PIX_IN[8786] NB2 NB1 CSA_VREF pixel
xPix8787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[87] VREF PIX_IN[8787] NB2 NB1 CSA_VREF pixel
xPix8788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[87] VREF PIX_IN[8788] NB2 NB1 CSA_VREF pixel
xPix8789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[87] VREF PIX_IN[8789] NB2 NB1 CSA_VREF pixel
xPix8790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[87] VREF PIX_IN[8790] NB2 NB1 CSA_VREF pixel
xPix8791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[87] VREF PIX_IN[8791] NB2 NB1 CSA_VREF pixel
xPix8792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[87] VREF PIX_IN[8792] NB2 NB1 CSA_VREF pixel
xPix8793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[87] VREF PIX_IN[8793] NB2 NB1 CSA_VREF pixel
xPix8794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[87] VREF PIX_IN[8794] NB2 NB1 CSA_VREF pixel
xPix8795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[87] VREF PIX_IN[8795] NB2 NB1 CSA_VREF pixel
xPix8796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[87] VREF PIX_IN[8796] NB2 NB1 CSA_VREF pixel
xPix8797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[87] VREF PIX_IN[8797] NB2 NB1 CSA_VREF pixel
xPix8798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[87] VREF PIX_IN[8798] NB2 NB1 CSA_VREF pixel
xPix8799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[87] VREF PIX_IN[8799] NB2 NB1 CSA_VREF pixel
xPix8800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[88] VREF PIX_IN[8800] NB2 NB1 CSA_VREF pixel
xPix8801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[88] VREF PIX_IN[8801] NB2 NB1 CSA_VREF pixel
xPix8802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[88] VREF PIX_IN[8802] NB2 NB1 CSA_VREF pixel
xPix8803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[88] VREF PIX_IN[8803] NB2 NB1 CSA_VREF pixel
xPix8804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[88] VREF PIX_IN[8804] NB2 NB1 CSA_VREF pixel
xPix8805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[88] VREF PIX_IN[8805] NB2 NB1 CSA_VREF pixel
xPix8806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[88] VREF PIX_IN[8806] NB2 NB1 CSA_VREF pixel
xPix8807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[88] VREF PIX_IN[8807] NB2 NB1 CSA_VREF pixel
xPix8808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[88] VREF PIX_IN[8808] NB2 NB1 CSA_VREF pixel
xPix8809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[88] VREF PIX_IN[8809] NB2 NB1 CSA_VREF pixel
xPix8810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[88] VREF PIX_IN[8810] NB2 NB1 CSA_VREF pixel
xPix8811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[88] VREF PIX_IN[8811] NB2 NB1 CSA_VREF pixel
xPix8812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[88] VREF PIX_IN[8812] NB2 NB1 CSA_VREF pixel
xPix8813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[88] VREF PIX_IN[8813] NB2 NB1 CSA_VREF pixel
xPix8814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[88] VREF PIX_IN[8814] NB2 NB1 CSA_VREF pixel
xPix8815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[88] VREF PIX_IN[8815] NB2 NB1 CSA_VREF pixel
xPix8816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[88] VREF PIX_IN[8816] NB2 NB1 CSA_VREF pixel
xPix8817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[88] VREF PIX_IN[8817] NB2 NB1 CSA_VREF pixel
xPix8818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[88] VREF PIX_IN[8818] NB2 NB1 CSA_VREF pixel
xPix8819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[88] VREF PIX_IN[8819] NB2 NB1 CSA_VREF pixel
xPix8820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[88] VREF PIX_IN[8820] NB2 NB1 CSA_VREF pixel
xPix8821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[88] VREF PIX_IN[8821] NB2 NB1 CSA_VREF pixel
xPix8822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[88] VREF PIX_IN[8822] NB2 NB1 CSA_VREF pixel
xPix8823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[88] VREF PIX_IN[8823] NB2 NB1 CSA_VREF pixel
xPix8824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[88] VREF PIX_IN[8824] NB2 NB1 CSA_VREF pixel
xPix8825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[88] VREF PIX_IN[8825] NB2 NB1 CSA_VREF pixel
xPix8826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[88] VREF PIX_IN[8826] NB2 NB1 CSA_VREF pixel
xPix8827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[88] VREF PIX_IN[8827] NB2 NB1 CSA_VREF pixel
xPix8828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[88] VREF PIX_IN[8828] NB2 NB1 CSA_VREF pixel
xPix8829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[88] VREF PIX_IN[8829] NB2 NB1 CSA_VREF pixel
xPix8830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[88] VREF PIX_IN[8830] NB2 NB1 CSA_VREF pixel
xPix8831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[88] VREF PIX_IN[8831] NB2 NB1 CSA_VREF pixel
xPix8832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[88] VREF PIX_IN[8832] NB2 NB1 CSA_VREF pixel
xPix8833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[88] VREF PIX_IN[8833] NB2 NB1 CSA_VREF pixel
xPix8834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[88] VREF PIX_IN[8834] NB2 NB1 CSA_VREF pixel
xPix8835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[88] VREF PIX_IN[8835] NB2 NB1 CSA_VREF pixel
xPix8836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[88] VREF PIX_IN[8836] NB2 NB1 CSA_VREF pixel
xPix8837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[88] VREF PIX_IN[8837] NB2 NB1 CSA_VREF pixel
xPix8838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[88] VREF PIX_IN[8838] NB2 NB1 CSA_VREF pixel
xPix8839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[88] VREF PIX_IN[8839] NB2 NB1 CSA_VREF pixel
xPix8840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[88] VREF PIX_IN[8840] NB2 NB1 CSA_VREF pixel
xPix8841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[88] VREF PIX_IN[8841] NB2 NB1 CSA_VREF pixel
xPix8842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[88] VREF PIX_IN[8842] NB2 NB1 CSA_VREF pixel
xPix8843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[88] VREF PIX_IN[8843] NB2 NB1 CSA_VREF pixel
xPix8844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[88] VREF PIX_IN[8844] NB2 NB1 CSA_VREF pixel
xPix8845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[88] VREF PIX_IN[8845] NB2 NB1 CSA_VREF pixel
xPix8846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[88] VREF PIX_IN[8846] NB2 NB1 CSA_VREF pixel
xPix8847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[88] VREF PIX_IN[8847] NB2 NB1 CSA_VREF pixel
xPix8848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[88] VREF PIX_IN[8848] NB2 NB1 CSA_VREF pixel
xPix8849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[88] VREF PIX_IN[8849] NB2 NB1 CSA_VREF pixel
xPix8850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[88] VREF PIX_IN[8850] NB2 NB1 CSA_VREF pixel
xPix8851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[88] VREF PIX_IN[8851] NB2 NB1 CSA_VREF pixel
xPix8852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[88] VREF PIX_IN[8852] NB2 NB1 CSA_VREF pixel
xPix8853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[88] VREF PIX_IN[8853] NB2 NB1 CSA_VREF pixel
xPix8854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[88] VREF PIX_IN[8854] NB2 NB1 CSA_VREF pixel
xPix8855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[88] VREF PIX_IN[8855] NB2 NB1 CSA_VREF pixel
xPix8856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[88] VREF PIX_IN[8856] NB2 NB1 CSA_VREF pixel
xPix8857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[88] VREF PIX_IN[8857] NB2 NB1 CSA_VREF pixel
xPix8858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[88] VREF PIX_IN[8858] NB2 NB1 CSA_VREF pixel
xPix8859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[88] VREF PIX_IN[8859] NB2 NB1 CSA_VREF pixel
xPix8860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[88] VREF PIX_IN[8860] NB2 NB1 CSA_VREF pixel
xPix8861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[88] VREF PIX_IN[8861] NB2 NB1 CSA_VREF pixel
xPix8862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[88] VREF PIX_IN[8862] NB2 NB1 CSA_VREF pixel
xPix8863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[88] VREF PIX_IN[8863] NB2 NB1 CSA_VREF pixel
xPix8864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[88] VREF PIX_IN[8864] NB2 NB1 CSA_VREF pixel
xPix8865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[88] VREF PIX_IN[8865] NB2 NB1 CSA_VREF pixel
xPix8866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[88] VREF PIX_IN[8866] NB2 NB1 CSA_VREF pixel
xPix8867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[88] VREF PIX_IN[8867] NB2 NB1 CSA_VREF pixel
xPix8868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[88] VREF PIX_IN[8868] NB2 NB1 CSA_VREF pixel
xPix8869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[88] VREF PIX_IN[8869] NB2 NB1 CSA_VREF pixel
xPix8870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[88] VREF PIX_IN[8870] NB2 NB1 CSA_VREF pixel
xPix8871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[88] VREF PIX_IN[8871] NB2 NB1 CSA_VREF pixel
xPix8872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[88] VREF PIX_IN[8872] NB2 NB1 CSA_VREF pixel
xPix8873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[88] VREF PIX_IN[8873] NB2 NB1 CSA_VREF pixel
xPix8874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[88] VREF PIX_IN[8874] NB2 NB1 CSA_VREF pixel
xPix8875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[88] VREF PIX_IN[8875] NB2 NB1 CSA_VREF pixel
xPix8876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[88] VREF PIX_IN[8876] NB2 NB1 CSA_VREF pixel
xPix8877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[88] VREF PIX_IN[8877] NB2 NB1 CSA_VREF pixel
xPix8878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[88] VREF PIX_IN[8878] NB2 NB1 CSA_VREF pixel
xPix8879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[88] VREF PIX_IN[8879] NB2 NB1 CSA_VREF pixel
xPix8880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[88] VREF PIX_IN[8880] NB2 NB1 CSA_VREF pixel
xPix8881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[88] VREF PIX_IN[8881] NB2 NB1 CSA_VREF pixel
xPix8882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[88] VREF PIX_IN[8882] NB2 NB1 CSA_VREF pixel
xPix8883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[88] VREF PIX_IN[8883] NB2 NB1 CSA_VREF pixel
xPix8884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[88] VREF PIX_IN[8884] NB2 NB1 CSA_VREF pixel
xPix8885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[88] VREF PIX_IN[8885] NB2 NB1 CSA_VREF pixel
xPix8886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[88] VREF PIX_IN[8886] NB2 NB1 CSA_VREF pixel
xPix8887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[88] VREF PIX_IN[8887] NB2 NB1 CSA_VREF pixel
xPix8888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[88] VREF PIX_IN[8888] NB2 NB1 CSA_VREF pixel
xPix8889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[88] VREF PIX_IN[8889] NB2 NB1 CSA_VREF pixel
xPix8890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[88] VREF PIX_IN[8890] NB2 NB1 CSA_VREF pixel
xPix8891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[88] VREF PIX_IN[8891] NB2 NB1 CSA_VREF pixel
xPix8892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[88] VREF PIX_IN[8892] NB2 NB1 CSA_VREF pixel
xPix8893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[88] VREF PIX_IN[8893] NB2 NB1 CSA_VREF pixel
xPix8894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[88] VREF PIX_IN[8894] NB2 NB1 CSA_VREF pixel
xPix8895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[88] VREF PIX_IN[8895] NB2 NB1 CSA_VREF pixel
xPix8896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[88] VREF PIX_IN[8896] NB2 NB1 CSA_VREF pixel
xPix8897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[88] VREF PIX_IN[8897] NB2 NB1 CSA_VREF pixel
xPix8898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[88] VREF PIX_IN[8898] NB2 NB1 CSA_VREF pixel
xPix8899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[88] VREF PIX_IN[8899] NB2 NB1 CSA_VREF pixel
xPix8900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[89] VREF PIX_IN[8900] NB2 NB1 CSA_VREF pixel
xPix8901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[89] VREF PIX_IN[8901] NB2 NB1 CSA_VREF pixel
xPix8902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[89] VREF PIX_IN[8902] NB2 NB1 CSA_VREF pixel
xPix8903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[89] VREF PIX_IN[8903] NB2 NB1 CSA_VREF pixel
xPix8904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[89] VREF PIX_IN[8904] NB2 NB1 CSA_VREF pixel
xPix8905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[89] VREF PIX_IN[8905] NB2 NB1 CSA_VREF pixel
xPix8906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[89] VREF PIX_IN[8906] NB2 NB1 CSA_VREF pixel
xPix8907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[89] VREF PIX_IN[8907] NB2 NB1 CSA_VREF pixel
xPix8908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[89] VREF PIX_IN[8908] NB2 NB1 CSA_VREF pixel
xPix8909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[89] VREF PIX_IN[8909] NB2 NB1 CSA_VREF pixel
xPix8910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[89] VREF PIX_IN[8910] NB2 NB1 CSA_VREF pixel
xPix8911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[89] VREF PIX_IN[8911] NB2 NB1 CSA_VREF pixel
xPix8912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[89] VREF PIX_IN[8912] NB2 NB1 CSA_VREF pixel
xPix8913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[89] VREF PIX_IN[8913] NB2 NB1 CSA_VREF pixel
xPix8914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[89] VREF PIX_IN[8914] NB2 NB1 CSA_VREF pixel
xPix8915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[89] VREF PIX_IN[8915] NB2 NB1 CSA_VREF pixel
xPix8916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[89] VREF PIX_IN[8916] NB2 NB1 CSA_VREF pixel
xPix8917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[89] VREF PIX_IN[8917] NB2 NB1 CSA_VREF pixel
xPix8918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[89] VREF PIX_IN[8918] NB2 NB1 CSA_VREF pixel
xPix8919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[89] VREF PIX_IN[8919] NB2 NB1 CSA_VREF pixel
xPix8920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[89] VREF PIX_IN[8920] NB2 NB1 CSA_VREF pixel
xPix8921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[89] VREF PIX_IN[8921] NB2 NB1 CSA_VREF pixel
xPix8922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[89] VREF PIX_IN[8922] NB2 NB1 CSA_VREF pixel
xPix8923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[89] VREF PIX_IN[8923] NB2 NB1 CSA_VREF pixel
xPix8924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[89] VREF PIX_IN[8924] NB2 NB1 CSA_VREF pixel
xPix8925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[89] VREF PIX_IN[8925] NB2 NB1 CSA_VREF pixel
xPix8926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[89] VREF PIX_IN[8926] NB2 NB1 CSA_VREF pixel
xPix8927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[89] VREF PIX_IN[8927] NB2 NB1 CSA_VREF pixel
xPix8928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[89] VREF PIX_IN[8928] NB2 NB1 CSA_VREF pixel
xPix8929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[89] VREF PIX_IN[8929] NB2 NB1 CSA_VREF pixel
xPix8930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[89] VREF PIX_IN[8930] NB2 NB1 CSA_VREF pixel
xPix8931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[89] VREF PIX_IN[8931] NB2 NB1 CSA_VREF pixel
xPix8932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[89] VREF PIX_IN[8932] NB2 NB1 CSA_VREF pixel
xPix8933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[89] VREF PIX_IN[8933] NB2 NB1 CSA_VREF pixel
xPix8934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[89] VREF PIX_IN[8934] NB2 NB1 CSA_VREF pixel
xPix8935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[89] VREF PIX_IN[8935] NB2 NB1 CSA_VREF pixel
xPix8936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[89] VREF PIX_IN[8936] NB2 NB1 CSA_VREF pixel
xPix8937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[89] VREF PIX_IN[8937] NB2 NB1 CSA_VREF pixel
xPix8938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[89] VREF PIX_IN[8938] NB2 NB1 CSA_VREF pixel
xPix8939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[89] VREF PIX_IN[8939] NB2 NB1 CSA_VREF pixel
xPix8940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[89] VREF PIX_IN[8940] NB2 NB1 CSA_VREF pixel
xPix8941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[89] VREF PIX_IN[8941] NB2 NB1 CSA_VREF pixel
xPix8942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[89] VREF PIX_IN[8942] NB2 NB1 CSA_VREF pixel
xPix8943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[89] VREF PIX_IN[8943] NB2 NB1 CSA_VREF pixel
xPix8944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[89] VREF PIX_IN[8944] NB2 NB1 CSA_VREF pixel
xPix8945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[89] VREF PIX_IN[8945] NB2 NB1 CSA_VREF pixel
xPix8946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[89] VREF PIX_IN[8946] NB2 NB1 CSA_VREF pixel
xPix8947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[89] VREF PIX_IN[8947] NB2 NB1 CSA_VREF pixel
xPix8948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[89] VREF PIX_IN[8948] NB2 NB1 CSA_VREF pixel
xPix8949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[89] VREF PIX_IN[8949] NB2 NB1 CSA_VREF pixel
xPix8950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[89] VREF PIX_IN[8950] NB2 NB1 CSA_VREF pixel
xPix8951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[89] VREF PIX_IN[8951] NB2 NB1 CSA_VREF pixel
xPix8952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[89] VREF PIX_IN[8952] NB2 NB1 CSA_VREF pixel
xPix8953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[89] VREF PIX_IN[8953] NB2 NB1 CSA_VREF pixel
xPix8954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[89] VREF PIX_IN[8954] NB2 NB1 CSA_VREF pixel
xPix8955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[89] VREF PIX_IN[8955] NB2 NB1 CSA_VREF pixel
xPix8956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[89] VREF PIX_IN[8956] NB2 NB1 CSA_VREF pixel
xPix8957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[89] VREF PIX_IN[8957] NB2 NB1 CSA_VREF pixel
xPix8958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[89] VREF PIX_IN[8958] NB2 NB1 CSA_VREF pixel
xPix8959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[89] VREF PIX_IN[8959] NB2 NB1 CSA_VREF pixel
xPix8960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[89] VREF PIX_IN[8960] NB2 NB1 CSA_VREF pixel
xPix8961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[89] VREF PIX_IN[8961] NB2 NB1 CSA_VREF pixel
xPix8962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[89] VREF PIX_IN[8962] NB2 NB1 CSA_VREF pixel
xPix8963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[89] VREF PIX_IN[8963] NB2 NB1 CSA_VREF pixel
xPix8964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[89] VREF PIX_IN[8964] NB2 NB1 CSA_VREF pixel
xPix8965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[89] VREF PIX_IN[8965] NB2 NB1 CSA_VREF pixel
xPix8966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[89] VREF PIX_IN[8966] NB2 NB1 CSA_VREF pixel
xPix8967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[89] VREF PIX_IN[8967] NB2 NB1 CSA_VREF pixel
xPix8968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[89] VREF PIX_IN[8968] NB2 NB1 CSA_VREF pixel
xPix8969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[89] VREF PIX_IN[8969] NB2 NB1 CSA_VREF pixel
xPix8970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[89] VREF PIX_IN[8970] NB2 NB1 CSA_VREF pixel
xPix8971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[89] VREF PIX_IN[8971] NB2 NB1 CSA_VREF pixel
xPix8972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[89] VREF PIX_IN[8972] NB2 NB1 CSA_VREF pixel
xPix8973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[89] VREF PIX_IN[8973] NB2 NB1 CSA_VREF pixel
xPix8974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[89] VREF PIX_IN[8974] NB2 NB1 CSA_VREF pixel
xPix8975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[89] VREF PIX_IN[8975] NB2 NB1 CSA_VREF pixel
xPix8976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[89] VREF PIX_IN[8976] NB2 NB1 CSA_VREF pixel
xPix8977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[89] VREF PIX_IN[8977] NB2 NB1 CSA_VREF pixel
xPix8978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[89] VREF PIX_IN[8978] NB2 NB1 CSA_VREF pixel
xPix8979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[89] VREF PIX_IN[8979] NB2 NB1 CSA_VREF pixel
xPix8980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[89] VREF PIX_IN[8980] NB2 NB1 CSA_VREF pixel
xPix8981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[89] VREF PIX_IN[8981] NB2 NB1 CSA_VREF pixel
xPix8982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[89] VREF PIX_IN[8982] NB2 NB1 CSA_VREF pixel
xPix8983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[89] VREF PIX_IN[8983] NB2 NB1 CSA_VREF pixel
xPix8984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[89] VREF PIX_IN[8984] NB2 NB1 CSA_VREF pixel
xPix8985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[89] VREF PIX_IN[8985] NB2 NB1 CSA_VREF pixel
xPix8986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[89] VREF PIX_IN[8986] NB2 NB1 CSA_VREF pixel
xPix8987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[89] VREF PIX_IN[8987] NB2 NB1 CSA_VREF pixel
xPix8988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[89] VREF PIX_IN[8988] NB2 NB1 CSA_VREF pixel
xPix8989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[89] VREF PIX_IN[8989] NB2 NB1 CSA_VREF pixel
xPix8990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[89] VREF PIX_IN[8990] NB2 NB1 CSA_VREF pixel
xPix8991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[89] VREF PIX_IN[8991] NB2 NB1 CSA_VREF pixel
xPix8992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[89] VREF PIX_IN[8992] NB2 NB1 CSA_VREF pixel
xPix8993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[89] VREF PIX_IN[8993] NB2 NB1 CSA_VREF pixel
xPix8994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[89] VREF PIX_IN[8994] NB2 NB1 CSA_VREF pixel
xPix8995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[89] VREF PIX_IN[8995] NB2 NB1 CSA_VREF pixel
xPix8996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[89] VREF PIX_IN[8996] NB2 NB1 CSA_VREF pixel
xPix8997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[89] VREF PIX_IN[8997] NB2 NB1 CSA_VREF pixel
xPix8998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[89] VREF PIX_IN[8998] NB2 NB1 CSA_VREF pixel
xPix8999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[89] VREF PIX_IN[8999] NB2 NB1 CSA_VREF pixel
xPix9000 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[90] VREF PIX_IN[9000] NB2 NB1 CSA_VREF pixel
xPix9001 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[90] VREF PIX_IN[9001] NB2 NB1 CSA_VREF pixel
xPix9002 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[90] VREF PIX_IN[9002] NB2 NB1 CSA_VREF pixel
xPix9003 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[90] VREF PIX_IN[9003] NB2 NB1 CSA_VREF pixel
xPix9004 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[90] VREF PIX_IN[9004] NB2 NB1 CSA_VREF pixel
xPix9005 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[90] VREF PIX_IN[9005] NB2 NB1 CSA_VREF pixel
xPix9006 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[90] VREF PIX_IN[9006] NB2 NB1 CSA_VREF pixel
xPix9007 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[90] VREF PIX_IN[9007] NB2 NB1 CSA_VREF pixel
xPix9008 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[90] VREF PIX_IN[9008] NB2 NB1 CSA_VREF pixel
xPix9009 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[90] VREF PIX_IN[9009] NB2 NB1 CSA_VREF pixel
xPix9010 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[90] VREF PIX_IN[9010] NB2 NB1 CSA_VREF pixel
xPix9011 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[90] VREF PIX_IN[9011] NB2 NB1 CSA_VREF pixel
xPix9012 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[90] VREF PIX_IN[9012] NB2 NB1 CSA_VREF pixel
xPix9013 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[90] VREF PIX_IN[9013] NB2 NB1 CSA_VREF pixel
xPix9014 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[90] VREF PIX_IN[9014] NB2 NB1 CSA_VREF pixel
xPix9015 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[90] VREF PIX_IN[9015] NB2 NB1 CSA_VREF pixel
xPix9016 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[90] VREF PIX_IN[9016] NB2 NB1 CSA_VREF pixel
xPix9017 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[90] VREF PIX_IN[9017] NB2 NB1 CSA_VREF pixel
xPix9018 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[90] VREF PIX_IN[9018] NB2 NB1 CSA_VREF pixel
xPix9019 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[90] VREF PIX_IN[9019] NB2 NB1 CSA_VREF pixel
xPix9020 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[90] VREF PIX_IN[9020] NB2 NB1 CSA_VREF pixel
xPix9021 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[90] VREF PIX_IN[9021] NB2 NB1 CSA_VREF pixel
xPix9022 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[90] VREF PIX_IN[9022] NB2 NB1 CSA_VREF pixel
xPix9023 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[90] VREF PIX_IN[9023] NB2 NB1 CSA_VREF pixel
xPix9024 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[90] VREF PIX_IN[9024] NB2 NB1 CSA_VREF pixel
xPix9025 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[90] VREF PIX_IN[9025] NB2 NB1 CSA_VREF pixel
xPix9026 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[90] VREF PIX_IN[9026] NB2 NB1 CSA_VREF pixel
xPix9027 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[90] VREF PIX_IN[9027] NB2 NB1 CSA_VREF pixel
xPix9028 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[90] VREF PIX_IN[9028] NB2 NB1 CSA_VREF pixel
xPix9029 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[90] VREF PIX_IN[9029] NB2 NB1 CSA_VREF pixel
xPix9030 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[90] VREF PIX_IN[9030] NB2 NB1 CSA_VREF pixel
xPix9031 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[90] VREF PIX_IN[9031] NB2 NB1 CSA_VREF pixel
xPix9032 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[90] VREF PIX_IN[9032] NB2 NB1 CSA_VREF pixel
xPix9033 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[90] VREF PIX_IN[9033] NB2 NB1 CSA_VREF pixel
xPix9034 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[90] VREF PIX_IN[9034] NB2 NB1 CSA_VREF pixel
xPix9035 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[90] VREF PIX_IN[9035] NB2 NB1 CSA_VREF pixel
xPix9036 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[90] VREF PIX_IN[9036] NB2 NB1 CSA_VREF pixel
xPix9037 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[90] VREF PIX_IN[9037] NB2 NB1 CSA_VREF pixel
xPix9038 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[90] VREF PIX_IN[9038] NB2 NB1 CSA_VREF pixel
xPix9039 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[90] VREF PIX_IN[9039] NB2 NB1 CSA_VREF pixel
xPix9040 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[90] VREF PIX_IN[9040] NB2 NB1 CSA_VREF pixel
xPix9041 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[90] VREF PIX_IN[9041] NB2 NB1 CSA_VREF pixel
xPix9042 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[90] VREF PIX_IN[9042] NB2 NB1 CSA_VREF pixel
xPix9043 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[90] VREF PIX_IN[9043] NB2 NB1 CSA_VREF pixel
xPix9044 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[90] VREF PIX_IN[9044] NB2 NB1 CSA_VREF pixel
xPix9045 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[90] VREF PIX_IN[9045] NB2 NB1 CSA_VREF pixel
xPix9046 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[90] VREF PIX_IN[9046] NB2 NB1 CSA_VREF pixel
xPix9047 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[90] VREF PIX_IN[9047] NB2 NB1 CSA_VREF pixel
xPix9048 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[90] VREF PIX_IN[9048] NB2 NB1 CSA_VREF pixel
xPix9049 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[90] VREF PIX_IN[9049] NB2 NB1 CSA_VREF pixel
xPix9050 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[90] VREF PIX_IN[9050] NB2 NB1 CSA_VREF pixel
xPix9051 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[90] VREF PIX_IN[9051] NB2 NB1 CSA_VREF pixel
xPix9052 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[90] VREF PIX_IN[9052] NB2 NB1 CSA_VREF pixel
xPix9053 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[90] VREF PIX_IN[9053] NB2 NB1 CSA_VREF pixel
xPix9054 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[90] VREF PIX_IN[9054] NB2 NB1 CSA_VREF pixel
xPix9055 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[90] VREF PIX_IN[9055] NB2 NB1 CSA_VREF pixel
xPix9056 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[90] VREF PIX_IN[9056] NB2 NB1 CSA_VREF pixel
xPix9057 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[90] VREF PIX_IN[9057] NB2 NB1 CSA_VREF pixel
xPix9058 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[90] VREF PIX_IN[9058] NB2 NB1 CSA_VREF pixel
xPix9059 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[90] VREF PIX_IN[9059] NB2 NB1 CSA_VREF pixel
xPix9060 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[90] VREF PIX_IN[9060] NB2 NB1 CSA_VREF pixel
xPix9061 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[90] VREF PIX_IN[9061] NB2 NB1 CSA_VREF pixel
xPix9062 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[90] VREF PIX_IN[9062] NB2 NB1 CSA_VREF pixel
xPix9063 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[90] VREF PIX_IN[9063] NB2 NB1 CSA_VREF pixel
xPix9064 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[90] VREF PIX_IN[9064] NB2 NB1 CSA_VREF pixel
xPix9065 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[90] VREF PIX_IN[9065] NB2 NB1 CSA_VREF pixel
xPix9066 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[90] VREF PIX_IN[9066] NB2 NB1 CSA_VREF pixel
xPix9067 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[90] VREF PIX_IN[9067] NB2 NB1 CSA_VREF pixel
xPix9068 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[90] VREF PIX_IN[9068] NB2 NB1 CSA_VREF pixel
xPix9069 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[90] VREF PIX_IN[9069] NB2 NB1 CSA_VREF pixel
xPix9070 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[90] VREF PIX_IN[9070] NB2 NB1 CSA_VREF pixel
xPix9071 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[90] VREF PIX_IN[9071] NB2 NB1 CSA_VREF pixel
xPix9072 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[90] VREF PIX_IN[9072] NB2 NB1 CSA_VREF pixel
xPix9073 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[90] VREF PIX_IN[9073] NB2 NB1 CSA_VREF pixel
xPix9074 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[90] VREF PIX_IN[9074] NB2 NB1 CSA_VREF pixel
xPix9075 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[90] VREF PIX_IN[9075] NB2 NB1 CSA_VREF pixel
xPix9076 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[90] VREF PIX_IN[9076] NB2 NB1 CSA_VREF pixel
xPix9077 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[90] VREF PIX_IN[9077] NB2 NB1 CSA_VREF pixel
xPix9078 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[90] VREF PIX_IN[9078] NB2 NB1 CSA_VREF pixel
xPix9079 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[90] VREF PIX_IN[9079] NB2 NB1 CSA_VREF pixel
xPix9080 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[90] VREF PIX_IN[9080] NB2 NB1 CSA_VREF pixel
xPix9081 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[90] VREF PIX_IN[9081] NB2 NB1 CSA_VREF pixel
xPix9082 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[90] VREF PIX_IN[9082] NB2 NB1 CSA_VREF pixel
xPix9083 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[90] VREF PIX_IN[9083] NB2 NB1 CSA_VREF pixel
xPix9084 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[90] VREF PIX_IN[9084] NB2 NB1 CSA_VREF pixel
xPix9085 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[90] VREF PIX_IN[9085] NB2 NB1 CSA_VREF pixel
xPix9086 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[90] VREF PIX_IN[9086] NB2 NB1 CSA_VREF pixel
xPix9087 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[90] VREF PIX_IN[9087] NB2 NB1 CSA_VREF pixel
xPix9088 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[90] VREF PIX_IN[9088] NB2 NB1 CSA_VREF pixel
xPix9089 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[90] VREF PIX_IN[9089] NB2 NB1 CSA_VREF pixel
xPix9090 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[90] VREF PIX_IN[9090] NB2 NB1 CSA_VREF pixel
xPix9091 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[90] VREF PIX_IN[9091] NB2 NB1 CSA_VREF pixel
xPix9092 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[90] VREF PIX_IN[9092] NB2 NB1 CSA_VREF pixel
xPix9093 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[90] VREF PIX_IN[9093] NB2 NB1 CSA_VREF pixel
xPix9094 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[90] VREF PIX_IN[9094] NB2 NB1 CSA_VREF pixel
xPix9095 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[90] VREF PIX_IN[9095] NB2 NB1 CSA_VREF pixel
xPix9096 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[90] VREF PIX_IN[9096] NB2 NB1 CSA_VREF pixel
xPix9097 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[90] VREF PIX_IN[9097] NB2 NB1 CSA_VREF pixel
xPix9098 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[90] VREF PIX_IN[9098] NB2 NB1 CSA_VREF pixel
xPix9099 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[90] VREF PIX_IN[9099] NB2 NB1 CSA_VREF pixel
xPix9100 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[91] VREF PIX_IN[9100] NB2 NB1 CSA_VREF pixel
xPix9101 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[91] VREF PIX_IN[9101] NB2 NB1 CSA_VREF pixel
xPix9102 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[91] VREF PIX_IN[9102] NB2 NB1 CSA_VREF pixel
xPix9103 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[91] VREF PIX_IN[9103] NB2 NB1 CSA_VREF pixel
xPix9104 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[91] VREF PIX_IN[9104] NB2 NB1 CSA_VREF pixel
xPix9105 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[91] VREF PIX_IN[9105] NB2 NB1 CSA_VREF pixel
xPix9106 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[91] VREF PIX_IN[9106] NB2 NB1 CSA_VREF pixel
xPix9107 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[91] VREF PIX_IN[9107] NB2 NB1 CSA_VREF pixel
xPix9108 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[91] VREF PIX_IN[9108] NB2 NB1 CSA_VREF pixel
xPix9109 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[91] VREF PIX_IN[9109] NB2 NB1 CSA_VREF pixel
xPix9110 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[91] VREF PIX_IN[9110] NB2 NB1 CSA_VREF pixel
xPix9111 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[91] VREF PIX_IN[9111] NB2 NB1 CSA_VREF pixel
xPix9112 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[91] VREF PIX_IN[9112] NB2 NB1 CSA_VREF pixel
xPix9113 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[91] VREF PIX_IN[9113] NB2 NB1 CSA_VREF pixel
xPix9114 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[91] VREF PIX_IN[9114] NB2 NB1 CSA_VREF pixel
xPix9115 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[91] VREF PIX_IN[9115] NB2 NB1 CSA_VREF pixel
xPix9116 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[91] VREF PIX_IN[9116] NB2 NB1 CSA_VREF pixel
xPix9117 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[91] VREF PIX_IN[9117] NB2 NB1 CSA_VREF pixel
xPix9118 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[91] VREF PIX_IN[9118] NB2 NB1 CSA_VREF pixel
xPix9119 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[91] VREF PIX_IN[9119] NB2 NB1 CSA_VREF pixel
xPix9120 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[91] VREF PIX_IN[9120] NB2 NB1 CSA_VREF pixel
xPix9121 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[91] VREF PIX_IN[9121] NB2 NB1 CSA_VREF pixel
xPix9122 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[91] VREF PIX_IN[9122] NB2 NB1 CSA_VREF pixel
xPix9123 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[91] VREF PIX_IN[9123] NB2 NB1 CSA_VREF pixel
xPix9124 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[91] VREF PIX_IN[9124] NB2 NB1 CSA_VREF pixel
xPix9125 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[91] VREF PIX_IN[9125] NB2 NB1 CSA_VREF pixel
xPix9126 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[91] VREF PIX_IN[9126] NB2 NB1 CSA_VREF pixel
xPix9127 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[91] VREF PIX_IN[9127] NB2 NB1 CSA_VREF pixel
xPix9128 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[91] VREF PIX_IN[9128] NB2 NB1 CSA_VREF pixel
xPix9129 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[91] VREF PIX_IN[9129] NB2 NB1 CSA_VREF pixel
xPix9130 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[91] VREF PIX_IN[9130] NB2 NB1 CSA_VREF pixel
xPix9131 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[91] VREF PIX_IN[9131] NB2 NB1 CSA_VREF pixel
xPix9132 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[91] VREF PIX_IN[9132] NB2 NB1 CSA_VREF pixel
xPix9133 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[91] VREF PIX_IN[9133] NB2 NB1 CSA_VREF pixel
xPix9134 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[91] VREF PIX_IN[9134] NB2 NB1 CSA_VREF pixel
xPix9135 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[91] VREF PIX_IN[9135] NB2 NB1 CSA_VREF pixel
xPix9136 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[91] VREF PIX_IN[9136] NB2 NB1 CSA_VREF pixel
xPix9137 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[91] VREF PIX_IN[9137] NB2 NB1 CSA_VREF pixel
xPix9138 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[91] VREF PIX_IN[9138] NB2 NB1 CSA_VREF pixel
xPix9139 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[91] VREF PIX_IN[9139] NB2 NB1 CSA_VREF pixel
xPix9140 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[91] VREF PIX_IN[9140] NB2 NB1 CSA_VREF pixel
xPix9141 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[91] VREF PIX_IN[9141] NB2 NB1 CSA_VREF pixel
xPix9142 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[91] VREF PIX_IN[9142] NB2 NB1 CSA_VREF pixel
xPix9143 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[91] VREF PIX_IN[9143] NB2 NB1 CSA_VREF pixel
xPix9144 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[91] VREF PIX_IN[9144] NB2 NB1 CSA_VREF pixel
xPix9145 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[91] VREF PIX_IN[9145] NB2 NB1 CSA_VREF pixel
xPix9146 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[91] VREF PIX_IN[9146] NB2 NB1 CSA_VREF pixel
xPix9147 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[91] VREF PIX_IN[9147] NB2 NB1 CSA_VREF pixel
xPix9148 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[91] VREF PIX_IN[9148] NB2 NB1 CSA_VREF pixel
xPix9149 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[91] VREF PIX_IN[9149] NB2 NB1 CSA_VREF pixel
xPix9150 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[91] VREF PIX_IN[9150] NB2 NB1 CSA_VREF pixel
xPix9151 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[91] VREF PIX_IN[9151] NB2 NB1 CSA_VREF pixel
xPix9152 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[91] VREF PIX_IN[9152] NB2 NB1 CSA_VREF pixel
xPix9153 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[91] VREF PIX_IN[9153] NB2 NB1 CSA_VREF pixel
xPix9154 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[91] VREF PIX_IN[9154] NB2 NB1 CSA_VREF pixel
xPix9155 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[91] VREF PIX_IN[9155] NB2 NB1 CSA_VREF pixel
xPix9156 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[91] VREF PIX_IN[9156] NB2 NB1 CSA_VREF pixel
xPix9157 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[91] VREF PIX_IN[9157] NB2 NB1 CSA_VREF pixel
xPix9158 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[91] VREF PIX_IN[9158] NB2 NB1 CSA_VREF pixel
xPix9159 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[91] VREF PIX_IN[9159] NB2 NB1 CSA_VREF pixel
xPix9160 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[91] VREF PIX_IN[9160] NB2 NB1 CSA_VREF pixel
xPix9161 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[91] VREF PIX_IN[9161] NB2 NB1 CSA_VREF pixel
xPix9162 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[91] VREF PIX_IN[9162] NB2 NB1 CSA_VREF pixel
xPix9163 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[91] VREF PIX_IN[9163] NB2 NB1 CSA_VREF pixel
xPix9164 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[91] VREF PIX_IN[9164] NB2 NB1 CSA_VREF pixel
xPix9165 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[91] VREF PIX_IN[9165] NB2 NB1 CSA_VREF pixel
xPix9166 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[91] VREF PIX_IN[9166] NB2 NB1 CSA_VREF pixel
xPix9167 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[91] VREF PIX_IN[9167] NB2 NB1 CSA_VREF pixel
xPix9168 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[91] VREF PIX_IN[9168] NB2 NB1 CSA_VREF pixel
xPix9169 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[91] VREF PIX_IN[9169] NB2 NB1 CSA_VREF pixel
xPix9170 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[91] VREF PIX_IN[9170] NB2 NB1 CSA_VREF pixel
xPix9171 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[91] VREF PIX_IN[9171] NB2 NB1 CSA_VREF pixel
xPix9172 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[91] VREF PIX_IN[9172] NB2 NB1 CSA_VREF pixel
xPix9173 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[91] VREF PIX_IN[9173] NB2 NB1 CSA_VREF pixel
xPix9174 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[91] VREF PIX_IN[9174] NB2 NB1 CSA_VREF pixel
xPix9175 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[91] VREF PIX_IN[9175] NB2 NB1 CSA_VREF pixel
xPix9176 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[91] VREF PIX_IN[9176] NB2 NB1 CSA_VREF pixel
xPix9177 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[91] VREF PIX_IN[9177] NB2 NB1 CSA_VREF pixel
xPix9178 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[91] VREF PIX_IN[9178] NB2 NB1 CSA_VREF pixel
xPix9179 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[91] VREF PIX_IN[9179] NB2 NB1 CSA_VREF pixel
xPix9180 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[91] VREF PIX_IN[9180] NB2 NB1 CSA_VREF pixel
xPix9181 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[91] VREF PIX_IN[9181] NB2 NB1 CSA_VREF pixel
xPix9182 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[91] VREF PIX_IN[9182] NB2 NB1 CSA_VREF pixel
xPix9183 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[91] VREF PIX_IN[9183] NB2 NB1 CSA_VREF pixel
xPix9184 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[91] VREF PIX_IN[9184] NB2 NB1 CSA_VREF pixel
xPix9185 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[91] VREF PIX_IN[9185] NB2 NB1 CSA_VREF pixel
xPix9186 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[91] VREF PIX_IN[9186] NB2 NB1 CSA_VREF pixel
xPix9187 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[91] VREF PIX_IN[9187] NB2 NB1 CSA_VREF pixel
xPix9188 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[91] VREF PIX_IN[9188] NB2 NB1 CSA_VREF pixel
xPix9189 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[91] VREF PIX_IN[9189] NB2 NB1 CSA_VREF pixel
xPix9190 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[91] VREF PIX_IN[9190] NB2 NB1 CSA_VREF pixel
xPix9191 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[91] VREF PIX_IN[9191] NB2 NB1 CSA_VREF pixel
xPix9192 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[91] VREF PIX_IN[9192] NB2 NB1 CSA_VREF pixel
xPix9193 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[91] VREF PIX_IN[9193] NB2 NB1 CSA_VREF pixel
xPix9194 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[91] VREF PIX_IN[9194] NB2 NB1 CSA_VREF pixel
xPix9195 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[91] VREF PIX_IN[9195] NB2 NB1 CSA_VREF pixel
xPix9196 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[91] VREF PIX_IN[9196] NB2 NB1 CSA_VREF pixel
xPix9197 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[91] VREF PIX_IN[9197] NB2 NB1 CSA_VREF pixel
xPix9198 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[91] VREF PIX_IN[9198] NB2 NB1 CSA_VREF pixel
xPix9199 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[91] VREF PIX_IN[9199] NB2 NB1 CSA_VREF pixel
xPix9200 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[92] VREF PIX_IN[9200] NB2 NB1 CSA_VREF pixel
xPix9201 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[92] VREF PIX_IN[9201] NB2 NB1 CSA_VREF pixel
xPix9202 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[92] VREF PIX_IN[9202] NB2 NB1 CSA_VREF pixel
xPix9203 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[92] VREF PIX_IN[9203] NB2 NB1 CSA_VREF pixel
xPix9204 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[92] VREF PIX_IN[9204] NB2 NB1 CSA_VREF pixel
xPix9205 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[92] VREF PIX_IN[9205] NB2 NB1 CSA_VREF pixel
xPix9206 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[92] VREF PIX_IN[9206] NB2 NB1 CSA_VREF pixel
xPix9207 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[92] VREF PIX_IN[9207] NB2 NB1 CSA_VREF pixel
xPix9208 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[92] VREF PIX_IN[9208] NB2 NB1 CSA_VREF pixel
xPix9209 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[92] VREF PIX_IN[9209] NB2 NB1 CSA_VREF pixel
xPix9210 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[92] VREF PIX_IN[9210] NB2 NB1 CSA_VREF pixel
xPix9211 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[92] VREF PIX_IN[9211] NB2 NB1 CSA_VREF pixel
xPix9212 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[92] VREF PIX_IN[9212] NB2 NB1 CSA_VREF pixel
xPix9213 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[92] VREF PIX_IN[9213] NB2 NB1 CSA_VREF pixel
xPix9214 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[92] VREF PIX_IN[9214] NB2 NB1 CSA_VREF pixel
xPix9215 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[92] VREF PIX_IN[9215] NB2 NB1 CSA_VREF pixel
xPix9216 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[92] VREF PIX_IN[9216] NB2 NB1 CSA_VREF pixel
xPix9217 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[92] VREF PIX_IN[9217] NB2 NB1 CSA_VREF pixel
xPix9218 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[92] VREF PIX_IN[9218] NB2 NB1 CSA_VREF pixel
xPix9219 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[92] VREF PIX_IN[9219] NB2 NB1 CSA_VREF pixel
xPix9220 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[92] VREF PIX_IN[9220] NB2 NB1 CSA_VREF pixel
xPix9221 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[92] VREF PIX_IN[9221] NB2 NB1 CSA_VREF pixel
xPix9222 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[92] VREF PIX_IN[9222] NB2 NB1 CSA_VREF pixel
xPix9223 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[92] VREF PIX_IN[9223] NB2 NB1 CSA_VREF pixel
xPix9224 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[92] VREF PIX_IN[9224] NB2 NB1 CSA_VREF pixel
xPix9225 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[92] VREF PIX_IN[9225] NB2 NB1 CSA_VREF pixel
xPix9226 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[92] VREF PIX_IN[9226] NB2 NB1 CSA_VREF pixel
xPix9227 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[92] VREF PIX_IN[9227] NB2 NB1 CSA_VREF pixel
xPix9228 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[92] VREF PIX_IN[9228] NB2 NB1 CSA_VREF pixel
xPix9229 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[92] VREF PIX_IN[9229] NB2 NB1 CSA_VREF pixel
xPix9230 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[92] VREF PIX_IN[9230] NB2 NB1 CSA_VREF pixel
xPix9231 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[92] VREF PIX_IN[9231] NB2 NB1 CSA_VREF pixel
xPix9232 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[92] VREF PIX_IN[9232] NB2 NB1 CSA_VREF pixel
xPix9233 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[92] VREF PIX_IN[9233] NB2 NB1 CSA_VREF pixel
xPix9234 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[92] VREF PIX_IN[9234] NB2 NB1 CSA_VREF pixel
xPix9235 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[92] VREF PIX_IN[9235] NB2 NB1 CSA_VREF pixel
xPix9236 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[92] VREF PIX_IN[9236] NB2 NB1 CSA_VREF pixel
xPix9237 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[92] VREF PIX_IN[9237] NB2 NB1 CSA_VREF pixel
xPix9238 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[92] VREF PIX_IN[9238] NB2 NB1 CSA_VREF pixel
xPix9239 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[92] VREF PIX_IN[9239] NB2 NB1 CSA_VREF pixel
xPix9240 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[92] VREF PIX_IN[9240] NB2 NB1 CSA_VREF pixel
xPix9241 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[92] VREF PIX_IN[9241] NB2 NB1 CSA_VREF pixel
xPix9242 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[92] VREF PIX_IN[9242] NB2 NB1 CSA_VREF pixel
xPix9243 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[92] VREF PIX_IN[9243] NB2 NB1 CSA_VREF pixel
xPix9244 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[92] VREF PIX_IN[9244] NB2 NB1 CSA_VREF pixel
xPix9245 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[92] VREF PIX_IN[9245] NB2 NB1 CSA_VREF pixel
xPix9246 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[92] VREF PIX_IN[9246] NB2 NB1 CSA_VREF pixel
xPix9247 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[92] VREF PIX_IN[9247] NB2 NB1 CSA_VREF pixel
xPix9248 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[92] VREF PIX_IN[9248] NB2 NB1 CSA_VREF pixel
xPix9249 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[92] VREF PIX_IN[9249] NB2 NB1 CSA_VREF pixel
xPix9250 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[92] VREF PIX_IN[9250] NB2 NB1 CSA_VREF pixel
xPix9251 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[92] VREF PIX_IN[9251] NB2 NB1 CSA_VREF pixel
xPix9252 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[92] VREF PIX_IN[9252] NB2 NB1 CSA_VREF pixel
xPix9253 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[92] VREF PIX_IN[9253] NB2 NB1 CSA_VREF pixel
xPix9254 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[92] VREF PIX_IN[9254] NB2 NB1 CSA_VREF pixel
xPix9255 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[92] VREF PIX_IN[9255] NB2 NB1 CSA_VREF pixel
xPix9256 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[92] VREF PIX_IN[9256] NB2 NB1 CSA_VREF pixel
xPix9257 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[92] VREF PIX_IN[9257] NB2 NB1 CSA_VREF pixel
xPix9258 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[92] VREF PIX_IN[9258] NB2 NB1 CSA_VREF pixel
xPix9259 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[92] VREF PIX_IN[9259] NB2 NB1 CSA_VREF pixel
xPix9260 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[92] VREF PIX_IN[9260] NB2 NB1 CSA_VREF pixel
xPix9261 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[92] VREF PIX_IN[9261] NB2 NB1 CSA_VREF pixel
xPix9262 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[92] VREF PIX_IN[9262] NB2 NB1 CSA_VREF pixel
xPix9263 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[92] VREF PIX_IN[9263] NB2 NB1 CSA_VREF pixel
xPix9264 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[92] VREF PIX_IN[9264] NB2 NB1 CSA_VREF pixel
xPix9265 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[92] VREF PIX_IN[9265] NB2 NB1 CSA_VREF pixel
xPix9266 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[92] VREF PIX_IN[9266] NB2 NB1 CSA_VREF pixel
xPix9267 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[92] VREF PIX_IN[9267] NB2 NB1 CSA_VREF pixel
xPix9268 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[92] VREF PIX_IN[9268] NB2 NB1 CSA_VREF pixel
xPix9269 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[92] VREF PIX_IN[9269] NB2 NB1 CSA_VREF pixel
xPix9270 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[92] VREF PIX_IN[9270] NB2 NB1 CSA_VREF pixel
xPix9271 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[92] VREF PIX_IN[9271] NB2 NB1 CSA_VREF pixel
xPix9272 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[92] VREF PIX_IN[9272] NB2 NB1 CSA_VREF pixel
xPix9273 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[92] VREF PIX_IN[9273] NB2 NB1 CSA_VREF pixel
xPix9274 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[92] VREF PIX_IN[9274] NB2 NB1 CSA_VREF pixel
xPix9275 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[92] VREF PIX_IN[9275] NB2 NB1 CSA_VREF pixel
xPix9276 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[92] VREF PIX_IN[9276] NB2 NB1 CSA_VREF pixel
xPix9277 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[92] VREF PIX_IN[9277] NB2 NB1 CSA_VREF pixel
xPix9278 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[92] VREF PIX_IN[9278] NB2 NB1 CSA_VREF pixel
xPix9279 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[92] VREF PIX_IN[9279] NB2 NB1 CSA_VREF pixel
xPix9280 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[92] VREF PIX_IN[9280] NB2 NB1 CSA_VREF pixel
xPix9281 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[92] VREF PIX_IN[9281] NB2 NB1 CSA_VREF pixel
xPix9282 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[92] VREF PIX_IN[9282] NB2 NB1 CSA_VREF pixel
xPix9283 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[92] VREF PIX_IN[9283] NB2 NB1 CSA_VREF pixel
xPix9284 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[92] VREF PIX_IN[9284] NB2 NB1 CSA_VREF pixel
xPix9285 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[92] VREF PIX_IN[9285] NB2 NB1 CSA_VREF pixel
xPix9286 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[92] VREF PIX_IN[9286] NB2 NB1 CSA_VREF pixel
xPix9287 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[92] VREF PIX_IN[9287] NB2 NB1 CSA_VREF pixel
xPix9288 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[92] VREF PIX_IN[9288] NB2 NB1 CSA_VREF pixel
xPix9289 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[92] VREF PIX_IN[9289] NB2 NB1 CSA_VREF pixel
xPix9290 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[92] VREF PIX_IN[9290] NB2 NB1 CSA_VREF pixel
xPix9291 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[92] VREF PIX_IN[9291] NB2 NB1 CSA_VREF pixel
xPix9292 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[92] VREF PIX_IN[9292] NB2 NB1 CSA_VREF pixel
xPix9293 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[92] VREF PIX_IN[9293] NB2 NB1 CSA_VREF pixel
xPix9294 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[92] VREF PIX_IN[9294] NB2 NB1 CSA_VREF pixel
xPix9295 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[92] VREF PIX_IN[9295] NB2 NB1 CSA_VREF pixel
xPix9296 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[92] VREF PIX_IN[9296] NB2 NB1 CSA_VREF pixel
xPix9297 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[92] VREF PIX_IN[9297] NB2 NB1 CSA_VREF pixel
xPix9298 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[92] VREF PIX_IN[9298] NB2 NB1 CSA_VREF pixel
xPix9299 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[92] VREF PIX_IN[9299] NB2 NB1 CSA_VREF pixel
xPix9300 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[93] VREF PIX_IN[9300] NB2 NB1 CSA_VREF pixel
xPix9301 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[93] VREF PIX_IN[9301] NB2 NB1 CSA_VREF pixel
xPix9302 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[93] VREF PIX_IN[9302] NB2 NB1 CSA_VREF pixel
xPix9303 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[93] VREF PIX_IN[9303] NB2 NB1 CSA_VREF pixel
xPix9304 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[93] VREF PIX_IN[9304] NB2 NB1 CSA_VREF pixel
xPix9305 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[93] VREF PIX_IN[9305] NB2 NB1 CSA_VREF pixel
xPix9306 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[93] VREF PIX_IN[9306] NB2 NB1 CSA_VREF pixel
xPix9307 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[93] VREF PIX_IN[9307] NB2 NB1 CSA_VREF pixel
xPix9308 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[93] VREF PIX_IN[9308] NB2 NB1 CSA_VREF pixel
xPix9309 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[93] VREF PIX_IN[9309] NB2 NB1 CSA_VREF pixel
xPix9310 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[93] VREF PIX_IN[9310] NB2 NB1 CSA_VREF pixel
xPix9311 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[93] VREF PIX_IN[9311] NB2 NB1 CSA_VREF pixel
xPix9312 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[93] VREF PIX_IN[9312] NB2 NB1 CSA_VREF pixel
xPix9313 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[93] VREF PIX_IN[9313] NB2 NB1 CSA_VREF pixel
xPix9314 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[93] VREF PIX_IN[9314] NB2 NB1 CSA_VREF pixel
xPix9315 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[93] VREF PIX_IN[9315] NB2 NB1 CSA_VREF pixel
xPix9316 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[93] VREF PIX_IN[9316] NB2 NB1 CSA_VREF pixel
xPix9317 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[93] VREF PIX_IN[9317] NB2 NB1 CSA_VREF pixel
xPix9318 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[93] VREF PIX_IN[9318] NB2 NB1 CSA_VREF pixel
xPix9319 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[93] VREF PIX_IN[9319] NB2 NB1 CSA_VREF pixel
xPix9320 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[93] VREF PIX_IN[9320] NB2 NB1 CSA_VREF pixel
xPix9321 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[93] VREF PIX_IN[9321] NB2 NB1 CSA_VREF pixel
xPix9322 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[93] VREF PIX_IN[9322] NB2 NB1 CSA_VREF pixel
xPix9323 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[93] VREF PIX_IN[9323] NB2 NB1 CSA_VREF pixel
xPix9324 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[93] VREF PIX_IN[9324] NB2 NB1 CSA_VREF pixel
xPix9325 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[93] VREF PIX_IN[9325] NB2 NB1 CSA_VREF pixel
xPix9326 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[93] VREF PIX_IN[9326] NB2 NB1 CSA_VREF pixel
xPix9327 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[93] VREF PIX_IN[9327] NB2 NB1 CSA_VREF pixel
xPix9328 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[93] VREF PIX_IN[9328] NB2 NB1 CSA_VREF pixel
xPix9329 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[93] VREF PIX_IN[9329] NB2 NB1 CSA_VREF pixel
xPix9330 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[93] VREF PIX_IN[9330] NB2 NB1 CSA_VREF pixel
xPix9331 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[93] VREF PIX_IN[9331] NB2 NB1 CSA_VREF pixel
xPix9332 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[93] VREF PIX_IN[9332] NB2 NB1 CSA_VREF pixel
xPix9333 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[93] VREF PIX_IN[9333] NB2 NB1 CSA_VREF pixel
xPix9334 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[93] VREF PIX_IN[9334] NB2 NB1 CSA_VREF pixel
xPix9335 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[93] VREF PIX_IN[9335] NB2 NB1 CSA_VREF pixel
xPix9336 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[93] VREF PIX_IN[9336] NB2 NB1 CSA_VREF pixel
xPix9337 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[93] VREF PIX_IN[9337] NB2 NB1 CSA_VREF pixel
xPix9338 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[93] VREF PIX_IN[9338] NB2 NB1 CSA_VREF pixel
xPix9339 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[93] VREF PIX_IN[9339] NB2 NB1 CSA_VREF pixel
xPix9340 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[93] VREF PIX_IN[9340] NB2 NB1 CSA_VREF pixel
xPix9341 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[93] VREF PIX_IN[9341] NB2 NB1 CSA_VREF pixel
xPix9342 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[93] VREF PIX_IN[9342] NB2 NB1 CSA_VREF pixel
xPix9343 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[93] VREF PIX_IN[9343] NB2 NB1 CSA_VREF pixel
xPix9344 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[93] VREF PIX_IN[9344] NB2 NB1 CSA_VREF pixel
xPix9345 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[93] VREF PIX_IN[9345] NB2 NB1 CSA_VREF pixel
xPix9346 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[93] VREF PIX_IN[9346] NB2 NB1 CSA_VREF pixel
xPix9347 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[93] VREF PIX_IN[9347] NB2 NB1 CSA_VREF pixel
xPix9348 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[93] VREF PIX_IN[9348] NB2 NB1 CSA_VREF pixel
xPix9349 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[93] VREF PIX_IN[9349] NB2 NB1 CSA_VREF pixel
xPix9350 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[93] VREF PIX_IN[9350] NB2 NB1 CSA_VREF pixel
xPix9351 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[93] VREF PIX_IN[9351] NB2 NB1 CSA_VREF pixel
xPix9352 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[93] VREF PIX_IN[9352] NB2 NB1 CSA_VREF pixel
xPix9353 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[93] VREF PIX_IN[9353] NB2 NB1 CSA_VREF pixel
xPix9354 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[93] VREF PIX_IN[9354] NB2 NB1 CSA_VREF pixel
xPix9355 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[93] VREF PIX_IN[9355] NB2 NB1 CSA_VREF pixel
xPix9356 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[93] VREF PIX_IN[9356] NB2 NB1 CSA_VREF pixel
xPix9357 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[93] VREF PIX_IN[9357] NB2 NB1 CSA_VREF pixel
xPix9358 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[93] VREF PIX_IN[9358] NB2 NB1 CSA_VREF pixel
xPix9359 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[93] VREF PIX_IN[9359] NB2 NB1 CSA_VREF pixel
xPix9360 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[93] VREF PIX_IN[9360] NB2 NB1 CSA_VREF pixel
xPix9361 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[93] VREF PIX_IN[9361] NB2 NB1 CSA_VREF pixel
xPix9362 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[93] VREF PIX_IN[9362] NB2 NB1 CSA_VREF pixel
xPix9363 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[93] VREF PIX_IN[9363] NB2 NB1 CSA_VREF pixel
xPix9364 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[93] VREF PIX_IN[9364] NB2 NB1 CSA_VREF pixel
xPix9365 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[93] VREF PIX_IN[9365] NB2 NB1 CSA_VREF pixel
xPix9366 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[93] VREF PIX_IN[9366] NB2 NB1 CSA_VREF pixel
xPix9367 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[93] VREF PIX_IN[9367] NB2 NB1 CSA_VREF pixel
xPix9368 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[93] VREF PIX_IN[9368] NB2 NB1 CSA_VREF pixel
xPix9369 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[93] VREF PIX_IN[9369] NB2 NB1 CSA_VREF pixel
xPix9370 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[93] VREF PIX_IN[9370] NB2 NB1 CSA_VREF pixel
xPix9371 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[93] VREF PIX_IN[9371] NB2 NB1 CSA_VREF pixel
xPix9372 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[93] VREF PIX_IN[9372] NB2 NB1 CSA_VREF pixel
xPix9373 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[93] VREF PIX_IN[9373] NB2 NB1 CSA_VREF pixel
xPix9374 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[93] VREF PIX_IN[9374] NB2 NB1 CSA_VREF pixel
xPix9375 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[93] VREF PIX_IN[9375] NB2 NB1 CSA_VREF pixel
xPix9376 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[93] VREF PIX_IN[9376] NB2 NB1 CSA_VREF pixel
xPix9377 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[93] VREF PIX_IN[9377] NB2 NB1 CSA_VREF pixel
xPix9378 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[93] VREF PIX_IN[9378] NB2 NB1 CSA_VREF pixel
xPix9379 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[93] VREF PIX_IN[9379] NB2 NB1 CSA_VREF pixel
xPix9380 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[93] VREF PIX_IN[9380] NB2 NB1 CSA_VREF pixel
xPix9381 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[93] VREF PIX_IN[9381] NB2 NB1 CSA_VREF pixel
xPix9382 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[93] VREF PIX_IN[9382] NB2 NB1 CSA_VREF pixel
xPix9383 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[93] VREF PIX_IN[9383] NB2 NB1 CSA_VREF pixel
xPix9384 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[93] VREF PIX_IN[9384] NB2 NB1 CSA_VREF pixel
xPix9385 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[93] VREF PIX_IN[9385] NB2 NB1 CSA_VREF pixel
xPix9386 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[93] VREF PIX_IN[9386] NB2 NB1 CSA_VREF pixel
xPix9387 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[93] VREF PIX_IN[9387] NB2 NB1 CSA_VREF pixel
xPix9388 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[93] VREF PIX_IN[9388] NB2 NB1 CSA_VREF pixel
xPix9389 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[93] VREF PIX_IN[9389] NB2 NB1 CSA_VREF pixel
xPix9390 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[93] VREF PIX_IN[9390] NB2 NB1 CSA_VREF pixel
xPix9391 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[93] VREF PIX_IN[9391] NB2 NB1 CSA_VREF pixel
xPix9392 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[93] VREF PIX_IN[9392] NB2 NB1 CSA_VREF pixel
xPix9393 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[93] VREF PIX_IN[9393] NB2 NB1 CSA_VREF pixel
xPix9394 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[93] VREF PIX_IN[9394] NB2 NB1 CSA_VREF pixel
xPix9395 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[93] VREF PIX_IN[9395] NB2 NB1 CSA_VREF pixel
xPix9396 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[93] VREF PIX_IN[9396] NB2 NB1 CSA_VREF pixel
xPix9397 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[93] VREF PIX_IN[9397] NB2 NB1 CSA_VREF pixel
xPix9398 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[93] VREF PIX_IN[9398] NB2 NB1 CSA_VREF pixel
xPix9399 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[93] VREF PIX_IN[9399] NB2 NB1 CSA_VREF pixel
xPix9400 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[94] VREF PIX_IN[9400] NB2 NB1 CSA_VREF pixel
xPix9401 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[94] VREF PIX_IN[9401] NB2 NB1 CSA_VREF pixel
xPix9402 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[94] VREF PIX_IN[9402] NB2 NB1 CSA_VREF pixel
xPix9403 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[94] VREF PIX_IN[9403] NB2 NB1 CSA_VREF pixel
xPix9404 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[94] VREF PIX_IN[9404] NB2 NB1 CSA_VREF pixel
xPix9405 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[94] VREF PIX_IN[9405] NB2 NB1 CSA_VREF pixel
xPix9406 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[94] VREF PIX_IN[9406] NB2 NB1 CSA_VREF pixel
xPix9407 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[94] VREF PIX_IN[9407] NB2 NB1 CSA_VREF pixel
xPix9408 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[94] VREF PIX_IN[9408] NB2 NB1 CSA_VREF pixel
xPix9409 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[94] VREF PIX_IN[9409] NB2 NB1 CSA_VREF pixel
xPix9410 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[94] VREF PIX_IN[9410] NB2 NB1 CSA_VREF pixel
xPix9411 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[94] VREF PIX_IN[9411] NB2 NB1 CSA_VREF pixel
xPix9412 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[94] VREF PIX_IN[9412] NB2 NB1 CSA_VREF pixel
xPix9413 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[94] VREF PIX_IN[9413] NB2 NB1 CSA_VREF pixel
xPix9414 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[94] VREF PIX_IN[9414] NB2 NB1 CSA_VREF pixel
xPix9415 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[94] VREF PIX_IN[9415] NB2 NB1 CSA_VREF pixel
xPix9416 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[94] VREF PIX_IN[9416] NB2 NB1 CSA_VREF pixel
xPix9417 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[94] VREF PIX_IN[9417] NB2 NB1 CSA_VREF pixel
xPix9418 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[94] VREF PIX_IN[9418] NB2 NB1 CSA_VREF pixel
xPix9419 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[94] VREF PIX_IN[9419] NB2 NB1 CSA_VREF pixel
xPix9420 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[94] VREF PIX_IN[9420] NB2 NB1 CSA_VREF pixel
xPix9421 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[94] VREF PIX_IN[9421] NB2 NB1 CSA_VREF pixel
xPix9422 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[94] VREF PIX_IN[9422] NB2 NB1 CSA_VREF pixel
xPix9423 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[94] VREF PIX_IN[9423] NB2 NB1 CSA_VREF pixel
xPix9424 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[94] VREF PIX_IN[9424] NB2 NB1 CSA_VREF pixel
xPix9425 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[94] VREF PIX_IN[9425] NB2 NB1 CSA_VREF pixel
xPix9426 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[94] VREF PIX_IN[9426] NB2 NB1 CSA_VREF pixel
xPix9427 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[94] VREF PIX_IN[9427] NB2 NB1 CSA_VREF pixel
xPix9428 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[94] VREF PIX_IN[9428] NB2 NB1 CSA_VREF pixel
xPix9429 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[94] VREF PIX_IN[9429] NB2 NB1 CSA_VREF pixel
xPix9430 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[94] VREF PIX_IN[9430] NB2 NB1 CSA_VREF pixel
xPix9431 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[94] VREF PIX_IN[9431] NB2 NB1 CSA_VREF pixel
xPix9432 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[94] VREF PIX_IN[9432] NB2 NB1 CSA_VREF pixel
xPix9433 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[94] VREF PIX_IN[9433] NB2 NB1 CSA_VREF pixel
xPix9434 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[94] VREF PIX_IN[9434] NB2 NB1 CSA_VREF pixel
xPix9435 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[94] VREF PIX_IN[9435] NB2 NB1 CSA_VREF pixel
xPix9436 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[94] VREF PIX_IN[9436] NB2 NB1 CSA_VREF pixel
xPix9437 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[94] VREF PIX_IN[9437] NB2 NB1 CSA_VREF pixel
xPix9438 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[94] VREF PIX_IN[9438] NB2 NB1 CSA_VREF pixel
xPix9439 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[94] VREF PIX_IN[9439] NB2 NB1 CSA_VREF pixel
xPix9440 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[94] VREF PIX_IN[9440] NB2 NB1 CSA_VREF pixel
xPix9441 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[94] VREF PIX_IN[9441] NB2 NB1 CSA_VREF pixel
xPix9442 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[94] VREF PIX_IN[9442] NB2 NB1 CSA_VREF pixel
xPix9443 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[94] VREF PIX_IN[9443] NB2 NB1 CSA_VREF pixel
xPix9444 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[94] VREF PIX_IN[9444] NB2 NB1 CSA_VREF pixel
xPix9445 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[94] VREF PIX_IN[9445] NB2 NB1 CSA_VREF pixel
xPix9446 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[94] VREF PIX_IN[9446] NB2 NB1 CSA_VREF pixel
xPix9447 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[94] VREF PIX_IN[9447] NB2 NB1 CSA_VREF pixel
xPix9448 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[94] VREF PIX_IN[9448] NB2 NB1 CSA_VREF pixel
xPix9449 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[94] VREF PIX_IN[9449] NB2 NB1 CSA_VREF pixel
xPix9450 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[94] VREF PIX_IN[9450] NB2 NB1 CSA_VREF pixel
xPix9451 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[94] VREF PIX_IN[9451] NB2 NB1 CSA_VREF pixel
xPix9452 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[94] VREF PIX_IN[9452] NB2 NB1 CSA_VREF pixel
xPix9453 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[94] VREF PIX_IN[9453] NB2 NB1 CSA_VREF pixel
xPix9454 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[94] VREF PIX_IN[9454] NB2 NB1 CSA_VREF pixel
xPix9455 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[94] VREF PIX_IN[9455] NB2 NB1 CSA_VREF pixel
xPix9456 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[94] VREF PIX_IN[9456] NB2 NB1 CSA_VREF pixel
xPix9457 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[94] VREF PIX_IN[9457] NB2 NB1 CSA_VREF pixel
xPix9458 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[94] VREF PIX_IN[9458] NB2 NB1 CSA_VREF pixel
xPix9459 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[94] VREF PIX_IN[9459] NB2 NB1 CSA_VREF pixel
xPix9460 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[94] VREF PIX_IN[9460] NB2 NB1 CSA_VREF pixel
xPix9461 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[94] VREF PIX_IN[9461] NB2 NB1 CSA_VREF pixel
xPix9462 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[94] VREF PIX_IN[9462] NB2 NB1 CSA_VREF pixel
xPix9463 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[94] VREF PIX_IN[9463] NB2 NB1 CSA_VREF pixel
xPix9464 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[94] VREF PIX_IN[9464] NB2 NB1 CSA_VREF pixel
xPix9465 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[94] VREF PIX_IN[9465] NB2 NB1 CSA_VREF pixel
xPix9466 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[94] VREF PIX_IN[9466] NB2 NB1 CSA_VREF pixel
xPix9467 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[94] VREF PIX_IN[9467] NB2 NB1 CSA_VREF pixel
xPix9468 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[94] VREF PIX_IN[9468] NB2 NB1 CSA_VREF pixel
xPix9469 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[94] VREF PIX_IN[9469] NB2 NB1 CSA_VREF pixel
xPix9470 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[94] VREF PIX_IN[9470] NB2 NB1 CSA_VREF pixel
xPix9471 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[94] VREF PIX_IN[9471] NB2 NB1 CSA_VREF pixel
xPix9472 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[94] VREF PIX_IN[9472] NB2 NB1 CSA_VREF pixel
xPix9473 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[94] VREF PIX_IN[9473] NB2 NB1 CSA_VREF pixel
xPix9474 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[94] VREF PIX_IN[9474] NB2 NB1 CSA_VREF pixel
xPix9475 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[94] VREF PIX_IN[9475] NB2 NB1 CSA_VREF pixel
xPix9476 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[94] VREF PIX_IN[9476] NB2 NB1 CSA_VREF pixel
xPix9477 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[94] VREF PIX_IN[9477] NB2 NB1 CSA_VREF pixel
xPix9478 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[94] VREF PIX_IN[9478] NB2 NB1 CSA_VREF pixel
xPix9479 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[94] VREF PIX_IN[9479] NB2 NB1 CSA_VREF pixel
xPix9480 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[94] VREF PIX_IN[9480] NB2 NB1 CSA_VREF pixel
xPix9481 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[94] VREF PIX_IN[9481] NB2 NB1 CSA_VREF pixel
xPix9482 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[94] VREF PIX_IN[9482] NB2 NB1 CSA_VREF pixel
xPix9483 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[94] VREF PIX_IN[9483] NB2 NB1 CSA_VREF pixel
xPix9484 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[94] VREF PIX_IN[9484] NB2 NB1 CSA_VREF pixel
xPix9485 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[94] VREF PIX_IN[9485] NB2 NB1 CSA_VREF pixel
xPix9486 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[94] VREF PIX_IN[9486] NB2 NB1 CSA_VREF pixel
xPix9487 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[94] VREF PIX_IN[9487] NB2 NB1 CSA_VREF pixel
xPix9488 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[94] VREF PIX_IN[9488] NB2 NB1 CSA_VREF pixel
xPix9489 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[94] VREF PIX_IN[9489] NB2 NB1 CSA_VREF pixel
xPix9490 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[94] VREF PIX_IN[9490] NB2 NB1 CSA_VREF pixel
xPix9491 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[94] VREF PIX_IN[9491] NB2 NB1 CSA_VREF pixel
xPix9492 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[94] VREF PIX_IN[9492] NB2 NB1 CSA_VREF pixel
xPix9493 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[94] VREF PIX_IN[9493] NB2 NB1 CSA_VREF pixel
xPix9494 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[94] VREF PIX_IN[9494] NB2 NB1 CSA_VREF pixel
xPix9495 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[94] VREF PIX_IN[9495] NB2 NB1 CSA_VREF pixel
xPix9496 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[94] VREF PIX_IN[9496] NB2 NB1 CSA_VREF pixel
xPix9497 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[94] VREF PIX_IN[9497] NB2 NB1 CSA_VREF pixel
xPix9498 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[94] VREF PIX_IN[9498] NB2 NB1 CSA_VREF pixel
xPix9499 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[94] VREF PIX_IN[9499] NB2 NB1 CSA_VREF pixel
xPix9500 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[95] VREF PIX_IN[9500] NB2 NB1 CSA_VREF pixel
xPix9501 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[95] VREF PIX_IN[9501] NB2 NB1 CSA_VREF pixel
xPix9502 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[95] VREF PIX_IN[9502] NB2 NB1 CSA_VREF pixel
xPix9503 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[95] VREF PIX_IN[9503] NB2 NB1 CSA_VREF pixel
xPix9504 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[95] VREF PIX_IN[9504] NB2 NB1 CSA_VREF pixel
xPix9505 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[95] VREF PIX_IN[9505] NB2 NB1 CSA_VREF pixel
xPix9506 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[95] VREF PIX_IN[9506] NB2 NB1 CSA_VREF pixel
xPix9507 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[95] VREF PIX_IN[9507] NB2 NB1 CSA_VREF pixel
xPix9508 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[95] VREF PIX_IN[9508] NB2 NB1 CSA_VREF pixel
xPix9509 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[95] VREF PIX_IN[9509] NB2 NB1 CSA_VREF pixel
xPix9510 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[95] VREF PIX_IN[9510] NB2 NB1 CSA_VREF pixel
xPix9511 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[95] VREF PIX_IN[9511] NB2 NB1 CSA_VREF pixel
xPix9512 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[95] VREF PIX_IN[9512] NB2 NB1 CSA_VREF pixel
xPix9513 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[95] VREF PIX_IN[9513] NB2 NB1 CSA_VREF pixel
xPix9514 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[95] VREF PIX_IN[9514] NB2 NB1 CSA_VREF pixel
xPix9515 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[95] VREF PIX_IN[9515] NB2 NB1 CSA_VREF pixel
xPix9516 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[95] VREF PIX_IN[9516] NB2 NB1 CSA_VREF pixel
xPix9517 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[95] VREF PIX_IN[9517] NB2 NB1 CSA_VREF pixel
xPix9518 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[95] VREF PIX_IN[9518] NB2 NB1 CSA_VREF pixel
xPix9519 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[95] VREF PIX_IN[9519] NB2 NB1 CSA_VREF pixel
xPix9520 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[95] VREF PIX_IN[9520] NB2 NB1 CSA_VREF pixel
xPix9521 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[95] VREF PIX_IN[9521] NB2 NB1 CSA_VREF pixel
xPix9522 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[95] VREF PIX_IN[9522] NB2 NB1 CSA_VREF pixel
xPix9523 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[95] VREF PIX_IN[9523] NB2 NB1 CSA_VREF pixel
xPix9524 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[95] VREF PIX_IN[9524] NB2 NB1 CSA_VREF pixel
xPix9525 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[95] VREF PIX_IN[9525] NB2 NB1 CSA_VREF pixel
xPix9526 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[95] VREF PIX_IN[9526] NB2 NB1 CSA_VREF pixel
xPix9527 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[95] VREF PIX_IN[9527] NB2 NB1 CSA_VREF pixel
xPix9528 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[95] VREF PIX_IN[9528] NB2 NB1 CSA_VREF pixel
xPix9529 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[95] VREF PIX_IN[9529] NB2 NB1 CSA_VREF pixel
xPix9530 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[95] VREF PIX_IN[9530] NB2 NB1 CSA_VREF pixel
xPix9531 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[95] VREF PIX_IN[9531] NB2 NB1 CSA_VREF pixel
xPix9532 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[95] VREF PIX_IN[9532] NB2 NB1 CSA_VREF pixel
xPix9533 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[95] VREF PIX_IN[9533] NB2 NB1 CSA_VREF pixel
xPix9534 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[95] VREF PIX_IN[9534] NB2 NB1 CSA_VREF pixel
xPix9535 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[95] VREF PIX_IN[9535] NB2 NB1 CSA_VREF pixel
xPix9536 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[95] VREF PIX_IN[9536] NB2 NB1 CSA_VREF pixel
xPix9537 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[95] VREF PIX_IN[9537] NB2 NB1 CSA_VREF pixel
xPix9538 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[95] VREF PIX_IN[9538] NB2 NB1 CSA_VREF pixel
xPix9539 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[95] VREF PIX_IN[9539] NB2 NB1 CSA_VREF pixel
xPix9540 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[95] VREF PIX_IN[9540] NB2 NB1 CSA_VREF pixel
xPix9541 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[95] VREF PIX_IN[9541] NB2 NB1 CSA_VREF pixel
xPix9542 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[95] VREF PIX_IN[9542] NB2 NB1 CSA_VREF pixel
xPix9543 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[95] VREF PIX_IN[9543] NB2 NB1 CSA_VREF pixel
xPix9544 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[95] VREF PIX_IN[9544] NB2 NB1 CSA_VREF pixel
xPix9545 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[95] VREF PIX_IN[9545] NB2 NB1 CSA_VREF pixel
xPix9546 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[95] VREF PIX_IN[9546] NB2 NB1 CSA_VREF pixel
xPix9547 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[95] VREF PIX_IN[9547] NB2 NB1 CSA_VREF pixel
xPix9548 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[95] VREF PIX_IN[9548] NB2 NB1 CSA_VREF pixel
xPix9549 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[95] VREF PIX_IN[9549] NB2 NB1 CSA_VREF pixel
xPix9550 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[95] VREF PIX_IN[9550] NB2 NB1 CSA_VREF pixel
xPix9551 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[95] VREF PIX_IN[9551] NB2 NB1 CSA_VREF pixel
xPix9552 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[95] VREF PIX_IN[9552] NB2 NB1 CSA_VREF pixel
xPix9553 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[95] VREF PIX_IN[9553] NB2 NB1 CSA_VREF pixel
xPix9554 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[95] VREF PIX_IN[9554] NB2 NB1 CSA_VREF pixel
xPix9555 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[95] VREF PIX_IN[9555] NB2 NB1 CSA_VREF pixel
xPix9556 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[95] VREF PIX_IN[9556] NB2 NB1 CSA_VREF pixel
xPix9557 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[95] VREF PIX_IN[9557] NB2 NB1 CSA_VREF pixel
xPix9558 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[95] VREF PIX_IN[9558] NB2 NB1 CSA_VREF pixel
xPix9559 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[95] VREF PIX_IN[9559] NB2 NB1 CSA_VREF pixel
xPix9560 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[95] VREF PIX_IN[9560] NB2 NB1 CSA_VREF pixel
xPix9561 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[95] VREF PIX_IN[9561] NB2 NB1 CSA_VREF pixel
xPix9562 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[95] VREF PIX_IN[9562] NB2 NB1 CSA_VREF pixel
xPix9563 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[95] VREF PIX_IN[9563] NB2 NB1 CSA_VREF pixel
xPix9564 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[95] VREF PIX_IN[9564] NB2 NB1 CSA_VREF pixel
xPix9565 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[95] VREF PIX_IN[9565] NB2 NB1 CSA_VREF pixel
xPix9566 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[95] VREF PIX_IN[9566] NB2 NB1 CSA_VREF pixel
xPix9567 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[95] VREF PIX_IN[9567] NB2 NB1 CSA_VREF pixel
xPix9568 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[95] VREF PIX_IN[9568] NB2 NB1 CSA_VREF pixel
xPix9569 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[95] VREF PIX_IN[9569] NB2 NB1 CSA_VREF pixel
xPix9570 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[95] VREF PIX_IN[9570] NB2 NB1 CSA_VREF pixel
xPix9571 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[95] VREF PIX_IN[9571] NB2 NB1 CSA_VREF pixel
xPix9572 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[95] VREF PIX_IN[9572] NB2 NB1 CSA_VREF pixel
xPix9573 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[95] VREF PIX_IN[9573] NB2 NB1 CSA_VREF pixel
xPix9574 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[95] VREF PIX_IN[9574] NB2 NB1 CSA_VREF pixel
xPix9575 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[95] VREF PIX_IN[9575] NB2 NB1 CSA_VREF pixel
xPix9576 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[95] VREF PIX_IN[9576] NB2 NB1 CSA_VREF pixel
xPix9577 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[95] VREF PIX_IN[9577] NB2 NB1 CSA_VREF pixel
xPix9578 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[95] VREF PIX_IN[9578] NB2 NB1 CSA_VREF pixel
xPix9579 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[95] VREF PIX_IN[9579] NB2 NB1 CSA_VREF pixel
xPix9580 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[95] VREF PIX_IN[9580] NB2 NB1 CSA_VREF pixel
xPix9581 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[95] VREF PIX_IN[9581] NB2 NB1 CSA_VREF pixel
xPix9582 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[95] VREF PIX_IN[9582] NB2 NB1 CSA_VREF pixel
xPix9583 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[95] VREF PIX_IN[9583] NB2 NB1 CSA_VREF pixel
xPix9584 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[95] VREF PIX_IN[9584] NB2 NB1 CSA_VREF pixel
xPix9585 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[95] VREF PIX_IN[9585] NB2 NB1 CSA_VREF pixel
xPix9586 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[95] VREF PIX_IN[9586] NB2 NB1 CSA_VREF pixel
xPix9587 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[95] VREF PIX_IN[9587] NB2 NB1 CSA_VREF pixel
xPix9588 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[95] VREF PIX_IN[9588] NB2 NB1 CSA_VREF pixel
xPix9589 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[95] VREF PIX_IN[9589] NB2 NB1 CSA_VREF pixel
xPix9590 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[95] VREF PIX_IN[9590] NB2 NB1 CSA_VREF pixel
xPix9591 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[95] VREF PIX_IN[9591] NB2 NB1 CSA_VREF pixel
xPix9592 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[95] VREF PIX_IN[9592] NB2 NB1 CSA_VREF pixel
xPix9593 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[95] VREF PIX_IN[9593] NB2 NB1 CSA_VREF pixel
xPix9594 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[95] VREF PIX_IN[9594] NB2 NB1 CSA_VREF pixel
xPix9595 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[95] VREF PIX_IN[9595] NB2 NB1 CSA_VREF pixel
xPix9596 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[95] VREF PIX_IN[9596] NB2 NB1 CSA_VREF pixel
xPix9597 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[95] VREF PIX_IN[9597] NB2 NB1 CSA_VREF pixel
xPix9598 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[95] VREF PIX_IN[9598] NB2 NB1 CSA_VREF pixel
xPix9599 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[95] VREF PIX_IN[9599] NB2 NB1 CSA_VREF pixel
xPix9600 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[96] VREF PIX_IN[9600] NB2 NB1 CSA_VREF pixel
xPix9601 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[96] VREF PIX_IN[9601] NB2 NB1 CSA_VREF pixel
xPix9602 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[96] VREF PIX_IN[9602] NB2 NB1 CSA_VREF pixel
xPix9603 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[96] VREF PIX_IN[9603] NB2 NB1 CSA_VREF pixel
xPix9604 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[96] VREF PIX_IN[9604] NB2 NB1 CSA_VREF pixel
xPix9605 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[96] VREF PIX_IN[9605] NB2 NB1 CSA_VREF pixel
xPix9606 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[96] VREF PIX_IN[9606] NB2 NB1 CSA_VREF pixel
xPix9607 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[96] VREF PIX_IN[9607] NB2 NB1 CSA_VREF pixel
xPix9608 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[96] VREF PIX_IN[9608] NB2 NB1 CSA_VREF pixel
xPix9609 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[96] VREF PIX_IN[9609] NB2 NB1 CSA_VREF pixel
xPix9610 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[96] VREF PIX_IN[9610] NB2 NB1 CSA_VREF pixel
xPix9611 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[96] VREF PIX_IN[9611] NB2 NB1 CSA_VREF pixel
xPix9612 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[96] VREF PIX_IN[9612] NB2 NB1 CSA_VREF pixel
xPix9613 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[96] VREF PIX_IN[9613] NB2 NB1 CSA_VREF pixel
xPix9614 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[96] VREF PIX_IN[9614] NB2 NB1 CSA_VREF pixel
xPix9615 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[96] VREF PIX_IN[9615] NB2 NB1 CSA_VREF pixel
xPix9616 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[96] VREF PIX_IN[9616] NB2 NB1 CSA_VREF pixel
xPix9617 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[96] VREF PIX_IN[9617] NB2 NB1 CSA_VREF pixel
xPix9618 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[96] VREF PIX_IN[9618] NB2 NB1 CSA_VREF pixel
xPix9619 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[96] VREF PIX_IN[9619] NB2 NB1 CSA_VREF pixel
xPix9620 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[96] VREF PIX_IN[9620] NB2 NB1 CSA_VREF pixel
xPix9621 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[96] VREF PIX_IN[9621] NB2 NB1 CSA_VREF pixel
xPix9622 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[96] VREF PIX_IN[9622] NB2 NB1 CSA_VREF pixel
xPix9623 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[96] VREF PIX_IN[9623] NB2 NB1 CSA_VREF pixel
xPix9624 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[96] VREF PIX_IN[9624] NB2 NB1 CSA_VREF pixel
xPix9625 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[96] VREF PIX_IN[9625] NB2 NB1 CSA_VREF pixel
xPix9626 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[96] VREF PIX_IN[9626] NB2 NB1 CSA_VREF pixel
xPix9627 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[96] VREF PIX_IN[9627] NB2 NB1 CSA_VREF pixel
xPix9628 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[96] VREF PIX_IN[9628] NB2 NB1 CSA_VREF pixel
xPix9629 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[96] VREF PIX_IN[9629] NB2 NB1 CSA_VREF pixel
xPix9630 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[96] VREF PIX_IN[9630] NB2 NB1 CSA_VREF pixel
xPix9631 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[96] VREF PIX_IN[9631] NB2 NB1 CSA_VREF pixel
xPix9632 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[96] VREF PIX_IN[9632] NB2 NB1 CSA_VREF pixel
xPix9633 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[96] VREF PIX_IN[9633] NB2 NB1 CSA_VREF pixel
xPix9634 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[96] VREF PIX_IN[9634] NB2 NB1 CSA_VREF pixel
xPix9635 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[96] VREF PIX_IN[9635] NB2 NB1 CSA_VREF pixel
xPix9636 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[96] VREF PIX_IN[9636] NB2 NB1 CSA_VREF pixel
xPix9637 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[96] VREF PIX_IN[9637] NB2 NB1 CSA_VREF pixel
xPix9638 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[96] VREF PIX_IN[9638] NB2 NB1 CSA_VREF pixel
xPix9639 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[96] VREF PIX_IN[9639] NB2 NB1 CSA_VREF pixel
xPix9640 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[96] VREF PIX_IN[9640] NB2 NB1 CSA_VREF pixel
xPix9641 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[96] VREF PIX_IN[9641] NB2 NB1 CSA_VREF pixel
xPix9642 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[96] VREF PIX_IN[9642] NB2 NB1 CSA_VREF pixel
xPix9643 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[96] VREF PIX_IN[9643] NB2 NB1 CSA_VREF pixel
xPix9644 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[96] VREF PIX_IN[9644] NB2 NB1 CSA_VREF pixel
xPix9645 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[96] VREF PIX_IN[9645] NB2 NB1 CSA_VREF pixel
xPix9646 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[96] VREF PIX_IN[9646] NB2 NB1 CSA_VREF pixel
xPix9647 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[96] VREF PIX_IN[9647] NB2 NB1 CSA_VREF pixel
xPix9648 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[96] VREF PIX_IN[9648] NB2 NB1 CSA_VREF pixel
xPix9649 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[96] VREF PIX_IN[9649] NB2 NB1 CSA_VREF pixel
xPix9650 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[96] VREF PIX_IN[9650] NB2 NB1 CSA_VREF pixel
xPix9651 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[96] VREF PIX_IN[9651] NB2 NB1 CSA_VREF pixel
xPix9652 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[96] VREF PIX_IN[9652] NB2 NB1 CSA_VREF pixel
xPix9653 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[96] VREF PIX_IN[9653] NB2 NB1 CSA_VREF pixel
xPix9654 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[96] VREF PIX_IN[9654] NB2 NB1 CSA_VREF pixel
xPix9655 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[96] VREF PIX_IN[9655] NB2 NB1 CSA_VREF pixel
xPix9656 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[96] VREF PIX_IN[9656] NB2 NB1 CSA_VREF pixel
xPix9657 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[96] VREF PIX_IN[9657] NB2 NB1 CSA_VREF pixel
xPix9658 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[96] VREF PIX_IN[9658] NB2 NB1 CSA_VREF pixel
xPix9659 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[96] VREF PIX_IN[9659] NB2 NB1 CSA_VREF pixel
xPix9660 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[96] VREF PIX_IN[9660] NB2 NB1 CSA_VREF pixel
xPix9661 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[96] VREF PIX_IN[9661] NB2 NB1 CSA_VREF pixel
xPix9662 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[96] VREF PIX_IN[9662] NB2 NB1 CSA_VREF pixel
xPix9663 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[96] VREF PIX_IN[9663] NB2 NB1 CSA_VREF pixel
xPix9664 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[96] VREF PIX_IN[9664] NB2 NB1 CSA_VREF pixel
xPix9665 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[96] VREF PIX_IN[9665] NB2 NB1 CSA_VREF pixel
xPix9666 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[96] VREF PIX_IN[9666] NB2 NB1 CSA_VREF pixel
xPix9667 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[96] VREF PIX_IN[9667] NB2 NB1 CSA_VREF pixel
xPix9668 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[96] VREF PIX_IN[9668] NB2 NB1 CSA_VREF pixel
xPix9669 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[96] VREF PIX_IN[9669] NB2 NB1 CSA_VREF pixel
xPix9670 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[96] VREF PIX_IN[9670] NB2 NB1 CSA_VREF pixel
xPix9671 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[96] VREF PIX_IN[9671] NB2 NB1 CSA_VREF pixel
xPix9672 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[96] VREF PIX_IN[9672] NB2 NB1 CSA_VREF pixel
xPix9673 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[96] VREF PIX_IN[9673] NB2 NB1 CSA_VREF pixel
xPix9674 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[96] VREF PIX_IN[9674] NB2 NB1 CSA_VREF pixel
xPix9675 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[96] VREF PIX_IN[9675] NB2 NB1 CSA_VREF pixel
xPix9676 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[96] VREF PIX_IN[9676] NB2 NB1 CSA_VREF pixel
xPix9677 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[96] VREF PIX_IN[9677] NB2 NB1 CSA_VREF pixel
xPix9678 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[96] VREF PIX_IN[9678] NB2 NB1 CSA_VREF pixel
xPix9679 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[96] VREF PIX_IN[9679] NB2 NB1 CSA_VREF pixel
xPix9680 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[96] VREF PIX_IN[9680] NB2 NB1 CSA_VREF pixel
xPix9681 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[96] VREF PIX_IN[9681] NB2 NB1 CSA_VREF pixel
xPix9682 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[96] VREF PIX_IN[9682] NB2 NB1 CSA_VREF pixel
xPix9683 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[96] VREF PIX_IN[9683] NB2 NB1 CSA_VREF pixel
xPix9684 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[96] VREF PIX_IN[9684] NB2 NB1 CSA_VREF pixel
xPix9685 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[96] VREF PIX_IN[9685] NB2 NB1 CSA_VREF pixel
xPix9686 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[96] VREF PIX_IN[9686] NB2 NB1 CSA_VREF pixel
xPix9687 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[96] VREF PIX_IN[9687] NB2 NB1 CSA_VREF pixel
xPix9688 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[96] VREF PIX_IN[9688] NB2 NB1 CSA_VREF pixel
xPix9689 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[96] VREF PIX_IN[9689] NB2 NB1 CSA_VREF pixel
xPix9690 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[96] VREF PIX_IN[9690] NB2 NB1 CSA_VREF pixel
xPix9691 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[96] VREF PIX_IN[9691] NB2 NB1 CSA_VREF pixel
xPix9692 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[96] VREF PIX_IN[9692] NB2 NB1 CSA_VREF pixel
xPix9693 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[96] VREF PIX_IN[9693] NB2 NB1 CSA_VREF pixel
xPix9694 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[96] VREF PIX_IN[9694] NB2 NB1 CSA_VREF pixel
xPix9695 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[96] VREF PIX_IN[9695] NB2 NB1 CSA_VREF pixel
xPix9696 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[96] VREF PIX_IN[9696] NB2 NB1 CSA_VREF pixel
xPix9697 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[96] VREF PIX_IN[9697] NB2 NB1 CSA_VREF pixel
xPix9698 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[96] VREF PIX_IN[9698] NB2 NB1 CSA_VREF pixel
xPix9699 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[96] VREF PIX_IN[9699] NB2 NB1 CSA_VREF pixel
xPix9700 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[97] VREF PIX_IN[9700] NB2 NB1 CSA_VREF pixel
xPix9701 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[97] VREF PIX_IN[9701] NB2 NB1 CSA_VREF pixel
xPix9702 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[97] VREF PIX_IN[9702] NB2 NB1 CSA_VREF pixel
xPix9703 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[97] VREF PIX_IN[9703] NB2 NB1 CSA_VREF pixel
xPix9704 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[97] VREF PIX_IN[9704] NB2 NB1 CSA_VREF pixel
xPix9705 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[97] VREF PIX_IN[9705] NB2 NB1 CSA_VREF pixel
xPix9706 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[97] VREF PIX_IN[9706] NB2 NB1 CSA_VREF pixel
xPix9707 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[97] VREF PIX_IN[9707] NB2 NB1 CSA_VREF pixel
xPix9708 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[97] VREF PIX_IN[9708] NB2 NB1 CSA_VREF pixel
xPix9709 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[97] VREF PIX_IN[9709] NB2 NB1 CSA_VREF pixel
xPix9710 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[97] VREF PIX_IN[9710] NB2 NB1 CSA_VREF pixel
xPix9711 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[97] VREF PIX_IN[9711] NB2 NB1 CSA_VREF pixel
xPix9712 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[97] VREF PIX_IN[9712] NB2 NB1 CSA_VREF pixel
xPix9713 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[97] VREF PIX_IN[9713] NB2 NB1 CSA_VREF pixel
xPix9714 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[97] VREF PIX_IN[9714] NB2 NB1 CSA_VREF pixel
xPix9715 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[97] VREF PIX_IN[9715] NB2 NB1 CSA_VREF pixel
xPix9716 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[97] VREF PIX_IN[9716] NB2 NB1 CSA_VREF pixel
xPix9717 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[97] VREF PIX_IN[9717] NB2 NB1 CSA_VREF pixel
xPix9718 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[97] VREF PIX_IN[9718] NB2 NB1 CSA_VREF pixel
xPix9719 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[97] VREF PIX_IN[9719] NB2 NB1 CSA_VREF pixel
xPix9720 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[97] VREF PIX_IN[9720] NB2 NB1 CSA_VREF pixel
xPix9721 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[97] VREF PIX_IN[9721] NB2 NB1 CSA_VREF pixel
xPix9722 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[97] VREF PIX_IN[9722] NB2 NB1 CSA_VREF pixel
xPix9723 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[97] VREF PIX_IN[9723] NB2 NB1 CSA_VREF pixel
xPix9724 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[97] VREF PIX_IN[9724] NB2 NB1 CSA_VREF pixel
xPix9725 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[97] VREF PIX_IN[9725] NB2 NB1 CSA_VREF pixel
xPix9726 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[97] VREF PIX_IN[9726] NB2 NB1 CSA_VREF pixel
xPix9727 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[97] VREF PIX_IN[9727] NB2 NB1 CSA_VREF pixel
xPix9728 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[97] VREF PIX_IN[9728] NB2 NB1 CSA_VREF pixel
xPix9729 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[97] VREF PIX_IN[9729] NB2 NB1 CSA_VREF pixel
xPix9730 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[97] VREF PIX_IN[9730] NB2 NB1 CSA_VREF pixel
xPix9731 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[97] VREF PIX_IN[9731] NB2 NB1 CSA_VREF pixel
xPix9732 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[97] VREF PIX_IN[9732] NB2 NB1 CSA_VREF pixel
xPix9733 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[97] VREF PIX_IN[9733] NB2 NB1 CSA_VREF pixel
xPix9734 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[97] VREF PIX_IN[9734] NB2 NB1 CSA_VREF pixel
xPix9735 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[97] VREF PIX_IN[9735] NB2 NB1 CSA_VREF pixel
xPix9736 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[97] VREF PIX_IN[9736] NB2 NB1 CSA_VREF pixel
xPix9737 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[97] VREF PIX_IN[9737] NB2 NB1 CSA_VREF pixel
xPix9738 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[97] VREF PIX_IN[9738] NB2 NB1 CSA_VREF pixel
xPix9739 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[97] VREF PIX_IN[9739] NB2 NB1 CSA_VREF pixel
xPix9740 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[97] VREF PIX_IN[9740] NB2 NB1 CSA_VREF pixel
xPix9741 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[97] VREF PIX_IN[9741] NB2 NB1 CSA_VREF pixel
xPix9742 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[97] VREF PIX_IN[9742] NB2 NB1 CSA_VREF pixel
xPix9743 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[97] VREF PIX_IN[9743] NB2 NB1 CSA_VREF pixel
xPix9744 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[97] VREF PIX_IN[9744] NB2 NB1 CSA_VREF pixel
xPix9745 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[97] VREF PIX_IN[9745] NB2 NB1 CSA_VREF pixel
xPix9746 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[97] VREF PIX_IN[9746] NB2 NB1 CSA_VREF pixel
xPix9747 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[97] VREF PIX_IN[9747] NB2 NB1 CSA_VREF pixel
xPix9748 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[97] VREF PIX_IN[9748] NB2 NB1 CSA_VREF pixel
xPix9749 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[97] VREF PIX_IN[9749] NB2 NB1 CSA_VREF pixel
xPix9750 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[97] VREF PIX_IN[9750] NB2 NB1 CSA_VREF pixel
xPix9751 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[97] VREF PIX_IN[9751] NB2 NB1 CSA_VREF pixel
xPix9752 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[97] VREF PIX_IN[9752] NB2 NB1 CSA_VREF pixel
xPix9753 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[97] VREF PIX_IN[9753] NB2 NB1 CSA_VREF pixel
xPix9754 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[97] VREF PIX_IN[9754] NB2 NB1 CSA_VREF pixel
xPix9755 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[97] VREF PIX_IN[9755] NB2 NB1 CSA_VREF pixel
xPix9756 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[97] VREF PIX_IN[9756] NB2 NB1 CSA_VREF pixel
xPix9757 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[97] VREF PIX_IN[9757] NB2 NB1 CSA_VREF pixel
xPix9758 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[97] VREF PIX_IN[9758] NB2 NB1 CSA_VREF pixel
xPix9759 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[97] VREF PIX_IN[9759] NB2 NB1 CSA_VREF pixel
xPix9760 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[97] VREF PIX_IN[9760] NB2 NB1 CSA_VREF pixel
xPix9761 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[97] VREF PIX_IN[9761] NB2 NB1 CSA_VREF pixel
xPix9762 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[97] VREF PIX_IN[9762] NB2 NB1 CSA_VREF pixel
xPix9763 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[97] VREF PIX_IN[9763] NB2 NB1 CSA_VREF pixel
xPix9764 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[97] VREF PIX_IN[9764] NB2 NB1 CSA_VREF pixel
xPix9765 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[97] VREF PIX_IN[9765] NB2 NB1 CSA_VREF pixel
xPix9766 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[97] VREF PIX_IN[9766] NB2 NB1 CSA_VREF pixel
xPix9767 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[97] VREF PIX_IN[9767] NB2 NB1 CSA_VREF pixel
xPix9768 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[97] VREF PIX_IN[9768] NB2 NB1 CSA_VREF pixel
xPix9769 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[97] VREF PIX_IN[9769] NB2 NB1 CSA_VREF pixel
xPix9770 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[97] VREF PIX_IN[9770] NB2 NB1 CSA_VREF pixel
xPix9771 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[97] VREF PIX_IN[9771] NB2 NB1 CSA_VREF pixel
xPix9772 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[97] VREF PIX_IN[9772] NB2 NB1 CSA_VREF pixel
xPix9773 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[97] VREF PIX_IN[9773] NB2 NB1 CSA_VREF pixel
xPix9774 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[97] VREF PIX_IN[9774] NB2 NB1 CSA_VREF pixel
xPix9775 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[97] VREF PIX_IN[9775] NB2 NB1 CSA_VREF pixel
xPix9776 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[97] VREF PIX_IN[9776] NB2 NB1 CSA_VREF pixel
xPix9777 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[97] VREF PIX_IN[9777] NB2 NB1 CSA_VREF pixel
xPix9778 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[97] VREF PIX_IN[9778] NB2 NB1 CSA_VREF pixel
xPix9779 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[97] VREF PIX_IN[9779] NB2 NB1 CSA_VREF pixel
xPix9780 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[97] VREF PIX_IN[9780] NB2 NB1 CSA_VREF pixel
xPix9781 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[97] VREF PIX_IN[9781] NB2 NB1 CSA_VREF pixel
xPix9782 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[97] VREF PIX_IN[9782] NB2 NB1 CSA_VREF pixel
xPix9783 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[97] VREF PIX_IN[9783] NB2 NB1 CSA_VREF pixel
xPix9784 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[97] VREF PIX_IN[9784] NB2 NB1 CSA_VREF pixel
xPix9785 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[97] VREF PIX_IN[9785] NB2 NB1 CSA_VREF pixel
xPix9786 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[97] VREF PIX_IN[9786] NB2 NB1 CSA_VREF pixel
xPix9787 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[97] VREF PIX_IN[9787] NB2 NB1 CSA_VREF pixel
xPix9788 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[97] VREF PIX_IN[9788] NB2 NB1 CSA_VREF pixel
xPix9789 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[97] VREF PIX_IN[9789] NB2 NB1 CSA_VREF pixel
xPix9790 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[97] VREF PIX_IN[9790] NB2 NB1 CSA_VREF pixel
xPix9791 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[97] VREF PIX_IN[9791] NB2 NB1 CSA_VREF pixel
xPix9792 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[97] VREF PIX_IN[9792] NB2 NB1 CSA_VREF pixel
xPix9793 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[97] VREF PIX_IN[9793] NB2 NB1 CSA_VREF pixel
xPix9794 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[97] VREF PIX_IN[9794] NB2 NB1 CSA_VREF pixel
xPix9795 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[97] VREF PIX_IN[9795] NB2 NB1 CSA_VREF pixel
xPix9796 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[97] VREF PIX_IN[9796] NB2 NB1 CSA_VREF pixel
xPix9797 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[97] VREF PIX_IN[9797] NB2 NB1 CSA_VREF pixel
xPix9798 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[97] VREF PIX_IN[9798] NB2 NB1 CSA_VREF pixel
xPix9799 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[97] VREF PIX_IN[9799] NB2 NB1 CSA_VREF pixel
xPix9800 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[98] VREF PIX_IN[9800] NB2 NB1 CSA_VREF pixel
xPix9801 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[98] VREF PIX_IN[9801] NB2 NB1 CSA_VREF pixel
xPix9802 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[98] VREF PIX_IN[9802] NB2 NB1 CSA_VREF pixel
xPix9803 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[98] VREF PIX_IN[9803] NB2 NB1 CSA_VREF pixel
xPix9804 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[98] VREF PIX_IN[9804] NB2 NB1 CSA_VREF pixel
xPix9805 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[98] VREF PIX_IN[9805] NB2 NB1 CSA_VREF pixel
xPix9806 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[98] VREF PIX_IN[9806] NB2 NB1 CSA_VREF pixel
xPix9807 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[98] VREF PIX_IN[9807] NB2 NB1 CSA_VREF pixel
xPix9808 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[98] VREF PIX_IN[9808] NB2 NB1 CSA_VREF pixel
xPix9809 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[98] VREF PIX_IN[9809] NB2 NB1 CSA_VREF pixel
xPix9810 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[98] VREF PIX_IN[9810] NB2 NB1 CSA_VREF pixel
xPix9811 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[98] VREF PIX_IN[9811] NB2 NB1 CSA_VREF pixel
xPix9812 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[98] VREF PIX_IN[9812] NB2 NB1 CSA_VREF pixel
xPix9813 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[98] VREF PIX_IN[9813] NB2 NB1 CSA_VREF pixel
xPix9814 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[98] VREF PIX_IN[9814] NB2 NB1 CSA_VREF pixel
xPix9815 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[98] VREF PIX_IN[9815] NB2 NB1 CSA_VREF pixel
xPix9816 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[98] VREF PIX_IN[9816] NB2 NB1 CSA_VREF pixel
xPix9817 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[98] VREF PIX_IN[9817] NB2 NB1 CSA_VREF pixel
xPix9818 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[98] VREF PIX_IN[9818] NB2 NB1 CSA_VREF pixel
xPix9819 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[98] VREF PIX_IN[9819] NB2 NB1 CSA_VREF pixel
xPix9820 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[98] VREF PIX_IN[9820] NB2 NB1 CSA_VREF pixel
xPix9821 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[98] VREF PIX_IN[9821] NB2 NB1 CSA_VREF pixel
xPix9822 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[98] VREF PIX_IN[9822] NB2 NB1 CSA_VREF pixel
xPix9823 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[98] VREF PIX_IN[9823] NB2 NB1 CSA_VREF pixel
xPix9824 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[98] VREF PIX_IN[9824] NB2 NB1 CSA_VREF pixel
xPix9825 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[98] VREF PIX_IN[9825] NB2 NB1 CSA_VREF pixel
xPix9826 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[98] VREF PIX_IN[9826] NB2 NB1 CSA_VREF pixel
xPix9827 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[98] VREF PIX_IN[9827] NB2 NB1 CSA_VREF pixel
xPix9828 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[98] VREF PIX_IN[9828] NB2 NB1 CSA_VREF pixel
xPix9829 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[98] VREF PIX_IN[9829] NB2 NB1 CSA_VREF pixel
xPix9830 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[98] VREF PIX_IN[9830] NB2 NB1 CSA_VREF pixel
xPix9831 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[98] VREF PIX_IN[9831] NB2 NB1 CSA_VREF pixel
xPix9832 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[98] VREF PIX_IN[9832] NB2 NB1 CSA_VREF pixel
xPix9833 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[98] VREF PIX_IN[9833] NB2 NB1 CSA_VREF pixel
xPix9834 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[98] VREF PIX_IN[9834] NB2 NB1 CSA_VREF pixel
xPix9835 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[98] VREF PIX_IN[9835] NB2 NB1 CSA_VREF pixel
xPix9836 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[98] VREF PIX_IN[9836] NB2 NB1 CSA_VREF pixel
xPix9837 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[98] VREF PIX_IN[9837] NB2 NB1 CSA_VREF pixel
xPix9838 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[98] VREF PIX_IN[9838] NB2 NB1 CSA_VREF pixel
xPix9839 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[98] VREF PIX_IN[9839] NB2 NB1 CSA_VREF pixel
xPix9840 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[98] VREF PIX_IN[9840] NB2 NB1 CSA_VREF pixel
xPix9841 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[98] VREF PIX_IN[9841] NB2 NB1 CSA_VREF pixel
xPix9842 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[98] VREF PIX_IN[9842] NB2 NB1 CSA_VREF pixel
xPix9843 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[98] VREF PIX_IN[9843] NB2 NB1 CSA_VREF pixel
xPix9844 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[98] VREF PIX_IN[9844] NB2 NB1 CSA_VREF pixel
xPix9845 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[98] VREF PIX_IN[9845] NB2 NB1 CSA_VREF pixel
xPix9846 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[98] VREF PIX_IN[9846] NB2 NB1 CSA_VREF pixel
xPix9847 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[98] VREF PIX_IN[9847] NB2 NB1 CSA_VREF pixel
xPix9848 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[98] VREF PIX_IN[9848] NB2 NB1 CSA_VREF pixel
xPix9849 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[98] VREF PIX_IN[9849] NB2 NB1 CSA_VREF pixel
xPix9850 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[98] VREF PIX_IN[9850] NB2 NB1 CSA_VREF pixel
xPix9851 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[98] VREF PIX_IN[9851] NB2 NB1 CSA_VREF pixel
xPix9852 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[98] VREF PIX_IN[9852] NB2 NB1 CSA_VREF pixel
xPix9853 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[98] VREF PIX_IN[9853] NB2 NB1 CSA_VREF pixel
xPix9854 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[98] VREF PIX_IN[9854] NB2 NB1 CSA_VREF pixel
xPix9855 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[98] VREF PIX_IN[9855] NB2 NB1 CSA_VREF pixel
xPix9856 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[98] VREF PIX_IN[9856] NB2 NB1 CSA_VREF pixel
xPix9857 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[98] VREF PIX_IN[9857] NB2 NB1 CSA_VREF pixel
xPix9858 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[98] VREF PIX_IN[9858] NB2 NB1 CSA_VREF pixel
xPix9859 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[98] VREF PIX_IN[9859] NB2 NB1 CSA_VREF pixel
xPix9860 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[98] VREF PIX_IN[9860] NB2 NB1 CSA_VREF pixel
xPix9861 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[98] VREF PIX_IN[9861] NB2 NB1 CSA_VREF pixel
xPix9862 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[98] VREF PIX_IN[9862] NB2 NB1 CSA_VREF pixel
xPix9863 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[98] VREF PIX_IN[9863] NB2 NB1 CSA_VREF pixel
xPix9864 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[98] VREF PIX_IN[9864] NB2 NB1 CSA_VREF pixel
xPix9865 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[98] VREF PIX_IN[9865] NB2 NB1 CSA_VREF pixel
xPix9866 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[98] VREF PIX_IN[9866] NB2 NB1 CSA_VREF pixel
xPix9867 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[98] VREF PIX_IN[9867] NB2 NB1 CSA_VREF pixel
xPix9868 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[98] VREF PIX_IN[9868] NB2 NB1 CSA_VREF pixel
xPix9869 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[98] VREF PIX_IN[9869] NB2 NB1 CSA_VREF pixel
xPix9870 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[98] VREF PIX_IN[9870] NB2 NB1 CSA_VREF pixel
xPix9871 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[98] VREF PIX_IN[9871] NB2 NB1 CSA_VREF pixel
xPix9872 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[98] VREF PIX_IN[9872] NB2 NB1 CSA_VREF pixel
xPix9873 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[98] VREF PIX_IN[9873] NB2 NB1 CSA_VREF pixel
xPix9874 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[98] VREF PIX_IN[9874] NB2 NB1 CSA_VREF pixel
xPix9875 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[98] VREF PIX_IN[9875] NB2 NB1 CSA_VREF pixel
xPix9876 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[98] VREF PIX_IN[9876] NB2 NB1 CSA_VREF pixel
xPix9877 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[98] VREF PIX_IN[9877] NB2 NB1 CSA_VREF pixel
xPix9878 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[98] VREF PIX_IN[9878] NB2 NB1 CSA_VREF pixel
xPix9879 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[98] VREF PIX_IN[9879] NB2 NB1 CSA_VREF pixel
xPix9880 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[98] VREF PIX_IN[9880] NB2 NB1 CSA_VREF pixel
xPix9881 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[98] VREF PIX_IN[9881] NB2 NB1 CSA_VREF pixel
xPix9882 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[98] VREF PIX_IN[9882] NB2 NB1 CSA_VREF pixel
xPix9883 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[98] VREF PIX_IN[9883] NB2 NB1 CSA_VREF pixel
xPix9884 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[98] VREF PIX_IN[9884] NB2 NB1 CSA_VREF pixel
xPix9885 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[98] VREF PIX_IN[9885] NB2 NB1 CSA_VREF pixel
xPix9886 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[98] VREF PIX_IN[9886] NB2 NB1 CSA_VREF pixel
xPix9887 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[98] VREF PIX_IN[9887] NB2 NB1 CSA_VREF pixel
xPix9888 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[98] VREF PIX_IN[9888] NB2 NB1 CSA_VREF pixel
xPix9889 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[98] VREF PIX_IN[9889] NB2 NB1 CSA_VREF pixel
xPix9890 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[98] VREF PIX_IN[9890] NB2 NB1 CSA_VREF pixel
xPix9891 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[98] VREF PIX_IN[9891] NB2 NB1 CSA_VREF pixel
xPix9892 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[98] VREF PIX_IN[9892] NB2 NB1 CSA_VREF pixel
xPix9893 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[98] VREF PIX_IN[9893] NB2 NB1 CSA_VREF pixel
xPix9894 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[98] VREF PIX_IN[9894] NB2 NB1 CSA_VREF pixel
xPix9895 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[98] VREF PIX_IN[9895] NB2 NB1 CSA_VREF pixel
xPix9896 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[98] VREF PIX_IN[9896] NB2 NB1 CSA_VREF pixel
xPix9897 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[98] VREF PIX_IN[9897] NB2 NB1 CSA_VREF pixel
xPix9898 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[98] VREF PIX_IN[9898] NB2 NB1 CSA_VREF pixel
xPix9899 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[98] VREF PIX_IN[9899] NB2 NB1 CSA_VREF pixel
xPix9900 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[99] VREF PIX_IN[9900] NB2 NB1 CSA_VREF pixel
xPix9901 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[99] VREF PIX_IN[9901] NB2 NB1 CSA_VREF pixel
xPix9902 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[99] VREF PIX_IN[9902] NB2 NB1 CSA_VREF pixel
xPix9903 VDD GND SF_IB gring VBIAS COL_OUT[3] ROW_SEL[99] VREF PIX_IN[9903] NB2 NB1 CSA_VREF pixel
xPix9904 VDD GND SF_IB gring VBIAS COL_OUT[4] ROW_SEL[99] VREF PIX_IN[9904] NB2 NB1 CSA_VREF pixel
xPix9905 VDD GND SF_IB gring VBIAS COL_OUT[5] ROW_SEL[99] VREF PIX_IN[9905] NB2 NB1 CSA_VREF pixel
xPix9906 VDD GND SF_IB gring VBIAS COL_OUT[6] ROW_SEL[99] VREF PIX_IN[9906] NB2 NB1 CSA_VREF pixel
xPix9907 VDD GND SF_IB gring VBIAS COL_OUT[7] ROW_SEL[99] VREF PIX_IN[9907] NB2 NB1 CSA_VREF pixel
xPix9908 VDD GND SF_IB gring VBIAS COL_OUT[8] ROW_SEL[99] VREF PIX_IN[9908] NB2 NB1 CSA_VREF pixel
xPix9909 VDD GND SF_IB gring VBIAS COL_OUT[9] ROW_SEL[99] VREF PIX_IN[9909] NB2 NB1 CSA_VREF pixel
xPix9910 VDD GND SF_IB gring VBIAS COL_OUT[10] ROW_SEL[99] VREF PIX_IN[9910] NB2 NB1 CSA_VREF pixel
xPix9911 VDD GND SF_IB gring VBIAS COL_OUT[11] ROW_SEL[99] VREF PIX_IN[9911] NB2 NB1 CSA_VREF pixel
xPix9912 VDD GND SF_IB gring VBIAS COL_OUT[12] ROW_SEL[99] VREF PIX_IN[9912] NB2 NB1 CSA_VREF pixel
xPix9913 VDD GND SF_IB gring VBIAS COL_OUT[13] ROW_SEL[99] VREF PIX_IN[9913] NB2 NB1 CSA_VREF pixel
xPix9914 VDD GND SF_IB gring VBIAS COL_OUT[14] ROW_SEL[99] VREF PIX_IN[9914] NB2 NB1 CSA_VREF pixel
xPix9915 VDD GND SF_IB gring VBIAS COL_OUT[15] ROW_SEL[99] VREF PIX_IN[9915] NB2 NB1 CSA_VREF pixel
xPix9916 VDD GND SF_IB gring VBIAS COL_OUT[16] ROW_SEL[99] VREF PIX_IN[9916] NB2 NB1 CSA_VREF pixel
xPix9917 VDD GND SF_IB gring VBIAS COL_OUT[17] ROW_SEL[99] VREF PIX_IN[9917] NB2 NB1 CSA_VREF pixel
xPix9918 VDD GND SF_IB gring VBIAS COL_OUT[18] ROW_SEL[99] VREF PIX_IN[9918] NB2 NB1 CSA_VREF pixel
xPix9919 VDD GND SF_IB gring VBIAS COL_OUT[19] ROW_SEL[99] VREF PIX_IN[9919] NB2 NB1 CSA_VREF pixel
xPix9920 VDD GND SF_IB gring VBIAS COL_OUT[20] ROW_SEL[99] VREF PIX_IN[9920] NB2 NB1 CSA_VREF pixel
xPix9921 VDD GND SF_IB gring VBIAS COL_OUT[21] ROW_SEL[99] VREF PIX_IN[9921] NB2 NB1 CSA_VREF pixel
xPix9922 VDD GND SF_IB gring VBIAS COL_OUT[22] ROW_SEL[99] VREF PIX_IN[9922] NB2 NB1 CSA_VREF pixel
xPix9923 VDD GND SF_IB gring VBIAS COL_OUT[23] ROW_SEL[99] VREF PIX_IN[9923] NB2 NB1 CSA_VREF pixel
xPix9924 VDD GND SF_IB gring VBIAS COL_OUT[24] ROW_SEL[99] VREF PIX_IN[9924] NB2 NB1 CSA_VREF pixel
xPix9925 VDD GND SF_IB gring VBIAS COL_OUT[25] ROW_SEL[99] VREF PIX_IN[9925] NB2 NB1 CSA_VREF pixel
xPix9926 VDD GND SF_IB gring VBIAS COL_OUT[26] ROW_SEL[99] VREF PIX_IN[9926] NB2 NB1 CSA_VREF pixel
xPix9927 VDD GND SF_IB gring VBIAS COL_OUT[27] ROW_SEL[99] VREF PIX_IN[9927] NB2 NB1 CSA_VREF pixel
xPix9928 VDD GND SF_IB gring VBIAS COL_OUT[28] ROW_SEL[99] VREF PIX_IN[9928] NB2 NB1 CSA_VREF pixel
xPix9929 VDD GND SF_IB gring VBIAS COL_OUT[29] ROW_SEL[99] VREF PIX_IN[9929] NB2 NB1 CSA_VREF pixel
xPix9930 VDD GND SF_IB gring VBIAS COL_OUT[30] ROW_SEL[99] VREF PIX_IN[9930] NB2 NB1 CSA_VREF pixel
xPix9931 VDD GND SF_IB gring VBIAS COL_OUT[31] ROW_SEL[99] VREF PIX_IN[9931] NB2 NB1 CSA_VREF pixel
xPix9932 VDD GND SF_IB gring VBIAS COL_OUT[32] ROW_SEL[99] VREF PIX_IN[9932] NB2 NB1 CSA_VREF pixel
xPix9933 VDD GND SF_IB gring VBIAS COL_OUT[33] ROW_SEL[99] VREF PIX_IN[9933] NB2 NB1 CSA_VREF pixel
xPix9934 VDD GND SF_IB gring VBIAS COL_OUT[34] ROW_SEL[99] VREF PIX_IN[9934] NB2 NB1 CSA_VREF pixel
xPix9935 VDD GND SF_IB gring VBIAS COL_OUT[35] ROW_SEL[99] VREF PIX_IN[9935] NB2 NB1 CSA_VREF pixel
xPix9936 VDD GND SF_IB gring VBIAS COL_OUT[36] ROW_SEL[99] VREF PIX_IN[9936] NB2 NB1 CSA_VREF pixel
xPix9937 VDD GND SF_IB gring VBIAS COL_OUT[37] ROW_SEL[99] VREF PIX_IN[9937] NB2 NB1 CSA_VREF pixel
xPix9938 VDD GND SF_IB gring VBIAS COL_OUT[38] ROW_SEL[99] VREF PIX_IN[9938] NB2 NB1 CSA_VREF pixel
xPix9939 VDD GND SF_IB gring VBIAS COL_OUT[39] ROW_SEL[99] VREF PIX_IN[9939] NB2 NB1 CSA_VREF pixel
xPix9940 VDD GND SF_IB gring VBIAS COL_OUT[40] ROW_SEL[99] VREF PIX_IN[9940] NB2 NB1 CSA_VREF pixel
xPix9941 VDD GND SF_IB gring VBIAS COL_OUT[41] ROW_SEL[99] VREF PIX_IN[9941] NB2 NB1 CSA_VREF pixel
xPix9942 VDD GND SF_IB gring VBIAS COL_OUT[42] ROW_SEL[99] VREF PIX_IN[9942] NB2 NB1 CSA_VREF pixel
xPix9943 VDD GND SF_IB gring VBIAS COL_OUT[43] ROW_SEL[99] VREF PIX_IN[9943] NB2 NB1 CSA_VREF pixel
xPix9944 VDD GND SF_IB gring VBIAS COL_OUT[44] ROW_SEL[99] VREF PIX_IN[9944] NB2 NB1 CSA_VREF pixel
xPix9945 VDD GND SF_IB gring VBIAS COL_OUT[45] ROW_SEL[99] VREF PIX_IN[9945] NB2 NB1 CSA_VREF pixel
xPix9946 VDD GND SF_IB gring VBIAS COL_OUT[46] ROW_SEL[99] VREF PIX_IN[9946] NB2 NB1 CSA_VREF pixel
xPix9947 VDD GND SF_IB gring VBIAS COL_OUT[47] ROW_SEL[99] VREF PIX_IN[9947] NB2 NB1 CSA_VREF pixel
xPix9948 VDD GND SF_IB gring VBIAS COL_OUT[48] ROW_SEL[99] VREF PIX_IN[9948] NB2 NB1 CSA_VREF pixel
xPix9949 VDD GND SF_IB gring VBIAS COL_OUT[49] ROW_SEL[99] VREF PIX_IN[9949] NB2 NB1 CSA_VREF pixel
xPix9950 VDD GND SF_IB gring VBIAS COL_OUT[50] ROW_SEL[99] VREF PIX_IN[9950] NB2 NB1 CSA_VREF pixel
xPix9951 VDD GND SF_IB gring VBIAS COL_OUT[51] ROW_SEL[99] VREF PIX_IN[9951] NB2 NB1 CSA_VREF pixel
xPix9952 VDD GND SF_IB gring VBIAS COL_OUT[52] ROW_SEL[99] VREF PIX_IN[9952] NB2 NB1 CSA_VREF pixel
xPix9953 VDD GND SF_IB gring VBIAS COL_OUT[53] ROW_SEL[99] VREF PIX_IN[9953] NB2 NB1 CSA_VREF pixel
xPix9954 VDD GND SF_IB gring VBIAS COL_OUT[54] ROW_SEL[99] VREF PIX_IN[9954] NB2 NB1 CSA_VREF pixel
xPix9955 VDD GND SF_IB gring VBIAS COL_OUT[55] ROW_SEL[99] VREF PIX_IN[9955] NB2 NB1 CSA_VREF pixel
xPix9956 VDD GND SF_IB gring VBIAS COL_OUT[56] ROW_SEL[99] VREF PIX_IN[9956] NB2 NB1 CSA_VREF pixel
xPix9957 VDD GND SF_IB gring VBIAS COL_OUT[57] ROW_SEL[99] VREF PIX_IN[9957] NB2 NB1 CSA_VREF pixel
xPix9958 VDD GND SF_IB gring VBIAS COL_OUT[58] ROW_SEL[99] VREF PIX_IN[9958] NB2 NB1 CSA_VREF pixel
xPix9959 VDD GND SF_IB gring VBIAS COL_OUT[59] ROW_SEL[99] VREF PIX_IN[9959] NB2 NB1 CSA_VREF pixel
xPix9960 VDD GND SF_IB gring VBIAS COL_OUT[60] ROW_SEL[99] VREF PIX_IN[9960] NB2 NB1 CSA_VREF pixel
xPix9961 VDD GND SF_IB gring VBIAS COL_OUT[61] ROW_SEL[99] VREF PIX_IN[9961] NB2 NB1 CSA_VREF pixel
xPix9962 VDD GND SF_IB gring VBIAS COL_OUT[62] ROW_SEL[99] VREF PIX_IN[9962] NB2 NB1 CSA_VREF pixel
xPix9963 VDD GND SF_IB gring VBIAS COL_OUT[63] ROW_SEL[99] VREF PIX_IN[9963] NB2 NB1 CSA_VREF pixel
xPix9964 VDD GND SF_IB gring VBIAS COL_OUT[64] ROW_SEL[99] VREF PIX_IN[9964] NB2 NB1 CSA_VREF pixel
xPix9965 VDD GND SF_IB gring VBIAS COL_OUT[65] ROW_SEL[99] VREF PIX_IN[9965] NB2 NB1 CSA_VREF pixel
xPix9966 VDD GND SF_IB gring VBIAS COL_OUT[66] ROW_SEL[99] VREF PIX_IN[9966] NB2 NB1 CSA_VREF pixel
xPix9967 VDD GND SF_IB gring VBIAS COL_OUT[67] ROW_SEL[99] VREF PIX_IN[9967] NB2 NB1 CSA_VREF pixel
xPix9968 VDD GND SF_IB gring VBIAS COL_OUT[68] ROW_SEL[99] VREF PIX_IN[9968] NB2 NB1 CSA_VREF pixel
xPix9969 VDD GND SF_IB gring VBIAS COL_OUT[69] ROW_SEL[99] VREF PIX_IN[9969] NB2 NB1 CSA_VREF pixel
xPix9970 VDD GND SF_IB gring VBIAS COL_OUT[70] ROW_SEL[99] VREF PIX_IN[9970] NB2 NB1 CSA_VREF pixel
xPix9971 VDD GND SF_IB gring VBIAS COL_OUT[71] ROW_SEL[99] VREF PIX_IN[9971] NB2 NB1 CSA_VREF pixel
xPix9972 VDD GND SF_IB gring VBIAS COL_OUT[72] ROW_SEL[99] VREF PIX_IN[9972] NB2 NB1 CSA_VREF pixel
xPix9973 VDD GND SF_IB gring VBIAS COL_OUT[73] ROW_SEL[99] VREF PIX_IN[9973] NB2 NB1 CSA_VREF pixel
xPix9974 VDD GND SF_IB gring VBIAS COL_OUT[74] ROW_SEL[99] VREF PIX_IN[9974] NB2 NB1 CSA_VREF pixel
xPix9975 VDD GND SF_IB gring VBIAS COL_OUT[75] ROW_SEL[99] VREF PIX_IN[9975] NB2 NB1 CSA_VREF pixel
xPix9976 VDD GND SF_IB gring VBIAS COL_OUT[76] ROW_SEL[99] VREF PIX_IN[9976] NB2 NB1 CSA_VREF pixel
xPix9977 VDD GND SF_IB gring VBIAS COL_OUT[77] ROW_SEL[99] VREF PIX_IN[9977] NB2 NB1 CSA_VREF pixel
xPix9978 VDD GND SF_IB gring VBIAS COL_OUT[78] ROW_SEL[99] VREF PIX_IN[9978] NB2 NB1 CSA_VREF pixel
xPix9979 VDD GND SF_IB gring VBIAS COL_OUT[79] ROW_SEL[99] VREF PIX_IN[9979] NB2 NB1 CSA_VREF pixel
xPix9980 VDD GND SF_IB gring VBIAS COL_OUT[80] ROW_SEL[99] VREF PIX_IN[9980] NB2 NB1 CSA_VREF pixel
xPix9981 VDD GND SF_IB gring VBIAS COL_OUT[81] ROW_SEL[99] VREF PIX_IN[9981] NB2 NB1 CSA_VREF pixel
xPix9982 VDD GND SF_IB gring VBIAS COL_OUT[82] ROW_SEL[99] VREF PIX_IN[9982] NB2 NB1 CSA_VREF pixel
xPix9983 VDD GND SF_IB gring VBIAS COL_OUT[83] ROW_SEL[99] VREF PIX_IN[9983] NB2 NB1 CSA_VREF pixel
xPix9984 VDD GND SF_IB gring VBIAS COL_OUT[84] ROW_SEL[99] VREF PIX_IN[9984] NB2 NB1 CSA_VREF pixel
xPix9985 VDD GND SF_IB gring VBIAS COL_OUT[85] ROW_SEL[99] VREF PIX_IN[9985] NB2 NB1 CSA_VREF pixel
xPix9986 VDD GND SF_IB gring VBIAS COL_OUT[86] ROW_SEL[99] VREF PIX_IN[9986] NB2 NB1 CSA_VREF pixel
xPix9987 VDD GND SF_IB gring VBIAS COL_OUT[87] ROW_SEL[99] VREF PIX_IN[9987] NB2 NB1 CSA_VREF pixel
xPix9988 VDD GND SF_IB gring VBIAS COL_OUT[88] ROW_SEL[99] VREF PIX_IN[9988] NB2 NB1 CSA_VREF pixel
xPix9989 VDD GND SF_IB gring VBIAS COL_OUT[89] ROW_SEL[99] VREF PIX_IN[9989] NB2 NB1 CSA_VREF pixel
xPix9990 VDD GND SF_IB gring VBIAS COL_OUT[90] ROW_SEL[99] VREF PIX_IN[9990] NB2 NB1 CSA_VREF pixel
xPix9991 VDD GND SF_IB gring VBIAS COL_OUT[91] ROW_SEL[99] VREF PIX_IN[9991] NB2 NB1 CSA_VREF pixel
xPix9992 VDD GND SF_IB gring VBIAS COL_OUT[92] ROW_SEL[99] VREF PIX_IN[9992] NB2 NB1 CSA_VREF pixel
xPix9993 VDD GND SF_IB gring VBIAS COL_OUT[93] ROW_SEL[99] VREF PIX_IN[9993] NB2 NB1 CSA_VREF pixel
xPix9994 VDD GND SF_IB gring VBIAS COL_OUT[94] ROW_SEL[99] VREF PIX_IN[9994] NB2 NB1 CSA_VREF pixel
xPix9995 VDD GND SF_IB gring VBIAS COL_OUT[95] ROW_SEL[99] VREF PIX_IN[9995] NB2 NB1 CSA_VREF pixel
xPix9996 VDD GND SF_IB gring VBIAS COL_OUT[96] ROW_SEL[99] VREF PIX_IN[9996] NB2 NB1 CSA_VREF pixel
xPix9997 VDD GND SF_IB gring VBIAS COL_OUT[97] ROW_SEL[99] VREF PIX_IN[9997] NB2 NB1 CSA_VREF pixel
xPix9998 VDD GND SF_IB gring VBIAS COL_OUT[98] ROW_SEL[99] VREF PIX_IN[9998] NB2 NB1 CSA_VREF pixel
xPix9999 VDD GND SF_IB gring VBIAS COL_OUT[99] ROW_SEL[99] VREF PIX_IN[9999] NB2 NB1 CSA_VREF pixel
XM0 COL_OUT[0] COL_SEL[0] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 COL_OUT[1] COL_SEL[1] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 COL_OUT[2] COL_SEL[2] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 COL_OUT[3] COL_SEL[3] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 COL_OUT[4] COL_SEL[4] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 COL_OUT[5] COL_SEL[5] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 COL_OUT[6] COL_SEL[6] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 COL_OUT[7] COL_SEL[7] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 COL_OUT[8] COL_SEL[8] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 COL_OUT[9] COL_SEL[9] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 COL_OUT[10] COL_SEL[10] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 COL_OUT[11] COL_SEL[11] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 COL_OUT[12] COL_SEL[12] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 COL_OUT[13] COL_SEL[13] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 COL_OUT[14] COL_SEL[14] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 COL_OUT[15] COL_SEL[15] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 COL_OUT[16] COL_SEL[16] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 COL_OUT[17] COL_SEL[17] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 COL_OUT[18] COL_SEL[18] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM19 COL_OUT[19] COL_SEL[19] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20 COL_OUT[20] COL_SEL[20] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21 COL_OUT[21] COL_SEL[21] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM22 COL_OUT[22] COL_SEL[22] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23 COL_OUT[23] COL_SEL[23] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 COL_OUT[24] COL_SEL[24] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM25 COL_OUT[25] COL_SEL[25] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM26 COL_OUT[26] COL_SEL[26] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM27 COL_OUT[27] COL_SEL[27] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM28 COL_OUT[28] COL_SEL[28] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM29 COL_OUT[29] COL_SEL[29] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM30 COL_OUT[30] COL_SEL[30] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM31 COL_OUT[31] COL_SEL[31] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM32 COL_OUT[32] COL_SEL[32] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM33 COL_OUT[33] COL_SEL[33] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM34 COL_OUT[34] COL_SEL[34] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM35 COL_OUT[35] COL_SEL[35] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM36 COL_OUT[36] COL_SEL[36] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM37 COL_OUT[37] COL_SEL[37] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM38 COL_OUT[38] COL_SEL[38] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM39 COL_OUT[39] COL_SEL[39] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM40 COL_OUT[40] COL_SEL[40] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM41 COL_OUT[41] COL_SEL[41] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM42 COL_OUT[42] COL_SEL[42] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM43 COL_OUT[43] COL_SEL[43] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM44 COL_OUT[44] COL_SEL[44] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM45 COL_OUT[45] COL_SEL[45] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM46 COL_OUT[46] COL_SEL[46] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM47 COL_OUT[47] COL_SEL[47] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM48 COL_OUT[48] COL_SEL[48] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM49 COL_OUT[49] COL_SEL[49] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM50 COL_OUT[50] COL_SEL[50] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM51 COL_OUT[51] COL_SEL[51] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM52 COL_OUT[52] COL_SEL[52] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM53 COL_OUT[53] COL_SEL[53] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM54 COL_OUT[54] COL_SEL[54] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM55 COL_OUT[55] COL_SEL[55] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM56 COL_OUT[56] COL_SEL[56] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM57 COL_OUT[57] COL_SEL[57] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM58 COL_OUT[58] COL_SEL[58] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM59 COL_OUT[59] COL_SEL[59] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM60 COL_OUT[60] COL_SEL[60] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM61 COL_OUT[61] COL_SEL[61] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM62 COL_OUT[62] COL_SEL[62] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM63 COL_OUT[63] COL_SEL[63] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM64 COL_OUT[64] COL_SEL[64] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM65 COL_OUT[65] COL_SEL[65] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM66 COL_OUT[66] COL_SEL[66] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM67 COL_OUT[67] COL_SEL[67] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM68 COL_OUT[68] COL_SEL[68] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM69 COL_OUT[69] COL_SEL[69] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM70 COL_OUT[70] COL_SEL[70] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM71 COL_OUT[71] COL_SEL[71] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM72 COL_OUT[72] COL_SEL[72] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM73 COL_OUT[73] COL_SEL[73] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM74 COL_OUT[74] COL_SEL[74] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM75 COL_OUT[75] COL_SEL[75] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM76 COL_OUT[76] COL_SEL[76] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM77 COL_OUT[77] COL_SEL[77] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM78 COL_OUT[78] COL_SEL[78] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM79 COL_OUT[79] COL_SEL[79] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM80 COL_OUT[80] COL_SEL[80] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM81 COL_OUT[81] COL_SEL[81] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM82 COL_OUT[82] COL_SEL[82] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM83 COL_OUT[83] COL_SEL[83] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM84 COL_OUT[84] COL_SEL[84] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM85 COL_OUT[85] COL_SEL[85] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM86 COL_OUT[86] COL_SEL[86] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM87 COL_OUT[87] COL_SEL[87] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM88 COL_OUT[88] COL_SEL[88] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM89 COL_OUT[89] COL_SEL[89] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM90 COL_OUT[90] COL_SEL[90] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM91 COL_OUT[91] COL_SEL[91] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM92 COL_OUT[92] COL_SEL[92] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM93 COL_OUT[93] COL_SEL[93] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM94 COL_OUT[94] COL_SEL[94] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM95 COL_OUT[95] COL_SEL[95] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM96 COL_OUT[96] COL_SEL[96] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM97 COL_OUT[97] COL_SEL[97] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM98 COL_OUT[98] COL_SEL[98] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM99 COL_OUT[99] COL_SEL[99] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  pixel/pixel.sym # of pins=12
** sym_path: /home/hni/TopmetalSe-Respin/xschem/pixel/pixel.sym
** sch_path: /home/hni/TopmetalSe-Respin/xschem/pixel/pixel.sch
.subckt pixel VDD GND SF_IB gring VBIAS pix_out ROW_SEL VREF AMP_IN NB2 NB1 CSA_VREF
*.PININFO pix_out:O SF_IB:I ROW_SEL:I VREF:I AMP_IN:I NB1:I CSA_VREF:I VBIAS:I NB2:I VDD:I GND:I gring:I
XM2 net2 ROW_SEL pix_out GND sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 GND AMP_OUT net1 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 SF_IB VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 VDD net1 net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 VDD net6 AMP_OUT GND sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net5 net5 net7 VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net8 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net7 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 AMP_OUT NB2 GND GND sky130_fd_pr__nfet_01v8_lvt L=1.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 net4 NB1 GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC3 AMP_IN AMP_OUT sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=1 m=1
XM4 net3 VREF net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 AMP_IN CSA_VREF AMP_OUT VDD sky130_fd_pr__pfet_01v8_lvt L=7.95 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net6 net5 net8 VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net5 VBIAS net3 GND sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net9 AMP_IN net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 net6 VBIAS net9 GND sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMD_4 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMD_1 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.65 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMD_2 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt L=3.35 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
