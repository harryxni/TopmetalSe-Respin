magic
tech sky130A
magscale 1 2
timestamp 1758069660
<< error_s >>
rect 39054 13636 39063 13637
rect 39341 13636 39350 13637
rect 115252 13636 115261 13637
rect 115539 13636 115548 13637
rect 191450 13636 191459 13637
rect 191737 13636 191746 13637
rect 267648 13636 267657 13637
rect 267935 13636 267944 13637
rect 39045 13619 39048 13628
rect 39054 13627 39110 13628
rect 39134 13627 39190 13628
rect 39214 13627 39270 13628
rect 39294 13627 39350 13628
rect 39356 13619 39359 13628
rect 115243 13619 115246 13628
rect 115252 13627 115308 13628
rect 115332 13627 115388 13628
rect 115412 13627 115468 13628
rect 115492 13627 115548 13628
rect 115554 13619 115557 13628
rect 191441 13619 191444 13628
rect 191450 13627 191506 13628
rect 191530 13627 191586 13628
rect 191610 13627 191666 13628
rect 191690 13627 191746 13628
rect 191752 13619 191755 13628
rect 267639 13619 267642 13628
rect 267648 13627 267704 13628
rect 267728 13627 267784 13628
rect 267808 13627 267864 13628
rect 267888 13627 267944 13628
rect 267950 13619 267953 13628
rect 207110 13568 207119 13569
rect 207157 13568 207166 13569
rect 208030 13568 208039 13569
rect 208077 13568 208086 13569
rect 207101 13559 207175 13560
rect 207101 13551 207110 13559
rect 207165 13557 207175 13559
rect 207166 13551 207175 13557
rect 208021 13559 208095 13560
rect 208021 13551 208030 13559
rect 208085 13551 208095 13559
rect 207165 13504 207166 13507
rect 208085 13504 208086 13551
rect 213274 13432 213276 13433
rect 213328 13432 213330 13433
rect 219806 13432 219815 13433
rect 219853 13432 219862 13433
rect 227074 13432 227083 13433
rect 227121 13432 227130 13433
rect 229190 13432 229192 13433
rect 229244 13432 229246 13433
rect 238114 13432 238123 13433
rect 238161 13432 238170 13433
rect 239494 13432 239496 13433
rect 239548 13432 239550 13433
rect 268934 13432 268943 13433
rect 268981 13432 268990 13433
rect 273166 13432 273175 13433
rect 273213 13432 273222 13433
rect 213265 13423 213339 13424
rect 213265 13415 213274 13423
rect 213329 13421 213339 13423
rect 213330 13415 213339 13421
rect 219797 13423 219871 13424
rect 219797 13415 219806 13423
rect 219861 13415 219871 13423
rect 227065 13423 227139 13424
rect 227065 13415 227074 13423
rect 227129 13421 227139 13423
rect 227130 13415 227139 13421
rect 229181 13423 229255 13424
rect 229181 13415 229190 13423
rect 229245 13415 229255 13423
rect 238105 13423 238179 13424
rect 238105 13415 238114 13423
rect 238169 13421 238179 13423
rect 238170 13415 238179 13421
rect 239485 13423 239559 13424
rect 239485 13415 239494 13423
rect 239549 13415 239559 13423
rect 268925 13423 268999 13424
rect 268925 13415 268934 13423
rect 268989 13421 268999 13423
rect 268990 13415 268999 13421
rect 273157 13423 273231 13424
rect 273157 13415 273166 13423
rect 273221 13415 273231 13423
rect 213329 13368 213330 13371
rect 219861 13368 219862 13415
rect 227129 13368 227130 13371
rect 229245 13368 229246 13415
rect 238169 13368 238170 13371
rect 239549 13368 239550 13415
rect 268989 13368 268990 13371
rect 273221 13368 273222 13415
rect 200854 13296 200863 13297
rect 200901 13296 200910 13297
rect 203430 13296 203439 13297
rect 203477 13296 203486 13297
rect 205546 13296 205555 13297
rect 205593 13296 205602 13297
rect 205730 13296 205739 13297
rect 205777 13296 205786 13297
rect 207202 13296 207204 13297
rect 207256 13296 207258 13297
rect 207938 13296 207940 13297
rect 207992 13296 207994 13297
rect 230386 13296 230388 13297
rect 230440 13296 230442 13297
rect 232134 13296 232143 13297
rect 232181 13296 232190 13297
rect 263414 13296 263423 13297
rect 263461 13296 263470 13297
rect 265530 13296 265539 13297
rect 265577 13296 265586 13297
rect 269026 13296 269035 13297
rect 269073 13296 269082 13297
rect 273258 13296 273260 13297
rect 273312 13296 273314 13297
rect 200845 13287 200919 13288
rect 200845 13279 200854 13287
rect 200909 13285 200919 13287
rect 200910 13279 200919 13285
rect 203421 13287 203495 13288
rect 203421 13279 203430 13287
rect 203485 13279 203495 13287
rect 205537 13287 205611 13288
rect 205537 13279 205546 13287
rect 205601 13285 205611 13287
rect 205602 13279 205611 13285
rect 205721 13287 205795 13288
rect 205721 13279 205730 13287
rect 205785 13279 205795 13287
rect 207193 13287 207267 13288
rect 207193 13279 207202 13287
rect 207257 13285 207267 13287
rect 207258 13279 207267 13285
rect 207929 13287 208003 13288
rect 207929 13279 207938 13287
rect 207993 13279 208003 13287
rect 230377 13287 230451 13288
rect 230377 13279 230386 13287
rect 230441 13285 230451 13287
rect 230442 13279 230451 13285
rect 232125 13287 232199 13288
rect 232125 13279 232134 13287
rect 232189 13279 232199 13287
rect 263405 13287 263479 13288
rect 263405 13279 263414 13287
rect 263469 13285 263479 13287
rect 263470 13279 263479 13285
rect 265521 13287 265595 13288
rect 265521 13279 265530 13287
rect 265585 13279 265595 13287
rect 269017 13287 269091 13288
rect 269017 13279 269026 13287
rect 269081 13285 269091 13287
rect 269082 13279 269091 13285
rect 273249 13287 273323 13288
rect 273249 13279 273258 13287
rect 273313 13279 273323 13287
rect 200909 13232 200910 13235
rect 203485 13232 203486 13279
rect 205601 13232 205602 13235
rect 205785 13232 205786 13279
rect 207257 13232 207258 13235
rect 207993 13232 207994 13279
rect 230441 13232 230442 13235
rect 232189 13232 232190 13279
rect 263469 13232 263470 13235
rect 265585 13232 265586 13279
rect 269081 13232 269082 13235
rect 273313 13232 273314 13279
rect 86958 13160 86967 13161
rect 87005 13160 87014 13161
rect 91834 13160 91843 13161
rect 91881 13160 91890 13161
rect 225418 13160 225420 13161
rect 225472 13160 225474 13161
rect 227074 13160 227076 13161
rect 227128 13160 227130 13161
rect 86949 13151 87023 13152
rect 86949 13143 86958 13151
rect 87013 13149 87023 13151
rect 87014 13143 87023 13149
rect 91825 13151 91899 13152
rect 91825 13143 91834 13151
rect 91889 13143 91899 13151
rect 225409 13151 225483 13152
rect 225409 13143 225418 13151
rect 225473 13149 225483 13151
rect 225474 13143 225483 13149
rect 227065 13151 227139 13152
rect 227065 13143 227074 13151
rect 227129 13143 227139 13151
rect 87013 13096 87014 13099
rect 91889 13096 91890 13143
rect 225473 13096 225474 13099
rect 227129 13096 227130 13143
rect 77154 13092 77163 13093
rect 77441 13092 77450 13093
rect 153352 13092 153361 13093
rect 153639 13092 153648 13093
rect 229550 13092 229559 13093
rect 229837 13092 229846 13093
rect 77145 13075 77148 13084
rect 77154 13083 77210 13084
rect 77234 13083 77290 13084
rect 77314 13083 77370 13084
rect 77394 13083 77450 13084
rect 77456 13075 77459 13084
rect 153343 13075 153346 13084
rect 153352 13083 153408 13084
rect 153432 13083 153488 13084
rect 153512 13083 153568 13084
rect 153592 13083 153648 13084
rect 153654 13075 153657 13084
rect 229541 13075 229544 13084
rect 229550 13083 229606 13084
rect 229630 13083 229686 13084
rect 229710 13083 229766 13084
rect 229790 13083 229846 13084
rect 229852 13075 229855 13084
rect 256606 13024 256615 13025
rect 256653 13024 256662 13025
rect 257986 13024 257995 13025
rect 258033 13024 258042 13025
rect 256597 13015 256671 13016
rect 256597 13007 256606 13015
rect 256661 13013 256671 13015
rect 256662 13007 256671 13013
rect 257977 13015 258051 13016
rect 257977 13007 257986 13015
rect 258041 13007 258051 13015
rect 256661 12960 256662 12963
rect 258041 12960 258042 13007
rect 155038 12888 155047 12889
rect 155085 12888 155094 12889
rect 194598 12888 194607 12889
rect 194645 12888 194654 12889
rect 195794 12888 195803 12889
rect 195841 12888 195850 12889
rect 197358 12888 197367 12889
rect 197405 12888 197414 12889
rect 299478 12888 299487 12889
rect 299525 12888 299534 12889
rect 155029 12879 155103 12880
rect 155029 12871 155038 12879
rect 155093 12877 155103 12879
rect 155094 12871 155103 12877
rect 194589 12879 194663 12880
rect 194589 12871 194598 12879
rect 194653 12877 194663 12879
rect 194654 12871 194663 12877
rect 195785 12879 195859 12880
rect 195785 12871 195794 12879
rect 195849 12871 195859 12879
rect 197349 12879 197423 12880
rect 197349 12871 197358 12879
rect 197413 12877 197423 12879
rect 197414 12871 197423 12877
rect 299469 12879 299543 12880
rect 299469 12871 299478 12879
rect 299533 12871 299543 12879
rect 155093 12824 155094 12827
rect 194653 12824 194654 12827
rect 195849 12824 195850 12871
rect 197413 12824 197414 12827
rect 299533 12824 299534 12871
rect 87786 12752 87795 12753
rect 87833 12752 87842 12753
rect 90730 12752 90739 12753
rect 90777 12752 90786 12753
rect 195058 12752 195067 12753
rect 195105 12752 195114 12753
rect 207846 12752 207855 12753
rect 207893 12752 207902 12753
rect 238298 12752 238307 12753
rect 238345 12752 238354 12753
rect 242162 12752 242171 12753
rect 242209 12752 242218 12753
rect 262310 12752 262312 12753
rect 262364 12752 262366 12753
rect 263506 12752 263515 12753
rect 263553 12752 263562 12753
rect 264334 12752 264343 12753
rect 264381 12752 264390 12753
rect 267094 12752 267103 12753
rect 267141 12752 267150 12753
rect 267646 12752 267655 12753
rect 267693 12752 267702 12753
rect 268106 12752 268115 12753
rect 268153 12752 268162 12753
rect 87777 12743 87851 12744
rect 87777 12735 87786 12743
rect 87841 12741 87851 12743
rect 87842 12735 87851 12741
rect 90721 12743 90795 12744
rect 90721 12735 90730 12743
rect 90785 12735 90795 12743
rect 195049 12743 195123 12744
rect 195049 12735 195058 12743
rect 195113 12741 195123 12743
rect 195114 12735 195123 12741
rect 207837 12743 207911 12744
rect 207837 12735 207846 12743
rect 207901 12735 207911 12743
rect 238289 12743 238363 12744
rect 238289 12735 238298 12743
rect 238353 12741 238363 12743
rect 238354 12735 238363 12741
rect 242153 12743 242227 12744
rect 242153 12735 242162 12743
rect 242217 12735 242227 12743
rect 262301 12743 262375 12744
rect 262301 12735 262310 12743
rect 262365 12741 262375 12743
rect 262366 12735 262375 12741
rect 263497 12743 263571 12744
rect 263497 12735 263506 12743
rect 263561 12735 263571 12743
rect 264325 12743 264399 12744
rect 264325 12735 264334 12743
rect 264389 12741 264399 12743
rect 264390 12735 264399 12741
rect 267085 12743 267159 12744
rect 267085 12735 267094 12743
rect 267149 12735 267159 12743
rect 267637 12743 267711 12744
rect 267637 12735 267646 12743
rect 267701 12741 267711 12743
rect 267702 12735 267711 12741
rect 268097 12743 268171 12744
rect 268097 12735 268106 12743
rect 268161 12735 268171 12743
rect 87841 12688 87842 12691
rect 90785 12688 90786 12735
rect 143305 12732 143306 12733
rect 143339 12722 143340 12733
rect 195113 12688 195114 12691
rect 207901 12688 207902 12735
rect 238353 12688 238354 12691
rect 242217 12688 242218 12735
rect 262365 12688 262366 12691
rect 263561 12688 263562 12735
rect 264389 12688 264390 12691
rect 267149 12688 267150 12735
rect 267701 12688 267702 12691
rect 268161 12688 268162 12735
rect 157890 12616 157892 12617
rect 157944 12616 157946 12617
rect 160282 12616 160284 12617
rect 160336 12616 160338 12617
rect 191838 12616 191847 12617
rect 191885 12616 191894 12617
rect 192206 12616 192215 12617
rect 192253 12616 192262 12617
rect 200394 12616 200403 12617
rect 200441 12616 200450 12617
rect 205270 12616 205272 12617
rect 205324 12616 205326 12617
rect 251914 12616 251916 12617
rect 251968 12616 251970 12617
rect 257066 12616 257075 12617
rect 257113 12616 257122 12617
rect 157881 12607 157955 12608
rect 157881 12599 157890 12607
rect 157945 12605 157955 12607
rect 157946 12599 157955 12605
rect 160273 12607 160347 12608
rect 160273 12599 160282 12607
rect 160337 12599 160347 12607
rect 191829 12607 191903 12608
rect 191829 12599 191838 12607
rect 191893 12605 191903 12607
rect 191894 12599 191903 12605
rect 192197 12607 192271 12608
rect 192197 12599 192206 12607
rect 192261 12599 192271 12607
rect 200385 12607 200459 12608
rect 200385 12599 200394 12607
rect 200449 12605 200459 12607
rect 200450 12599 200459 12605
rect 205261 12607 205335 12608
rect 205261 12599 205270 12607
rect 205325 12599 205335 12607
rect 251905 12607 251979 12608
rect 251905 12599 251914 12607
rect 251969 12605 251979 12607
rect 251970 12599 251979 12605
rect 257057 12607 257131 12608
rect 257057 12599 257066 12607
rect 257121 12599 257131 12607
rect 157945 12552 157946 12555
rect 160337 12552 160338 12599
rect 191893 12552 191894 12555
rect 192261 12552 192262 12599
rect 200449 12552 200450 12555
rect 205325 12552 205326 12599
rect 251969 12552 251970 12555
rect 257121 12552 257122 12599
rect 39054 12548 39063 12549
rect 39341 12548 39350 12549
rect 115252 12548 115261 12549
rect 115539 12548 115548 12549
rect 191450 12548 191459 12549
rect 191737 12548 191746 12549
rect 267648 12548 267657 12549
rect 267935 12548 267944 12549
rect 39045 12531 39048 12540
rect 39054 12539 39110 12540
rect 39134 12539 39190 12540
rect 39214 12539 39270 12540
rect 39294 12539 39350 12540
rect 39356 12531 39359 12540
rect 115243 12531 115246 12540
rect 115252 12539 115308 12540
rect 115332 12539 115388 12540
rect 115412 12539 115468 12540
rect 115492 12539 115548 12540
rect 115554 12531 115557 12540
rect 191441 12531 191444 12540
rect 191450 12539 191506 12540
rect 191530 12539 191586 12540
rect 191610 12539 191666 12540
rect 191690 12539 191746 12540
rect 191752 12531 191755 12540
rect 267639 12531 267642 12540
rect 267648 12539 267704 12540
rect 267728 12539 267784 12540
rect 267808 12539 267864 12540
rect 267888 12539 267944 12540
rect 267950 12531 267953 12540
rect 251822 12480 251831 12481
rect 251869 12480 251878 12481
rect 257158 12480 257167 12481
rect 257205 12480 257214 12481
rect 251813 12471 251887 12472
rect 251813 12463 251822 12471
rect 251877 12469 251887 12471
rect 251878 12463 251887 12469
rect 257149 12471 257223 12472
rect 257149 12463 257158 12471
rect 257213 12463 257223 12471
rect 251877 12416 251878 12419
rect 257213 12416 257214 12463
rect 88154 12344 88163 12345
rect 88201 12344 88210 12345
rect 89902 12344 89911 12345
rect 89949 12344 89958 12345
rect 163594 12344 163603 12345
rect 163641 12344 163650 12345
rect 193034 12344 193043 12345
rect 193081 12344 193090 12345
rect 88145 12335 88219 12336
rect 88145 12327 88154 12335
rect 88209 12333 88219 12335
rect 88210 12327 88219 12333
rect 89893 12335 89967 12336
rect 89893 12327 89902 12335
rect 89957 12327 89967 12335
rect 163585 12335 163659 12336
rect 163585 12327 163594 12335
rect 163649 12333 163659 12335
rect 163650 12327 163659 12333
rect 193025 12335 193099 12336
rect 193025 12327 193034 12335
rect 193089 12327 193099 12335
rect 88209 12280 88210 12283
rect 89957 12280 89958 12327
rect 163649 12280 163650 12283
rect 193089 12280 193090 12327
rect 29366 12208 29368 12209
rect 29420 12208 29422 12209
rect 30746 12208 30755 12209
rect 30793 12208 30802 12209
rect 31390 12208 31399 12209
rect 31437 12208 31446 12209
rect 40590 12208 40592 12209
rect 40644 12208 40646 12209
rect 42430 12208 42439 12209
rect 42477 12208 42486 12209
rect 29357 12199 29431 12200
rect 29357 12191 29366 12199
rect 29421 12197 29431 12199
rect 29422 12191 29431 12197
rect 30737 12199 30811 12200
rect 30737 12191 30746 12199
rect 30801 12197 30811 12199
rect 30802 12191 30811 12197
rect 31381 12199 31455 12200
rect 31381 12191 31390 12199
rect 31445 12191 31455 12199
rect 40581 12199 40655 12200
rect 40581 12191 40590 12199
rect 40645 12197 40655 12199
rect 40646 12191 40655 12197
rect 42421 12199 42495 12200
rect 42421 12191 42430 12199
rect 42485 12191 42495 12199
rect 29421 12144 29422 12147
rect 30801 12144 30802 12147
rect 31445 12144 31446 12191
rect 40645 12144 40646 12147
rect 42485 12144 42486 12191
rect 77154 12004 77163 12005
rect 77441 12004 77450 12005
rect 153352 12004 153361 12005
rect 153639 12004 153648 12005
rect 229550 12004 229559 12005
rect 229837 12004 229846 12005
rect 77145 11987 77148 11996
rect 77154 11995 77210 11996
rect 77234 11995 77290 11996
rect 77314 11995 77370 11996
rect 77394 11995 77450 11996
rect 77456 11987 77459 11996
rect 153343 11987 153346 11996
rect 153352 11995 153408 11996
rect 153432 11995 153488 11996
rect 153512 11995 153568 11996
rect 153592 11995 153648 11996
rect 153654 11987 153657 11996
rect 229541 11987 229544 11996
rect 229550 11995 229606 11996
rect 229630 11995 229686 11996
rect 229710 11995 229766 11996
rect 229790 11995 229846 11996
rect 229852 11987 229855 11996
rect 189630 11800 189639 11801
rect 189677 11800 189686 11801
rect 193034 11800 193043 11801
rect 193081 11800 193090 11801
rect 189621 11791 189695 11792
rect 189621 11783 189630 11791
rect 189685 11789 189695 11791
rect 189686 11783 189695 11789
rect 193025 11791 193099 11792
rect 193025 11783 193034 11791
rect 193089 11783 193099 11791
rect 189685 11736 189686 11739
rect 193089 11736 193090 11783
rect 231006 11703 231007 11753
rect 231040 11712 231041 11746
rect 39054 11460 39063 11461
rect 39341 11460 39350 11461
rect 115252 11460 115261 11461
rect 115539 11460 115548 11461
rect 191450 11460 191459 11461
rect 191737 11460 191746 11461
rect 267648 11460 267657 11461
rect 267935 11460 267944 11461
rect 39045 11443 39048 11452
rect 39054 11451 39110 11452
rect 39134 11451 39190 11452
rect 39214 11451 39270 11452
rect 39294 11451 39350 11452
rect 39356 11443 39359 11452
rect 115243 11443 115246 11452
rect 115252 11451 115308 11452
rect 115332 11451 115388 11452
rect 115412 11451 115468 11452
rect 115492 11451 115548 11452
rect 115554 11443 115557 11452
rect 191441 11443 191444 11452
rect 191450 11451 191506 11452
rect 191530 11451 191586 11452
rect 191610 11451 191666 11452
rect 191690 11451 191746 11452
rect 191752 11443 191755 11452
rect 267639 11443 267642 11452
rect 267648 11451 267704 11452
rect 267728 11451 267784 11452
rect 267808 11451 267864 11452
rect 267888 11451 267944 11452
rect 267950 11443 267953 11452
rect 190894 11095 190895 11145
rect 190928 11100 190929 11134
rect 140420 11032 140454 11033
rect 156060 11032 156094 11033
rect 140409 10998 140470 10999
rect 156049 10998 156110 10999
rect 77154 10916 77163 10917
rect 77441 10916 77450 10917
rect 153352 10916 153361 10917
rect 153639 10916 153648 10917
rect 229550 10916 229559 10917
rect 229837 10916 229846 10917
rect 77145 10899 77148 10908
rect 77154 10907 77210 10908
rect 77234 10907 77290 10908
rect 77314 10907 77370 10908
rect 77394 10907 77450 10908
rect 77456 10899 77459 10908
rect 153343 10899 153346 10908
rect 153352 10907 153408 10908
rect 153432 10907 153488 10908
rect 153512 10907 153568 10908
rect 153592 10907 153648 10908
rect 153654 10899 153657 10908
rect 229541 10899 229544 10908
rect 229550 10907 229606 10908
rect 229630 10907 229686 10908
rect 229710 10907 229766 10908
rect 229790 10907 229846 10908
rect 229852 10899 229855 10908
rect 269186 10615 269187 10665
rect 269220 10624 269221 10658
rect 187490 10522 187501 10557
rect 187524 10556 187535 10557
rect 39054 10372 39063 10373
rect 39341 10372 39350 10373
rect 115252 10372 115261 10373
rect 115539 10372 115548 10373
rect 191450 10372 191459 10373
rect 191737 10372 191746 10373
rect 267648 10372 267657 10373
rect 267935 10372 267944 10373
rect 39045 10355 39048 10364
rect 39054 10363 39110 10364
rect 39134 10363 39190 10364
rect 39214 10363 39270 10364
rect 39294 10363 39350 10364
rect 39356 10355 39359 10364
rect 115243 10355 115246 10364
rect 115252 10363 115308 10364
rect 115332 10363 115388 10364
rect 115412 10363 115468 10364
rect 115492 10363 115548 10364
rect 115554 10355 115557 10364
rect 191441 10355 191444 10364
rect 191450 10363 191506 10364
rect 191530 10363 191586 10364
rect 191610 10363 191666 10364
rect 191690 10363 191746 10364
rect 191752 10355 191755 10364
rect 267639 10355 267642 10364
rect 267648 10363 267704 10364
rect 267728 10363 267784 10364
rect 267808 10363 267864 10364
rect 267888 10363 267944 10364
rect 267950 10355 267953 10364
rect 304446 10032 304448 10033
rect 304500 10032 304502 10033
rect 304437 10023 304511 10024
rect 304437 10015 304446 10023
rect 304501 10021 304511 10023
rect 304502 10015 304511 10021
rect 304501 9968 304502 9971
rect 77154 9828 77163 9829
rect 77441 9828 77450 9829
rect 153352 9828 153361 9829
rect 153639 9828 153648 9829
rect 229550 9828 229559 9829
rect 229837 9828 229846 9829
rect 77145 9811 77148 9820
rect 77154 9819 77210 9820
rect 77234 9819 77290 9820
rect 77314 9819 77370 9820
rect 77394 9819 77450 9820
rect 77456 9811 77459 9820
rect 153343 9811 153346 9820
rect 153352 9819 153408 9820
rect 153432 9819 153488 9820
rect 153512 9819 153568 9820
rect 153592 9819 153648 9820
rect 153654 9811 153657 9820
rect 229541 9811 229544 9820
rect 229550 9819 229606 9820
rect 229630 9819 229686 9820
rect 229710 9819 229766 9820
rect 229790 9819 229846 9820
rect 229852 9811 229855 9820
rect 39054 9284 39063 9285
rect 39341 9284 39350 9285
rect 115252 9284 115261 9285
rect 115539 9284 115548 9285
rect 191450 9284 191459 9285
rect 191737 9284 191746 9285
rect 267648 9284 267657 9285
rect 267935 9284 267944 9285
rect 39045 9267 39048 9276
rect 39054 9275 39110 9276
rect 39134 9275 39190 9276
rect 39214 9275 39270 9276
rect 39294 9275 39350 9276
rect 39356 9267 39359 9276
rect 115243 9267 115246 9276
rect 115252 9275 115308 9276
rect 115332 9275 115388 9276
rect 115412 9275 115468 9276
rect 115492 9275 115548 9276
rect 115554 9267 115557 9276
rect 191441 9267 191444 9276
rect 191450 9275 191506 9276
rect 191530 9275 191586 9276
rect 191610 9275 191666 9276
rect 191690 9275 191746 9276
rect 191752 9267 191755 9276
rect 267639 9267 267642 9276
rect 267648 9275 267704 9276
rect 267728 9275 267784 9276
rect 267808 9275 267864 9276
rect 267888 9275 267944 9276
rect 267950 9267 267953 9276
rect 77154 8740 77163 8741
rect 77441 8740 77450 8741
rect 153352 8740 153361 8741
rect 153639 8740 153648 8741
rect 229550 8740 229559 8741
rect 229837 8740 229846 8741
rect 77145 8723 77148 8732
rect 77154 8731 77210 8732
rect 77234 8731 77290 8732
rect 77314 8731 77370 8732
rect 77394 8731 77450 8732
rect 77456 8723 77459 8732
rect 153343 8723 153346 8732
rect 153352 8731 153408 8732
rect 153432 8731 153488 8732
rect 153512 8731 153568 8732
rect 153592 8731 153648 8732
rect 153654 8723 153657 8732
rect 229541 8723 229544 8732
rect 229550 8731 229606 8732
rect 229630 8731 229686 8732
rect 229710 8731 229766 8732
rect 229790 8731 229846 8732
rect 229852 8723 229855 8732
rect 39054 8196 39063 8197
rect 39341 8196 39350 8197
rect 115252 8196 115261 8197
rect 115539 8196 115548 8197
rect 191450 8196 191459 8197
rect 191737 8196 191746 8197
rect 267648 8196 267657 8197
rect 267935 8196 267944 8197
rect 39045 8179 39048 8188
rect 39054 8187 39110 8188
rect 39134 8187 39190 8188
rect 39214 8187 39270 8188
rect 39294 8187 39350 8188
rect 39356 8179 39359 8188
rect 115243 8179 115246 8188
rect 115252 8187 115308 8188
rect 115332 8187 115388 8188
rect 115412 8187 115468 8188
rect 115492 8187 115548 8188
rect 115554 8179 115557 8188
rect 191441 8179 191444 8188
rect 191450 8187 191506 8188
rect 191530 8187 191586 8188
rect 191610 8187 191666 8188
rect 191690 8187 191746 8188
rect 191752 8179 191755 8188
rect 267639 8179 267642 8188
rect 267648 8187 267704 8188
rect 267728 8187 267784 8188
rect 267808 8187 267864 8188
rect 267888 8187 267944 8188
rect 267950 8179 267953 8188
rect 77154 7652 77163 7653
rect 77441 7652 77450 7653
rect 153352 7652 153361 7653
rect 153639 7652 153648 7653
rect 229550 7652 229559 7653
rect 229837 7652 229846 7653
rect 77145 7635 77148 7644
rect 77154 7643 77210 7644
rect 77234 7643 77290 7644
rect 77314 7643 77370 7644
rect 77394 7643 77450 7644
rect 77456 7635 77459 7644
rect 153343 7635 153346 7644
rect 153352 7643 153408 7644
rect 153432 7643 153488 7644
rect 153512 7643 153568 7644
rect 153592 7643 153648 7644
rect 153654 7635 153657 7644
rect 229541 7635 229544 7644
rect 229550 7643 229606 7644
rect 229630 7643 229686 7644
rect 229710 7643 229766 7644
rect 229790 7643 229846 7644
rect 229852 7635 229855 7644
rect 39054 7108 39063 7109
rect 39341 7108 39350 7109
rect 115252 7108 115261 7109
rect 115539 7108 115548 7109
rect 191450 7108 191459 7109
rect 191737 7108 191746 7109
rect 267648 7108 267657 7109
rect 267935 7108 267944 7109
rect 39045 7091 39048 7100
rect 39054 7099 39110 7100
rect 39134 7099 39190 7100
rect 39214 7099 39270 7100
rect 39294 7099 39350 7100
rect 39356 7091 39359 7100
rect 115243 7091 115246 7100
rect 115252 7099 115308 7100
rect 115332 7099 115388 7100
rect 115412 7099 115468 7100
rect 115492 7099 115548 7100
rect 115554 7091 115557 7100
rect 191441 7091 191444 7100
rect 191450 7099 191506 7100
rect 191530 7099 191586 7100
rect 191610 7099 191666 7100
rect 191690 7099 191746 7100
rect 191752 7091 191755 7100
rect 267639 7091 267642 7100
rect 267648 7099 267704 7100
rect 267728 7099 267784 7100
rect 267808 7099 267864 7100
rect 267888 7099 267944 7100
rect 267950 7091 267953 7100
rect 77154 6564 77163 6565
rect 77441 6564 77450 6565
rect 153352 6564 153361 6565
rect 153639 6564 153648 6565
rect 229550 6564 229559 6565
rect 229837 6564 229846 6565
rect 77145 6547 77148 6556
rect 77154 6555 77210 6556
rect 77234 6555 77290 6556
rect 77314 6555 77370 6556
rect 77394 6555 77450 6556
rect 77456 6547 77459 6556
rect 153343 6547 153346 6556
rect 153352 6555 153408 6556
rect 153432 6555 153488 6556
rect 153512 6555 153568 6556
rect 153592 6555 153648 6556
rect 153654 6547 153657 6556
rect 229541 6547 229544 6556
rect 229550 6555 229606 6556
rect 229630 6555 229686 6556
rect 229710 6555 229766 6556
rect 229790 6555 229846 6556
rect 229852 6547 229855 6556
rect 304238 6170 304249 6205
rect 304272 6204 304283 6205
rect 39054 6020 39063 6021
rect 39341 6020 39350 6021
rect 115252 6020 115261 6021
rect 115539 6020 115548 6021
rect 191450 6020 191459 6021
rect 191737 6020 191746 6021
rect 267648 6020 267657 6021
rect 267935 6020 267944 6021
rect 39045 6003 39048 6012
rect 39054 6011 39110 6012
rect 39134 6011 39190 6012
rect 39214 6011 39270 6012
rect 39294 6011 39350 6012
rect 39356 6003 39359 6012
rect 115243 6003 115246 6012
rect 115252 6011 115308 6012
rect 115332 6011 115388 6012
rect 115412 6011 115468 6012
rect 115492 6011 115548 6012
rect 115554 6003 115557 6012
rect 191441 6003 191444 6012
rect 191450 6011 191506 6012
rect 191530 6011 191586 6012
rect 191610 6011 191666 6012
rect 191690 6011 191746 6012
rect 191752 6003 191755 6012
rect 267639 6003 267642 6012
rect 267648 6011 267704 6012
rect 267728 6011 267784 6012
rect 267808 6011 267864 6012
rect 267888 6011 267944 6012
rect 267950 6003 267953 6012
rect 303986 5952 303995 5953
rect 304033 5952 304042 5953
rect 303977 5943 304051 5944
rect 303977 5935 303986 5943
rect 304041 5941 304051 5943
rect 304042 5935 304051 5941
rect 304041 5888 304042 5891
rect 77154 5476 77163 5477
rect 77441 5476 77450 5477
rect 153352 5476 153361 5477
rect 153639 5476 153648 5477
rect 229550 5476 229559 5477
rect 229837 5476 229846 5477
rect 77145 5459 77148 5468
rect 77154 5467 77210 5468
rect 77234 5467 77290 5468
rect 77314 5467 77370 5468
rect 77394 5467 77450 5468
rect 77456 5459 77459 5468
rect 153343 5459 153346 5468
rect 153352 5467 153408 5468
rect 153432 5467 153488 5468
rect 153512 5467 153568 5468
rect 153592 5467 153648 5468
rect 153654 5459 153657 5468
rect 229541 5459 229544 5468
rect 229550 5467 229606 5468
rect 229630 5467 229686 5468
rect 229710 5467 229766 5468
rect 229790 5467 229846 5468
rect 229852 5459 229855 5468
rect 39054 4932 39063 4933
rect 39341 4932 39350 4933
rect 115252 4932 115261 4933
rect 115539 4932 115548 4933
rect 191450 4932 191459 4933
rect 191737 4932 191746 4933
rect 267648 4932 267657 4933
rect 267935 4932 267944 4933
rect 39045 4915 39048 4924
rect 39054 4923 39110 4924
rect 39134 4923 39190 4924
rect 39214 4923 39270 4924
rect 39294 4923 39350 4924
rect 39356 4915 39359 4924
rect 115243 4915 115246 4924
rect 115252 4923 115308 4924
rect 115332 4923 115388 4924
rect 115412 4923 115468 4924
rect 115492 4923 115548 4924
rect 115554 4915 115557 4924
rect 191441 4915 191444 4924
rect 191450 4923 191506 4924
rect 191530 4923 191586 4924
rect 191610 4923 191666 4924
rect 191690 4923 191746 4924
rect 191752 4915 191755 4924
rect 267639 4915 267642 4924
rect 267648 4923 267704 4924
rect 267728 4923 267784 4924
rect 267808 4923 267864 4924
rect 267888 4923 267944 4924
rect 267950 4915 267953 4924
rect 77154 4388 77163 4389
rect 77441 4388 77450 4389
rect 153352 4388 153361 4389
rect 153639 4388 153648 4389
rect 229550 4388 229559 4389
rect 229837 4388 229846 4389
rect 77145 4371 77148 4380
rect 77154 4379 77210 4380
rect 77234 4379 77290 4380
rect 77314 4379 77370 4380
rect 77394 4379 77450 4380
rect 77456 4371 77459 4380
rect 153343 4371 153346 4380
rect 153352 4379 153408 4380
rect 153432 4379 153488 4380
rect 153512 4379 153568 4380
rect 153592 4379 153648 4380
rect 153654 4371 153657 4380
rect 229541 4371 229544 4380
rect 229550 4379 229606 4380
rect 229630 4379 229686 4380
rect 229710 4379 229766 4380
rect 229790 4379 229846 4380
rect 229852 4371 229855 4380
rect 39054 3844 39063 3845
rect 39341 3844 39350 3845
rect 115252 3844 115261 3845
rect 115539 3844 115548 3845
rect 191450 3844 191459 3845
rect 191737 3844 191746 3845
rect 267648 3844 267657 3845
rect 267935 3844 267944 3845
rect 39045 3827 39048 3836
rect 39054 3835 39110 3836
rect 39134 3835 39190 3836
rect 39214 3835 39270 3836
rect 39294 3835 39350 3836
rect 39356 3827 39359 3836
rect 115243 3827 115246 3836
rect 115252 3835 115308 3836
rect 115332 3835 115388 3836
rect 115412 3835 115468 3836
rect 115492 3835 115548 3836
rect 115554 3827 115557 3836
rect 191441 3827 191444 3836
rect 191450 3835 191506 3836
rect 191530 3835 191586 3836
rect 191610 3835 191666 3836
rect 191690 3835 191746 3836
rect 191752 3827 191755 3836
rect 267639 3827 267642 3836
rect 267648 3835 267704 3836
rect 267728 3835 267784 3836
rect 267808 3835 267864 3836
rect 267888 3835 267944 3836
rect 267950 3827 267953 3836
rect 77154 3300 77163 3301
rect 77441 3300 77450 3301
rect 153352 3300 153361 3301
rect 153639 3300 153648 3301
rect 229550 3300 229559 3301
rect 229837 3300 229846 3301
rect 77145 3283 77148 3292
rect 77154 3291 77210 3292
rect 77234 3291 77290 3292
rect 77314 3291 77370 3292
rect 77394 3291 77450 3292
rect 77456 3283 77459 3292
rect 153343 3283 153346 3292
rect 153352 3291 153408 3292
rect 153432 3291 153488 3292
rect 153512 3291 153568 3292
rect 153592 3291 153648 3292
rect 153654 3283 153657 3292
rect 229541 3283 229544 3292
rect 229550 3291 229606 3292
rect 229630 3291 229686 3292
rect 229710 3291 229766 3292
rect 229790 3291 229846 3292
rect 229852 3283 229855 3292
rect 39054 2756 39063 2757
rect 39341 2756 39350 2757
rect 115252 2756 115261 2757
rect 115539 2756 115548 2757
rect 191450 2756 191459 2757
rect 191737 2756 191746 2757
rect 267648 2756 267657 2757
rect 267935 2756 267944 2757
rect 39045 2739 39048 2748
rect 39054 2747 39110 2748
rect 39134 2747 39190 2748
rect 39214 2747 39270 2748
rect 39294 2747 39350 2748
rect 39356 2739 39359 2748
rect 115243 2739 115246 2748
rect 115252 2747 115308 2748
rect 115332 2747 115388 2748
rect 115412 2747 115468 2748
rect 115492 2747 115548 2748
rect 115554 2739 115557 2748
rect 191441 2739 191444 2748
rect 191450 2747 191506 2748
rect 191530 2747 191586 2748
rect 191610 2747 191666 2748
rect 191690 2747 191746 2748
rect 191752 2739 191755 2748
rect 267639 2739 267642 2748
rect 267648 2747 267704 2748
rect 267728 2747 267784 2748
rect 267808 2747 267864 2748
rect 267888 2747 267944 2748
rect 267950 2739 267953 2748
rect 77154 2212 77163 2213
rect 77441 2212 77450 2213
rect 153352 2212 153361 2213
rect 153639 2212 153648 2213
rect 229550 2212 229559 2213
rect 229837 2212 229846 2213
rect 77145 2195 77148 2204
rect 77154 2203 77210 2204
rect 77234 2203 77290 2204
rect 77314 2203 77370 2204
rect 77394 2203 77450 2204
rect 77456 2195 77459 2204
rect 153343 2195 153346 2204
rect 153352 2203 153408 2204
rect 153432 2203 153488 2204
rect 153512 2203 153568 2204
rect 153592 2203 153648 2204
rect 153654 2195 153657 2204
rect 229541 2195 229544 2204
rect 229550 2203 229606 2204
rect 229630 2203 229686 2204
rect 229710 2203 229766 2204
rect 229790 2203 229846 2204
rect 229852 2195 229855 2204
rect 302238 2008 302247 2009
rect 302285 2008 302294 2009
rect 302229 1999 302303 2000
rect 302229 1991 302238 1999
rect 302293 1997 302303 1999
rect 302294 1991 302303 1997
rect 302293 1944 302294 1947
<< viali >>
rect 1592 13480 1626 13514
rect 4628 13480 4662 13514
rect 7664 13480 7698 13514
rect 10792 13480 10826 13514
rect 14104 13480 14138 13514
rect 16864 13480 16898 13514
rect 19992 13480 20026 13514
rect 23028 13480 23062 13514
rect 25696 13480 25730 13514
rect 29008 13480 29042 13514
rect 31584 13480 31618 13514
rect 47592 13480 47626 13514
rect 50352 13480 50386 13514
rect 50996 13480 51030 13514
rect 142904 13480 142938 13514
rect 144744 13480 144778 13514
rect 148320 13480 148354 13514
rect 157624 13480 157658 13514
rect 182740 13480 182774 13514
rect 185776 13480 185810 13514
rect 210340 13480 210374 13514
rect 213376 13480 213410 13514
rect 269392 13480 269426 13514
rect 274280 13480 274314 13514
rect 274924 13480 274958 13514
rect 277868 13480 277902 13514
rect 280904 13480 280938 13514
rect 284584 13480 284618 13514
rect 287160 13480 287194 13514
rect 290104 13480 290138 13514
rect 293232 13480 293266 13514
rect 296268 13480 296302 13514
rect 299304 13480 299338 13514
rect 301420 13480 301454 13514
rect 301788 13480 301822 13514
rect 302156 13480 302190 13514
rect 302984 13480 303018 13514
rect 303352 13480 303386 13514
rect 44280 13412 44314 13446
rect 60472 13412 60506 13446
rect 63048 13412 63082 13446
rect 75376 13412 75410 13446
rect 93960 13412 93994 13446
rect 101136 13412 101170 13446
rect 109416 13412 109450 13446
rect 111256 13412 111290 13446
rect 121284 13412 121318 13446
rect 124136 13412 124170 13446
rect 136648 13412 136682 13446
rect 140328 13412 140362 13446
rect 155784 13412 155818 13446
rect 170412 13412 170446 13446
rect 173080 13412 173114 13446
rect 173816 13412 173850 13446
rect 175840 13412 175874 13446
rect 178140 13412 178174 13446
rect 181544 13412 181578 13446
rect 199852 13412 199886 13446
rect 203900 13412 203934 13446
rect 216412 13412 216446 13446
rect 220184 13412 220218 13446
rect 226624 13412 226658 13446
rect 229660 13412 229694 13446
rect 239964 13412 239998 13446
rect 247140 13412 247174 13446
rect 249532 13412 249566 13446
rect 252844 13412 252878 13446
rect 255420 13412 255454 13446
rect 259468 13412 259502 13446
rect 262688 13412 262722 13446
rect 266000 13412 266034 13446
rect 26340 13344 26374 13378
rect 27260 13344 27294 13378
rect 34712 13344 34746 13378
rect 37564 13344 37598 13378
rect 45568 13344 45602 13378
rect 51640 13344 51674 13378
rect 72708 13344 72742 13378
rect 73628 13344 73662 13378
rect 78504 13344 78538 13378
rect 80252 13344 80286 13378
rect 81540 13344 81574 13378
rect 81632 13344 81666 13378
rect 98008 13344 98042 13378
rect 98192 13344 98226 13378
rect 112268 13344 112302 13378
rect 120272 13344 120306 13378
rect 125700 13344 125734 13378
rect 126712 13344 126746 13378
rect 130300 13344 130334 13378
rect 132600 13344 132634 13378
rect 148056 13344 148090 13378
rect 150908 13344 150942 13378
rect 153484 13344 153518 13378
rect 160936 13344 160970 13378
rect 166640 13344 166674 13378
rect 167560 13344 167594 13378
rect 174276 13344 174310 13378
rect 174368 13344 174402 13378
rect 178968 13344 179002 13378
rect 182096 13344 182130 13378
rect 188536 13344 188570 13378
rect 189824 13344 189858 13378
rect 198748 13344 198782 13378
rect 201140 13344 201174 13378
rect 204728 13344 204762 13378
rect 207856 13344 207890 13378
rect 224324 13344 224358 13378
rect 227084 13344 227118 13378
rect 227176 13344 227210 13378
rect 230488 13344 230522 13378
rect 232236 13344 232270 13378
rect 237204 13344 237238 13378
rect 237296 13344 237330 13378
rect 240792 13344 240826 13378
rect 243368 13344 243402 13378
rect 245116 13344 245150 13378
rect 250176 13344 250210 13378
rect 262044 13344 262078 13378
rect 263240 13344 263274 13378
rect 266552 13344 266586 13378
rect 269128 13344 269162 13378
rect 271704 13344 271738 13378
rect 304456 13344 304490 13378
rect 304916 13344 304950 13378
rect 305376 13344 305410 13378
rect 1776 13276 1810 13310
rect 4812 13276 4846 13310
rect 7848 13276 7882 13310
rect 10976 13276 11010 13310
rect 14288 13276 14322 13310
rect 17048 13276 17082 13310
rect 20176 13276 20210 13310
rect 23212 13276 23246 13310
rect 26064 13276 26098 13310
rect 29836 13276 29870 13310
rect 32412 13276 32446 13310
rect 40140 13276 40174 13310
rect 42532 13276 42566 13310
rect 47776 13276 47810 13310
rect 50536 13276 50570 13310
rect 51364 13276 51398 13310
rect 53020 13276 53054 13310
rect 55596 13276 55630 13310
rect 57896 13276 57930 13310
rect 60656 13276 60690 13310
rect 63232 13276 63266 13310
rect 66176 13276 66210 13310
rect 69304 13276 69338 13310
rect 72524 13276 72558 13310
rect 76204 13276 76238 13310
rect 82460 13276 82494 13310
rect 83104 13276 83138 13310
rect 83932 13276 83966 13310
rect 86508 13276 86542 13310
rect 88808 13276 88842 13310
rect 94144 13276 94178 13310
rect 96904 13276 96938 13310
rect 99388 13276 99422 13310
rect 101964 13276 101998 13310
rect 104264 13276 104298 13310
rect 109600 13276 109634 13310
rect 111440 13276 111474 13310
rect 114844 13276 114878 13310
rect 117420 13276 117454 13310
rect 120180 13276 120214 13310
rect 121468 13276 121502 13310
rect 124320 13276 124354 13310
rect 126620 13276 126654 13310
rect 127540 13276 127574 13310
rect 136832 13276 136866 13310
rect 140512 13276 140546 13310
rect 143088 13276 143122 13310
rect 144928 13276 144962 13310
rect 145756 13276 145790 13310
rect 155968 13276 156002 13310
rect 156428 13276 156462 13310
rect 157808 13276 157842 13310
rect 158636 13276 158670 13310
rect 163512 13276 163546 13310
rect 170596 13276 170630 13310
rect 173264 13276 173298 13310
rect 174184 13276 174218 13310
rect 175656 13276 175690 13310
rect 176392 13276 176426 13310
rect 182004 13276 182038 13310
rect 182924 13276 182958 13310
rect 185960 13276 185994 13310
rect 187340 13276 187374 13310
rect 188444 13276 188478 13310
rect 189548 13276 189582 13310
rect 191848 13276 191882 13310
rect 194424 13276 194458 13310
rect 200036 13276 200070 13310
rect 202152 13276 202186 13310
rect 207672 13276 207706 13310
rect 210524 13276 210558 13310
rect 213560 13276 213594 13310
rect 216596 13276 216630 13310
rect 220368 13276 220402 13310
rect 222944 13276 222978 13310
rect 225888 13276 225922 13310
rect 227912 13276 227946 13310
rect 233064 13276 233098 13310
rect 233892 13276 233926 13310
rect 235088 13276 235122 13310
rect 237112 13276 237146 13310
rect 238216 13276 238250 13310
rect 247324 13276 247358 13310
rect 249992 13276 250026 13310
rect 251096 13276 251130 13310
rect 253672 13276 253706 13310
rect 256248 13276 256282 13310
rect 259652 13276 259686 13310
rect 264252 13276 264286 13310
rect 268576 13276 268610 13310
rect 274464 13276 274498 13310
rect 275108 13276 275142 13310
rect 278052 13276 278086 13310
rect 281088 13276 281122 13310
rect 284768 13276 284802 13310
rect 287344 13276 287378 13310
rect 290288 13276 290322 13310
rect 293416 13276 293450 13310
rect 296452 13276 296486 13310
rect 299488 13276 299522 13310
rect 303720 13276 303754 13310
rect 27536 13208 27570 13242
rect 30112 13208 30146 13242
rect 32688 13208 32722 13242
rect 34988 13208 35022 13242
rect 37840 13208 37874 13242
rect 40416 13208 40450 13242
rect 42808 13208 42842 13242
rect 45476 13208 45510 13242
rect 53296 13208 53330 13242
rect 55872 13208 55906 13242
rect 58172 13208 58206 13242
rect 73904 13208 73938 13242
rect 76480 13208 76514 13242
rect 78780 13208 78814 13242
rect 84208 13208 84242 13242
rect 86784 13208 86818 13242
rect 89084 13208 89118 13242
rect 91844 13208 91878 13242
rect 92028 13208 92062 13242
rect 99664 13208 99698 13242
rect 102240 13208 102274 13242
rect 104540 13208 104574 13242
rect 112544 13208 112578 13242
rect 115120 13208 115154 13242
rect 117696 13208 117730 13242
rect 120088 13208 120122 13242
rect 125516 13208 125550 13242
rect 127816 13208 127850 13242
rect 130576 13208 130610 13242
rect 132876 13208 132910 13242
rect 146032 13208 146066 13242
rect 150080 13208 150114 13242
rect 151184 13208 151218 13242
rect 153760 13208 153794 13242
rect 156520 13208 156554 13242
rect 158912 13208 158946 13242
rect 161212 13208 161246 13242
rect 163788 13208 163822 13242
rect 166548 13208 166582 13242
rect 167376 13208 167410 13242
rect 176668 13208 176702 13242
rect 179244 13208 179278 13242
rect 181912 13208 181946 13242
rect 187432 13208 187466 13242
rect 192124 13208 192158 13242
rect 193872 13208 193906 13242
rect 194700 13208 194734 13242
rect 196448 13208 196482 13242
rect 197828 13208 197862 13242
rect 198656 13208 198690 13242
rect 202428 13208 202462 13242
rect 205004 13208 205038 13242
rect 228188 13208 228222 13242
rect 230764 13208 230798 13242
rect 238492 13208 238526 13242
rect 241068 13208 241102 13242
rect 243644 13208 243678 13242
rect 251372 13208 251406 13242
rect 253948 13208 253982 13242
rect 256524 13208 256558 13242
rect 261860 13208 261894 13242
rect 263056 13208 263090 13242
rect 264528 13208 264562 13242
rect 266828 13208 266862 13242
rect 271980 13208 272014 13242
rect 26156 13140 26190 13174
rect 34160 13140 34194 13174
rect 36460 13140 36494 13174
rect 39312 13140 39346 13174
rect 41888 13140 41922 13174
rect 45016 13140 45050 13174
rect 45384 13140 45418 13174
rect 51456 13140 51490 13174
rect 54768 13140 54802 13174
rect 57344 13140 57378 13174
rect 59644 13140 59678 13174
rect 65992 13140 66026 13174
rect 69120 13140 69154 13174
rect 72064 13140 72098 13174
rect 72432 13140 72466 13174
rect 77952 13140 77986 13174
rect 81080 13140 81114 13174
rect 81448 13140 81482 13174
rect 82276 13140 82310 13174
rect 82920 13140 82954 13174
rect 85680 13140 85714 13174
rect 88256 13140 88290 13174
rect 90556 13140 90590 13174
rect 96720 13140 96754 13174
rect 97548 13140 97582 13174
rect 97916 13140 97950 13174
rect 103712 13140 103746 13174
rect 106012 13140 106046 13174
rect 114016 13140 114050 13174
rect 116592 13140 116626 13174
rect 119168 13140 119202 13174
rect 119720 13140 119754 13174
rect 126160 13140 126194 13174
rect 126528 13140 126562 13174
rect 129288 13140 129322 13174
rect 132048 13140 132082 13174
rect 134348 13140 134382 13174
rect 147504 13140 147538 13174
rect 152656 13140 152690 13174
rect 155232 13140 155266 13174
rect 160384 13140 160418 13174
rect 162684 13140 162718 13174
rect 165260 13140 165294 13174
rect 166088 13140 166122 13174
rect 166456 13140 166490 13174
rect 180716 13140 180750 13174
rect 187984 13140 188018 13174
rect 188352 13140 188386 13174
rect 191296 13140 191330 13174
rect 198196 13140 198230 13174
rect 198564 13140 198598 13174
rect 200496 13140 200530 13174
rect 200864 13140 200898 13174
rect 200956 13140 200990 13174
rect 206476 13140 206510 13174
rect 207304 13140 207338 13174
rect 207764 13140 207798 13174
rect 222760 13140 222794 13174
rect 223680 13140 223714 13174
rect 224048 13140 224082 13174
rect 224140 13140 224174 13174
rect 225704 13140 225738 13174
rect 226992 13140 227026 13174
rect 233156 13140 233190 13174
rect 233708 13140 233742 13174
rect 234904 13140 234938 13174
rect 236744 13140 236778 13174
rect 242540 13140 242574 13174
rect 249900 13140 249934 13174
rect 257996 13140 258030 13174
rect 263148 13140 263182 13174
rect 270876 13140 270910 13174
rect 273452 13140 273486 13174
rect 295900 13140 295934 13174
rect 26064 12936 26098 12970
rect 27444 12936 27478 12970
rect 33884 12936 33918 12970
rect 34804 12936 34838 12970
rect 35540 12936 35574 12970
rect 36644 12936 36678 12970
rect 42532 12936 42566 12970
rect 43452 12936 43486 12970
rect 44556 12936 44590 12970
rect 52008 12936 52042 12970
rect 53572 12936 53606 12970
rect 53940 12936 53974 12970
rect 58540 12936 58574 12970
rect 72156 12936 72190 12970
rect 89544 12936 89578 12970
rect 91108 12936 91142 12970
rect 112268 12936 112302 12970
rect 118248 12936 118282 12970
rect 118708 12936 118742 12970
rect 126712 12936 126746 12970
rect 128092 12936 128126 12970
rect 128736 12936 128770 12970
rect 129196 12936 129230 12970
rect 130300 12936 130334 12970
rect 133520 12936 133554 12970
rect 134348 12936 134382 12970
rect 145480 12936 145514 12970
rect 151460 12936 151494 12970
rect 152748 12936 152782 12970
rect 153116 12936 153150 12970
rect 153484 12936 153518 12970
rect 153852 12936 153886 12970
rect 154220 12936 154254 12970
rect 154956 12936 154990 12970
rect 156060 12936 156094 12970
rect 156428 12936 156462 12970
rect 156796 12936 156830 12970
rect 157164 12936 157198 12970
rect 163604 12936 163638 12970
rect 164432 12936 164466 12970
rect 167836 12936 167870 12970
rect 175012 12936 175046 12970
rect 175656 12936 175690 12970
rect 180808 12936 180842 12970
rect 192308 12936 192342 12970
rect 195988 12936 196022 12970
rect 206568 12936 206602 12970
rect 252384 12936 252418 12970
rect 264620 12936 264654 12970
rect 302616 12936 302650 12970
rect 304456 12936 304490 12970
rect 29008 12868 29042 12902
rect 36552 12868 36586 12902
rect 37380 12868 37414 12902
rect 38484 12868 38518 12902
rect 39772 12868 39806 12902
rect 58632 12868 58666 12902
rect 77860 12868 77894 12902
rect 78596 12868 78630 12902
rect 99480 12868 99514 12902
rect 104632 12868 104666 12902
rect 104724 12868 104758 12902
rect 112360 12868 112394 12902
rect 114016 12868 114050 12902
rect 115672 12868 115706 12902
rect 133612 12868 133646 12902
rect 145940 12868 145974 12902
rect 159280 12868 159314 12902
rect 164524 12868 164558 12902
rect 181636 12868 181670 12902
rect 189548 12868 189582 12902
rect 190928 12868 190962 12902
rect 193320 12868 193354 12902
rect 195896 12868 195930 12902
rect 231040 12868 231074 12902
rect 238768 12868 238802 12902
rect 240976 12868 241010 12902
rect 245300 12868 245334 12902
rect 251372 12868 251406 12902
rect 252476 12868 252510 12902
rect 261768 12868 261802 12902
rect 263240 12868 263274 12902
rect 263424 12868 263458 12902
rect 265540 12868 265574 12902
rect 271796 12868 271830 12902
rect 272900 12868 272934 12902
rect 305008 12868 305042 12902
rect 305468 12868 305502 12902
rect 26248 12800 26282 12834
rect 27812 12800 27846 12834
rect 34712 12800 34746 12834
rect 35724 12800 35758 12834
rect 38392 12800 38426 12834
rect 41704 12800 41738 12834
rect 42440 12800 42474 12834
rect 44740 12800 44774 12834
rect 52192 12800 52226 12834
rect 52928 12800 52962 12834
rect 54032 12800 54066 12834
rect 54768 12800 54802 12834
rect 57068 12800 57102 12834
rect 72340 12800 72374 12834
rect 75100 12800 75134 12834
rect 75560 12800 75594 12834
rect 77768 12800 77802 12834
rect 78504 12800 78538 12834
rect 79332 12800 79366 12834
rect 79792 12800 79826 12834
rect 86232 12800 86266 12834
rect 90464 12800 90498 12834
rect 91292 12800 91326 12834
rect 98560 12800 98594 12834
rect 106104 12800 106138 12834
rect 113096 12800 113130 12834
rect 113832 12800 113866 12834
rect 114660 12800 114694 12834
rect 118892 12800 118926 12834
rect 126896 12800 126930 12834
rect 127448 12800 127482 12834
rect 128276 12800 128310 12834
rect 129104 12800 129138 12834
rect 130208 12800 130242 12834
rect 130852 12800 130886 12834
rect 134532 12800 134566 12834
rect 135360 12800 135394 12834
rect 142996 12800 143030 12834
rect 145848 12800 145882 12834
rect 147044 12800 147078 12834
rect 149896 12800 149930 12834
rect 154864 12800 154898 12834
rect 159188 12800 159222 12834
rect 160016 12800 160050 12834
rect 161212 12800 161246 12834
rect 161856 12800 161890 12834
rect 165352 12800 165386 12834
rect 166548 12800 166582 12834
rect 167376 12800 167410 12834
rect 168020 12800 168054 12834
rect 175196 12800 175230 12834
rect 175840 12800 175874 12834
rect 176392 12800 176426 12834
rect 178600 12800 178634 12834
rect 180992 12800 181026 12834
rect 181544 12800 181578 12834
rect 182188 12800 182222 12834
rect 188076 12800 188110 12834
rect 188628 12800 188662 12834
rect 189364 12800 189398 12834
rect 191020 12800 191054 12834
rect 192216 12800 192250 12834
rect 195068 12800 195102 12834
rect 197368 12800 197402 12834
rect 197460 12800 197494 12834
rect 198380 12800 198414 12834
rect 200496 12800 200530 12834
rect 201324 12800 201358 12834
rect 204820 12800 204854 12834
rect 207488 12800 207522 12834
rect 226716 12800 226750 12834
rect 227360 12800 227394 12834
rect 227912 12800 227946 12834
rect 230304 12800 230338 12834
rect 230764 12800 230798 12834
rect 233064 12800 233098 12834
rect 237020 12800 237054 12834
rect 237664 12800 237698 12834
rect 238492 12800 238526 12834
rect 240700 12800 240734 12834
rect 243828 12800 243862 12834
rect 244564 12800 244598 12834
rect 244748 12800 244782 12834
rect 245208 12800 245242 12834
rect 250360 12800 250394 12834
rect 251556 12800 251590 12834
rect 256248 12800 256282 12834
rect 257076 12800 257110 12834
rect 262504 12800 262538 12834
rect 264160 12800 264194 12834
rect 264804 12800 264838 12834
rect 265264 12800 265298 12834
rect 267840 12800 267874 12834
rect 269128 12800 269162 12834
rect 271704 12800 271738 12834
rect 302800 12800 302834 12834
rect 304640 12800 304674 12834
rect 27904 12732 27938 12766
rect 28088 12732 28122 12766
rect 29100 12732 29134 12766
rect 29284 12732 29318 12766
rect 29836 12732 29870 12766
rect 30112 12732 30146 12766
rect 32136 12732 32170 12766
rect 32412 12732 32446 12766
rect 34896 12732 34930 12766
rect 37564 12732 37598 12766
rect 38576 12732 38610 12766
rect 39496 12732 39530 12766
rect 43544 12732 43578 12766
rect 43728 12732 43762 12766
rect 54124 12732 54158 12766
rect 55044 12732 55078 12766
rect 58724 12732 58758 12766
rect 75836 12732 75870 12766
rect 80068 12732 80102 12766
rect 84024 12732 84058 12766
rect 84300 12732 84334 12766
rect 86508 12732 86542 12766
rect 89636 12732 89670 12766
rect 89820 12732 89854 12766
rect 99204 12732 99238 12766
rect 101412 12732 101446 12766
rect 101688 12732 101722 12766
rect 104816 12732 104850 12766
rect 112544 12732 112578 12766
rect 113188 12732 113222 12766
rect 115764 12732 115798 12766
rect 115856 12732 115890 12766
rect 116500 12732 116534 12766
rect 116776 12732 116810 12766
rect 129380 12732 129414 12766
rect 131128 12732 131162 12766
rect 132600 12732 132634 12766
rect 133796 12732 133830 12766
rect 143272 12732 143306 12766
rect 146124 12732 146158 12766
rect 147504 12732 147538 12766
rect 147780 12732 147814 12766
rect 149252 12732 149286 12766
rect 151552 12732 151586 12766
rect 151736 12732 151770 12766
rect 155048 12732 155082 12766
rect 159464 12732 159498 12766
rect 162132 12732 162166 12766
rect 164616 12732 164650 12766
rect 176668 12732 176702 12766
rect 178876 12732 178910 12766
rect 191204 12732 191238 12766
rect 192400 12732 192434 12766
rect 193044 12732 193078 12766
rect 196172 12732 196206 12766
rect 197644 12732 197678 12766
rect 198104 12732 198138 12766
rect 200588 12732 200622 12766
rect 202612 12732 202646 12766
rect 202888 12732 202922 12766
rect 205096 12732 205130 12766
rect 228188 12732 228222 12766
rect 233156 12732 233190 12766
rect 252568 12732 252602 12766
rect 253672 12732 253706 12766
rect 253948 12732 253982 12766
rect 255420 12732 255454 12766
rect 256340 12732 256374 12766
rect 256432 12732 256466 12766
rect 267932 12732 267966 12766
rect 268024 12732 268058 12766
rect 269404 12732 269438 12766
rect 271980 12732 272014 12766
rect 272992 12732 273026 12766
rect 273084 12732 273118 12766
rect 74916 12664 74950 12698
rect 79148 12664 79182 12698
rect 81540 12664 81574 12698
rect 100952 12664 100986 12698
rect 105920 12664 105954 12698
rect 135544 12664 135578 12698
rect 152380 12664 152414 12698
rect 154496 12664 154530 12698
rect 158820 12664 158854 12698
rect 160200 12664 160234 12698
rect 167192 12664 167226 12698
rect 187892 12664 187926 12698
rect 207304 12664 207338 12698
rect 227176 12664 227210 12698
rect 237480 12664 237514 12698
rect 250176 12664 250210 12698
rect 255880 12664 255914 12698
rect 262688 12664 262722 12698
rect 28640 12596 28674 12630
rect 31584 12596 31618 12630
rect 34344 12596 34378 12630
rect 38024 12596 38058 12630
rect 41244 12596 41278 12630
rect 41796 12596 41830 12630
rect 43084 12596 43118 12630
rect 53020 12596 53054 12630
rect 56516 12596 56550 12630
rect 57160 12596 57194 12630
rect 58172 12596 58206 12630
rect 77308 12596 77342 12630
rect 85772 12596 85806 12630
rect 87980 12596 88014 12630
rect 89176 12596 89210 12630
rect 90556 12596 90590 12630
rect 98376 12596 98410 12630
rect 103160 12596 103194 12630
rect 104264 12596 104298 12630
rect 111900 12596 111934 12630
rect 114752 12596 114786 12630
rect 115304 12596 115338 12630
rect 127540 12596 127574 12630
rect 133152 12596 133186 12630
rect 146860 12596 146894 12630
rect 149988 12596 150022 12630
rect 151092 12596 151126 12630
rect 161304 12596 161338 12630
rect 164064 12596 164098 12630
rect 165444 12596 165478 12630
rect 166640 12596 166674 12630
rect 178140 12596 178174 12630
rect 180348 12596 180382 12630
rect 182280 12596 182314 12630
rect 188720 12596 188754 12630
rect 190560 12596 190594 12630
rect 191848 12596 191882 12630
rect 195528 12596 195562 12630
rect 197000 12596 197034 12630
rect 198196 12596 198230 12630
rect 201140 12596 201174 12630
rect 204360 12596 204394 12630
rect 226532 12596 226566 12630
rect 229660 12596 229694 12630
rect 230120 12596 230154 12630
rect 232512 12596 232546 12630
rect 236836 12596 236870 12630
rect 240240 12596 240274 12630
rect 242448 12596 242482 12630
rect 243920 12596 243954 12630
rect 252016 12596 252050 12630
rect 257168 12596 257202 12630
rect 261860 12596 261894 12630
rect 263976 12596 264010 12630
rect 267012 12596 267046 12630
rect 267472 12596 267506 12630
rect 270876 12596 270910 12630
rect 271336 12596 271370 12630
rect 272532 12596 272566 12630
rect 31308 12392 31342 12426
rect 33976 12392 34010 12426
rect 34804 12392 34838 12426
rect 37196 12392 37230 12426
rect 38484 12392 38518 12426
rect 39220 12392 39254 12426
rect 43176 12392 43210 12426
rect 43820 12392 43854 12426
rect 54124 12392 54158 12426
rect 54676 12392 54710 12426
rect 57344 12392 57378 12426
rect 57988 12392 58022 12426
rect 75192 12392 75226 12426
rect 79332 12392 79366 12426
rect 80252 12392 80286 12426
rect 85588 12392 85622 12426
rect 86416 12392 86450 12426
rect 88900 12392 88934 12426
rect 90188 12392 90222 12426
rect 99112 12392 99146 12426
rect 99848 12392 99882 12426
rect 103896 12392 103930 12426
rect 105184 12392 105218 12426
rect 113096 12392 113130 12426
rect 113740 12392 113774 12426
rect 118432 12392 118466 12426
rect 127724 12392 127758 12426
rect 130852 12392 130886 12426
rect 132692 12392 132726 12426
rect 147320 12392 147354 12426
rect 152564 12392 152598 12426
rect 154128 12392 154162 12426
rect 165352 12392 165386 12426
rect 175932 12392 175966 12426
rect 181360 12392 181394 12426
rect 188536 12392 188570 12426
rect 190192 12392 190226 12426
rect 201692 12392 201726 12426
rect 206476 12392 206510 12426
rect 227808 12392 227842 12426
rect 232236 12392 232270 12426
rect 239964 12392 239998 12426
rect 243552 12392 243586 12426
rect 244196 12392 244230 12426
rect 251096 12392 251130 12426
rect 256892 12392 256926 12426
rect 262504 12392 262538 12426
rect 264620 12392 264654 12426
rect 271060 12392 271094 12426
rect 305468 12392 305502 12426
rect 77492 12324 77526 12358
rect 89452 12324 89486 12358
rect 148424 12324 148458 12358
rect 153300 12324 153334 12358
rect 160016 12324 160050 12358
rect 166088 12324 166122 12358
rect 180900 12324 180934 12358
rect 192584 12324 192618 12358
rect 201140 12324 201174 12358
rect 229752 12324 229786 12358
rect 238768 12324 238802 12358
rect 242356 12324 242390 12358
rect 252108 12324 252142 12358
rect 254316 12324 254350 12358
rect 256340 12324 256374 12358
rect 264068 12324 264102 12358
rect 271704 12324 271738 12358
rect 27720 12256 27754 12290
rect 28732 12256 28766 12290
rect 28916 12256 28950 12290
rect 29560 12256 29594 12290
rect 31768 12256 31802 12290
rect 40876 12256 40910 12290
rect 52376 12256 52410 12290
rect 55688 12256 55722 12290
rect 56700 12256 56734 12290
rect 76756 12256 76790 12290
rect 76940 12256 76974 12290
rect 78136 12256 78170 12290
rect 84484 12256 84518 12290
rect 84668 12256 84702 12290
rect 87060 12256 87094 12290
rect 88164 12256 88198 12290
rect 100952 12256 100986 12290
rect 103160 12256 103194 12290
rect 104540 12256 104574 12290
rect 114384 12256 114418 12290
rect 117788 12256 117822 12290
rect 131864 12256 131898 12290
rect 152104 12256 152138 12290
rect 152196 12256 152230 12290
rect 153944 12256 153978 12290
rect 161304 12256 161338 12290
rect 161488 12256 161522 12290
rect 162500 12256 162534 12290
rect 162684 12256 162718 12290
rect 163604 12256 163638 12290
rect 177036 12256 177070 12290
rect 177128 12256 177162 12290
rect 190836 12256 190870 12290
rect 193688 12256 193722 12290
rect 197552 12256 197586 12290
rect 203532 12256 203566 12290
rect 204728 12256 204762 12290
rect 231592 12256 231626 12290
rect 239320 12256 239354 12290
rect 241436 12256 241470 12290
rect 242816 12256 242850 12290
rect 242908 12256 242942 12290
rect 252568 12256 252602 12290
rect 255328 12256 255362 12290
rect 265724 12256 265758 12290
rect 265908 12256 265942 12290
rect 268760 12256 268794 12290
rect 272256 12256 272290 12290
rect 27444 12188 27478 12222
rect 28640 12188 28674 12222
rect 34160 12188 34194 12222
rect 34712 12188 34746 12222
rect 35356 12188 35390 12222
rect 36368 12188 36402 12222
rect 37104 12188 37138 12222
rect 38668 12188 38702 12222
rect 39128 12188 39162 12222
rect 40600 12188 40634 12222
rect 41428 12188 41462 12222
rect 43728 12188 43762 12222
rect 54584 12188 54618 12222
rect 56608 12188 56642 12222
rect 57528 12188 57562 12222
rect 58172 12188 58206 12222
rect 75376 12188 75410 12222
rect 76664 12188 76698 12222
rect 77952 12188 77986 12222
rect 79240 12188 79274 12222
rect 80160 12188 80194 12222
rect 84392 12188 84426 12222
rect 85496 12188 85530 12222
rect 86876 12188 86910 12222
rect 87980 12188 88014 12222
rect 88808 12188 88842 12222
rect 89636 12188 89670 12222
rect 90096 12188 90130 12222
rect 99296 12188 99330 12222
rect 99756 12188 99790 12222
rect 102976 12188 103010 12222
rect 103804 12188 103838 12222
rect 104448 12188 104482 12222
rect 105092 12188 105126 12222
rect 113280 12188 113314 12222
rect 113924 12188 113958 12222
rect 117604 12188 117638 12222
rect 118340 12188 118374 12222
rect 127908 12188 127942 12222
rect 128644 12188 128678 12222
rect 129104 12188 129138 12222
rect 131680 12188 131714 12222
rect 132600 12188 132634 12222
rect 137752 12188 137786 12222
rect 147504 12188 147538 12222
rect 148332 12188 148366 12222
rect 149436 12188 149470 12222
rect 152472 12188 152506 12222
rect 154312 12188 154346 12222
rect 160200 12188 160234 12222
rect 161212 12188 161246 12222
rect 176116 12188 176150 12222
rect 176944 12188 176978 12222
rect 179152 12188 179186 12222
rect 181544 12188 181578 12222
rect 188720 12188 188754 12222
rect 189548 12188 189582 12222
rect 190376 12188 190410 12222
rect 194424 12188 194458 12222
rect 196448 12188 196482 12222
rect 196724 12188 196758 12222
rect 197460 12188 197494 12222
rect 201048 12188 201082 12222
rect 201876 12188 201910 12222
rect 203256 12188 203290 12222
rect 227544 12188 227578 12222
rect 229936 12188 229970 12222
rect 232144 12188 232178 12222
rect 238032 12188 238066 12222
rect 239136 12188 239170 12222
rect 239228 12188 239262 12222
rect 240148 12188 240182 12222
rect 241252 12188 241286 12222
rect 243736 12188 243770 12222
rect 244380 12188 244414 12222
rect 251280 12188 251314 12222
rect 251924 12188 251958 12222
rect 255144 12188 255178 12222
rect 256248 12188 256282 12222
rect 257076 12188 257110 12222
rect 262688 12188 262722 12222
rect 263976 12188 264010 12222
rect 264804 12188 264838 12222
rect 266552 12188 266586 12222
rect 270968 12188 271002 12222
rect 272072 12188 272106 12222
rect 29836 12120 29870 12154
rect 32044 12120 32078 12154
rect 35448 12120 35482 12154
rect 41704 12120 41738 12154
rect 52652 12120 52686 12154
rect 55504 12120 55538 12154
rect 100768 12120 100802 12154
rect 100860 12120 100894 12154
rect 101964 12120 101998 12154
rect 102148 12120 102182 12154
rect 114660 12120 114694 12154
rect 117512 12120 117546 12154
rect 129380 12120 129414 12154
rect 138028 12120 138062 12154
rect 145848 12120 145882 12154
rect 146216 12120 146250 12154
rect 153668 12120 153702 12154
rect 163880 12120 163914 12154
rect 165904 12120 165938 12154
rect 177956 12120 177990 12154
rect 179428 12120 179462 12154
rect 191112 12120 191146 12154
rect 193412 12120 193446 12154
rect 194700 12120 194734 12154
rect 205004 12120 205038 12154
rect 249072 12120 249106 12154
rect 249256 12120 249290 12154
rect 252844 12120 252878 12154
rect 265632 12120 265666 12154
rect 266828 12120 266862 12154
rect 269036 12120 269070 12154
rect 27076 12052 27110 12086
rect 27536 12052 27570 12086
rect 28272 12052 28306 12086
rect 33516 12052 33550 12086
rect 36460 12052 36494 12086
rect 40232 12052 40266 12086
rect 40692 12052 40726 12086
rect 56056 12052 56090 12086
rect 56148 12052 56182 12086
rect 56516 12052 56550 12086
rect 76296 12052 76330 12086
rect 77860 12052 77894 12086
rect 84024 12052 84058 12086
rect 86784 12052 86818 12086
rect 87612 12052 87646 12086
rect 88072 12052 88106 12086
rect 100400 12052 100434 12086
rect 102608 12052 102642 12086
rect 103068 12052 103102 12086
rect 116132 12052 116166 12086
rect 117144 12052 117178 12086
rect 128460 12052 128494 12086
rect 131312 12052 131346 12086
rect 131772 12052 131806 12086
rect 150724 12052 150758 12086
rect 151644 12052 151678 12086
rect 152012 12052 152046 12086
rect 153760 12052 153794 12086
rect 160844 12052 160878 12086
rect 162040 12052 162074 12086
rect 162408 12052 162442 12086
rect 176576 12052 176610 12086
rect 178048 12052 178082 12086
rect 189640 12052 189674 12086
rect 193044 12052 193078 12086
rect 193504 12052 193538 12086
rect 196816 12052 196850 12086
rect 197000 12052 197034 12086
rect 197368 12052 197402 12086
rect 202888 12052 202922 12086
rect 203348 12052 203382 12086
rect 229292 12052 229326 12086
rect 230948 12052 230982 12086
rect 231316 12052 231350 12086
rect 231408 12052 231442 12086
rect 238216 12052 238250 12086
rect 240884 12052 240918 12086
rect 241344 12052 241378 12086
rect 242724 12052 242758 12086
rect 254776 12052 254810 12086
rect 255236 12052 255270 12086
rect 265264 12052 265298 12086
rect 268300 12052 268334 12086
rect 270508 12052 270542 12086
rect 272164 12052 272198 12086
rect 27812 11848 27846 11882
rect 32596 11848 32630 11882
rect 33792 11848 33826 11882
rect 34436 11848 34470 11882
rect 34988 11848 35022 11882
rect 38392 11848 38426 11882
rect 39036 11848 39070 11882
rect 39680 11848 39714 11882
rect 40140 11848 40174 11882
rect 41152 11848 41186 11882
rect 41704 11848 41738 11882
rect 52836 11848 52870 11882
rect 53664 11848 53698 11882
rect 54400 11848 54434 11882
rect 55320 11848 55354 11882
rect 56516 11848 56550 11882
rect 57160 11848 57194 11882
rect 75560 11848 75594 11882
rect 76020 11848 76054 11882
rect 76940 11848 76974 11882
rect 77860 11848 77894 11882
rect 78504 11848 78538 11882
rect 84392 11848 84426 11882
rect 86048 11848 86082 11882
rect 87152 11848 87186 11882
rect 87888 11848 87922 11882
rect 88900 11848 88934 11882
rect 100216 11848 100250 11882
rect 100952 11848 100986 11882
rect 101872 11848 101906 11882
rect 113832 11848 113866 11882
rect 115028 11848 115062 11882
rect 116224 11848 116258 11882
rect 116960 11848 116994 11882
rect 117604 11848 117638 11882
rect 129380 11848 129414 11882
rect 130484 11848 130518 11882
rect 130944 11848 130978 11882
rect 132416 11848 132450 11882
rect 151092 11848 151126 11882
rect 152012 11848 152046 11882
rect 152748 11848 152782 11882
rect 162316 11848 162350 11882
rect 162960 11848 162994 11882
rect 163512 11848 163546 11882
rect 164248 11848 164282 11882
rect 164892 11848 164926 11882
rect 176484 11848 176518 11882
rect 177588 11848 177622 11882
rect 178048 11848 178082 11882
rect 179152 11848 179186 11882
rect 180072 11848 180106 11882
rect 190836 11848 190870 11882
rect 196264 11848 196298 11882
rect 202888 11848 202922 11882
rect 204084 11848 204118 11882
rect 205188 11848 205222 11882
rect 228280 11848 228314 11882
rect 229476 11848 229510 11882
rect 230396 11848 230430 11882
rect 231592 11848 231626 11882
rect 238768 11848 238802 11882
rect 240332 11848 240366 11882
rect 241068 11848 241102 11882
rect 241804 11848 241838 11882
rect 251832 11848 251866 11882
rect 254132 11848 254166 11882
rect 254960 11848 254994 11882
rect 255604 11848 255638 11882
rect 264988 11848 265022 11882
rect 267380 11848 267414 11882
rect 268208 11848 268242 11882
rect 271428 11848 271462 11882
rect 28824 11780 28858 11814
rect 40048 11780 40082 11814
rect 202336 11780 202370 11814
rect 203992 11780 204026 11814
rect 205280 11780 205314 11814
rect 228372 11780 228406 11814
rect 229568 11780 229602 11814
rect 238676 11780 238710 11814
rect 254040 11780 254074 11814
rect 264436 11780 264470 11814
rect 27996 11712 28030 11746
rect 29652 11712 29686 11746
rect 32504 11712 32538 11746
rect 33700 11712 33734 11746
rect 34344 11712 34378 11746
rect 35172 11712 35206 11746
rect 38576 11712 38610 11746
rect 39220 11712 39254 11746
rect 41060 11712 41094 11746
rect 41888 11712 41922 11746
rect 42900 11712 42934 11746
rect 53020 11712 53054 11746
rect 53848 11712 53882 11746
rect 54308 11712 54342 11746
rect 56424 11712 56458 11746
rect 57068 11712 57102 11746
rect 75928 11712 75962 11746
rect 77124 11712 77158 11746
rect 77768 11712 77802 11746
rect 78688 11712 78722 11746
rect 84576 11712 84610 11746
rect 85220 11712 85254 11746
rect 86140 11712 86174 11746
rect 86968 11712 87002 11746
rect 87796 11712 87830 11746
rect 88808 11712 88842 11746
rect 100400 11712 100434 11746
rect 100860 11712 100894 11746
rect 103160 11712 103194 11746
rect 114016 11712 114050 11746
rect 115120 11712 115154 11746
rect 116408 11712 116442 11746
rect 116868 11712 116902 11746
rect 117512 11712 117546 11746
rect 129288 11712 129322 11746
rect 130852 11712 130886 11746
rect 131680 11712 131714 11746
rect 132600 11712 132634 11746
rect 147780 11712 147814 11746
rect 151276 11712 151310 11746
rect 152196 11712 152230 11746
rect 152656 11712 152690 11746
rect 161120 11712 161154 11746
rect 161764 11712 161798 11746
rect 162224 11712 162258 11746
rect 162868 11712 162902 11746
rect 163696 11712 163730 11746
rect 164156 11712 164190 11746
rect 164800 11712 164834 11746
rect 176668 11712 176702 11746
rect 177956 11712 177990 11746
rect 179244 11712 179278 11746
rect 179980 11712 180014 11746
rect 189640 11712 189674 11746
rect 190100 11712 190134 11746
rect 190744 11712 190778 11746
rect 191848 11712 191882 11746
rect 194056 11712 194090 11746
rect 196448 11712 196482 11746
rect 202244 11712 202278 11746
rect 203072 11712 203106 11746
rect 230304 11712 230338 11746
rect 230948 11712 230982 11746
rect 231040 11712 231074 11746
rect 231776 11712 231810 11746
rect 240240 11712 240274 11746
rect 241252 11712 241286 11746
rect 241712 11712 241746 11746
rect 242540 11712 242574 11746
rect 252016 11712 252050 11746
rect 252384 11712 252418 11746
rect 252752 11712 252786 11746
rect 254868 11712 254902 11746
rect 255512 11712 255546 11746
rect 264344 11712 264378 11746
rect 265172 11712 265206 11746
rect 265632 11712 265666 11746
rect 269128 11712 269162 11746
rect 271336 11712 271370 11746
rect 28916 11644 28950 11678
rect 29100 11644 29134 11678
rect 29928 11644 29962 11678
rect 32688 11644 32722 11678
rect 40232 11644 40266 11678
rect 43084 11644 43118 11678
rect 55412 11644 55446 11678
rect 55596 11644 55630 11678
rect 76204 11644 76238 11678
rect 86324 11644 86358 11678
rect 101964 11644 101998 11678
rect 102056 11644 102090 11678
rect 115304 11644 115338 11678
rect 131036 11644 131070 11678
rect 148332 11644 148366 11678
rect 148608 11644 148642 11678
rect 178140 11644 178174 11678
rect 179336 11644 179370 11678
rect 192124 11644 192158 11678
rect 194332 11644 194366 11678
rect 195804 11644 195838 11678
rect 204268 11644 204302 11678
rect 205464 11644 205498 11678
rect 228464 11644 228498 11678
rect 229752 11644 229786 11678
rect 240424 11644 240458 11678
rect 254224 11644 254258 11678
rect 265908 11644 265942 11678
rect 268300 11644 268334 11678
rect 268392 11644 268426 11678
rect 269404 11644 269438 11678
rect 270876 11644 270910 11678
rect 43452 11576 43486 11610
rect 147596 11576 147630 11610
rect 160936 11576 160970 11610
rect 161580 11576 161614 11610
rect 178784 11576 178818 11610
rect 190192 11576 190226 11610
rect 227912 11576 227946 11610
rect 239872 11576 239906 11610
rect 252936 11576 252970 11610
rect 28456 11508 28490 11542
rect 31400 11508 31434 11542
rect 32136 11508 32170 11542
rect 54952 11508 54986 11542
rect 85036 11508 85070 11542
rect 85680 11508 85714 11542
rect 101504 11508 101538 11542
rect 102976 11508 103010 11542
rect 114660 11508 114694 11542
rect 131864 11508 131898 11542
rect 150080 11508 150114 11542
rect 189456 11508 189490 11542
rect 193596 11508 193630 11542
rect 203624 11508 203658 11542
rect 204820 11508 204854 11542
rect 229108 11508 229142 11542
rect 242356 11508 242390 11542
rect 253672 11508 253706 11542
rect 267840 11508 267874 11542
rect 28824 11304 28858 11338
rect 33608 11304 33642 11338
rect 40324 11304 40358 11338
rect 41060 11304 41094 11338
rect 41612 11304 41646 11338
rect 55320 11304 55354 11338
rect 56240 11304 56274 11338
rect 76480 11304 76514 11338
rect 78228 11304 78262 11338
rect 86232 11304 86266 11338
rect 86968 11304 87002 11338
rect 88256 11304 88290 11338
rect 102884 11304 102918 11338
rect 116040 11304 116074 11338
rect 117144 11304 117178 11338
rect 130484 11304 130518 11338
rect 131220 11304 131254 11338
rect 131772 11304 131806 11338
rect 148056 11304 148090 11338
rect 150816 11304 150850 11338
rect 157348 11304 157382 11338
rect 162040 11304 162074 11338
rect 162684 11304 162718 11338
rect 163604 11304 163638 11338
rect 239964 11304 239998 11338
rect 240884 11304 240918 11338
rect 241436 11304 241470 11338
rect 242172 11304 242206 11338
rect 252568 11304 252602 11338
rect 253120 11304 253154 11338
rect 253764 11304 253798 11338
rect 265540 11304 265574 11338
rect 268024 11304 268058 11338
rect 42256 11236 42290 11270
rect 87612 11236 87646 11270
rect 103528 11236 103562 11270
rect 115396 11236 115430 11270
rect 149896 11236 149930 11270
rect 254408 11236 254442 11270
rect 266828 11236 266862 11270
rect 29652 11168 29686 11202
rect 32320 11168 32354 11202
rect 32504 11168 32538 11202
rect 102332 11168 102366 11202
rect 148516 11168 148550 11202
rect 148700 11168 148734 11202
rect 177588 11168 177622 11202
rect 178232 11168 178266 11202
rect 190284 11168 190318 11202
rect 192032 11168 192066 11202
rect 193780 11168 193814 11202
rect 194976 11168 195010 11202
rect 202888 11168 202922 11202
rect 264988 11168 265022 11202
rect 267472 11168 267506 11202
rect 268576 11168 268610 11202
rect 269404 11168 269438 11202
rect 270600 11168 270634 11202
rect 29008 11100 29042 11134
rect 32228 11100 32262 11134
rect 33516 11100 33550 11134
rect 40508 11100 40542 11134
rect 40968 11100 41002 11134
rect 41796 11100 41830 11134
rect 42440 11100 42474 11134
rect 55504 11100 55538 11134
rect 56424 11100 56458 11134
rect 76664 11100 76698 11134
rect 78412 11100 78446 11134
rect 86416 11100 86450 11134
rect 86876 11100 86910 11134
rect 87796 11100 87830 11134
rect 88440 11100 88474 11134
rect 102148 11100 102182 11134
rect 103068 11100 103102 11134
rect 103712 11100 103746 11134
rect 115304 11100 115338 11134
rect 116224 11100 116258 11134
rect 117328 11100 117362 11134
rect 130668 11100 130702 11134
rect 131128 11100 131162 11134
rect 131956 11100 131990 11134
rect 142076 11100 142110 11134
rect 151000 11100 151034 11134
rect 162224 11100 162258 11134
rect 162868 11100 162902 11134
rect 163512 11100 163546 11134
rect 177496 11100 177530 11134
rect 178140 11100 178174 11134
rect 179152 11100 179186 11134
rect 190192 11100 190226 11134
rect 190836 11100 190870 11134
rect 190928 11100 190962 11134
rect 194792 11100 194826 11134
rect 195804 11100 195838 11134
rect 202336 11100 202370 11134
rect 202796 11100 202830 11134
rect 203440 11100 203474 11134
rect 204912 11100 204946 11134
rect 229384 11100 229418 11134
rect 239872 11100 239906 11134
rect 240792 11100 240826 11134
rect 241620 11100 241654 11134
rect 242080 11100 242114 11134
rect 252476 11100 252510 11134
rect 253304 11100 253338 11134
rect 253948 11100 253982 11134
rect 254592 11100 254626 11134
rect 264896 11100 264930 11134
rect 265724 11100 265758 11134
rect 267196 11100 267230 11134
rect 268208 11100 268242 11134
rect 270416 11100 270450 11134
rect 270508 11100 270542 11134
rect 29928 11032 29962 11066
rect 140420 11032 140454 11066
rect 149620 11032 149654 11066
rect 156060 11032 156094 11066
rect 192308 11032 192342 11066
rect 267288 11032 267322 11066
rect 269220 11032 269254 11066
rect 269312 11032 269346 11066
rect 31400 10964 31434 10998
rect 31860 10964 31894 10998
rect 148424 10964 148458 10998
rect 178968 10964 179002 10998
rect 194424 10964 194458 10998
rect 194884 10964 194918 10998
rect 195620 10964 195654 10998
rect 202152 10964 202186 10998
rect 203532 10964 203566 10998
rect 204728 10964 204762 10998
rect 229200 10964 229234 10998
rect 268852 10964 268886 10998
rect 270048 10964 270082 10998
rect 29652 10760 29686 10794
rect 30664 10760 30698 10794
rect 30756 10760 30790 10794
rect 32136 10760 32170 10794
rect 32780 10760 32814 10794
rect 33424 10760 33458 10794
rect 101688 10760 101722 10794
rect 130484 10760 130518 10794
rect 141984 10760 142018 10794
rect 148884 10760 148918 10794
rect 150724 10760 150758 10794
rect 191848 10760 191882 10794
rect 194240 10760 194274 10794
rect 202888 10760 202922 10794
rect 253672 10760 253706 10794
rect 266552 10760 266586 10794
rect 267748 10760 267782 10794
rect 268392 10760 268426 10794
rect 140696 10692 140730 10726
rect 156152 10692 156186 10726
rect 193504 10692 193538 10726
rect 29836 10624 29870 10658
rect 32320 10624 32354 10658
rect 32964 10624 32998 10658
rect 33608 10624 33642 10658
rect 101872 10624 101906 10658
rect 130392 10624 130426 10658
rect 149068 10624 149102 10658
rect 150632 10624 150666 10658
rect 187248 10624 187282 10658
rect 191296 10624 191330 10658
rect 192032 10624 192066 10658
rect 192676 10624 192710 10658
rect 194148 10624 194182 10658
rect 203072 10624 203106 10658
rect 253856 10624 253890 10658
rect 266000 10624 266034 10658
rect 266460 10624 266494 10658
rect 267104 10624 267138 10658
rect 267932 10624 267966 10658
rect 268576 10624 268610 10658
rect 269128 10624 269162 10658
rect 269220 10624 269254 10658
rect 30848 10556 30882 10590
rect 187524 10556 187558 10590
rect 30296 10488 30330 10522
rect 191112 10488 191146 10522
rect 192860 10488 192894 10522
rect 193688 10488 193722 10522
rect 267196 10488 267230 10522
rect 157624 10420 157658 10454
rect 265816 10420 265850 10454
rect 30940 10216 30974 10250
rect 31676 10216 31710 10250
rect 32872 10216 32906 10250
rect 33608 10216 33642 10250
rect 191848 10216 191882 10250
rect 193136 10216 193170 10250
rect 267748 10216 267782 10250
rect 269036 10216 269070 10250
rect 30296 10148 30330 10182
rect 32320 10148 32354 10182
rect 267104 10148 267138 10182
rect 268484 10148 268518 10182
rect 157808 10080 157842 10114
rect 30480 10012 30514 10046
rect 31124 10012 31158 10046
rect 31584 10012 31618 10046
rect 32228 10012 32262 10046
rect 33056 10012 33090 10046
rect 33516 10012 33550 10046
rect 140420 10012 140454 10046
rect 156060 10012 156094 10046
rect 192032 10012 192066 10046
rect 192676 10012 192710 10046
rect 193320 10012 193354 10046
rect 267288 10012 267322 10046
rect 267932 10012 267966 10046
rect 268392 10012 268426 10046
rect 269220 10012 269254 10046
rect 304456 10012 304490 10046
rect 304824 9944 304858 9978
rect 141708 9876 141742 9910
rect 192492 9876 192526 9910
rect 32872 9604 32906 9638
rect 140696 9604 140730 9638
rect 156152 9604 156186 9638
rect 157900 9604 157934 9638
rect 193044 9604 193078 9638
rect 267932 9604 267966 9638
rect 31308 9536 31342 9570
rect 32136 9536 32170 9570
rect 32780 9536 32814 9570
rect 192492 9536 192526 9570
rect 192952 9536 192986 9570
rect 267840 9536 267874 9570
rect 32228 9468 32262 9502
rect 31124 9400 31158 9434
rect 192308 9400 192342 9434
rect 141984 9332 142018 9366
rect 1592 8448 1626 8482
rect 1408 8312 1442 8346
rect 1960 8312 1994 8346
rect 2328 8312 2362 8346
rect 2696 8312 2730 8346
rect 3064 8312 3098 8346
rect 303996 6272 304030 6306
rect 304272 6204 304306 6238
<< metal1 >>
rect 189902 13852 189908 13864
rect 72344 13824 75500 13852
rect 28994 13744 29000 13796
rect 29052 13784 29058 13796
rect 32950 13784 32956 13796
rect 29052 13756 32956 13784
rect 29052 13744 29058 13756
rect 32950 13744 32956 13756
rect 33008 13744 33014 13796
rect 46198 13744 46204 13796
rect 46256 13784 46262 13796
rect 63402 13784 63408 13796
rect 46256 13756 63408 13784
rect 46256 13744 46262 13756
rect 63402 13744 63408 13756
rect 63460 13744 63466 13796
rect 69290 13744 69296 13796
rect 69348 13784 69354 13796
rect 72344 13784 72372 13824
rect 75362 13784 75368 13796
rect 69348 13756 72372 13784
rect 72436 13756 75368 13784
rect 69348 13744 69354 13756
rect 72436 13728 72464 13756
rect 75362 13744 75368 13756
rect 75420 13744 75426 13796
rect 75472 13784 75500 13824
rect 189276 13824 189908 13852
rect 76006 13784 76012 13796
rect 75472 13756 76012 13784
rect 76006 13744 76012 13756
rect 76064 13744 76070 13796
rect 90634 13744 90640 13796
rect 90692 13784 90698 13796
rect 102410 13784 102416 13796
rect 90692 13756 102416 13784
rect 90692 13744 90698 13756
rect 102410 13744 102416 13756
rect 102468 13744 102474 13796
rect 113818 13744 113824 13796
rect 113876 13784 113882 13796
rect 125502 13784 125508 13796
rect 113876 13756 125508 13784
rect 113876 13744 113882 13756
rect 125502 13744 125508 13756
rect 125560 13784 125566 13796
rect 131850 13784 131856 13796
rect 125560 13756 131856 13784
rect 125560 13744 125566 13756
rect 131850 13744 131856 13756
rect 131908 13744 131914 13796
rect 161658 13744 161664 13796
rect 161716 13784 161722 13796
rect 166074 13784 166080 13796
rect 161716 13756 166080 13784
rect 161716 13744 161722 13756
rect 166074 13744 166080 13756
rect 166132 13784 166138 13796
rect 167362 13784 167368 13796
rect 166132 13756 167368 13784
rect 166132 13744 166138 13756
rect 167362 13744 167368 13756
rect 167420 13744 167426 13796
rect 174170 13744 174176 13796
rect 174228 13784 174234 13796
rect 177758 13784 177764 13796
rect 174228 13756 177764 13784
rect 174228 13744 174234 13756
rect 177758 13744 177764 13756
rect 177816 13744 177822 13796
rect 181898 13744 181904 13796
rect 181956 13784 181962 13796
rect 189276 13784 189304 13824
rect 189902 13812 189908 13824
rect 189960 13812 189966 13864
rect 181956 13756 189304 13784
rect 181956 13744 181962 13756
rect 189350 13744 189356 13796
rect 189408 13784 189414 13796
rect 193214 13784 193220 13796
rect 189408 13756 193220 13784
rect 189408 13744 189414 13756
rect 193214 13744 193220 13756
rect 193272 13744 193278 13796
rect 195974 13744 195980 13796
rect 196032 13784 196038 13796
rect 302786 13784 302792 13796
rect 196032 13756 302792 13784
rect 196032 13744 196038 13756
rect 302786 13744 302792 13756
rect 302844 13744 302850 13796
rect 27154 13676 27160 13728
rect 27212 13716 27218 13728
rect 36538 13716 36544 13728
rect 27212 13688 36544 13716
rect 27212 13676 27218 13688
rect 36538 13676 36544 13688
rect 36596 13676 36602 13728
rect 42518 13676 42524 13728
rect 42576 13716 42582 13728
rect 47854 13716 47860 13728
rect 42576 13688 47860 13716
rect 42576 13676 42582 13688
rect 47854 13676 47860 13688
rect 47912 13676 47918 13728
rect 51626 13676 51632 13728
rect 51684 13716 51690 13728
rect 54110 13716 54116 13728
rect 51684 13688 54116 13716
rect 51684 13676 51690 13688
rect 54110 13676 54116 13688
rect 54168 13676 54174 13728
rect 66162 13676 66168 13728
rect 66220 13716 66226 13728
rect 72418 13716 72424 13728
rect 66220 13688 72424 13716
rect 66220 13676 66226 13688
rect 72418 13676 72424 13688
rect 72476 13676 72482 13728
rect 73890 13676 73896 13728
rect 73948 13716 73954 13728
rect 76374 13716 76380 13728
rect 73948 13688 76380 13716
rect 73948 13676 73954 13688
rect 76374 13676 76380 13688
rect 76432 13676 76438 13728
rect 83090 13676 83096 13728
rect 83148 13716 83154 13728
rect 86402 13716 86408 13728
rect 83148 13688 86408 13716
rect 83148 13676 83154 13688
rect 86402 13676 86408 13688
rect 86460 13676 86466 13728
rect 91830 13676 91836 13728
rect 91888 13716 91894 13728
rect 101950 13716 101956 13728
rect 91888 13688 101956 13716
rect 91888 13676 91894 13688
rect 101950 13676 101956 13688
rect 102008 13676 102014 13728
rect 114646 13676 114652 13728
rect 114704 13716 114710 13728
rect 127434 13716 127440 13728
rect 114704 13688 127440 13716
rect 114704 13676 114710 13688
rect 127434 13676 127440 13688
rect 127492 13676 127498 13728
rect 127526 13676 127532 13728
rect 127584 13716 127590 13728
rect 129734 13716 129740 13728
rect 127584 13688 129740 13716
rect 127584 13676 127590 13688
rect 129734 13676 129740 13688
rect 129792 13676 129798 13728
rect 133598 13676 133604 13728
rect 133656 13716 133662 13728
rect 136818 13716 136824 13728
rect 133656 13688 136824 13716
rect 133656 13676 133662 13688
rect 136818 13676 136824 13688
rect 136876 13676 136882 13728
rect 148134 13676 148140 13728
rect 148192 13716 148198 13728
rect 150434 13716 150440 13728
rect 148192 13688 150440 13716
rect 148192 13676 148198 13688
rect 150434 13676 150440 13688
rect 150492 13676 150498 13728
rect 157150 13676 157156 13728
rect 157208 13716 157214 13728
rect 301406 13716 301412 13728
rect 157208 13688 301412 13716
rect 157208 13676 157214 13688
rect 301406 13676 301412 13688
rect 301464 13676 301470 13728
rect 1104 13626 305808 13648
rect 1104 13574 39048 13626
rect 39100 13574 39112 13626
rect 39164 13574 39176 13626
rect 39228 13574 39240 13626
rect 39292 13574 39304 13626
rect 39356 13574 115246 13626
rect 115298 13574 115310 13626
rect 115362 13574 115374 13626
rect 115426 13574 115438 13626
rect 115490 13574 115502 13626
rect 115554 13574 191444 13626
rect 191496 13574 191508 13626
rect 191560 13574 191572 13626
rect 191624 13574 191636 13626
rect 191688 13574 191700 13626
rect 191752 13574 267642 13626
rect 267694 13574 267706 13626
rect 267758 13574 267770 13626
rect 267822 13574 267834 13626
rect 267886 13574 267898 13626
rect 267950 13574 305808 13626
rect 1104 13552 305808 13574
rect 1578 13512 1584 13524
rect 1538 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 4614 13512 4620 13524
rect 4574 13484 4620 13512
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 7650 13512 7656 13524
rect 7610 13484 7656 13512
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 10778 13512 10784 13524
rect 10738 13484 10784 13512
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14092 13514 14150 13520
rect 14092 13512 14104 13514
rect 13872 13484 14104 13512
rect 13872 13472 13878 13484
rect 14092 13480 14104 13484
rect 14138 13480 14150 13514
rect 16850 13512 16856 13524
rect 16810 13484 16856 13512
rect 14092 13474 14150 13480
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 19978 13512 19984 13524
rect 19938 13484 19984 13512
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 23014 13512 23020 13524
rect 22974 13484 23020 13512
rect 23014 13472 23020 13484
rect 23072 13472 23078 13524
rect 25684 13514 25742 13520
rect 25684 13480 25696 13514
rect 25730 13512 25742 13514
rect 27614 13512 27620 13524
rect 25730 13484 27620 13512
rect 25730 13480 25742 13484
rect 25684 13474 25742 13480
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 27706 13472 27712 13524
rect 27764 13512 27770 13524
rect 28996 13514 29054 13520
rect 28996 13512 29008 13514
rect 27764 13484 29008 13512
rect 27764 13472 27770 13484
rect 28996 13480 29008 13484
rect 29042 13480 29054 13514
rect 28996 13474 29054 13480
rect 30466 13472 30472 13524
rect 30524 13512 30530 13524
rect 31572 13514 31630 13520
rect 31572 13512 31584 13514
rect 30524 13484 31584 13512
rect 30524 13472 30530 13484
rect 31572 13480 31584 13484
rect 31618 13480 31630 13514
rect 31572 13474 31630 13480
rect 36538 13472 36544 13524
rect 36596 13512 36602 13524
rect 46198 13512 46204 13524
rect 36596 13484 46204 13512
rect 36596 13472 36602 13484
rect 46198 13472 46204 13484
rect 46256 13472 46262 13524
rect 47578 13512 47584 13524
rect 47538 13484 47584 13512
rect 47578 13472 47584 13484
rect 47636 13472 47642 13524
rect 50340 13514 50398 13520
rect 50340 13480 50352 13514
rect 50386 13512 50398 13514
rect 50522 13512 50528 13524
rect 50386 13484 50528 13512
rect 50386 13480 50398 13484
rect 50340 13474 50398 13480
rect 50522 13472 50528 13484
rect 50580 13472 50586 13524
rect 50984 13514 51042 13520
rect 50984 13480 50996 13514
rect 51030 13512 51042 13514
rect 53006 13512 53012 13524
rect 51030 13484 53012 13512
rect 51030 13480 51042 13484
rect 50984 13474 51042 13480
rect 53006 13472 53012 13484
rect 53064 13472 53070 13524
rect 55582 13472 55588 13524
rect 55640 13512 55646 13524
rect 57882 13512 57888 13524
rect 55640 13484 57888 13512
rect 55640 13472 55646 13484
rect 57882 13472 57888 13484
rect 57940 13512 57946 13524
rect 61746 13512 61752 13524
rect 57940 13484 61752 13512
rect 57940 13472 57946 13484
rect 61746 13472 61752 13484
rect 61804 13472 61810 13524
rect 63402 13472 63408 13524
rect 63460 13512 63466 13524
rect 142890 13512 142896 13524
rect 63460 13484 142154 13512
rect 142850 13484 142896 13512
rect 63460 13472 63466 13484
rect 27154 13444 27160 13456
rect 6886 13416 27160 13444
rect 6886 13376 6914 13416
rect 27154 13404 27160 13416
rect 27212 13404 27218 13456
rect 44174 13404 44180 13456
rect 44232 13404 44238 13456
rect 44268 13446 44326 13452
rect 44268 13412 44280 13446
rect 44314 13412 44326 13446
rect 44268 13406 44326 13412
rect 26328 13378 26386 13384
rect 1780 13348 6914 13376
rect 10980 13348 26096 13376
rect 1780 13316 1808 13348
rect 1764 13310 1822 13316
rect 1764 13276 1776 13310
rect 1810 13276 1822 13310
rect 4798 13308 4804 13320
rect 4758 13280 4804 13308
rect 1764 13270 1822 13276
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 10980 13316 11008 13348
rect 7836 13310 7894 13316
rect 7836 13276 7848 13310
rect 7882 13276 7894 13310
rect 7836 13270 7894 13276
rect 10964 13310 11022 13316
rect 10964 13276 10976 13310
rect 11010 13276 11022 13310
rect 14274 13308 14280 13320
rect 14234 13280 14280 13308
rect 10964 13270 11022 13276
rect 7852 13240 7880 13270
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 17034 13308 17040 13320
rect 16994 13280 17040 13308
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 20162 13308 20168 13320
rect 20122 13280 20168 13308
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 23198 13308 23204 13320
rect 23158 13280 23204 13308
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 26068 13316 26096 13348
rect 26328 13344 26340 13378
rect 26374 13376 26386 13378
rect 26970 13376 26976 13388
rect 26374 13348 26976 13376
rect 26374 13344 26386 13348
rect 26328 13338 26386 13344
rect 26970 13336 26976 13348
rect 27028 13336 27034 13388
rect 27248 13378 27306 13384
rect 27248 13344 27260 13378
rect 27294 13376 27306 13378
rect 34700 13378 34758 13384
rect 34700 13376 34712 13378
rect 27294 13348 34712 13376
rect 27294 13344 27306 13348
rect 27248 13338 27306 13344
rect 34700 13344 34712 13348
rect 34746 13376 34758 13378
rect 37552 13378 37610 13384
rect 34746 13348 37044 13376
rect 34746 13344 34758 13348
rect 34700 13338 34758 13344
rect 26052 13310 26110 13316
rect 26052 13276 26064 13310
rect 26098 13276 26110 13310
rect 29822 13308 29828 13320
rect 29782 13280 29828 13308
rect 26052 13270 26110 13276
rect 26068 13240 26096 13270
rect 29822 13268 29828 13280
rect 29880 13268 29886 13320
rect 32398 13308 32404 13320
rect 32358 13280 32404 13308
rect 32398 13268 32404 13280
rect 32456 13268 32462 13320
rect 33778 13268 33784 13320
rect 33836 13268 33842 13320
rect 37016 13308 37044 13348
rect 37552 13344 37564 13378
rect 37598 13376 37610 13378
rect 44192 13376 44220 13404
rect 37598 13348 44220 13376
rect 37598 13344 37610 13348
rect 37552 13338 37610 13344
rect 44284 13320 44312 13406
rect 44358 13404 44364 13456
rect 44416 13444 44422 13456
rect 44416 13416 51856 13444
rect 44416 13404 44422 13416
rect 45554 13336 45560 13388
rect 45612 13376 45618 13388
rect 51626 13376 51632 13388
rect 45612 13348 45656 13376
rect 51586 13348 51632 13376
rect 45612 13336 45618 13348
rect 51626 13336 51632 13348
rect 51684 13336 51690 13388
rect 51828 13376 51856 13416
rect 59814 13404 59820 13456
rect 59872 13444 59878 13456
rect 60460 13446 60518 13452
rect 60460 13444 60472 13446
rect 59872 13416 60472 13444
rect 59872 13404 59878 13416
rect 60460 13412 60472 13416
rect 60506 13412 60518 13446
rect 63034 13444 63040 13456
rect 62994 13416 63040 13444
rect 60460 13406 60518 13412
rect 63034 13404 63040 13416
rect 63092 13404 63098 13456
rect 75362 13444 75368 13456
rect 63144 13416 73660 13444
rect 75322 13416 75368 13444
rect 63144 13376 63172 13416
rect 72694 13376 72700 13388
rect 51828 13348 63172 13376
rect 64846 13348 69428 13376
rect 72654 13348 72700 13376
rect 37016 13280 37596 13308
rect 27522 13240 27528 13252
rect 7852 13212 22094 13240
rect 26068 13212 27384 13240
rect 27482 13212 27528 13240
rect 22066 13172 22094 13212
rect 26144 13174 26202 13180
rect 26144 13172 26156 13174
rect 22066 13144 26156 13172
rect 26144 13140 26156 13144
rect 26190 13172 26202 13174
rect 27246 13172 27252 13184
rect 26190 13144 27252 13172
rect 26190 13140 26202 13144
rect 26144 13134 26202 13140
rect 27246 13132 27252 13144
rect 27304 13132 27310 13184
rect 27356 13172 27384 13212
rect 27522 13200 27528 13212
rect 27580 13200 27586 13252
rect 30100 13242 30158 13248
rect 28750 13212 29224 13240
rect 27706 13172 27712 13184
rect 27356 13144 27712 13172
rect 27706 13132 27712 13144
rect 27764 13132 27770 13184
rect 29196 13172 29224 13212
rect 30100 13208 30112 13242
rect 30146 13240 30158 13242
rect 30190 13240 30196 13252
rect 30146 13212 30196 13240
rect 30146 13208 30158 13212
rect 30100 13202 30158 13208
rect 30190 13200 30196 13212
rect 30248 13200 30254 13252
rect 32674 13240 32680 13252
rect 31326 13212 31754 13240
rect 32634 13212 32680 13240
rect 30466 13172 30472 13184
rect 29196 13144 30472 13172
rect 30466 13132 30472 13144
rect 30524 13132 30530 13184
rect 31726 13172 31754 13212
rect 32674 13200 32680 13212
rect 32732 13200 32738 13252
rect 34514 13200 34520 13252
rect 34572 13240 34578 13252
rect 34976 13242 35034 13248
rect 34976 13240 34988 13242
rect 34572 13212 34988 13240
rect 34572 13200 34578 13212
rect 34976 13208 34988 13212
rect 35022 13208 35034 13242
rect 34976 13202 35034 13208
rect 35986 13200 35992 13252
rect 36044 13200 36050 13252
rect 33594 13172 33600 13184
rect 31726 13144 33600 13172
rect 33594 13132 33600 13144
rect 33652 13132 33658 13184
rect 34146 13172 34152 13184
rect 34106 13144 34152 13172
rect 34146 13132 34152 13144
rect 34204 13132 34210 13184
rect 34330 13132 34336 13184
rect 34388 13172 34394 13184
rect 36448 13174 36506 13180
rect 36448 13172 36460 13174
rect 34388 13144 36460 13172
rect 34388 13132 34394 13144
rect 36448 13140 36460 13144
rect 36494 13172 36506 13174
rect 37458 13172 37464 13184
rect 36494 13144 37464 13172
rect 36494 13140 36506 13144
rect 36448 13134 36506 13140
rect 37458 13132 37464 13144
rect 37516 13132 37522 13184
rect 37568 13172 37596 13280
rect 38930 13268 38936 13320
rect 38988 13268 38994 13320
rect 40128 13310 40186 13316
rect 40128 13308 40140 13310
rect 39132 13280 40140 13308
rect 37826 13240 37832 13252
rect 37786 13212 37832 13240
rect 37826 13200 37832 13212
rect 37884 13200 37890 13252
rect 39132 13172 39160 13280
rect 40128 13276 40140 13280
rect 40174 13276 40186 13310
rect 42518 13308 42524 13320
rect 42478 13280 42524 13308
rect 40128 13270 40186 13276
rect 39298 13172 39304 13184
rect 37568 13144 39160 13172
rect 39258 13144 39304 13172
rect 39298 13132 39304 13144
rect 39356 13172 39362 13184
rect 39942 13172 39948 13184
rect 39356 13144 39948 13172
rect 39356 13132 39362 13144
rect 39942 13132 39948 13144
rect 40000 13132 40006 13184
rect 40144 13172 40172 13270
rect 42518 13268 42524 13280
rect 42576 13268 42582 13320
rect 44266 13268 44272 13320
rect 44324 13308 44330 13320
rect 47764 13310 47822 13316
rect 47764 13308 47776 13310
rect 44324 13280 47776 13308
rect 44324 13268 44330 13280
rect 47764 13276 47776 13280
rect 47810 13276 47822 13310
rect 47764 13270 47822 13276
rect 50524 13310 50582 13316
rect 50524 13276 50536 13310
rect 50570 13308 50582 13310
rect 51350 13308 51356 13320
rect 50570 13280 51356 13308
rect 50570 13276 50582 13280
rect 50524 13270 50582 13276
rect 40402 13240 40408 13252
rect 40362 13212 40408 13240
rect 40402 13200 40408 13212
rect 40460 13200 40466 13252
rect 41414 13200 41420 13252
rect 41472 13200 41478 13252
rect 42536 13240 42564 13268
rect 41800 13212 42564 13240
rect 42796 13242 42854 13248
rect 41800 13172 41828 13212
rect 42796 13208 42808 13242
rect 42842 13240 42854 13242
rect 42886 13240 42892 13252
rect 42842 13212 42892 13240
rect 42842 13208 42854 13212
rect 42796 13202 42854 13208
rect 42886 13200 42892 13212
rect 42944 13200 42950 13252
rect 43254 13200 43260 13252
rect 43312 13200 43318 13252
rect 45464 13242 45522 13248
rect 45464 13240 45476 13242
rect 44468 13212 45476 13240
rect 40144 13144 41828 13172
rect 41876 13174 41934 13180
rect 41876 13140 41888 13174
rect 41922 13172 41934 13174
rect 42426 13172 42432 13184
rect 41922 13144 42432 13172
rect 41922 13140 41934 13144
rect 41876 13134 41934 13140
rect 42426 13132 42432 13144
rect 42484 13172 42490 13184
rect 44468 13172 44496 13212
rect 45464 13208 45476 13212
rect 45510 13208 45522 13242
rect 45464 13202 45522 13208
rect 45002 13172 45008 13184
rect 42484 13144 44496 13172
rect 44962 13144 45008 13172
rect 42484 13132 42490 13144
rect 45002 13132 45008 13144
rect 45060 13132 45066 13184
rect 45370 13172 45376 13184
rect 45330 13144 45376 13172
rect 45370 13132 45376 13144
rect 45428 13132 45434 13184
rect 47780 13172 47808 13270
rect 51350 13268 51356 13280
rect 51408 13268 51414 13320
rect 53008 13310 53066 13316
rect 53008 13276 53020 13310
rect 53054 13276 53066 13310
rect 53008 13270 53066 13276
rect 47854 13200 47860 13252
rect 47912 13240 47918 13252
rect 53024 13240 53052 13270
rect 54386 13268 54392 13320
rect 54444 13268 54450 13320
rect 54754 13268 54760 13320
rect 54812 13308 54818 13320
rect 55582 13308 55588 13320
rect 54812 13280 55588 13308
rect 54812 13268 54818 13280
rect 55582 13268 55588 13280
rect 55640 13268 55646 13320
rect 57882 13308 57888 13320
rect 57842 13280 57888 13308
rect 57882 13268 57888 13280
rect 57940 13268 57946 13320
rect 60642 13308 60648 13320
rect 60602 13280 60648 13308
rect 60642 13268 60648 13280
rect 60700 13268 60706 13320
rect 63220 13310 63278 13316
rect 63220 13308 63232 13310
rect 61580 13280 63232 13308
rect 53282 13240 53288 13252
rect 47912 13212 53052 13240
rect 53242 13212 53288 13240
rect 47912 13200 47918 13212
rect 51444 13174 51502 13180
rect 51444 13172 51456 13174
rect 47780 13144 51456 13172
rect 51444 13140 51456 13144
rect 51490 13140 51502 13174
rect 53024 13172 53052 13212
rect 53282 13200 53288 13212
rect 53340 13200 53346 13252
rect 55858 13240 55864 13252
rect 54588 13212 54984 13240
rect 55818 13212 55864 13240
rect 54588 13172 54616 13212
rect 53024 13144 54616 13172
rect 51444 13134 51502 13140
rect 54662 13132 54668 13184
rect 54720 13172 54726 13184
rect 54756 13174 54814 13180
rect 54756 13172 54768 13174
rect 54720 13144 54768 13172
rect 54720 13132 54726 13144
rect 54756 13140 54768 13144
rect 54802 13140 54814 13174
rect 54956 13172 54984 13212
rect 55858 13200 55864 13212
rect 55916 13200 55922 13252
rect 56594 13200 56600 13252
rect 56652 13200 56658 13252
rect 57164 13212 57468 13240
rect 57164 13172 57192 13212
rect 57330 13172 57336 13184
rect 54956 13144 57192 13172
rect 57290 13144 57336 13172
rect 54756 13134 54814 13140
rect 57330 13132 57336 13144
rect 57388 13132 57394 13184
rect 57440 13172 57468 13212
rect 57698 13200 57704 13252
rect 57756 13240 57762 13252
rect 58160 13242 58218 13248
rect 58160 13240 58172 13242
rect 57756 13212 58172 13240
rect 57756 13200 57762 13212
rect 58160 13208 58172 13212
rect 58206 13208 58218 13242
rect 58160 13202 58218 13208
rect 58618 13200 58624 13252
rect 58676 13200 58682 13252
rect 61470 13240 61476 13252
rect 59464 13212 61476 13240
rect 59464 13172 59492 13212
rect 61470 13200 61476 13212
rect 61528 13200 61534 13252
rect 59630 13172 59636 13184
rect 57440 13144 59492 13172
rect 59590 13144 59636 13172
rect 59630 13132 59636 13144
rect 59688 13172 59694 13184
rect 61580 13172 61608 13280
rect 63220 13276 63232 13280
rect 63266 13308 63278 13310
rect 64846 13308 64874 13348
rect 66162 13308 66168 13320
rect 63266 13304 63356 13308
rect 63420 13304 64874 13308
rect 63266 13280 64874 13304
rect 66122 13280 66168 13308
rect 63266 13276 63278 13280
rect 63328 13276 63448 13280
rect 63220 13270 63278 13276
rect 66162 13268 66168 13280
rect 66220 13268 66226 13320
rect 69290 13308 69296 13320
rect 69250 13280 69296 13308
rect 69290 13268 69296 13280
rect 69348 13268 69354 13320
rect 69400 13308 69428 13348
rect 72694 13336 72700 13348
rect 72752 13336 72758 13388
rect 73632 13384 73660 13416
rect 75362 13404 75368 13416
rect 75420 13444 75426 13456
rect 75638 13444 75644 13456
rect 75420 13416 75644 13444
rect 75420 13404 75426 13416
rect 75638 13404 75644 13416
rect 75696 13404 75702 13456
rect 80026 13416 82492 13444
rect 73616 13378 73674 13384
rect 73616 13344 73628 13378
rect 73662 13376 73674 13378
rect 78492 13378 78550 13384
rect 78492 13376 78504 13378
rect 73662 13348 78504 13376
rect 73662 13344 73674 13348
rect 73616 13338 73674 13344
rect 78492 13344 78504 13348
rect 78538 13376 78550 13378
rect 80026 13376 80054 13416
rect 80238 13376 80244 13388
rect 78538 13348 80054 13376
rect 80150 13348 80244 13376
rect 78538 13344 78550 13348
rect 78492 13338 78550 13344
rect 80238 13336 80244 13348
rect 80296 13376 80302 13388
rect 81528 13378 81586 13384
rect 81528 13376 81540 13378
rect 80296 13348 81540 13376
rect 80296 13336 80302 13348
rect 81528 13344 81540 13348
rect 81574 13344 81586 13378
rect 81528 13338 81586 13344
rect 81618 13336 81624 13388
rect 81676 13376 81682 13388
rect 82464 13376 82492 13416
rect 93854 13404 93860 13456
rect 93912 13444 93918 13456
rect 93948 13446 94006 13452
rect 93948 13444 93960 13446
rect 93912 13416 93960 13444
rect 93912 13404 93918 13416
rect 93948 13412 93960 13416
rect 93994 13412 94006 13446
rect 93948 13406 94006 13412
rect 94516 13416 99374 13444
rect 94516 13376 94544 13416
rect 97996 13378 98054 13384
rect 97996 13376 98008 13378
rect 81676 13348 81720 13376
rect 82464 13348 94544 13376
rect 94608 13348 98008 13376
rect 81676 13336 81682 13348
rect 72512 13310 72570 13316
rect 72512 13308 72524 13310
rect 69400 13280 72524 13308
rect 72512 13276 72524 13280
rect 72558 13276 72570 13310
rect 72512 13270 72570 13276
rect 76192 13310 76250 13316
rect 76192 13276 76204 13310
rect 76238 13276 76250 13310
rect 78398 13308 78404 13320
rect 77602 13280 78404 13308
rect 76192 13270 76250 13276
rect 61746 13200 61752 13252
rect 61804 13240 61810 13252
rect 61804 13212 73844 13240
rect 61804 13200 61810 13212
rect 59688 13144 61608 13172
rect 59688 13132 59694 13144
rect 61654 13132 61660 13184
rect 61712 13172 61718 13184
rect 65886 13172 65892 13184
rect 61712 13144 65892 13172
rect 61712 13132 61718 13144
rect 65886 13132 65892 13144
rect 65944 13132 65950 13184
rect 65978 13132 65984 13184
rect 66036 13172 66042 13184
rect 69106 13172 69112 13184
rect 66036 13144 66080 13172
rect 69066 13144 69112 13172
rect 66036 13132 66042 13144
rect 69106 13132 69112 13144
rect 69164 13132 69170 13184
rect 72052 13174 72110 13180
rect 72052 13140 72064 13174
rect 72098 13172 72110 13174
rect 72326 13172 72332 13184
rect 72098 13144 72332 13172
rect 72098 13140 72110 13144
rect 72052 13134 72110 13140
rect 72326 13132 72332 13144
rect 72384 13132 72390 13184
rect 72418 13132 72424 13184
rect 72476 13172 72482 13184
rect 73816 13172 73844 13212
rect 73890 13200 73896 13252
rect 73948 13240 73954 13252
rect 75178 13240 75184 13252
rect 73948 13212 73992 13240
rect 75118 13212 75184 13240
rect 73948 13200 73954 13212
rect 75178 13200 75184 13212
rect 75236 13200 75242 13252
rect 76208 13172 76236 13270
rect 78398 13268 78404 13280
rect 78456 13268 78462 13320
rect 81434 13268 81440 13320
rect 81492 13268 81498 13320
rect 82448 13310 82506 13316
rect 82448 13276 82460 13310
rect 82494 13276 82506 13310
rect 83090 13308 83096 13320
rect 83050 13280 83096 13308
rect 82448 13270 82506 13276
rect 76466 13240 76472 13252
rect 76426 13212 76472 13240
rect 76466 13200 76472 13212
rect 76524 13200 76530 13252
rect 78766 13240 78772 13252
rect 77864 13212 78168 13240
rect 78726 13212 78772 13240
rect 77864 13172 77892 13212
rect 72476 13144 72520 13172
rect 73816 13144 77892 13172
rect 72476 13132 72482 13144
rect 77938 13132 77944 13184
rect 77996 13172 78002 13184
rect 78140 13172 78168 13212
rect 78766 13200 78772 13212
rect 78824 13200 78830 13252
rect 79318 13200 79324 13252
rect 79376 13200 79382 13252
rect 80054 13200 80060 13252
rect 80112 13240 80118 13252
rect 81452 13240 81480 13268
rect 82464 13240 82492 13270
rect 83090 13268 83096 13280
rect 83148 13268 83154 13320
rect 83918 13308 83924 13320
rect 83878 13280 83924 13308
rect 83918 13268 83924 13280
rect 83976 13268 83982 13320
rect 86496 13310 86554 13316
rect 86496 13308 86508 13310
rect 85592 13280 86508 13308
rect 83826 13240 83832 13252
rect 80112 13212 81112 13240
rect 81452 13212 82308 13240
rect 82464 13212 83832 13240
rect 80112 13200 80118 13212
rect 80790 13172 80796 13184
rect 77996 13144 78040 13172
rect 78140 13144 80796 13172
rect 77996 13132 78002 13144
rect 80790 13132 80796 13144
rect 80848 13132 80854 13184
rect 81084 13180 81112 13212
rect 81068 13174 81126 13180
rect 81068 13140 81080 13174
rect 81114 13140 81126 13174
rect 81434 13172 81440 13184
rect 81394 13144 81440 13172
rect 81068 13134 81126 13140
rect 81434 13132 81440 13144
rect 81492 13132 81498 13184
rect 82280 13180 82308 13212
rect 83826 13200 83832 13212
rect 83884 13200 83890 13252
rect 84196 13242 84254 13248
rect 84196 13208 84208 13242
rect 84242 13240 84254 13242
rect 84470 13240 84476 13252
rect 84242 13212 84476 13240
rect 84242 13208 84254 13212
rect 84196 13202 84254 13208
rect 84470 13200 84476 13212
rect 84528 13200 84534 13252
rect 85482 13240 85488 13252
rect 85422 13212 85488 13240
rect 85482 13200 85488 13212
rect 85540 13200 85546 13252
rect 82264 13174 82322 13180
rect 82264 13140 82276 13174
rect 82310 13140 82322 13174
rect 82906 13172 82912 13184
rect 82866 13144 82912 13172
rect 82264 13134 82322 13140
rect 82906 13132 82912 13144
rect 82964 13132 82970 13184
rect 83918 13132 83924 13184
rect 83976 13172 83982 13184
rect 85592 13172 85620 13280
rect 86496 13276 86508 13280
rect 86542 13276 86554 13310
rect 86496 13270 86554 13276
rect 83976 13144 85620 13172
rect 85668 13174 85726 13180
rect 83976 13132 83982 13144
rect 85668 13140 85680 13174
rect 85714 13172 85726 13174
rect 86034 13172 86040 13184
rect 85714 13144 86040 13172
rect 85714 13140 85726 13144
rect 85668 13134 85726 13140
rect 86034 13132 86040 13144
rect 86092 13132 86098 13184
rect 86512 13172 86540 13270
rect 87874 13268 87880 13320
rect 87932 13268 87938 13320
rect 88796 13310 88854 13316
rect 88796 13308 88808 13310
rect 88076 13280 88808 13308
rect 86770 13240 86776 13252
rect 86730 13212 86776 13240
rect 86770 13200 86776 13212
rect 86828 13200 86834 13252
rect 88076 13172 88104 13280
rect 88796 13276 88808 13280
rect 88842 13276 88854 13310
rect 94132 13310 94190 13316
rect 94132 13308 94144 13310
rect 88796 13270 88854 13276
rect 93136 13280 94144 13308
rect 88242 13172 88248 13184
rect 86512 13144 88104 13172
rect 88202 13144 88248 13172
rect 88242 13132 88248 13144
rect 88300 13132 88306 13184
rect 88812 13172 88840 13270
rect 89070 13240 89076 13252
rect 89030 13212 89076 13240
rect 89070 13200 89076 13212
rect 89128 13200 89134 13252
rect 89530 13200 89536 13252
rect 89588 13200 89594 13252
rect 91646 13240 91652 13252
rect 90468 13212 91652 13240
rect 90468 13172 90496 13212
rect 91646 13200 91652 13212
rect 91704 13200 91710 13252
rect 91830 13240 91836 13252
rect 91790 13212 91836 13240
rect 91830 13200 91836 13212
rect 91888 13200 91894 13252
rect 92014 13240 92020 13252
rect 91974 13212 92020 13240
rect 92014 13200 92020 13212
rect 92072 13200 92078 13252
rect 88812 13144 90496 13172
rect 90542 13132 90548 13184
rect 90600 13172 90606 13184
rect 93136 13172 93164 13280
rect 94132 13276 94144 13280
rect 94178 13308 94190 13310
rect 94608 13308 94636 13348
rect 97996 13344 98008 13348
rect 98042 13344 98054 13378
rect 97996 13338 98054 13344
rect 98180 13378 98238 13384
rect 98180 13344 98192 13378
rect 98226 13376 98238 13378
rect 99098 13376 99104 13388
rect 98226 13348 99104 13376
rect 98226 13344 98238 13348
rect 98180 13338 98238 13344
rect 99098 13336 99104 13348
rect 99156 13336 99162 13388
rect 99346 13376 99374 13416
rect 100754 13404 100760 13456
rect 100812 13444 100818 13456
rect 101124 13446 101182 13452
rect 101124 13444 101136 13446
rect 100812 13416 101136 13444
rect 100812 13404 100818 13416
rect 101124 13412 101136 13416
rect 101170 13412 101182 13446
rect 101124 13406 101182 13412
rect 109034 13404 109040 13456
rect 109092 13444 109098 13456
rect 109404 13446 109462 13452
rect 109404 13444 109416 13446
rect 109092 13416 109416 13444
rect 109092 13404 109098 13416
rect 109404 13412 109416 13416
rect 109450 13412 109462 13446
rect 109404 13406 109462 13412
rect 111244 13446 111302 13452
rect 111244 13412 111256 13446
rect 111290 13444 111302 13446
rect 111702 13444 111708 13456
rect 111290 13416 111708 13444
rect 111290 13412 111302 13416
rect 111244 13406 111302 13412
rect 111702 13404 111708 13416
rect 111760 13404 111766 13456
rect 118878 13404 118884 13456
rect 118936 13444 118942 13456
rect 121270 13444 121276 13456
rect 118936 13416 120304 13444
rect 121230 13416 121276 13444
rect 118936 13404 118942 13416
rect 112256 13378 112314 13384
rect 112256 13376 112268 13378
rect 99346 13348 112268 13376
rect 112256 13344 112268 13348
rect 112302 13376 112314 13378
rect 112302 13348 114876 13376
rect 112302 13344 112314 13348
rect 112256 13338 112314 13344
rect 114848 13320 114876 13348
rect 118234 13336 118240 13388
rect 118292 13376 118298 13388
rect 120276 13384 120304 13416
rect 121270 13404 121276 13416
rect 121328 13404 121334 13456
rect 124122 13444 124128 13456
rect 124082 13416 124128 13444
rect 124122 13404 124128 13416
rect 124180 13404 124186 13456
rect 127526 13444 127532 13456
rect 126716 13416 127532 13444
rect 126716 13384 126744 13416
rect 127526 13404 127532 13416
rect 127584 13404 127590 13456
rect 136634 13444 136640 13456
rect 136594 13416 136640 13444
rect 136634 13404 136640 13416
rect 136692 13404 136698 13456
rect 139578 13404 139584 13456
rect 139636 13444 139642 13456
rect 140316 13446 140374 13452
rect 140316 13444 140328 13446
rect 139636 13416 140328 13444
rect 139636 13404 139642 13416
rect 140316 13412 140328 13416
rect 140362 13412 140374 13446
rect 142126 13444 142154 13484
rect 142890 13472 142896 13484
rect 142948 13472 142954 13524
rect 144732 13514 144790 13520
rect 144732 13480 144744 13514
rect 144778 13512 144790 13514
rect 145742 13512 145748 13524
rect 144778 13484 145748 13512
rect 144778 13480 144790 13484
rect 144732 13474 144790 13480
rect 145742 13472 145748 13484
rect 145800 13472 145806 13524
rect 148134 13512 148140 13524
rect 145852 13484 148140 13512
rect 145852 13444 145880 13484
rect 148134 13472 148140 13484
rect 148192 13472 148198 13524
rect 148308 13514 148366 13520
rect 148308 13480 148320 13514
rect 148354 13512 148366 13514
rect 150802 13512 150808 13524
rect 148354 13484 150808 13512
rect 148354 13480 148366 13484
rect 148308 13474 148366 13480
rect 150802 13472 150808 13484
rect 150860 13472 150866 13524
rect 157242 13512 157248 13524
rect 152200 13484 157248 13512
rect 142126 13416 145880 13444
rect 140316 13406 140374 13412
rect 120260 13378 120318 13384
rect 118292 13348 120212 13376
rect 118292 13336 118298 13348
rect 94178 13280 94636 13308
rect 96892 13310 96950 13316
rect 94178 13276 94190 13280
rect 94132 13270 94190 13276
rect 96892 13276 96904 13310
rect 96938 13308 96950 13310
rect 99376 13310 99434 13316
rect 96938 13280 97948 13308
rect 96938 13276 96950 13280
rect 96892 13270 96950 13276
rect 96706 13172 96712 13184
rect 90600 13144 93164 13172
rect 96666 13144 96712 13172
rect 90600 13132 90606 13144
rect 96706 13132 96712 13144
rect 96764 13132 96770 13184
rect 97534 13172 97540 13184
rect 97494 13144 97540 13172
rect 97534 13132 97540 13144
rect 97592 13132 97598 13184
rect 97920 13180 97948 13280
rect 99376 13276 99388 13310
rect 99422 13276 99434 13310
rect 99376 13270 99434 13276
rect 97994 13200 98000 13252
rect 98052 13240 98058 13252
rect 99190 13240 99196 13252
rect 98052 13212 99196 13240
rect 98052 13200 98058 13212
rect 99190 13200 99196 13212
rect 99248 13240 99254 13252
rect 99392 13240 99420 13270
rect 101398 13268 101404 13320
rect 101456 13308 101462 13320
rect 101952 13310 102010 13316
rect 101952 13308 101964 13310
rect 101456 13280 101964 13308
rect 101456 13268 101462 13280
rect 101952 13276 101964 13280
rect 101998 13276 102010 13310
rect 101952 13270 102010 13276
rect 99650 13240 99656 13252
rect 99248 13212 99420 13240
rect 99610 13212 99656 13240
rect 99248 13200 99254 13212
rect 99650 13200 99656 13212
rect 99708 13200 99714 13252
rect 100938 13240 100944 13252
rect 100878 13212 100944 13240
rect 100938 13200 100944 13212
rect 100996 13200 101002 13252
rect 97904 13174 97962 13180
rect 97904 13140 97916 13174
rect 97950 13172 97962 13174
rect 101030 13172 101036 13184
rect 97950 13144 101036 13172
rect 97950 13140 97962 13144
rect 97904 13134 97962 13140
rect 101030 13132 101036 13144
rect 101088 13132 101094 13184
rect 101968 13172 101996 13270
rect 103330 13268 103336 13320
rect 103388 13268 103394 13320
rect 104250 13308 104256 13320
rect 103532 13280 104256 13308
rect 102226 13240 102232 13252
rect 102186 13212 102232 13240
rect 102226 13200 102232 13212
rect 102284 13200 102290 13252
rect 103532 13172 103560 13280
rect 104250 13268 104256 13280
rect 104308 13268 104314 13320
rect 109586 13308 109592 13320
rect 109546 13280 109592 13308
rect 109586 13268 109592 13280
rect 109644 13268 109650 13320
rect 111426 13308 111432 13320
rect 111386 13280 111432 13308
rect 111426 13268 111432 13280
rect 111484 13268 111490 13320
rect 114830 13308 114836 13320
rect 114790 13280 114836 13308
rect 114830 13268 114836 13280
rect 114888 13268 114894 13320
rect 117406 13308 117412 13320
rect 117366 13280 117412 13308
rect 117406 13268 117412 13280
rect 117464 13268 117470 13320
rect 118786 13268 118792 13320
rect 118844 13268 118850 13320
rect 120184 13316 120212 13348
rect 120260 13344 120272 13378
rect 120306 13344 120318 13378
rect 120260 13338 120318 13344
rect 125688 13378 125746 13384
rect 125688 13344 125700 13378
rect 125734 13376 125746 13378
rect 126700 13378 126758 13384
rect 126700 13376 126712 13378
rect 125734 13348 126712 13376
rect 125734 13344 125746 13348
rect 125688 13338 125746 13344
rect 126700 13344 126712 13348
rect 126746 13344 126758 13378
rect 130286 13376 130292 13388
rect 126700 13338 126758 13344
rect 127544 13348 130292 13376
rect 127544 13320 127572 13348
rect 130286 13336 130292 13348
rect 130344 13376 130350 13388
rect 132588 13378 132646 13384
rect 132588 13376 132600 13378
rect 130344 13348 132600 13376
rect 130344 13336 130350 13348
rect 132588 13344 132600 13348
rect 132634 13376 132646 13378
rect 142062 13376 142068 13388
rect 132634 13348 142068 13376
rect 132634 13344 132646 13348
rect 132588 13338 132646 13344
rect 142062 13336 142068 13348
rect 142120 13336 142126 13388
rect 148044 13378 148102 13384
rect 144932 13348 147674 13376
rect 120168 13310 120226 13316
rect 120168 13276 120180 13310
rect 120214 13308 120226 13310
rect 121456 13310 121514 13316
rect 121456 13308 121468 13310
rect 120214 13280 121468 13308
rect 120214 13276 120226 13280
rect 120168 13270 120226 13276
rect 121456 13276 121468 13280
rect 121502 13276 121514 13310
rect 124308 13310 124366 13316
rect 124308 13308 124320 13310
rect 121456 13270 121514 13276
rect 122806 13280 124320 13308
rect 104066 13200 104072 13252
rect 104124 13240 104130 13252
rect 104528 13242 104586 13248
rect 104528 13240 104540 13242
rect 104124 13212 104540 13240
rect 104124 13200 104130 13212
rect 104528 13208 104540 13212
rect 104574 13208 104586 13242
rect 104528 13202 104586 13208
rect 104986 13200 104992 13252
rect 105044 13200 105050 13252
rect 112530 13240 112536 13252
rect 112490 13212 112536 13240
rect 112530 13200 112536 13212
rect 112588 13200 112594 13252
rect 114186 13240 114192 13252
rect 113758 13212 114192 13240
rect 114186 13200 114192 13212
rect 114244 13200 114250 13252
rect 115106 13240 115112 13252
rect 115066 13212 115112 13240
rect 115106 13200 115112 13212
rect 115164 13200 115170 13252
rect 116946 13240 116952 13252
rect 116334 13212 116952 13240
rect 116946 13200 116952 13212
rect 117004 13200 117010 13252
rect 117682 13240 117688 13252
rect 117642 13212 117688 13240
rect 117682 13200 117688 13212
rect 117740 13200 117746 13252
rect 120076 13242 120134 13248
rect 120076 13240 120088 13242
rect 119172 13212 120088 13240
rect 101968 13144 103560 13172
rect 103698 13132 103704 13184
rect 103756 13172 103762 13184
rect 104434 13172 104440 13184
rect 103756 13144 104440 13172
rect 103756 13132 103762 13144
rect 104434 13132 104440 13144
rect 104492 13132 104498 13184
rect 104618 13132 104624 13184
rect 104676 13172 104682 13184
rect 106000 13174 106058 13180
rect 106000 13172 106012 13174
rect 104676 13144 106012 13172
rect 104676 13132 104682 13144
rect 106000 13140 106012 13144
rect 106046 13172 106058 13174
rect 109586 13172 109592 13184
rect 106046 13144 109592 13172
rect 106046 13140 106058 13144
rect 106000 13134 106058 13140
rect 109586 13132 109592 13144
rect 109644 13132 109650 13184
rect 114004 13174 114062 13180
rect 114004 13140 114016 13174
rect 114050 13172 114062 13174
rect 114554 13172 114560 13184
rect 114050 13144 114560 13172
rect 114050 13140 114062 13144
rect 114004 13134 114062 13140
rect 114554 13132 114560 13144
rect 114612 13172 114618 13184
rect 114922 13172 114928 13184
rect 114612 13144 114928 13172
rect 114612 13132 114618 13144
rect 114922 13132 114928 13144
rect 114980 13132 114986 13184
rect 115750 13132 115756 13184
rect 115808 13172 115814 13184
rect 116580 13174 116638 13180
rect 116580 13172 116592 13174
rect 115808 13144 116592 13172
rect 115808 13132 115814 13144
rect 116580 13140 116592 13144
rect 116626 13172 116638 13174
rect 118050 13172 118056 13184
rect 116626 13144 118056 13172
rect 116626 13140 116638 13144
rect 116580 13134 116638 13140
rect 118050 13132 118056 13144
rect 118108 13132 118114 13184
rect 119172 13180 119200 13212
rect 120076 13208 120088 13212
rect 120122 13240 120134 13242
rect 122806 13240 122834 13280
rect 124308 13276 124320 13280
rect 124354 13308 124366 13310
rect 126608 13310 126666 13316
rect 126608 13308 126620 13310
rect 124354 13280 126620 13308
rect 124354 13276 124366 13280
rect 124308 13270 124366 13276
rect 126608 13276 126620 13280
rect 126654 13276 126666 13310
rect 127526 13308 127532 13320
rect 127486 13280 127532 13308
rect 126608 13270 126666 13276
rect 127526 13268 127532 13280
rect 127584 13268 127590 13320
rect 129366 13308 129372 13320
rect 128938 13280 129372 13308
rect 129366 13268 129372 13280
rect 129424 13268 129430 13320
rect 136818 13308 136824 13320
rect 136778 13280 136824 13308
rect 136818 13268 136824 13280
rect 136876 13268 136882 13320
rect 140500 13310 140558 13316
rect 140500 13276 140512 13310
rect 140546 13276 140558 13310
rect 143074 13308 143080 13320
rect 143034 13280 143080 13308
rect 140500 13270 140558 13276
rect 125502 13240 125508 13252
rect 120122 13212 122834 13240
rect 125462 13212 125508 13240
rect 120122 13208 120134 13212
rect 120076 13202 120134 13208
rect 125502 13200 125508 13212
rect 125560 13200 125566 13252
rect 127802 13240 127808 13252
rect 127762 13212 127808 13240
rect 127802 13200 127808 13212
rect 127860 13200 127866 13252
rect 130564 13242 130622 13248
rect 130564 13240 130576 13242
rect 129108 13212 130576 13240
rect 119156 13174 119214 13180
rect 119156 13140 119168 13174
rect 119202 13140 119214 13174
rect 119706 13172 119712 13184
rect 119666 13144 119712 13172
rect 119156 13134 119214 13140
rect 119706 13132 119712 13144
rect 119764 13132 119770 13184
rect 126146 13172 126152 13184
rect 126106 13144 126152 13172
rect 126146 13132 126152 13144
rect 126204 13132 126210 13184
rect 126514 13172 126520 13184
rect 126474 13144 126520 13172
rect 126514 13132 126520 13144
rect 126572 13132 126578 13184
rect 128078 13132 128084 13184
rect 128136 13172 128142 13184
rect 129108 13172 129136 13212
rect 130564 13208 130576 13212
rect 130610 13208 130622 13242
rect 130564 13202 130622 13208
rect 131206 13200 131212 13252
rect 131264 13200 131270 13252
rect 132862 13240 132868 13252
rect 132822 13212 132868 13240
rect 132862 13200 132868 13212
rect 132920 13200 132926 13252
rect 133322 13200 133328 13252
rect 133380 13200 133386 13252
rect 140516 13240 140544 13270
rect 143074 13268 143080 13280
rect 143132 13268 143138 13320
rect 144932 13316 144960 13348
rect 144916 13310 144974 13316
rect 144916 13276 144928 13310
rect 144962 13276 144974 13310
rect 145742 13308 145748 13320
rect 145702 13280 145748 13308
rect 144916 13270 144974 13276
rect 145742 13268 145748 13280
rect 145800 13268 145806 13320
rect 147646 13308 147674 13348
rect 148044 13344 148056 13378
rect 148090 13376 148102 13378
rect 150896 13378 150954 13384
rect 150896 13376 150908 13378
rect 148090 13348 150908 13376
rect 148090 13344 148102 13348
rect 148044 13338 148102 13344
rect 150896 13344 150908 13348
rect 150942 13376 150954 13378
rect 152200 13376 152228 13484
rect 157242 13472 157248 13484
rect 157300 13472 157306 13524
rect 157612 13514 157670 13520
rect 157612 13480 157624 13514
rect 157658 13512 157670 13514
rect 157978 13512 157984 13524
rect 157658 13484 157984 13512
rect 157658 13480 157670 13484
rect 157612 13474 157670 13480
rect 157978 13472 157984 13484
rect 158036 13472 158042 13524
rect 159450 13472 159456 13524
rect 159508 13512 159514 13524
rect 161566 13512 161572 13524
rect 159508 13484 161572 13512
rect 159508 13472 159514 13484
rect 161566 13472 161572 13484
rect 161624 13512 161630 13524
rect 162670 13512 162676 13524
rect 161624 13484 162676 13512
rect 161624 13472 161630 13484
rect 162670 13472 162676 13484
rect 162728 13472 162734 13524
rect 163498 13472 163504 13524
rect 163556 13512 163562 13524
rect 176378 13512 176384 13524
rect 163556 13484 176384 13512
rect 163556 13472 163562 13484
rect 176378 13472 176384 13484
rect 176436 13472 176442 13524
rect 182726 13512 182732 13524
rect 176488 13484 182588 13512
rect 182686 13484 182732 13512
rect 154942 13404 154948 13456
rect 155000 13444 155006 13456
rect 155772 13446 155830 13452
rect 155772 13444 155784 13446
rect 155000 13416 155784 13444
rect 155000 13404 155006 13416
rect 155772 13412 155784 13416
rect 155818 13412 155830 13446
rect 155772 13406 155830 13412
rect 166442 13404 166448 13456
rect 166500 13444 166506 13456
rect 170398 13444 170404 13456
rect 166500 13416 170260 13444
rect 170358 13416 170404 13444
rect 166500 13404 166506 13416
rect 150942 13348 152228 13376
rect 153472 13378 153530 13384
rect 150942 13344 150954 13348
rect 150896 13338 150954 13344
rect 153472 13344 153484 13378
rect 153518 13376 153530 13378
rect 160922 13376 160928 13388
rect 153518 13348 158668 13376
rect 160834 13348 160928 13376
rect 153518 13344 153530 13348
rect 153472 13338 153530 13344
rect 158640 13320 158668 13348
rect 160922 13336 160928 13348
rect 160980 13376 160986 13388
rect 160980 13348 165108 13376
rect 160980 13336 160986 13348
rect 165080 13324 165108 13348
rect 165246 13336 165252 13388
rect 165304 13376 165310 13388
rect 166628 13378 166686 13384
rect 166628 13376 166640 13378
rect 165304 13348 166640 13376
rect 165304 13336 165310 13348
rect 166628 13344 166640 13348
rect 166674 13376 166686 13378
rect 167548 13378 167606 13384
rect 167548 13376 167560 13378
rect 166674 13348 167560 13376
rect 166674 13344 166686 13348
rect 166628 13338 166686 13344
rect 167548 13344 167560 13348
rect 167594 13344 167606 13378
rect 167548 13338 167606 13344
rect 147646 13280 148088 13308
rect 145926 13240 145932 13252
rect 134352 13212 145932 13240
rect 128136 13144 129136 13172
rect 128136 13132 128142 13144
rect 129182 13132 129188 13184
rect 129240 13172 129246 13184
rect 129276 13174 129334 13180
rect 129276 13172 129288 13174
rect 129240 13144 129288 13172
rect 129240 13132 129246 13144
rect 129276 13140 129288 13144
rect 129322 13140 129334 13174
rect 129276 13134 129334 13140
rect 131574 13132 131580 13184
rect 131632 13172 131638 13184
rect 132036 13174 132094 13180
rect 132036 13172 132048 13174
rect 131632 13144 132048 13172
rect 131632 13132 131638 13144
rect 132036 13140 132048 13144
rect 132082 13172 132094 13174
rect 133690 13172 133696 13184
rect 132082 13144 133696 13172
rect 132082 13140 132094 13144
rect 132036 13134 132094 13140
rect 133690 13132 133696 13144
rect 133748 13132 133754 13184
rect 134150 13132 134156 13184
rect 134208 13172 134214 13184
rect 134352 13180 134380 13212
rect 145926 13200 145932 13212
rect 145984 13200 145990 13252
rect 146018 13200 146024 13252
rect 146076 13240 146082 13252
rect 147582 13240 147588 13252
rect 146076 13212 146120 13240
rect 147246 13212 147588 13240
rect 146076 13200 146082 13212
rect 147582 13200 147588 13212
rect 147640 13200 147646 13252
rect 134336 13174 134394 13180
rect 134336 13172 134348 13174
rect 134208 13144 134348 13172
rect 134208 13132 134214 13144
rect 134336 13140 134348 13144
rect 134382 13140 134394 13174
rect 134336 13134 134394 13140
rect 145834 13132 145840 13184
rect 145892 13172 145898 13184
rect 147490 13172 147496 13184
rect 145892 13144 147496 13172
rect 145892 13132 145898 13144
rect 147490 13132 147496 13144
rect 147548 13132 147554 13184
rect 148060 13172 148088 13280
rect 155218 13268 155224 13320
rect 155276 13308 155282 13320
rect 155862 13308 155868 13320
rect 155276 13280 155868 13308
rect 155276 13268 155282 13280
rect 155862 13268 155868 13280
rect 155920 13308 155926 13320
rect 155956 13310 156014 13316
rect 155956 13308 155968 13310
rect 155920 13280 155968 13308
rect 155920 13268 155926 13280
rect 155956 13276 155968 13280
rect 156002 13276 156014 13310
rect 156414 13308 156420 13320
rect 156374 13280 156420 13308
rect 155956 13270 156014 13276
rect 156414 13268 156420 13280
rect 156472 13268 156478 13320
rect 157794 13308 157800 13320
rect 157754 13280 157800 13308
rect 157794 13268 157800 13280
rect 157852 13268 157858 13320
rect 158622 13308 158628 13320
rect 158582 13280 158628 13308
rect 158622 13268 158628 13280
rect 158680 13268 158686 13320
rect 162670 13268 162676 13320
rect 162728 13308 162734 13320
rect 163498 13308 163504 13320
rect 162728 13280 163360 13308
rect 163458 13280 163504 13308
rect 162728 13268 162734 13280
rect 150068 13242 150126 13248
rect 149546 13212 150020 13240
rect 149238 13172 149244 13184
rect 148060 13144 149244 13172
rect 149238 13132 149244 13144
rect 149296 13132 149302 13184
rect 149992 13172 150020 13212
rect 150068 13208 150080 13242
rect 150114 13240 150126 13242
rect 150434 13240 150440 13252
rect 150114 13212 150440 13240
rect 150114 13208 150126 13212
rect 150068 13202 150126 13208
rect 150434 13200 150440 13212
rect 150492 13200 150498 13252
rect 151078 13200 151084 13252
rect 151136 13240 151142 13252
rect 151172 13242 151230 13248
rect 151172 13240 151184 13242
rect 151136 13212 151184 13240
rect 151136 13200 151142 13212
rect 151172 13208 151184 13212
rect 151218 13208 151230 13242
rect 152458 13240 152464 13252
rect 152398 13212 152464 13240
rect 151172 13202 151230 13208
rect 152458 13200 152464 13212
rect 152516 13200 152522 13252
rect 153746 13240 153752 13252
rect 152568 13212 152872 13240
rect 153706 13212 153752 13240
rect 152568 13172 152596 13212
rect 149992 13144 152596 13172
rect 152642 13132 152648 13184
rect 152700 13172 152706 13184
rect 152844 13172 152872 13212
rect 153746 13200 153752 13212
rect 153804 13200 153810 13252
rect 154206 13200 154212 13252
rect 154264 13200 154270 13252
rect 156508 13242 156566 13248
rect 156508 13240 156520 13242
rect 155052 13212 156520 13240
rect 155052 13172 155080 13212
rect 156508 13208 156520 13212
rect 156554 13208 156566 13242
rect 156508 13202 156566 13208
rect 156598 13200 156604 13252
rect 156656 13240 156662 13252
rect 158898 13240 158904 13252
rect 156656 13212 157334 13240
rect 158858 13212 158904 13240
rect 156656 13200 156662 13212
rect 155218 13172 155224 13184
rect 152700 13144 152744 13172
rect 152844 13144 155080 13172
rect 155178 13144 155224 13172
rect 152700 13132 152706 13144
rect 155218 13132 155224 13144
rect 155276 13132 155282 13184
rect 157306 13172 157334 13212
rect 158898 13200 158904 13212
rect 158956 13200 158962 13252
rect 161198 13240 161204 13252
rect 160126 13212 160692 13240
rect 161158 13212 161204 13240
rect 159542 13172 159548 13184
rect 157306 13144 159548 13172
rect 159542 13132 159548 13144
rect 159600 13132 159606 13184
rect 160370 13172 160376 13184
rect 160330 13144 160376 13172
rect 160370 13132 160376 13144
rect 160428 13132 160434 13184
rect 160664 13172 160692 13212
rect 161198 13200 161204 13212
rect 161256 13200 161262 13252
rect 162762 13240 162768 13252
rect 162426 13212 162768 13240
rect 162762 13200 162768 13212
rect 162820 13200 162826 13252
rect 162026 13172 162032 13184
rect 160664 13144 162032 13172
rect 162026 13132 162032 13144
rect 162084 13132 162090 13184
rect 162486 13132 162492 13184
rect 162544 13172 162550 13184
rect 162672 13174 162730 13180
rect 162672 13172 162684 13174
rect 162544 13144 162684 13172
rect 162544 13132 162550 13144
rect 162672 13140 162684 13144
rect 162718 13140 162730 13174
rect 163332 13172 163360 13280
rect 163498 13268 163504 13280
rect 163556 13268 163562 13320
rect 164878 13268 164884 13320
rect 164936 13268 164942 13320
rect 165080 13308 165200 13324
rect 170232 13308 170260 13416
rect 170398 13404 170404 13416
rect 170456 13404 170462 13456
rect 173066 13444 173072 13456
rect 173026 13416 173072 13444
rect 173066 13404 173072 13416
rect 173124 13404 173130 13456
rect 173802 13444 173808 13456
rect 173762 13416 173808 13444
rect 173802 13404 173808 13416
rect 173860 13404 173866 13456
rect 175828 13446 175886 13452
rect 175828 13444 175840 13446
rect 174372 13416 175840 13444
rect 174372 13384 174400 13416
rect 175828 13412 175840 13416
rect 175874 13444 175886 13446
rect 175918 13444 175924 13456
rect 175874 13416 175924 13444
rect 175874 13412 175886 13416
rect 175828 13406 175886 13412
rect 175918 13404 175924 13416
rect 175976 13404 175982 13456
rect 176010 13404 176016 13456
rect 176068 13444 176074 13456
rect 176488 13444 176516 13484
rect 176068 13416 176516 13444
rect 176068 13404 176074 13416
rect 177758 13404 177764 13456
rect 177816 13444 177822 13456
rect 178128 13446 178186 13452
rect 178128 13444 178140 13446
rect 177816 13416 178140 13444
rect 177816 13404 177822 13416
rect 178128 13412 178140 13416
rect 178174 13412 178186 13446
rect 178128 13406 178186 13412
rect 180426 13404 180432 13456
rect 180484 13444 180490 13456
rect 181532 13446 181590 13452
rect 181532 13444 181544 13446
rect 180484 13416 181544 13444
rect 180484 13404 180490 13416
rect 181532 13412 181544 13416
rect 181578 13412 181590 13446
rect 181532 13406 181590 13412
rect 174264 13378 174322 13384
rect 174264 13376 174276 13378
rect 170600 13348 174276 13376
rect 170600 13316 170628 13348
rect 174264 13344 174276 13348
rect 174310 13344 174322 13378
rect 174264 13338 174322 13344
rect 174356 13378 174414 13384
rect 174356 13344 174368 13378
rect 174402 13344 174414 13378
rect 178956 13378 179014 13384
rect 178956 13376 178968 13378
rect 174356 13338 174414 13344
rect 174464 13348 175964 13376
rect 170584 13310 170642 13316
rect 170584 13308 170596 13310
rect 165080 13296 170168 13308
rect 165172 13280 170168 13296
rect 170232 13280 170596 13308
rect 163774 13240 163780 13252
rect 163734 13212 163780 13240
rect 163774 13200 163780 13212
rect 163832 13200 163838 13252
rect 165154 13240 165160 13252
rect 165080 13212 165160 13240
rect 164602 13172 164608 13184
rect 163332 13144 164608 13172
rect 162672 13134 162730 13140
rect 164602 13132 164608 13144
rect 164660 13172 164666 13184
rect 165080 13172 165108 13212
rect 165154 13200 165160 13212
rect 165212 13200 165218 13252
rect 166536 13242 166594 13248
rect 166536 13240 166548 13242
rect 165264 13212 166548 13240
rect 165264 13184 165292 13212
rect 166536 13208 166548 13212
rect 166582 13208 166594 13242
rect 167362 13240 167368 13252
rect 167274 13212 167368 13240
rect 166536 13202 166594 13208
rect 167362 13200 167368 13212
rect 167420 13200 167426 13252
rect 170140 13240 170168 13280
rect 170584 13276 170596 13280
rect 170630 13276 170642 13310
rect 170584 13270 170642 13276
rect 173252 13310 173310 13316
rect 173252 13276 173264 13310
rect 173298 13308 173310 13310
rect 174170 13308 174176 13320
rect 173298 13280 174176 13308
rect 173298 13276 173310 13280
rect 173252 13270 173310 13276
rect 174170 13268 174176 13280
rect 174228 13268 174234 13320
rect 174464 13240 174492 13348
rect 175644 13310 175702 13316
rect 175644 13308 175656 13310
rect 170140 13212 174492 13240
rect 174556 13280 175656 13308
rect 165246 13172 165252 13184
rect 164660 13144 165108 13172
rect 165206 13144 165252 13172
rect 164660 13132 164666 13144
rect 165246 13132 165252 13144
rect 165304 13132 165310 13184
rect 165338 13132 165344 13184
rect 165396 13172 165402 13184
rect 166076 13174 166134 13180
rect 166076 13172 166088 13174
rect 165396 13144 166088 13172
rect 165396 13132 165402 13144
rect 166076 13140 166088 13144
rect 166122 13140 166134 13174
rect 166442 13172 166448 13184
rect 166402 13144 166448 13172
rect 166076 13134 166134 13140
rect 166442 13132 166448 13144
rect 166500 13132 166506 13184
rect 167380 13172 167408 13200
rect 174556 13172 174584 13280
rect 175644 13276 175656 13280
rect 175690 13308 175702 13310
rect 175826 13308 175832 13320
rect 175690 13280 175832 13308
rect 175690 13276 175702 13280
rect 175644 13270 175702 13276
rect 175826 13268 175832 13280
rect 175884 13268 175890 13320
rect 175936 13304 175964 13348
rect 176120 13348 178968 13376
rect 176120 13304 176148 13348
rect 178956 13344 178968 13348
rect 179002 13376 179014 13378
rect 181898 13376 181904 13388
rect 179002 13348 181904 13376
rect 179002 13344 179014 13348
rect 178956 13338 179014 13344
rect 181898 13336 181904 13348
rect 181956 13336 181962 13388
rect 182082 13336 182088 13388
rect 182140 13376 182146 13388
rect 182560 13376 182588 13484
rect 182726 13472 182732 13484
rect 182784 13472 182790 13524
rect 185762 13512 185768 13524
rect 185722 13484 185768 13512
rect 185762 13472 185768 13484
rect 185820 13472 185826 13524
rect 189350 13512 189356 13524
rect 185872 13484 189356 13512
rect 185872 13376 185900 13484
rect 189350 13472 189356 13484
rect 189408 13472 189414 13524
rect 189460 13484 190868 13512
rect 188798 13404 188804 13456
rect 188856 13444 188862 13456
rect 189460 13444 189488 13484
rect 188856 13416 189488 13444
rect 188856 13404 188862 13416
rect 189534 13404 189540 13456
rect 189592 13444 189598 13456
rect 190840 13444 190868 13484
rect 190914 13472 190920 13524
rect 190972 13512 190978 13524
rect 193490 13512 193496 13524
rect 190972 13484 193496 13512
rect 190972 13472 190978 13484
rect 193490 13472 193496 13484
rect 193548 13472 193554 13524
rect 207106 13512 207112 13524
rect 197372 13484 207112 13512
rect 191834 13444 191840 13456
rect 189592 13416 189672 13444
rect 190840 13416 191840 13444
rect 189592 13404 189598 13416
rect 188522 13376 188528 13388
rect 182140 13348 182184 13376
rect 182560 13348 185900 13376
rect 185964 13348 187464 13376
rect 188482 13348 188528 13376
rect 182140 13336 182146 13348
rect 176378 13308 176384 13320
rect 175936 13276 176148 13304
rect 176338 13280 176384 13308
rect 176378 13268 176384 13280
rect 176436 13268 176442 13320
rect 180610 13268 180616 13320
rect 180668 13308 180674 13320
rect 185964 13316 185992 13348
rect 181992 13310 182050 13316
rect 181992 13308 182004 13310
rect 180668 13280 182004 13308
rect 180668 13268 180674 13280
rect 181992 13276 182004 13280
rect 182038 13308 182050 13310
rect 182912 13310 182970 13316
rect 182912 13308 182924 13310
rect 182038 13280 182924 13308
rect 182038 13276 182050 13280
rect 181992 13270 182050 13276
rect 182912 13276 182924 13280
rect 182958 13276 182970 13310
rect 182912 13270 182970 13276
rect 185948 13310 186006 13316
rect 185948 13276 185960 13310
rect 185994 13276 186006 13310
rect 185948 13270 186006 13276
rect 187328 13310 187386 13316
rect 187328 13276 187340 13310
rect 187374 13276 187386 13310
rect 187436 13308 187464 13348
rect 188522 13336 188528 13348
rect 188580 13336 188586 13388
rect 189644 13376 189672 13416
rect 191834 13404 191840 13416
rect 191892 13404 191898 13456
rect 197372 13444 197400 13484
rect 207106 13472 207112 13484
rect 207164 13472 207170 13524
rect 210326 13512 210332 13524
rect 207216 13484 207980 13512
rect 210286 13484 210332 13512
rect 195716 13416 197400 13444
rect 199840 13446 199898 13452
rect 189812 13378 189870 13384
rect 189812 13376 189824 13378
rect 189644 13348 189824 13376
rect 189812 13344 189824 13348
rect 189858 13344 189870 13378
rect 189812 13338 189870 13344
rect 189902 13336 189908 13388
rect 189960 13376 189966 13388
rect 195716 13376 195744 13416
rect 199840 13412 199852 13446
rect 199886 13444 199898 13446
rect 201954 13444 201960 13456
rect 199886 13416 201960 13444
rect 199886 13412 199898 13416
rect 199840 13406 199898 13412
rect 201954 13404 201960 13416
rect 202012 13404 202018 13456
rect 203426 13404 203432 13456
rect 203484 13444 203490 13456
rect 203888 13446 203946 13452
rect 203888 13444 203900 13446
rect 203484 13416 203900 13444
rect 203484 13404 203490 13416
rect 203888 13412 203900 13416
rect 203934 13412 203946 13446
rect 203888 13406 203946 13412
rect 206002 13404 206008 13456
rect 206060 13444 206066 13456
rect 207216 13444 207244 13484
rect 206060 13416 207244 13444
rect 206060 13404 206066 13416
rect 207750 13404 207756 13456
rect 207808 13444 207814 13456
rect 207808 13416 207888 13444
rect 207808 13404 207814 13416
rect 189960 13348 195744 13376
rect 189960 13336 189966 13348
rect 197630 13336 197636 13388
rect 197688 13376 197694 13388
rect 198736 13378 198794 13384
rect 198736 13376 198748 13378
rect 197688 13348 198748 13376
rect 197688 13336 197694 13348
rect 198736 13344 198748 13348
rect 198782 13344 198794 13378
rect 198736 13338 198794 13344
rect 201128 13378 201186 13384
rect 201128 13344 201140 13378
rect 201174 13376 201186 13378
rect 202046 13376 202052 13388
rect 201174 13348 202052 13376
rect 201174 13344 201186 13348
rect 201128 13338 201186 13344
rect 202046 13336 202052 13348
rect 202104 13336 202110 13388
rect 207860 13384 207888 13416
rect 204716 13378 204774 13384
rect 204716 13376 204728 13378
rect 202156 13348 204728 13376
rect 202156 13320 202184 13348
rect 204716 13344 204728 13348
rect 204762 13376 204774 13378
rect 207844 13378 207902 13384
rect 204762 13348 207796 13376
rect 204762 13344 204774 13348
rect 204716 13338 204774 13344
rect 188432 13310 188490 13316
rect 188432 13308 188444 13310
rect 187436 13280 188444 13308
rect 187328 13270 187386 13276
rect 188432 13276 188444 13280
rect 188478 13276 188490 13310
rect 189534 13308 189540 13320
rect 189494 13280 189540 13308
rect 188432 13270 188490 13276
rect 175734 13200 175740 13252
rect 175792 13240 175798 13252
rect 176656 13242 176714 13248
rect 176656 13240 176668 13242
rect 175792 13212 176668 13240
rect 175792 13200 175798 13212
rect 176656 13208 176668 13212
rect 176702 13208 176714 13242
rect 176656 13202 176714 13208
rect 177666 13200 177672 13252
rect 177724 13200 177730 13252
rect 179232 13242 179290 13248
rect 179232 13240 179244 13242
rect 177960 13212 179244 13240
rect 167380 13144 174584 13172
rect 174998 13132 175004 13184
rect 175056 13172 175062 13184
rect 177960 13172 177988 13212
rect 179232 13208 179244 13212
rect 179278 13208 179290 13242
rect 179232 13202 179290 13208
rect 179966 13200 179972 13252
rect 180024 13200 180030 13252
rect 180886 13200 180892 13252
rect 180944 13240 180950 13252
rect 181900 13242 181958 13248
rect 181900 13240 181912 13242
rect 180944 13212 181912 13240
rect 180944 13200 180950 13212
rect 181900 13208 181912 13212
rect 181946 13240 181958 13242
rect 185964 13240 185992 13270
rect 181946 13212 185992 13240
rect 181946 13208 181958 13212
rect 181900 13202 181958 13208
rect 180702 13172 180708 13184
rect 175056 13144 177988 13172
rect 180662 13144 180708 13172
rect 175056 13132 175062 13144
rect 180702 13132 180708 13144
rect 180760 13132 180766 13184
rect 187344 13172 187372 13270
rect 189534 13268 189540 13280
rect 189592 13268 189598 13320
rect 191836 13310 191894 13316
rect 191836 13276 191848 13310
rect 191882 13276 191894 13310
rect 191836 13270 191894 13276
rect 194412 13310 194470 13316
rect 194412 13276 194424 13310
rect 194458 13276 194470 13310
rect 194412 13270 194470 13276
rect 200024 13310 200082 13316
rect 200024 13276 200036 13310
rect 200070 13308 200082 13310
rect 201494 13308 201500 13320
rect 200070 13280 201500 13308
rect 200070 13276 200082 13280
rect 200024 13270 200082 13276
rect 187420 13242 187478 13248
rect 187420 13208 187432 13242
rect 187466 13240 187478 13242
rect 191852 13240 191880 13270
rect 187466 13212 190302 13240
rect 191208 13212 191880 13240
rect 187466 13208 187478 13212
rect 187420 13202 187478 13208
rect 187786 13172 187792 13184
rect 187344 13144 187792 13172
rect 187786 13132 187792 13144
rect 187844 13132 187850 13184
rect 187970 13172 187976 13184
rect 187930 13144 187976 13172
rect 187970 13132 187976 13144
rect 188028 13132 188034 13184
rect 188338 13172 188344 13184
rect 188298 13144 188344 13172
rect 188338 13132 188344 13144
rect 188396 13132 188402 13184
rect 189534 13132 189540 13184
rect 189592 13172 189598 13184
rect 191208 13172 191236 13212
rect 189592 13144 191236 13172
rect 191284 13174 191342 13180
rect 189592 13132 189598 13144
rect 191284 13140 191296 13174
rect 191330 13172 191342 13174
rect 191374 13172 191380 13184
rect 191330 13144 191380 13172
rect 191330 13140 191342 13144
rect 191284 13134 191342 13140
rect 191374 13132 191380 13144
rect 191432 13132 191438 13184
rect 191852 13172 191880 13212
rect 192112 13242 192170 13248
rect 192112 13208 192124 13242
rect 192158 13240 192170 13242
rect 192386 13240 192392 13252
rect 192158 13212 192392 13240
rect 192158 13208 192170 13212
rect 192112 13202 192170 13208
rect 192386 13200 192392 13212
rect 192444 13200 192450 13252
rect 193398 13240 193404 13252
rect 193338 13212 193404 13240
rect 193398 13200 193404 13212
rect 193456 13200 193462 13252
rect 193860 13242 193918 13248
rect 193860 13208 193872 13242
rect 193906 13240 193918 13242
rect 193950 13240 193956 13252
rect 193906 13212 193956 13240
rect 193906 13208 193918 13212
rect 193860 13202 193918 13208
rect 193950 13200 193956 13212
rect 194008 13200 194014 13252
rect 194428 13172 194456 13270
rect 201494 13268 201500 13280
rect 201552 13268 201558 13320
rect 202138 13308 202144 13320
rect 202098 13280 202144 13308
rect 202138 13268 202144 13280
rect 202196 13268 202202 13320
rect 207198 13308 207204 13320
rect 206296 13280 207204 13308
rect 194594 13200 194600 13252
rect 194652 13240 194658 13252
rect 194688 13242 194746 13248
rect 194688 13240 194700 13242
rect 194652 13212 194700 13240
rect 194652 13200 194658 13212
rect 194688 13208 194700 13212
rect 194734 13208 194746 13242
rect 194688 13202 194746 13208
rect 194778 13200 194784 13252
rect 194836 13240 194842 13252
rect 196434 13240 196440 13252
rect 194836 13212 195178 13240
rect 196346 13212 196440 13240
rect 194836 13200 194842 13212
rect 196434 13200 196440 13212
rect 196492 13240 196498 13252
rect 197354 13240 197360 13252
rect 196492 13212 197360 13240
rect 196492 13200 196498 13212
rect 197354 13200 197360 13212
rect 197412 13200 197418 13252
rect 197816 13242 197874 13248
rect 197816 13208 197828 13242
rect 197862 13240 197874 13242
rect 198644 13242 198702 13248
rect 197862 13212 198596 13240
rect 197862 13208 197874 13212
rect 197816 13202 197874 13208
rect 198568 13184 198596 13212
rect 198644 13208 198656 13242
rect 198690 13240 198702 13242
rect 202414 13240 202420 13252
rect 198690 13212 202184 13240
rect 202374 13212 202420 13240
rect 198690 13208 198702 13212
rect 198644 13202 198702 13208
rect 197722 13172 197728 13184
rect 191852 13144 197728 13172
rect 197722 13132 197728 13144
rect 197780 13132 197786 13184
rect 197906 13132 197912 13184
rect 197964 13172 197970 13184
rect 198184 13174 198242 13180
rect 198184 13172 198196 13174
rect 197964 13144 198196 13172
rect 197964 13132 197970 13144
rect 198184 13140 198196 13144
rect 198230 13140 198242 13174
rect 198550 13172 198556 13184
rect 198510 13144 198556 13172
rect 198184 13134 198242 13140
rect 198550 13132 198556 13144
rect 198608 13132 198614 13184
rect 200482 13172 200488 13184
rect 200442 13144 200488 13172
rect 200482 13132 200488 13144
rect 200540 13132 200546 13184
rect 200850 13172 200856 13184
rect 200810 13144 200856 13172
rect 200850 13132 200856 13144
rect 200908 13132 200914 13184
rect 200944 13174 201002 13180
rect 200944 13140 200956 13174
rect 200990 13172 201002 13174
rect 201310 13172 201316 13184
rect 200990 13144 201316 13172
rect 200990 13140 201002 13144
rect 200944 13134 201002 13140
rect 201310 13132 201316 13144
rect 201368 13132 201374 13184
rect 202156 13172 202184 13212
rect 202414 13200 202420 13212
rect 202472 13200 202478 13252
rect 203150 13200 203156 13252
rect 203208 13200 203214 13252
rect 203812 13212 204024 13240
rect 203812 13172 203840 13212
rect 202156 13144 203840 13172
rect 203996 13172 204024 13212
rect 204254 13200 204260 13252
rect 204312 13240 204318 13252
rect 204992 13242 205050 13248
rect 204992 13240 205004 13242
rect 204312 13212 205004 13240
rect 204312 13200 204318 13212
rect 204992 13208 205004 13212
rect 205038 13208 205050 13242
rect 204992 13202 205050 13208
rect 205450 13200 205456 13252
rect 205508 13200 205514 13252
rect 205634 13172 205640 13184
rect 203996 13144 205640 13172
rect 205634 13132 205640 13144
rect 205692 13132 205698 13184
rect 205726 13132 205732 13184
rect 205784 13172 205790 13184
rect 206296 13172 206324 13280
rect 207198 13268 207204 13280
rect 207256 13268 207262 13320
rect 207660 13310 207718 13316
rect 207660 13308 207672 13310
rect 207584 13280 207672 13308
rect 207584 13252 207612 13280
rect 207660 13276 207672 13280
rect 207706 13276 207718 13310
rect 207660 13270 207718 13276
rect 206370 13200 206376 13252
rect 206428 13240 206434 13252
rect 206428 13212 206876 13240
rect 206428 13200 206434 13212
rect 206464 13174 206522 13180
rect 206464 13172 206476 13174
rect 205784 13144 206476 13172
rect 205784 13132 205790 13144
rect 206464 13140 206476 13144
rect 206510 13140 206522 13174
rect 206848 13172 206876 13212
rect 207566 13200 207572 13252
rect 207624 13200 207630 13252
rect 207768 13240 207796 13348
rect 207844 13344 207856 13378
rect 207890 13344 207902 13378
rect 207952 13376 207980 13484
rect 210326 13472 210332 13484
rect 210384 13472 210390 13524
rect 213362 13512 213368 13524
rect 213322 13484 213368 13512
rect 213362 13472 213368 13484
rect 213420 13472 213426 13524
rect 268930 13512 268936 13524
rect 213472 13484 268936 13512
rect 208026 13404 208032 13456
rect 208084 13444 208090 13456
rect 213270 13444 213276 13456
rect 208084 13416 213276 13444
rect 208084 13404 208090 13416
rect 213270 13404 213276 13416
rect 213328 13404 213334 13456
rect 213472 13376 213500 13484
rect 268930 13472 268936 13484
rect 268988 13472 268994 13524
rect 269380 13514 269438 13520
rect 269380 13480 269392 13514
rect 269426 13512 269438 13514
rect 269574 13512 269580 13524
rect 269426 13484 269580 13512
rect 269426 13480 269438 13484
rect 269380 13474 269438 13480
rect 269574 13472 269580 13484
rect 269632 13472 269638 13524
rect 271782 13472 271788 13524
rect 271840 13512 271846 13524
rect 274268 13514 274326 13520
rect 274268 13512 274280 13514
rect 271840 13484 274280 13512
rect 271840 13472 271846 13484
rect 274268 13480 274280 13484
rect 274314 13480 274326 13514
rect 274910 13512 274916 13524
rect 274870 13484 274916 13512
rect 274268 13474 274326 13480
rect 274910 13472 274916 13484
rect 274968 13472 274974 13524
rect 277854 13512 277860 13524
rect 277814 13484 277860 13512
rect 277854 13472 277860 13484
rect 277912 13472 277918 13524
rect 280890 13512 280896 13524
rect 280850 13484 280896 13512
rect 280890 13472 280896 13484
rect 280948 13472 280954 13524
rect 284294 13472 284300 13524
rect 284352 13512 284358 13524
rect 284572 13514 284630 13520
rect 284572 13512 284584 13514
rect 284352 13484 284584 13512
rect 284352 13472 284358 13484
rect 284572 13480 284584 13484
rect 284618 13480 284630 13514
rect 284572 13474 284630 13480
rect 287054 13472 287060 13524
rect 287112 13512 287118 13524
rect 287148 13514 287206 13520
rect 287148 13512 287160 13514
rect 287112 13484 287160 13512
rect 287112 13472 287118 13484
rect 287148 13480 287160 13484
rect 287194 13480 287206 13514
rect 290090 13512 290096 13524
rect 290050 13484 290096 13512
rect 287148 13474 287206 13480
rect 290090 13472 290096 13484
rect 290148 13472 290154 13524
rect 293218 13512 293224 13524
rect 293178 13484 293224 13512
rect 293218 13472 293224 13484
rect 293276 13472 293282 13524
rect 296254 13512 296260 13524
rect 296214 13484 296260 13512
rect 296254 13472 296260 13484
rect 296312 13472 296318 13524
rect 299290 13512 299296 13524
rect 299250 13484 299296 13512
rect 299290 13472 299296 13484
rect 299348 13472 299354 13524
rect 301406 13512 301412 13524
rect 301366 13484 301412 13512
rect 301406 13472 301412 13484
rect 301464 13512 301470 13524
rect 301776 13514 301834 13520
rect 301776 13512 301788 13514
rect 301464 13484 301788 13512
rect 301464 13472 301470 13484
rect 301776 13480 301788 13484
rect 301822 13512 301834 13514
rect 302144 13514 302202 13520
rect 302144 13512 302156 13514
rect 301822 13484 302156 13512
rect 301822 13480 301834 13484
rect 301776 13474 301834 13480
rect 302144 13480 302156 13484
rect 302190 13512 302202 13514
rect 302972 13514 303030 13520
rect 302972 13512 302984 13514
rect 302190 13484 302984 13512
rect 302190 13480 302202 13484
rect 302144 13474 302202 13480
rect 302972 13480 302984 13484
rect 303018 13512 303030 13514
rect 303340 13514 303398 13520
rect 303340 13512 303352 13514
rect 303018 13484 303352 13512
rect 303018 13480 303030 13484
rect 302972 13474 303030 13480
rect 303340 13480 303352 13484
rect 303386 13480 303398 13514
rect 303340 13474 303398 13480
rect 216398 13444 216404 13456
rect 216358 13416 216404 13444
rect 216398 13404 216404 13416
rect 216456 13404 216462 13456
rect 219434 13404 219440 13456
rect 219492 13444 219498 13456
rect 220172 13446 220230 13452
rect 220172 13444 220184 13446
rect 219492 13416 220184 13444
rect 219492 13404 219498 13416
rect 220172 13412 220184 13416
rect 220218 13412 220230 13446
rect 224126 13444 224132 13456
rect 220172 13406 220230 13412
rect 220280 13416 224132 13444
rect 207952 13348 213500 13376
rect 207844 13338 207902 13344
rect 207934 13268 207940 13320
rect 207992 13308 207998 13320
rect 210512 13310 210570 13316
rect 210512 13308 210524 13310
rect 207992 13280 210524 13308
rect 207992 13268 207998 13280
rect 210512 13276 210524 13280
rect 210558 13276 210570 13310
rect 213546 13308 213552 13320
rect 213506 13280 213552 13308
rect 210512 13270 210570 13276
rect 213546 13268 213552 13280
rect 213604 13268 213610 13320
rect 216582 13308 216588 13320
rect 216494 13280 216588 13308
rect 216582 13268 216588 13280
rect 216640 13308 216646 13320
rect 220280 13308 220308 13416
rect 224126 13404 224132 13416
rect 224184 13404 224190 13456
rect 226426 13444 226432 13456
rect 224328 13416 226432 13444
rect 224034 13376 224040 13388
rect 220372 13348 224040 13376
rect 220372 13316 220400 13348
rect 224034 13336 224040 13348
rect 224092 13336 224098 13388
rect 224328 13384 224356 13416
rect 226426 13404 226432 13416
rect 226484 13404 226490 13456
rect 226610 13404 226616 13456
rect 226668 13444 226674 13456
rect 226668 13416 226712 13444
rect 226668 13404 226674 13416
rect 226886 13404 226892 13456
rect 226944 13444 226950 13456
rect 227898 13444 227904 13456
rect 226944 13416 227904 13444
rect 226944 13404 226950 13416
rect 227898 13404 227904 13416
rect 227956 13404 227962 13456
rect 229186 13404 229192 13456
rect 229244 13444 229250 13456
rect 229648 13446 229706 13452
rect 229648 13444 229660 13446
rect 229244 13416 229660 13444
rect 229244 13404 229250 13416
rect 229648 13412 229660 13416
rect 229694 13412 229706 13446
rect 229648 13406 229706 13412
rect 231780 13416 238340 13444
rect 224312 13378 224370 13384
rect 224312 13344 224324 13378
rect 224358 13344 224370 13378
rect 224312 13338 224370 13344
rect 224402 13336 224408 13388
rect 224460 13376 224466 13388
rect 227070 13376 227076 13388
rect 224460 13348 227076 13376
rect 224460 13336 224466 13348
rect 227070 13336 227076 13348
rect 227128 13336 227134 13388
rect 227162 13336 227168 13388
rect 227220 13376 227226 13388
rect 230476 13378 230534 13384
rect 230476 13376 230488 13378
rect 227220 13348 227264 13376
rect 227824 13348 230488 13376
rect 227220 13336 227226 13348
rect 216640 13280 220308 13308
rect 220356 13310 220414 13316
rect 216640 13268 216646 13280
rect 220356 13276 220368 13310
rect 220402 13276 220414 13310
rect 220356 13270 220414 13276
rect 222932 13310 222990 13316
rect 225876 13310 225934 13316
rect 222932 13276 222944 13310
rect 222978 13308 222990 13310
rect 225616 13308 225736 13310
rect 222978 13280 224356 13308
rect 222978 13276 222990 13280
rect 222932 13270 222990 13276
rect 224218 13240 224224 13252
rect 207768 13212 224224 13240
rect 224218 13200 224224 13212
rect 224276 13200 224282 13252
rect 207292 13174 207350 13180
rect 207292 13172 207304 13174
rect 206848 13144 207304 13172
rect 206464 13134 206522 13140
rect 207292 13140 207304 13144
rect 207338 13140 207350 13174
rect 207292 13134 207350 13140
rect 207382 13132 207388 13184
rect 207440 13172 207446 13184
rect 207752 13174 207810 13180
rect 207752 13172 207764 13174
rect 207440 13144 207764 13172
rect 207440 13132 207446 13144
rect 207752 13140 207764 13144
rect 207798 13172 207810 13174
rect 213546 13172 213552 13184
rect 207798 13144 213552 13172
rect 207798 13140 207810 13144
rect 207752 13134 207810 13140
rect 213546 13132 213552 13144
rect 213604 13132 213610 13184
rect 222746 13172 222752 13184
rect 222706 13144 222752 13172
rect 222746 13132 222752 13144
rect 222804 13132 222810 13184
rect 223666 13172 223672 13184
rect 223626 13144 223672 13172
rect 223666 13132 223672 13144
rect 223724 13132 223730 13184
rect 224034 13172 224040 13184
rect 223994 13144 224040 13172
rect 224034 13132 224040 13144
rect 224092 13132 224098 13184
rect 224126 13132 224132 13184
rect 224184 13172 224190 13184
rect 224328 13172 224356 13280
rect 225432 13282 225828 13308
rect 225432 13280 225644 13282
rect 225708 13280 225828 13282
rect 224402 13200 224408 13252
rect 224460 13240 224466 13252
rect 225432 13240 225460 13280
rect 224460 13212 225460 13240
rect 225800 13240 225828 13280
rect 225876 13276 225888 13310
rect 225922 13308 225934 13310
rect 227714 13308 227720 13320
rect 225922 13280 227720 13308
rect 225922 13276 225934 13280
rect 225876 13270 225934 13276
rect 227714 13268 227720 13280
rect 227772 13268 227778 13320
rect 227824 13240 227852 13348
rect 230476 13344 230488 13348
rect 230522 13376 230534 13378
rect 231780 13376 231808 13416
rect 230522 13348 231808 13376
rect 230522 13344 230534 13348
rect 230476 13338 230534 13344
rect 231946 13336 231952 13388
rect 232004 13376 232010 13388
rect 232224 13378 232282 13384
rect 232224 13376 232236 13378
rect 232004 13348 232236 13376
rect 232004 13336 232010 13348
rect 232224 13344 232236 13348
rect 232270 13344 232282 13378
rect 233142 13376 233148 13388
rect 232224 13338 232282 13344
rect 232700 13348 233148 13376
rect 227900 13310 227958 13316
rect 227900 13276 227912 13310
rect 227946 13276 227958 13310
rect 230382 13308 230388 13320
rect 229310 13280 230388 13308
rect 227900 13270 227958 13276
rect 225800 13212 227852 13240
rect 224460 13200 224466 13212
rect 227916 13184 227944 13270
rect 230382 13268 230388 13280
rect 230440 13268 230446 13320
rect 231854 13268 231860 13320
rect 231912 13268 231918 13320
rect 232038 13268 232044 13320
rect 232096 13308 232102 13320
rect 232700 13308 232728 13348
rect 233142 13336 233148 13348
rect 233200 13336 233206 13388
rect 233326 13336 233332 13388
rect 233384 13376 233390 13388
rect 237192 13378 237250 13384
rect 237192 13376 237204 13378
rect 233384 13348 237204 13376
rect 233384 13336 233390 13348
rect 233050 13308 233056 13320
rect 232096 13280 232728 13308
rect 233010 13280 233056 13308
rect 232096 13268 232102 13280
rect 233050 13268 233056 13280
rect 233108 13268 233114 13320
rect 233880 13310 233938 13316
rect 233160 13284 233740 13308
rect 233160 13280 233832 13284
rect 228082 13200 228088 13252
rect 228140 13240 228146 13252
rect 228176 13242 228234 13248
rect 228176 13240 228188 13242
rect 228140 13212 228188 13240
rect 228140 13200 228146 13212
rect 228176 13208 228188 13212
rect 228222 13208 228234 13242
rect 230750 13240 230756 13252
rect 230710 13212 230756 13240
rect 228176 13202 228234 13208
rect 230750 13200 230756 13212
rect 230808 13200 230814 13252
rect 233160 13240 233188 13280
rect 233712 13256 233832 13280
rect 233880 13276 233892 13310
rect 233926 13308 233938 13310
rect 233988 13308 234016 13348
rect 237192 13344 237204 13348
rect 237238 13344 237250 13378
rect 237192 13338 237250 13344
rect 237284 13378 237342 13384
rect 237284 13344 237296 13378
rect 237330 13376 237342 13378
rect 237926 13376 237932 13388
rect 237330 13348 237932 13376
rect 237330 13344 237342 13348
rect 237284 13338 237342 13344
rect 237926 13336 237932 13348
rect 237984 13336 237990 13388
rect 238110 13376 238116 13388
rect 238036 13348 238116 13376
rect 233926 13280 234016 13308
rect 235076 13310 235134 13316
rect 233926 13276 233938 13280
rect 233880 13270 233938 13276
rect 235076 13276 235088 13310
rect 235122 13308 235134 13310
rect 237100 13310 237158 13316
rect 237100 13308 237112 13310
rect 235122 13280 237112 13308
rect 235122 13276 235134 13280
rect 235076 13270 235134 13276
rect 237100 13276 237112 13280
rect 237146 13308 237158 13310
rect 238036 13308 238064 13348
rect 238110 13336 238116 13348
rect 238168 13336 238174 13388
rect 238312 13376 238340 13416
rect 239490 13404 239496 13456
rect 239548 13444 239554 13456
rect 239952 13446 240010 13452
rect 239952 13444 239964 13446
rect 239548 13416 239964 13444
rect 239548 13404 239554 13416
rect 239952 13412 239964 13416
rect 239998 13412 240010 13446
rect 239952 13406 240010 13412
rect 244642 13404 244648 13456
rect 244700 13444 244706 13456
rect 245378 13444 245384 13456
rect 244700 13416 245384 13444
rect 244700 13404 244706 13416
rect 245378 13404 245384 13416
rect 245436 13404 245442 13456
rect 247126 13444 247132 13456
rect 247086 13416 247132 13444
rect 247126 13404 247132 13416
rect 247184 13404 247190 13456
rect 249520 13446 249578 13452
rect 249520 13412 249532 13446
rect 249566 13444 249578 13446
rect 251082 13444 251088 13456
rect 249566 13416 251088 13444
rect 249566 13412 249578 13416
rect 249520 13406 249578 13412
rect 251082 13404 251088 13416
rect 251140 13404 251146 13456
rect 252462 13404 252468 13456
rect 252520 13444 252526 13456
rect 252832 13446 252890 13452
rect 252832 13444 252844 13446
rect 252520 13416 252844 13444
rect 252520 13404 252526 13416
rect 252832 13412 252844 13416
rect 252878 13412 252890 13446
rect 252832 13406 252890 13412
rect 254946 13404 254952 13456
rect 255004 13444 255010 13456
rect 255408 13446 255466 13452
rect 255408 13444 255420 13446
rect 255004 13416 255420 13444
rect 255004 13404 255010 13416
rect 255408 13412 255420 13416
rect 255454 13412 255466 13446
rect 259454 13444 259460 13456
rect 259414 13416 259460 13444
rect 255408 13406 255466 13412
rect 259454 13404 259460 13416
rect 259512 13404 259518 13456
rect 262676 13446 262734 13452
rect 262676 13412 262688 13446
rect 262722 13444 262734 13446
rect 263502 13444 263508 13456
rect 262722 13416 263508 13444
rect 262722 13412 262734 13416
rect 262676 13406 262734 13412
rect 263502 13404 263508 13416
rect 263560 13404 263566 13456
rect 265526 13404 265532 13456
rect 265584 13444 265590 13456
rect 265988 13446 266046 13452
rect 265988 13444 266000 13446
rect 265584 13416 266000 13444
rect 265584 13404 265590 13416
rect 265988 13412 266000 13416
rect 266034 13412 266046 13446
rect 265988 13406 266046 13412
rect 270402 13404 270408 13456
rect 270460 13444 270466 13456
rect 270460 13416 271828 13444
rect 270460 13404 270466 13416
rect 240780 13378 240838 13384
rect 240780 13376 240792 13378
rect 238312 13348 240792 13376
rect 240780 13344 240792 13348
rect 240826 13376 240838 13378
rect 243356 13378 243414 13384
rect 243356 13376 243368 13378
rect 240826 13348 243368 13376
rect 240826 13344 240838 13348
rect 240780 13338 240838 13344
rect 243356 13344 243368 13348
rect 243402 13344 243414 13378
rect 243356 13338 243414 13344
rect 244090 13336 244096 13388
rect 244148 13376 244154 13388
rect 245104 13378 245162 13384
rect 245104 13376 245116 13378
rect 244148 13348 245116 13376
rect 244148 13336 244154 13348
rect 245104 13344 245116 13348
rect 245150 13344 245162 13378
rect 245104 13338 245162 13344
rect 250164 13378 250222 13384
rect 250164 13344 250176 13378
rect 250210 13376 250222 13378
rect 250990 13376 250996 13388
rect 250210 13348 250996 13376
rect 250210 13344 250222 13348
rect 250164 13338 250222 13344
rect 238202 13308 238208 13320
rect 237146 13280 238064 13308
rect 238162 13280 238208 13308
rect 237146 13276 237158 13280
rect 237100 13270 237158 13276
rect 238202 13268 238208 13280
rect 238260 13268 238266 13320
rect 239766 13308 239772 13320
rect 239614 13280 239772 13308
rect 239766 13268 239772 13280
rect 239824 13268 239830 13320
rect 245120 13308 245148 13338
rect 250990 13336 250996 13348
rect 251048 13336 251054 13388
rect 262032 13378 262090 13384
rect 251100 13348 259776 13376
rect 251100 13320 251128 13348
rect 247312 13310 247370 13316
rect 247312 13308 247324 13310
rect 245120 13280 247324 13308
rect 247312 13276 247324 13280
rect 247358 13308 247370 13310
rect 249980 13310 250038 13316
rect 249980 13308 249992 13310
rect 247358 13280 249992 13308
rect 247358 13276 247370 13280
rect 247312 13270 247370 13276
rect 249980 13276 249992 13280
rect 250026 13276 250038 13310
rect 251082 13308 251088 13320
rect 251042 13280 251088 13308
rect 249980 13270 250038 13276
rect 251082 13268 251088 13280
rect 251140 13268 251146 13320
rect 253660 13310 253718 13316
rect 253660 13308 253672 13310
rect 252940 13280 253672 13308
rect 232056 13212 233188 13240
rect 233804 13240 233832 13256
rect 233804 13212 238432 13240
rect 225414 13172 225420 13184
rect 224184 13144 224228 13172
rect 224328 13144 225420 13172
rect 224184 13132 224190 13144
rect 225414 13132 225420 13144
rect 225472 13132 225478 13184
rect 225690 13172 225696 13184
rect 225650 13144 225696 13172
rect 225690 13132 225696 13144
rect 225748 13132 225754 13184
rect 226980 13174 227038 13180
rect 226980 13140 226992 13174
rect 227026 13172 227038 13174
rect 227070 13172 227076 13184
rect 227026 13144 227076 13172
rect 227026 13140 227038 13144
rect 226980 13134 227038 13140
rect 227070 13132 227076 13144
rect 227128 13172 227134 13184
rect 227622 13172 227628 13184
rect 227128 13144 227628 13172
rect 227128 13132 227134 13144
rect 227622 13132 227628 13144
rect 227680 13132 227686 13184
rect 227898 13172 227904 13184
rect 227810 13144 227904 13172
rect 227898 13132 227904 13144
rect 227956 13172 227962 13184
rect 232056 13172 232084 13212
rect 227956 13144 232084 13172
rect 227956 13132 227962 13144
rect 232130 13132 232136 13184
rect 232188 13172 232194 13184
rect 233144 13174 233202 13180
rect 233144 13172 233156 13174
rect 232188 13144 233156 13172
rect 232188 13132 232194 13144
rect 233144 13140 233156 13144
rect 233190 13140 233202 13174
rect 233144 13134 233202 13140
rect 233234 13132 233240 13184
rect 233292 13172 233298 13184
rect 233696 13174 233754 13180
rect 233696 13172 233708 13174
rect 233292 13144 233708 13172
rect 233292 13132 233298 13144
rect 233696 13140 233708 13144
rect 233742 13140 233754 13174
rect 234890 13172 234896 13184
rect 234850 13144 234896 13172
rect 233696 13134 233754 13140
rect 234890 13132 234896 13144
rect 234948 13132 234954 13184
rect 236732 13174 236790 13180
rect 236732 13140 236744 13174
rect 236778 13172 236790 13174
rect 237006 13172 237012 13184
rect 236778 13144 237012 13172
rect 236778 13140 236790 13144
rect 236732 13134 236790 13140
rect 237006 13132 237012 13144
rect 237064 13132 237070 13184
rect 238404 13172 238432 13212
rect 238478 13200 238484 13252
rect 238536 13240 238542 13252
rect 241054 13240 241060 13252
rect 238536 13212 238580 13240
rect 239784 13212 240088 13240
rect 241014 13212 241060 13240
rect 238536 13200 238542 13212
rect 239784 13172 239812 13212
rect 238404 13144 239812 13172
rect 240060 13172 240088 13212
rect 241054 13200 241060 13212
rect 241112 13200 241118 13252
rect 241790 13200 241796 13252
rect 241848 13200 241854 13252
rect 243630 13240 243636 13252
rect 242360 13212 242664 13240
rect 243590 13212 243636 13240
rect 242360 13172 242388 13212
rect 242526 13172 242532 13184
rect 240060 13144 242388 13172
rect 242486 13144 242532 13172
rect 242526 13132 242532 13144
rect 242584 13132 242590 13184
rect 242636 13172 242664 13212
rect 243630 13200 243636 13212
rect 243688 13200 243694 13252
rect 244918 13240 244924 13252
rect 244858 13212 244924 13240
rect 244918 13200 244924 13212
rect 244976 13200 244982 13252
rect 249720 13212 251312 13240
rect 249720 13172 249748 13212
rect 242636 13144 249748 13172
rect 249888 13174 249946 13180
rect 249888 13140 249900 13174
rect 249934 13172 249946 13174
rect 251174 13172 251180 13184
rect 249934 13144 251180 13172
rect 249934 13140 249946 13144
rect 249888 13134 249946 13140
rect 251174 13132 251180 13144
rect 251232 13132 251238 13184
rect 251284 13172 251312 13212
rect 251358 13200 251364 13252
rect 251416 13240 251422 13252
rect 251416 13212 251460 13240
rect 251416 13200 251422 13212
rect 252370 13200 252376 13252
rect 252428 13200 252434 13252
rect 252940 13172 252968 13280
rect 253660 13276 253672 13280
rect 253706 13276 253718 13310
rect 256234 13308 256240 13320
rect 253660 13270 253718 13276
rect 255240 13280 256240 13308
rect 253014 13200 253020 13252
rect 253072 13240 253078 13252
rect 253936 13242 253994 13248
rect 253936 13240 253948 13242
rect 253072 13212 253948 13240
rect 253072 13200 253078 13212
rect 253936 13208 253948 13212
rect 253982 13208 253994 13242
rect 253936 13202 253994 13208
rect 254946 13200 254952 13252
rect 255004 13200 255010 13252
rect 253474 13172 253480 13184
rect 251284 13144 253480 13172
rect 253474 13132 253480 13144
rect 253532 13172 253538 13184
rect 255240 13172 255268 13280
rect 256234 13268 256240 13280
rect 256292 13268 256298 13320
rect 259640 13310 259698 13316
rect 259640 13308 259652 13310
rect 257816 13280 259652 13308
rect 255314 13200 255320 13252
rect 255372 13240 255378 13252
rect 256512 13242 256570 13248
rect 256512 13240 256524 13242
rect 255372 13212 256524 13240
rect 255372 13200 255378 13212
rect 256512 13208 256524 13212
rect 256558 13208 256570 13242
rect 256512 13202 256570 13208
rect 256970 13200 256976 13252
rect 257028 13200 257034 13252
rect 253532 13144 255268 13172
rect 253532 13132 253538 13144
rect 256326 13132 256332 13184
rect 256384 13172 256390 13184
rect 257816 13172 257844 13280
rect 259640 13276 259652 13280
rect 259686 13276 259698 13310
rect 259748 13308 259776 13348
rect 262032 13344 262044 13378
rect 262078 13376 262090 13378
rect 263228 13378 263286 13384
rect 263228 13376 263240 13378
rect 262078 13348 263240 13376
rect 262078 13344 262090 13348
rect 262032 13338 262090 13344
rect 263228 13344 263240 13348
rect 263274 13376 263286 13378
rect 264146 13376 264152 13388
rect 263274 13348 264152 13376
rect 263274 13344 263286 13348
rect 263228 13338 263286 13344
rect 264146 13336 264152 13348
rect 264204 13336 264210 13388
rect 266540 13378 266598 13384
rect 266540 13376 266552 13378
rect 264256 13348 266552 13376
rect 264256 13316 264284 13348
rect 266540 13344 266552 13348
rect 266586 13376 266598 13378
rect 269116 13378 269174 13384
rect 269116 13376 269128 13378
rect 266586 13348 269128 13376
rect 266586 13344 266598 13348
rect 266540 13338 266598 13344
rect 269116 13344 269128 13348
rect 269162 13376 269174 13378
rect 271692 13378 271750 13384
rect 271692 13376 271704 13378
rect 269162 13348 271704 13376
rect 269162 13344 269174 13348
rect 269116 13338 269174 13344
rect 271692 13344 271704 13348
rect 271738 13344 271750 13378
rect 271800 13376 271828 13416
rect 272978 13404 272984 13456
rect 273036 13444 273042 13456
rect 273036 13416 278084 13444
rect 273036 13404 273042 13416
rect 271800 13348 273116 13376
rect 271692 13338 271750 13344
rect 264240 13310 264298 13316
rect 264240 13308 264252 13310
rect 259748 13280 264252 13308
rect 259640 13270 259698 13276
rect 264240 13276 264252 13280
rect 264286 13276 264298 13310
rect 264240 13270 264298 13276
rect 268564 13310 268622 13316
rect 268564 13276 268576 13310
rect 268610 13308 268622 13310
rect 268930 13308 268936 13320
rect 268610 13280 268936 13308
rect 268610 13276 268622 13280
rect 268564 13270 268622 13276
rect 268930 13268 268936 13280
rect 268988 13268 268994 13320
rect 273088 13294 273116 13348
rect 273162 13336 273168 13388
rect 273220 13376 273226 13388
rect 273220 13348 277992 13376
rect 273220 13336 273226 13348
rect 273254 13268 273260 13320
rect 273312 13308 273318 13320
rect 274452 13310 274510 13316
rect 274452 13308 274464 13310
rect 273312 13280 274464 13308
rect 273312 13268 273318 13280
rect 274452 13276 274464 13280
rect 274498 13276 274510 13310
rect 275094 13308 275100 13320
rect 275054 13280 275100 13308
rect 274452 13270 274510 13276
rect 275094 13268 275100 13280
rect 275152 13268 275158 13320
rect 261846 13240 261852 13252
rect 261806 13212 261852 13240
rect 261846 13200 261852 13212
rect 261904 13200 261910 13252
rect 263044 13242 263102 13248
rect 263044 13208 263056 13242
rect 263090 13240 263102 13242
rect 263410 13240 263416 13252
rect 263090 13212 263416 13240
rect 263090 13208 263102 13212
rect 263044 13202 263102 13208
rect 263410 13200 263416 13212
rect 263468 13200 263474 13252
rect 263502 13200 263508 13252
rect 263560 13240 263566 13252
rect 264422 13240 264428 13252
rect 263560 13212 264428 13240
rect 263560 13200 263566 13212
rect 264422 13200 264428 13212
rect 264480 13200 264486 13252
rect 264516 13242 264574 13248
rect 264516 13208 264528 13242
rect 264562 13240 264574 13242
rect 264606 13240 264612 13252
rect 264562 13212 264612 13240
rect 264562 13208 264574 13212
rect 264516 13202 264574 13208
rect 264606 13200 264612 13212
rect 264664 13200 264670 13252
rect 264974 13200 264980 13252
rect 265032 13200 265038 13252
rect 266816 13242 266874 13248
rect 265912 13212 266768 13240
rect 256384 13144 257844 13172
rect 256384 13132 256390 13144
rect 257982 13132 257988 13184
rect 258040 13172 258046 13184
rect 262950 13172 262956 13184
rect 258040 13144 262956 13172
rect 258040 13132 258046 13144
rect 262950 13132 262956 13144
rect 263008 13172 263014 13184
rect 263136 13174 263194 13180
rect 263136 13172 263148 13174
rect 263008 13144 263148 13172
rect 263008 13132 263014 13144
rect 263136 13140 263148 13144
rect 263182 13140 263194 13174
rect 263136 13134 263194 13140
rect 263318 13132 263324 13184
rect 263376 13172 263382 13184
rect 265912 13172 265940 13212
rect 263376 13144 265940 13172
rect 266740 13172 266768 13212
rect 266816 13208 266828 13242
rect 266862 13240 266874 13242
rect 266906 13240 266912 13252
rect 266862 13212 266912 13240
rect 266862 13208 266874 13212
rect 266816 13202 266874 13208
rect 266906 13200 266912 13212
rect 266964 13200 266970 13252
rect 268042 13212 268516 13240
rect 267642 13172 267648 13184
rect 266740 13144 267648 13172
rect 263376 13132 263382 13144
rect 267642 13132 267648 13144
rect 267700 13132 267706 13184
rect 268488 13172 268516 13212
rect 268746 13200 268752 13252
rect 268804 13240 268810 13252
rect 268804 13212 269882 13240
rect 268804 13200 268810 13212
rect 270678 13200 270684 13252
rect 270736 13240 270742 13252
rect 270736 13212 270908 13240
rect 270736 13200 270742 13212
rect 270770 13172 270776 13184
rect 268488 13144 270776 13172
rect 270770 13132 270776 13144
rect 270828 13132 270834 13184
rect 270880 13180 270908 13212
rect 270954 13200 270960 13252
rect 271012 13240 271018 13252
rect 271968 13242 272026 13248
rect 271968 13240 271980 13242
rect 271012 13212 271980 13240
rect 271012 13200 271018 13212
rect 271968 13208 271980 13212
rect 272014 13208 272026 13242
rect 277964 13240 277992 13348
rect 278056 13316 278084 13416
rect 303356 13376 303384 13474
rect 304444 13378 304502 13384
rect 304444 13376 304456 13378
rect 278148 13348 293448 13376
rect 303356 13348 304456 13376
rect 278040 13310 278098 13316
rect 278040 13276 278052 13310
rect 278086 13276 278098 13310
rect 278040 13270 278098 13276
rect 278148 13240 278176 13348
rect 281074 13308 281080 13320
rect 281034 13280 281080 13308
rect 281074 13268 281080 13280
rect 281132 13268 281138 13320
rect 284754 13308 284760 13320
rect 284714 13280 284760 13308
rect 284754 13268 284760 13280
rect 284812 13268 284818 13320
rect 287332 13310 287390 13316
rect 287332 13308 287344 13310
rect 287026 13280 287344 13308
rect 287026 13240 287054 13280
rect 287332 13276 287344 13280
rect 287378 13276 287390 13310
rect 290274 13308 290280 13320
rect 290234 13280 290280 13308
rect 287332 13270 287390 13276
rect 290274 13268 290280 13280
rect 290332 13268 290338 13320
rect 293420 13316 293448 13348
rect 304444 13344 304456 13348
rect 304490 13376 304502 13378
rect 304904 13378 304962 13384
rect 304904 13376 304916 13378
rect 304490 13348 304916 13376
rect 304490 13344 304502 13348
rect 304444 13338 304502 13344
rect 304904 13344 304916 13348
rect 304950 13376 304962 13378
rect 304994 13376 305000 13388
rect 304950 13348 305000 13376
rect 304950 13344 304962 13348
rect 304904 13338 304962 13344
rect 304994 13336 305000 13348
rect 305052 13376 305058 13388
rect 305364 13378 305422 13384
rect 305364 13376 305376 13378
rect 305052 13348 305376 13376
rect 305052 13336 305058 13348
rect 305364 13344 305376 13348
rect 305410 13344 305422 13378
rect 305364 13338 305422 13344
rect 293404 13310 293462 13316
rect 293404 13276 293416 13310
rect 293450 13276 293462 13310
rect 296440 13310 296498 13316
rect 296440 13308 296452 13310
rect 293404 13270 293462 13276
rect 295904 13280 296452 13308
rect 277964 13212 278176 13240
rect 282886 13212 287054 13240
rect 271968 13202 272026 13208
rect 270864 13174 270922 13180
rect 270864 13140 270876 13174
rect 270910 13172 270922 13174
rect 271782 13172 271788 13184
rect 270910 13144 271788 13172
rect 270910 13140 270922 13144
rect 270864 13134 270922 13140
rect 271782 13132 271788 13144
rect 271840 13132 271846 13184
rect 272886 13132 272892 13184
rect 272944 13172 272950 13184
rect 273440 13174 273498 13180
rect 273440 13172 273452 13174
rect 272944 13144 273452 13172
rect 272944 13132 272950 13144
rect 273440 13140 273452 13144
rect 273486 13172 273498 13174
rect 282886 13172 282914 13212
rect 295904 13184 295932 13280
rect 296440 13276 296452 13280
rect 296486 13276 296498 13310
rect 299474 13308 299480 13320
rect 299434 13280 299480 13308
rect 296440 13270 296498 13276
rect 299474 13268 299480 13280
rect 299532 13268 299538 13320
rect 303522 13268 303528 13320
rect 303580 13308 303586 13320
rect 303708 13310 303766 13316
rect 303708 13308 303720 13310
rect 303580 13280 303720 13308
rect 303580 13268 303586 13280
rect 303708 13276 303720 13280
rect 303754 13276 303766 13310
rect 303708 13270 303766 13276
rect 295886 13172 295892 13184
rect 273486 13144 282914 13172
rect 295846 13144 295892 13172
rect 273486 13140 273498 13144
rect 273440 13134 273498 13140
rect 295886 13132 295892 13144
rect 295944 13132 295950 13184
rect 1104 13082 305808 13104
rect 1104 13030 77148 13082
rect 77200 13030 77212 13082
rect 77264 13030 77276 13082
rect 77328 13030 77340 13082
rect 77392 13030 77404 13082
rect 77456 13030 153346 13082
rect 153398 13030 153410 13082
rect 153462 13030 153474 13082
rect 153526 13030 153538 13082
rect 153590 13030 153602 13082
rect 153654 13030 229544 13082
rect 229596 13030 229608 13082
rect 229660 13030 229672 13082
rect 229724 13030 229736 13082
rect 229788 13030 229800 13082
rect 229852 13030 305808 13082
rect 1104 13008 305808 13030
rect 26050 12968 26056 12980
rect 26010 12940 26056 12968
rect 26050 12928 26056 12940
rect 26108 12928 26114 12980
rect 27432 12970 27490 12976
rect 27432 12936 27444 12970
rect 27478 12936 27490 12970
rect 32214 12968 32220 12980
rect 27432 12930 27490 12936
rect 27632 12940 32220 12968
rect 20162 12860 20168 12912
rect 20220 12900 20226 12912
rect 20220 12872 22094 12900
rect 20220 12860 20226 12872
rect 22066 12628 22094 12872
rect 27338 12860 27344 12912
rect 27396 12900 27402 12912
rect 27448 12900 27476 12930
rect 27396 12872 27476 12900
rect 27396 12860 27402 12872
rect 26236 12834 26294 12840
rect 26236 12800 26248 12834
rect 26282 12832 26294 12834
rect 27632 12832 27660 12940
rect 32214 12928 32220 12940
rect 32272 12968 32278 12980
rect 33872 12970 33930 12976
rect 33872 12968 33884 12970
rect 32272 12940 33884 12968
rect 32272 12928 32278 12940
rect 33872 12936 33884 12940
rect 33918 12936 33930 12970
rect 33872 12930 33930 12936
rect 34146 12928 34152 12980
rect 34204 12968 34210 12980
rect 34792 12970 34850 12976
rect 34792 12968 34804 12970
rect 34204 12940 34804 12968
rect 34204 12928 34210 12940
rect 34792 12936 34804 12940
rect 34838 12936 34850 12970
rect 35526 12968 35532 12980
rect 35486 12940 35532 12968
rect 34792 12930 34850 12936
rect 35526 12928 35532 12940
rect 35584 12928 35590 12980
rect 36632 12970 36690 12976
rect 36632 12968 36644 12970
rect 35636 12940 36644 12968
rect 28994 12900 29000 12912
rect 26282 12804 27660 12832
rect 27724 12872 29000 12900
rect 26282 12800 26294 12804
rect 26236 12794 26294 12800
rect 23198 12724 23204 12776
rect 23256 12764 23262 12776
rect 27724 12764 27752 12872
rect 28994 12860 29000 12872
rect 29052 12860 29058 12912
rect 30374 12900 30380 12912
rect 29104 12872 30380 12900
rect 27800 12834 27858 12840
rect 27800 12800 27812 12834
rect 27846 12832 27858 12834
rect 27982 12832 27988 12844
rect 27846 12804 27988 12832
rect 27846 12800 27858 12804
rect 27800 12794 27858 12800
rect 27982 12792 27988 12804
rect 28040 12792 28046 12844
rect 23256 12736 27752 12764
rect 27892 12766 27950 12772
rect 23256 12724 23262 12736
rect 27892 12732 27904 12766
rect 27938 12732 27950 12766
rect 28074 12764 28080 12776
rect 28034 12736 28080 12764
rect 27892 12726 27950 12732
rect 27154 12656 27160 12708
rect 27212 12696 27218 12708
rect 27908 12696 27936 12726
rect 28074 12724 28080 12736
rect 28132 12724 28138 12776
rect 29104 12772 29132 12872
rect 30374 12860 30380 12872
rect 30432 12860 30438 12912
rect 31570 12900 31576 12912
rect 31326 12872 31576 12900
rect 31570 12860 31576 12872
rect 31628 12860 31634 12912
rect 34422 12900 34428 12912
rect 33626 12872 34428 12900
rect 34422 12860 34428 12872
rect 34480 12860 34486 12912
rect 35636 12900 35664 12940
rect 36632 12936 36644 12940
rect 36678 12936 36690 12970
rect 42520 12970 42578 12976
rect 36632 12930 36690 12936
rect 37384 12940 41414 12968
rect 37384 12908 37412 12940
rect 34532 12872 35664 12900
rect 36540 12902 36598 12908
rect 33686 12792 33692 12844
rect 33744 12832 33750 12844
rect 34532 12832 34560 12872
rect 36540 12868 36552 12902
rect 36586 12900 36598 12902
rect 37368 12902 37426 12908
rect 37368 12900 37380 12902
rect 36586 12872 37380 12900
rect 36586 12868 36598 12872
rect 36540 12862 36598 12868
rect 37368 12868 37380 12872
rect 37414 12868 37426 12902
rect 37368 12862 37426 12868
rect 37458 12860 37464 12912
rect 37516 12900 37522 12912
rect 38472 12902 38530 12908
rect 38472 12900 38484 12902
rect 37516 12872 38484 12900
rect 37516 12860 37522 12872
rect 38472 12868 38484 12872
rect 38518 12868 38530 12902
rect 38472 12862 38530 12868
rect 39666 12860 39672 12912
rect 39724 12900 39730 12912
rect 39760 12902 39818 12908
rect 39760 12900 39772 12902
rect 39724 12872 39772 12900
rect 39724 12860 39730 12872
rect 39760 12868 39772 12872
rect 39806 12868 39818 12902
rect 41046 12900 41052 12912
rect 40986 12872 41052 12900
rect 39760 12862 39818 12868
rect 41046 12860 41052 12872
rect 41104 12860 41110 12912
rect 41386 12900 41414 12940
rect 42520 12936 42532 12970
rect 42566 12968 42578 12970
rect 43254 12968 43260 12980
rect 42566 12940 43260 12968
rect 42566 12936 42578 12940
rect 42520 12930 42578 12936
rect 43254 12928 43260 12940
rect 43312 12928 43318 12980
rect 43440 12970 43498 12976
rect 43440 12936 43452 12970
rect 43486 12968 43498 12970
rect 44266 12968 44272 12980
rect 43486 12940 44272 12968
rect 43486 12936 43498 12940
rect 43440 12930 43498 12936
rect 44266 12928 44272 12940
rect 44324 12928 44330 12980
rect 44542 12968 44548 12980
rect 44502 12940 44548 12968
rect 44542 12928 44548 12940
rect 44600 12928 44606 12980
rect 51996 12970 52054 12976
rect 51996 12936 52008 12970
rect 52042 12968 52054 12970
rect 53282 12968 53288 12980
rect 52042 12940 53288 12968
rect 52042 12936 52054 12940
rect 51996 12930 52054 12936
rect 53282 12928 53288 12940
rect 53340 12928 53346 12980
rect 53560 12970 53618 12976
rect 53560 12936 53572 12970
rect 53606 12936 53618 12970
rect 53560 12930 53618 12936
rect 53928 12970 53986 12976
rect 53928 12936 53940 12970
rect 53974 12968 53986 12970
rect 54662 12968 54668 12980
rect 53974 12940 54668 12968
rect 53974 12936 53986 12940
rect 53928 12930 53986 12936
rect 42978 12900 42984 12912
rect 41386 12872 42984 12900
rect 42978 12860 42984 12872
rect 43036 12860 43042 12912
rect 53576 12900 53604 12930
rect 54662 12928 54668 12940
rect 54720 12928 54726 12980
rect 55858 12928 55864 12980
rect 55916 12968 55922 12980
rect 57974 12968 57980 12980
rect 55916 12940 57980 12968
rect 55916 12928 55922 12940
rect 57974 12928 57980 12940
rect 58032 12928 58038 12980
rect 58528 12970 58586 12976
rect 58528 12936 58540 12970
rect 58574 12968 58586 12970
rect 59630 12968 59636 12980
rect 58574 12940 59636 12968
rect 58574 12936 58586 12940
rect 58528 12930 58586 12936
rect 59630 12928 59636 12940
rect 59688 12928 59694 12980
rect 72142 12968 72148 12980
rect 72102 12940 72148 12968
rect 72142 12928 72148 12940
rect 72200 12928 72206 12980
rect 72326 12928 72332 12980
rect 72384 12968 72390 12980
rect 74718 12968 74724 12980
rect 72384 12940 74724 12968
rect 72384 12928 72390 12940
rect 74718 12928 74724 12940
rect 74776 12928 74782 12980
rect 83918 12968 83924 12980
rect 75564 12940 83924 12968
rect 52196 12872 53604 12900
rect 33744 12804 34560 12832
rect 34700 12834 34758 12840
rect 33744 12792 33750 12804
rect 34700 12800 34712 12834
rect 34746 12800 34758 12834
rect 34700 12794 34758 12800
rect 35712 12834 35770 12840
rect 35712 12800 35724 12834
rect 35758 12832 35770 12834
rect 38380 12834 38438 12840
rect 38380 12832 38392 12834
rect 35758 12804 38392 12832
rect 35758 12800 35770 12804
rect 35712 12794 35770 12800
rect 38380 12800 38392 12804
rect 38426 12832 38438 12834
rect 39298 12832 39304 12844
rect 38426 12804 39304 12832
rect 38426 12800 38438 12804
rect 38380 12794 38438 12800
rect 29088 12766 29146 12772
rect 29088 12764 29100 12766
rect 28276 12736 29100 12764
rect 27212 12668 27936 12696
rect 27212 12656 27218 12668
rect 28276 12628 28304 12736
rect 29088 12732 29100 12736
rect 29134 12732 29146 12766
rect 29088 12726 29146 12732
rect 29272 12766 29330 12772
rect 29272 12732 29284 12766
rect 29318 12764 29330 12766
rect 29638 12764 29644 12776
rect 29318 12736 29644 12764
rect 29318 12732 29330 12736
rect 29272 12726 29330 12732
rect 29638 12724 29644 12736
rect 29696 12724 29702 12776
rect 29822 12764 29828 12776
rect 29734 12736 29828 12764
rect 29822 12724 29828 12736
rect 29880 12724 29886 12776
rect 30098 12764 30104 12776
rect 30058 12736 30104 12764
rect 30098 12724 30104 12736
rect 30156 12724 30162 12776
rect 32124 12766 32182 12772
rect 32124 12732 32136 12766
rect 32170 12732 32182 12766
rect 32124 12726 32182 12732
rect 32400 12766 32458 12772
rect 32400 12732 32412 12766
rect 32446 12764 32458 12766
rect 33042 12764 33048 12776
rect 32446 12736 33048 12764
rect 32446 12732 32458 12736
rect 32400 12726 32458 12732
rect 22066 12600 28304 12628
rect 28628 12630 28686 12636
rect 28628 12596 28640 12630
rect 28674 12628 28686 12630
rect 28902 12628 28908 12640
rect 28674 12600 28908 12628
rect 28674 12596 28686 12600
rect 28628 12590 28686 12596
rect 28902 12588 28908 12600
rect 28960 12588 28966 12640
rect 29840 12628 29868 12724
rect 32140 12696 32168 12726
rect 33042 12724 33048 12736
rect 33100 12724 33106 12776
rect 33410 12724 33416 12776
rect 33468 12764 33474 12776
rect 34330 12764 34336 12776
rect 33468 12736 34336 12764
rect 33468 12724 33474 12736
rect 34330 12724 34336 12736
rect 34388 12764 34394 12776
rect 34716 12764 34744 12794
rect 39298 12792 39304 12804
rect 39356 12792 39362 12844
rect 41506 12792 41512 12844
rect 41564 12832 41570 12844
rect 41692 12834 41750 12840
rect 41692 12832 41704 12834
rect 41564 12804 41704 12832
rect 41564 12792 41570 12804
rect 41692 12800 41704 12804
rect 41738 12832 41750 12834
rect 42428 12834 42486 12840
rect 42428 12832 42440 12834
rect 41738 12804 42440 12832
rect 41738 12800 41750 12804
rect 41692 12794 41750 12800
rect 42428 12800 42440 12804
rect 42474 12800 42486 12834
rect 44728 12834 44786 12840
rect 44728 12832 44740 12834
rect 42428 12794 42486 12800
rect 43548 12804 44740 12832
rect 34388 12736 34744 12764
rect 34388 12724 34394 12736
rect 34882 12724 34888 12776
rect 34940 12764 34946 12776
rect 34940 12736 34984 12764
rect 34940 12724 34946 12736
rect 35342 12724 35348 12776
rect 35400 12764 35406 12776
rect 37552 12766 37610 12772
rect 37552 12764 37564 12766
rect 35400 12736 37564 12764
rect 35400 12724 35406 12736
rect 37552 12732 37564 12736
rect 37598 12732 37610 12766
rect 37552 12726 37610 12732
rect 38564 12766 38622 12772
rect 38564 12732 38576 12766
rect 38610 12764 38622 12766
rect 39390 12764 39396 12776
rect 38610 12736 39396 12764
rect 38610 12732 38622 12736
rect 38564 12726 38622 12732
rect 39390 12724 39396 12736
rect 39448 12724 39454 12776
rect 39484 12766 39542 12772
rect 39484 12732 39496 12766
rect 39530 12732 39542 12766
rect 39484 12726 39542 12732
rect 39500 12696 39528 12726
rect 40954 12724 40960 12776
rect 41012 12764 41018 12776
rect 43070 12764 43076 12776
rect 41012 12736 43076 12764
rect 41012 12724 41018 12736
rect 43070 12724 43076 12736
rect 43128 12724 43134 12776
rect 43162 12724 43168 12776
rect 43220 12764 43226 12776
rect 43548 12772 43576 12804
rect 44728 12800 44740 12804
rect 44774 12832 44786 12834
rect 45370 12832 45376 12844
rect 44774 12804 45376 12832
rect 44774 12800 44786 12804
rect 44728 12794 44786 12800
rect 45370 12792 45376 12804
rect 45428 12792 45434 12844
rect 52196 12840 52224 12872
rect 55490 12860 55496 12912
rect 55548 12860 55554 12912
rect 57330 12860 57336 12912
rect 57388 12900 57394 12912
rect 58620 12902 58678 12908
rect 58620 12900 58632 12902
rect 57388 12872 58632 12900
rect 57388 12860 57394 12872
rect 58620 12868 58632 12872
rect 58666 12900 58678 12902
rect 60642 12900 60648 12912
rect 58666 12872 60648 12900
rect 58666 12868 58678 12872
rect 58620 12862 58678 12868
rect 60642 12860 60648 12872
rect 60700 12860 60706 12912
rect 65886 12860 65892 12912
rect 65944 12900 65950 12912
rect 75564 12900 75592 12940
rect 77848 12902 77906 12908
rect 77848 12900 77860 12902
rect 65944 12872 75592 12900
rect 77050 12872 77860 12900
rect 65944 12860 65950 12872
rect 52180 12834 52238 12840
rect 52180 12800 52192 12834
rect 52226 12800 52238 12834
rect 52180 12794 52238 12800
rect 52916 12834 52974 12840
rect 52916 12800 52928 12834
rect 52962 12832 52974 12834
rect 53742 12832 53748 12844
rect 52962 12804 53748 12832
rect 52962 12800 52974 12804
rect 52916 12794 52974 12800
rect 53742 12792 53748 12804
rect 53800 12792 53806 12844
rect 54018 12838 54024 12844
rect 53944 12832 54024 12838
rect 53852 12804 54024 12832
rect 43532 12766 43590 12772
rect 43532 12764 43544 12766
rect 43220 12736 43544 12764
rect 43220 12724 43226 12736
rect 43532 12732 43544 12736
rect 43578 12732 43590 12766
rect 43532 12726 43590 12732
rect 43716 12766 43774 12772
rect 43716 12732 43728 12766
rect 43762 12764 43774 12766
rect 43806 12764 43812 12776
rect 43762 12736 43812 12764
rect 43762 12732 43774 12736
rect 43716 12726 43774 12732
rect 43806 12724 43812 12736
rect 43864 12764 43870 12776
rect 45462 12764 45468 12776
rect 43864 12736 45468 12764
rect 43864 12724 43870 12736
rect 45462 12724 45468 12736
rect 45520 12724 45526 12776
rect 51350 12724 51356 12776
rect 51408 12764 51414 12776
rect 53852 12764 53880 12804
rect 54018 12792 54024 12804
rect 54076 12792 54082 12844
rect 54754 12836 54760 12844
rect 54680 12832 54760 12836
rect 54666 12804 54760 12832
rect 54110 12764 54116 12776
rect 51408 12736 53880 12764
rect 54070 12736 54116 12764
rect 51408 12724 51414 12736
rect 54110 12724 54116 12736
rect 54168 12724 54174 12776
rect 54680 12696 54708 12804
rect 54754 12792 54760 12804
rect 54812 12792 54818 12844
rect 57056 12834 57114 12840
rect 57056 12800 57068 12834
rect 57102 12832 57114 12834
rect 57422 12832 57428 12844
rect 57102 12804 57428 12832
rect 57102 12800 57114 12804
rect 57056 12794 57114 12800
rect 57422 12792 57428 12804
rect 57480 12792 57486 12844
rect 72328 12834 72386 12840
rect 72328 12800 72340 12834
rect 72374 12832 72386 12834
rect 74810 12832 74816 12844
rect 72374 12804 74816 12832
rect 72374 12800 72386 12804
rect 72328 12794 72386 12800
rect 74810 12792 74816 12804
rect 74868 12792 74874 12844
rect 75088 12834 75146 12840
rect 75088 12800 75100 12834
rect 75134 12832 75146 12834
rect 75454 12832 75460 12844
rect 75134 12804 75460 12832
rect 75134 12800 75146 12804
rect 75088 12794 75146 12800
rect 75454 12792 75460 12804
rect 75512 12792 75518 12844
rect 75564 12840 75592 12872
rect 77848 12868 77860 12872
rect 77894 12868 77906 12902
rect 77848 12862 77906 12868
rect 78398 12860 78404 12912
rect 78456 12900 78462 12912
rect 78584 12902 78642 12908
rect 78584 12900 78596 12902
rect 78456 12872 78596 12900
rect 78456 12860 78462 12872
rect 78584 12868 78596 12872
rect 78630 12868 78642 12902
rect 78584 12862 78642 12868
rect 75548 12834 75606 12840
rect 75548 12800 75560 12834
rect 75594 12800 75606 12834
rect 75548 12794 75606 12800
rect 77756 12834 77814 12840
rect 77756 12800 77768 12834
rect 77802 12832 77814 12834
rect 78492 12834 78550 12840
rect 78492 12832 78504 12834
rect 77802 12804 78504 12832
rect 77802 12800 77814 12804
rect 77756 12794 77814 12800
rect 78492 12800 78504 12804
rect 78538 12832 78550 12834
rect 79320 12834 79378 12840
rect 78538 12804 78628 12832
rect 78538 12800 78550 12804
rect 78492 12794 78550 12800
rect 78600 12776 78628 12804
rect 79320 12800 79332 12834
rect 79366 12832 79378 12834
rect 79686 12832 79692 12844
rect 79366 12804 79692 12832
rect 79366 12800 79378 12804
rect 79320 12794 79378 12800
rect 79686 12792 79692 12804
rect 79744 12792 79750 12844
rect 79796 12840 79824 12940
rect 83918 12928 83924 12940
rect 83976 12928 83982 12980
rect 86494 12968 86500 12980
rect 84672 12940 86500 12968
rect 80514 12860 80520 12912
rect 80572 12860 80578 12912
rect 82906 12860 82912 12912
rect 82964 12900 82970 12912
rect 84672 12900 84700 12940
rect 86494 12928 86500 12940
rect 86552 12928 86558 12980
rect 87138 12968 87144 12980
rect 86880 12940 87144 12968
rect 86880 12900 86908 12940
rect 87138 12928 87144 12940
rect 87196 12928 87202 12980
rect 89532 12970 89590 12976
rect 89532 12936 89544 12970
rect 89578 12968 89590 12970
rect 89578 12940 89714 12968
rect 89578 12936 89590 12940
rect 89532 12930 89590 12936
rect 89686 12900 89714 12940
rect 90450 12928 90456 12980
rect 90508 12968 90514 12980
rect 91096 12970 91154 12976
rect 91096 12968 91108 12970
rect 90508 12940 91108 12968
rect 90508 12928 90514 12940
rect 91096 12936 91108 12940
rect 91142 12936 91154 12970
rect 91096 12930 91154 12936
rect 91646 12928 91652 12980
rect 91704 12968 91710 12980
rect 97994 12968 98000 12980
rect 91704 12940 98000 12968
rect 91704 12928 91710 12940
rect 97994 12928 98000 12940
rect 98052 12928 98058 12980
rect 99346 12940 108344 12968
rect 90542 12900 90548 12912
rect 82964 12872 84700 12900
rect 85514 12872 86908 12900
rect 87722 12872 89576 12900
rect 89686 12872 90548 12900
rect 82964 12860 82970 12872
rect 79780 12834 79838 12840
rect 79780 12800 79792 12834
rect 79826 12800 79838 12834
rect 86220 12834 86278 12840
rect 86220 12832 86232 12834
rect 79780 12794 79838 12800
rect 85500 12804 86232 12832
rect 55030 12764 55036 12776
rect 54990 12736 55036 12764
rect 55030 12724 55036 12736
rect 55088 12724 55094 12776
rect 58712 12766 58770 12772
rect 58712 12732 58724 12766
rect 58758 12732 58770 12766
rect 75824 12766 75882 12772
rect 75824 12764 75836 12766
rect 58712 12726 58770 12732
rect 74920 12736 75836 12764
rect 58728 12696 58756 12726
rect 74920 12704 74948 12736
rect 75824 12732 75836 12736
rect 75870 12732 75882 12766
rect 75824 12726 75882 12732
rect 78582 12724 78588 12776
rect 78640 12724 78646 12776
rect 80056 12766 80114 12772
rect 80056 12764 80068 12766
rect 79152 12736 80068 12764
rect 31128 12668 32168 12696
rect 31128 12628 31156 12668
rect 29840 12600 31156 12628
rect 31386 12588 31392 12640
rect 31444 12628 31450 12640
rect 31572 12630 31630 12636
rect 31572 12628 31584 12630
rect 31444 12600 31584 12628
rect 31444 12588 31450 12600
rect 31572 12596 31584 12600
rect 31618 12596 31630 12630
rect 32140 12628 32168 12668
rect 33428 12668 39528 12696
rect 32398 12628 32404 12640
rect 32140 12600 32404 12628
rect 31572 12590 31630 12596
rect 32398 12588 32404 12600
rect 32456 12628 32462 12640
rect 33428 12628 33456 12668
rect 32456 12600 33456 12628
rect 32456 12588 32462 12600
rect 34146 12588 34152 12640
rect 34204 12628 34210 12640
rect 34332 12630 34390 12636
rect 34332 12628 34344 12630
rect 34204 12600 34344 12628
rect 34204 12588 34210 12600
rect 34332 12596 34344 12600
rect 34378 12596 34390 12630
rect 38010 12628 38016 12640
rect 37970 12600 38016 12628
rect 34332 12590 34390 12596
rect 38010 12588 38016 12600
rect 38068 12588 38074 12640
rect 39500 12628 39528 12668
rect 40788 12668 54708 12696
rect 56336 12668 58756 12696
rect 74904 12698 74962 12704
rect 40788 12628 40816 12668
rect 56336 12640 56364 12668
rect 41230 12628 41236 12640
rect 39500 12600 40816 12628
rect 41190 12600 41236 12628
rect 41230 12588 41236 12600
rect 41288 12588 41294 12640
rect 41782 12628 41788 12640
rect 41742 12600 41788 12628
rect 41782 12588 41788 12600
rect 41840 12588 41846 12640
rect 42794 12588 42800 12640
rect 42852 12628 42858 12640
rect 43072 12630 43130 12636
rect 43072 12628 43084 12630
rect 42852 12600 43084 12628
rect 42852 12588 42858 12600
rect 43072 12596 43084 12600
rect 43118 12596 43130 12630
rect 43072 12590 43130 12596
rect 43254 12588 43260 12640
rect 43312 12628 43318 12640
rect 43806 12628 43812 12640
rect 43312 12600 43812 12628
rect 43312 12588 43318 12600
rect 43806 12588 43812 12600
rect 43864 12588 43870 12640
rect 53008 12630 53066 12636
rect 53008 12596 53020 12630
rect 53054 12628 53066 12630
rect 53098 12628 53104 12640
rect 53054 12600 53104 12628
rect 53054 12596 53066 12600
rect 53008 12590 53066 12596
rect 53098 12588 53104 12600
rect 53156 12588 53162 12640
rect 54110 12588 54116 12640
rect 54168 12628 54174 12640
rect 55582 12628 55588 12640
rect 54168 12600 55588 12628
rect 54168 12588 54174 12600
rect 55582 12588 55588 12600
rect 55640 12628 55646 12640
rect 56318 12628 56324 12640
rect 55640 12600 56324 12628
rect 55640 12588 55646 12600
rect 56318 12588 56324 12600
rect 56376 12588 56382 12640
rect 56502 12628 56508 12640
rect 56462 12600 56508 12628
rect 56502 12588 56508 12600
rect 56560 12588 56566 12640
rect 57164 12636 57192 12668
rect 74904 12664 74916 12698
rect 74950 12664 74962 12698
rect 77846 12696 77852 12708
rect 74904 12658 74962 12664
rect 76852 12668 77852 12696
rect 57148 12630 57206 12636
rect 57148 12596 57160 12630
rect 57194 12596 57206 12630
rect 57148 12590 57206 12596
rect 57238 12588 57244 12640
rect 57296 12628 57302 12640
rect 58160 12630 58218 12636
rect 58160 12628 58172 12630
rect 57296 12600 58172 12628
rect 57296 12588 57302 12600
rect 58160 12596 58172 12600
rect 58206 12596 58218 12630
rect 58160 12590 58218 12596
rect 72694 12588 72700 12640
rect 72752 12628 72758 12640
rect 74994 12628 75000 12640
rect 72752 12600 75000 12628
rect 72752 12588 72758 12600
rect 74994 12588 75000 12600
rect 75052 12588 75058 12640
rect 75178 12588 75184 12640
rect 75236 12628 75242 12640
rect 76852 12628 76880 12668
rect 77846 12656 77852 12668
rect 77904 12656 77910 12708
rect 78122 12656 78128 12708
rect 78180 12696 78186 12708
rect 79152 12704 79180 12736
rect 80056 12732 80068 12736
rect 80102 12732 80114 12766
rect 80056 12726 80114 12732
rect 80790 12724 80796 12776
rect 80848 12764 80854 12776
rect 84012 12766 84070 12772
rect 84012 12764 84024 12766
rect 80848 12736 84024 12764
rect 80848 12724 80854 12736
rect 84012 12732 84024 12736
rect 84058 12732 84070 12766
rect 84012 12726 84070 12732
rect 84288 12766 84346 12772
rect 84288 12732 84300 12766
rect 84334 12764 84346 12766
rect 84838 12764 84844 12776
rect 84334 12736 84844 12764
rect 84334 12732 84346 12736
rect 84288 12726 84346 12732
rect 79136 12698 79194 12704
rect 78180 12668 78720 12696
rect 78180 12656 78186 12668
rect 75236 12600 76880 12628
rect 75236 12588 75242 12600
rect 77202 12588 77208 12640
rect 77260 12628 77266 12640
rect 77296 12630 77354 12636
rect 77296 12628 77308 12630
rect 77260 12600 77308 12628
rect 77260 12588 77266 12600
rect 77296 12596 77308 12600
rect 77342 12596 77354 12630
rect 78692 12628 78720 12668
rect 79136 12664 79148 12698
rect 79182 12664 79194 12698
rect 79136 12658 79194 12664
rect 81434 12656 81440 12708
rect 81492 12696 81498 12708
rect 81528 12698 81586 12704
rect 81528 12696 81540 12698
rect 81492 12668 81540 12696
rect 81492 12656 81498 12668
rect 81528 12664 81540 12668
rect 81574 12664 81586 12698
rect 81528 12658 81586 12664
rect 81618 12628 81624 12640
rect 78692 12600 81624 12628
rect 77296 12590 77354 12596
rect 81618 12588 81624 12600
rect 81676 12588 81682 12640
rect 84028 12628 84056 12726
rect 84838 12724 84844 12736
rect 84896 12724 84902 12776
rect 85500 12764 85528 12804
rect 85316 12736 85528 12764
rect 85316 12628 85344 12736
rect 85758 12628 85764 12640
rect 84028 12600 85344 12628
rect 85718 12600 85764 12628
rect 85758 12588 85764 12600
rect 85816 12588 85822 12640
rect 86144 12628 86172 12804
rect 86220 12800 86232 12804
rect 86266 12800 86278 12834
rect 89548 12832 89576 12872
rect 90542 12860 90548 12872
rect 90600 12860 90606 12912
rect 90726 12860 90732 12912
rect 90784 12900 90790 12912
rect 99346 12900 99374 12940
rect 99466 12900 99472 12912
rect 90784 12872 99374 12900
rect 99426 12872 99472 12900
rect 90784 12860 90790 12872
rect 99466 12860 99472 12872
rect 99524 12860 99530 12912
rect 99926 12860 99932 12912
rect 99984 12860 99990 12912
rect 104618 12900 104624 12912
rect 104578 12872 104624 12900
rect 104618 12860 104624 12872
rect 104676 12860 104682 12912
rect 104710 12860 104716 12912
rect 104768 12900 104774 12912
rect 104768 12872 106136 12900
rect 104768 12860 104774 12872
rect 90174 12832 90180 12844
rect 89548 12804 90180 12832
rect 86220 12794 86278 12800
rect 90174 12792 90180 12804
rect 90232 12792 90238 12844
rect 90450 12832 90456 12844
rect 90362 12804 90456 12832
rect 90450 12792 90456 12804
rect 90508 12832 90514 12844
rect 90634 12832 90640 12844
rect 90508 12804 90640 12832
rect 90508 12792 90514 12804
rect 90634 12792 90640 12804
rect 90692 12792 90698 12844
rect 91280 12834 91338 12840
rect 91280 12800 91292 12834
rect 91326 12800 91338 12834
rect 91280 12794 91338 12800
rect 98548 12834 98606 12840
rect 98548 12800 98560 12834
rect 98594 12800 98606 12834
rect 105170 12832 105176 12844
rect 102810 12804 105176 12832
rect 98548 12794 98606 12800
rect 86494 12764 86500 12776
rect 86454 12736 86500 12764
rect 86494 12724 86500 12736
rect 86552 12724 86558 12776
rect 88242 12724 88248 12776
rect 88300 12764 88306 12776
rect 89624 12766 89682 12772
rect 89624 12764 89636 12766
rect 88300 12736 89636 12764
rect 88300 12724 88306 12736
rect 89624 12732 89636 12736
rect 89670 12764 89682 12766
rect 89714 12764 89720 12776
rect 89670 12736 89720 12764
rect 89670 12732 89682 12736
rect 89624 12726 89682 12732
rect 89714 12724 89720 12736
rect 89772 12724 89778 12776
rect 89808 12766 89866 12772
rect 89808 12732 89820 12766
rect 89854 12764 89866 12766
rect 89854 12736 89944 12764
rect 89854 12732 89866 12736
rect 89808 12726 89866 12732
rect 89916 12640 89944 12736
rect 90082 12724 90088 12776
rect 90140 12764 90146 12776
rect 91296 12764 91324 12794
rect 90140 12736 91324 12764
rect 90140 12724 90146 12736
rect 98564 12696 98592 12794
rect 105170 12792 105176 12804
rect 105228 12792 105234 12844
rect 106108 12840 106136 12872
rect 106092 12834 106150 12840
rect 106092 12800 106104 12834
rect 106138 12800 106150 12834
rect 106092 12794 106150 12800
rect 99190 12764 99196 12776
rect 99102 12736 99196 12764
rect 99190 12724 99196 12736
rect 99248 12764 99254 12776
rect 101398 12764 101404 12776
rect 99248 12736 101404 12764
rect 99248 12724 99254 12736
rect 101398 12724 101404 12736
rect 101456 12724 101462 12776
rect 101674 12764 101680 12776
rect 101634 12736 101680 12764
rect 101674 12724 101680 12736
rect 101732 12724 101738 12776
rect 104804 12766 104862 12772
rect 104804 12732 104816 12766
rect 104850 12732 104862 12766
rect 104804 12726 104862 12732
rect 100940 12698 100998 12704
rect 98564 12668 99328 12696
rect 87782 12628 87788 12640
rect 86144 12600 87788 12628
rect 87782 12588 87788 12600
rect 87840 12588 87846 12640
rect 87966 12628 87972 12640
rect 87926 12600 87972 12628
rect 87966 12588 87972 12600
rect 88024 12588 88030 12640
rect 88426 12588 88432 12640
rect 88484 12628 88490 12640
rect 89164 12630 89222 12636
rect 89164 12628 89176 12630
rect 88484 12600 89176 12628
rect 88484 12588 88490 12600
rect 89164 12596 89176 12600
rect 89210 12596 89222 12630
rect 89898 12628 89904 12640
rect 89810 12600 89904 12628
rect 89164 12590 89222 12596
rect 89898 12588 89904 12600
rect 89956 12628 89962 12640
rect 90544 12630 90602 12636
rect 90544 12628 90556 12630
rect 89956 12600 90556 12628
rect 89956 12588 89962 12600
rect 90544 12596 90556 12600
rect 90590 12596 90602 12630
rect 90544 12590 90602 12596
rect 98364 12630 98422 12636
rect 98364 12596 98376 12630
rect 98410 12628 98422 12630
rect 99190 12628 99196 12640
rect 98410 12600 99196 12628
rect 98410 12596 98422 12600
rect 98364 12590 98422 12596
rect 99190 12588 99196 12600
rect 99248 12588 99254 12640
rect 99300 12628 99328 12668
rect 100940 12664 100952 12698
rect 100986 12696 100998 12698
rect 101030 12696 101036 12708
rect 100986 12668 101036 12696
rect 100986 12664 100998 12668
rect 100940 12658 100998 12664
rect 101030 12656 101036 12668
rect 101088 12656 101094 12708
rect 103238 12656 103244 12708
rect 103296 12696 103302 12708
rect 104820 12696 104848 12726
rect 105906 12696 105912 12708
rect 103296 12668 104848 12696
rect 105866 12668 105912 12696
rect 103296 12656 103302 12668
rect 105906 12656 105912 12668
rect 105964 12656 105970 12708
rect 108316 12696 108344 12940
rect 111426 12928 111432 12980
rect 111484 12968 111490 12980
rect 112256 12970 112314 12976
rect 112256 12968 112268 12970
rect 111484 12940 112268 12968
rect 111484 12928 111490 12940
rect 112256 12936 112268 12940
rect 112302 12968 112314 12970
rect 114554 12968 114560 12980
rect 112302 12940 114560 12968
rect 112302 12936 112314 12940
rect 112256 12930 112314 12936
rect 114554 12928 114560 12940
rect 114612 12928 114618 12980
rect 114738 12928 114744 12980
rect 114796 12968 114802 12980
rect 117406 12968 117412 12980
rect 114796 12940 117412 12968
rect 114796 12928 114802 12940
rect 117406 12928 117412 12940
rect 117464 12928 117470 12980
rect 118234 12968 118240 12980
rect 118194 12940 118240 12968
rect 118234 12928 118240 12940
rect 118292 12928 118298 12980
rect 118694 12968 118700 12980
rect 118654 12940 118700 12968
rect 118694 12928 118700 12940
rect 118752 12928 118758 12980
rect 126700 12970 126758 12976
rect 126700 12936 126712 12970
rect 126746 12968 126758 12970
rect 126882 12968 126888 12980
rect 126746 12940 126888 12968
rect 126746 12936 126758 12940
rect 126700 12930 126758 12936
rect 126882 12928 126888 12940
rect 126940 12928 126946 12980
rect 128078 12968 128084 12980
rect 128038 12940 128084 12968
rect 128078 12928 128084 12940
rect 128136 12928 128142 12980
rect 128630 12928 128636 12980
rect 128688 12968 128694 12980
rect 128724 12970 128782 12976
rect 128724 12968 128736 12970
rect 128688 12940 128736 12968
rect 128688 12928 128694 12940
rect 128724 12936 128736 12940
rect 128770 12936 128782 12970
rect 129182 12968 129188 12980
rect 129142 12940 129188 12968
rect 128724 12930 128782 12936
rect 129182 12928 129188 12940
rect 129240 12928 129246 12980
rect 130288 12970 130346 12976
rect 130288 12936 130300 12970
rect 130334 12968 130346 12970
rect 133322 12968 133328 12980
rect 130334 12940 133328 12968
rect 130334 12936 130346 12940
rect 130288 12930 130346 12936
rect 133322 12928 133328 12940
rect 133380 12928 133386 12980
rect 133508 12970 133566 12976
rect 133508 12936 133520 12970
rect 133554 12968 133566 12970
rect 133554 12940 133828 12968
rect 133554 12936 133566 12940
rect 133508 12930 133566 12936
rect 109586 12860 109592 12912
rect 109644 12900 109650 12912
rect 112348 12902 112406 12908
rect 112348 12900 112360 12902
rect 109644 12872 112360 12900
rect 109644 12860 109650 12872
rect 112348 12868 112360 12872
rect 112394 12868 112406 12902
rect 114004 12902 114062 12908
rect 114004 12900 114016 12902
rect 112348 12862 112406 12868
rect 112548 12872 114016 12900
rect 112548 12772 112576 12872
rect 114004 12868 114016 12872
rect 114050 12900 114062 12902
rect 115660 12902 115718 12908
rect 114050 12872 115612 12900
rect 114050 12868 114062 12872
rect 114004 12862 114062 12868
rect 113082 12832 113088 12844
rect 113042 12804 113088 12832
rect 113082 12792 113088 12804
rect 113140 12792 113146 12844
rect 113818 12832 113824 12844
rect 113778 12804 113824 12832
rect 113818 12792 113824 12804
rect 113876 12792 113882 12844
rect 114646 12792 114652 12844
rect 114704 12832 114710 12844
rect 115584 12832 115612 12872
rect 115660 12868 115672 12902
rect 115706 12900 115718 12902
rect 115750 12900 115756 12912
rect 115706 12872 115756 12900
rect 115706 12868 115718 12872
rect 115660 12862 115718 12868
rect 115750 12860 115756 12872
rect 115808 12860 115814 12912
rect 117314 12860 117320 12912
rect 117372 12860 117378 12912
rect 126514 12860 126520 12912
rect 126572 12900 126578 12912
rect 129200 12900 129228 12928
rect 132402 12900 132408 12912
rect 126572 12872 129228 12900
rect 132342 12872 132408 12900
rect 126572 12860 126578 12872
rect 114704 12804 114748 12832
rect 115584 12804 115888 12832
rect 114704 12792 114710 12804
rect 115860 12776 115888 12804
rect 118050 12792 118056 12844
rect 118108 12832 118114 12844
rect 126900 12840 126928 12872
rect 132402 12860 132408 12872
rect 132460 12860 132466 12912
rect 133598 12900 133604 12912
rect 133558 12872 133604 12900
rect 133598 12860 133604 12872
rect 133656 12860 133662 12912
rect 133800 12900 133828 12940
rect 133874 12928 133880 12980
rect 133932 12968 133938 12980
rect 134336 12970 134394 12976
rect 134336 12968 134348 12970
rect 133932 12940 134348 12968
rect 133932 12928 133938 12940
rect 134336 12936 134348 12940
rect 134382 12936 134394 12970
rect 134336 12930 134394 12936
rect 145468 12970 145526 12976
rect 145468 12936 145480 12970
rect 145514 12968 145526 12970
rect 147674 12968 147680 12980
rect 145514 12940 147680 12968
rect 145514 12936 145526 12940
rect 145468 12930 145526 12936
rect 147674 12928 147680 12940
rect 147732 12928 147738 12980
rect 151448 12970 151506 12976
rect 148152 12940 149836 12968
rect 134150 12900 134156 12912
rect 133800 12872 134156 12900
rect 134150 12860 134156 12872
rect 134208 12860 134214 12912
rect 143074 12860 143080 12912
rect 143132 12900 143138 12912
rect 145926 12900 145932 12912
rect 143132 12872 145788 12900
rect 145886 12872 145932 12900
rect 143132 12860 143138 12872
rect 118880 12834 118938 12840
rect 118880 12832 118892 12834
rect 118108 12804 118892 12832
rect 118108 12792 118114 12804
rect 118880 12800 118892 12804
rect 118926 12800 118938 12834
rect 118880 12794 118938 12800
rect 126884 12834 126942 12840
rect 126884 12800 126896 12834
rect 126930 12800 126942 12834
rect 127434 12832 127440 12844
rect 127394 12804 127440 12832
rect 126884 12794 126942 12800
rect 127434 12792 127440 12804
rect 127492 12832 127498 12844
rect 128264 12834 128322 12840
rect 127492 12804 128216 12832
rect 127492 12792 127498 12804
rect 112532 12766 112590 12772
rect 112532 12732 112544 12766
rect 112578 12732 112590 12766
rect 112532 12726 112590 12732
rect 113176 12766 113234 12772
rect 113176 12732 113188 12766
rect 113222 12764 113234 12766
rect 113910 12764 113916 12776
rect 113222 12736 113916 12764
rect 113222 12732 113234 12736
rect 113176 12726 113234 12732
rect 113910 12724 113916 12736
rect 113968 12724 113974 12776
rect 114738 12724 114744 12776
rect 114796 12724 114802 12776
rect 115658 12724 115664 12776
rect 115716 12764 115722 12776
rect 115752 12766 115810 12772
rect 115752 12764 115764 12766
rect 115716 12736 115764 12764
rect 115716 12724 115722 12736
rect 115752 12732 115764 12736
rect 115798 12732 115810 12766
rect 115752 12726 115810 12732
rect 115842 12724 115848 12776
rect 115900 12764 115906 12776
rect 116488 12766 116546 12772
rect 115900 12736 115944 12764
rect 115900 12724 115906 12736
rect 116488 12732 116500 12766
rect 116534 12732 116546 12766
rect 116762 12764 116768 12776
rect 116722 12736 116768 12764
rect 116488 12726 116546 12732
rect 114756 12696 114784 12724
rect 108316 12668 114784 12696
rect 114830 12656 114836 12708
rect 114888 12696 114894 12708
rect 116504 12696 116532 12726
rect 116762 12724 116768 12736
rect 116820 12724 116826 12776
rect 127526 12764 127532 12776
rect 117792 12736 127532 12764
rect 114888 12668 116532 12696
rect 114888 12656 114894 12668
rect 100754 12628 100760 12640
rect 99300 12600 100760 12628
rect 100754 12588 100760 12600
rect 100812 12588 100818 12640
rect 103054 12588 103060 12640
rect 103112 12628 103118 12640
rect 103148 12630 103206 12636
rect 103148 12628 103160 12630
rect 103112 12600 103160 12628
rect 103112 12588 103118 12600
rect 103148 12596 103160 12600
rect 103194 12596 103206 12630
rect 103148 12590 103206 12596
rect 103606 12588 103612 12640
rect 103664 12628 103670 12640
rect 104252 12630 104310 12636
rect 104252 12628 104264 12630
rect 103664 12600 104264 12628
rect 103664 12588 103670 12600
rect 104252 12596 104264 12600
rect 104298 12596 104310 12630
rect 111886 12628 111892 12640
rect 111846 12600 111892 12628
rect 104252 12590 104310 12596
rect 111886 12588 111892 12600
rect 111944 12588 111950 12640
rect 113082 12588 113088 12640
rect 113140 12628 113146 12640
rect 114738 12628 114744 12640
rect 113140 12600 114744 12628
rect 113140 12588 113146 12600
rect 114738 12588 114744 12600
rect 114796 12588 114802 12640
rect 115292 12630 115350 12636
rect 115292 12596 115304 12630
rect 115338 12628 115350 12630
rect 115842 12628 115848 12640
rect 115338 12600 115848 12628
rect 115338 12596 115350 12600
rect 115292 12590 115350 12596
rect 115842 12588 115848 12600
rect 115900 12588 115906 12640
rect 116504 12628 116532 12668
rect 117792 12628 117820 12736
rect 127526 12724 127532 12736
rect 127584 12724 127590 12776
rect 116504 12600 117820 12628
rect 127528 12630 127586 12636
rect 127528 12596 127540 12630
rect 127574 12628 127586 12630
rect 128078 12628 128084 12640
rect 127574 12600 128084 12628
rect 127574 12596 127586 12600
rect 127528 12590 127586 12596
rect 128078 12588 128084 12600
rect 128136 12588 128142 12640
rect 128188 12628 128216 12804
rect 128264 12800 128276 12834
rect 128310 12800 128322 12834
rect 129090 12832 129096 12844
rect 129050 12804 129096 12832
rect 128264 12794 128322 12800
rect 128280 12696 128308 12794
rect 129090 12792 129096 12804
rect 129148 12792 129154 12844
rect 130196 12834 130254 12840
rect 130196 12832 130208 12834
rect 129200 12804 130208 12832
rect 128354 12724 128360 12776
rect 128412 12764 128418 12776
rect 129200 12764 129228 12804
rect 130196 12800 130208 12804
rect 130242 12800 130254 12834
rect 130196 12794 130254 12800
rect 130286 12792 130292 12844
rect 130344 12832 130350 12844
rect 130840 12834 130898 12840
rect 130840 12832 130852 12834
rect 130344 12804 130852 12832
rect 130344 12792 130350 12804
rect 130840 12800 130852 12804
rect 130886 12800 130898 12834
rect 130840 12794 130898 12800
rect 128412 12736 129228 12764
rect 129368 12766 129426 12772
rect 128412 12724 128418 12736
rect 129368 12732 129380 12766
rect 129414 12764 129426 12766
rect 129734 12764 129740 12776
rect 129414 12736 129740 12764
rect 129414 12732 129426 12736
rect 129368 12726 129426 12732
rect 129734 12724 129740 12736
rect 129792 12724 129798 12776
rect 131114 12764 131120 12776
rect 131074 12736 131120 12764
rect 131114 12724 131120 12736
rect 131172 12724 131178 12776
rect 132586 12724 132592 12776
rect 132644 12764 132650 12776
rect 133616 12764 133644 12860
rect 133690 12792 133696 12844
rect 133748 12836 133754 12844
rect 133748 12832 133828 12836
rect 134520 12834 134578 12840
rect 134520 12832 134532 12834
rect 133748 12808 134532 12832
rect 133748 12792 133754 12808
rect 133800 12804 134532 12808
rect 134520 12800 134532 12804
rect 134566 12800 134578 12834
rect 134520 12794 134578 12800
rect 135348 12834 135406 12840
rect 135348 12800 135360 12834
rect 135394 12832 135406 12834
rect 142984 12834 143042 12840
rect 142984 12832 142996 12834
rect 135394 12804 142996 12832
rect 135394 12800 135406 12804
rect 135348 12794 135406 12800
rect 142984 12800 142996 12804
rect 143030 12832 143042 12834
rect 145760 12832 145788 12872
rect 145926 12860 145932 12872
rect 145984 12860 145990 12912
rect 148152 12900 148180 12940
rect 146036 12872 148180 12900
rect 149808 12900 149836 12940
rect 151448 12936 151460 12970
rect 151494 12968 151506 12970
rect 152642 12968 152648 12980
rect 151494 12940 152648 12968
rect 151494 12936 151506 12940
rect 151448 12930 151506 12936
rect 152642 12928 152648 12940
rect 152700 12928 152706 12980
rect 152736 12970 152794 12976
rect 152736 12936 152748 12970
rect 152782 12968 152794 12970
rect 152826 12968 152832 12980
rect 152782 12940 152832 12968
rect 152782 12936 152794 12940
rect 152736 12930 152794 12936
rect 152826 12928 152832 12940
rect 152884 12968 152890 12980
rect 153104 12970 153162 12976
rect 153104 12968 153116 12970
rect 152884 12940 153116 12968
rect 152884 12928 152890 12940
rect 153104 12936 153116 12940
rect 153150 12968 153162 12970
rect 153472 12970 153530 12976
rect 153472 12968 153484 12970
rect 153150 12940 153484 12968
rect 153150 12936 153162 12940
rect 153104 12930 153162 12936
rect 153472 12936 153484 12940
rect 153518 12968 153530 12970
rect 153840 12970 153898 12976
rect 153840 12968 153852 12970
rect 153518 12940 153852 12968
rect 153518 12936 153530 12940
rect 153472 12930 153530 12936
rect 153840 12936 153852 12940
rect 153886 12968 153898 12970
rect 154208 12970 154266 12976
rect 154208 12968 154220 12970
rect 153886 12940 154220 12968
rect 153886 12936 153898 12940
rect 153840 12930 153898 12936
rect 154208 12936 154220 12940
rect 154254 12968 154266 12970
rect 154944 12970 155002 12976
rect 154944 12968 154956 12970
rect 154254 12940 154956 12968
rect 154254 12936 154266 12940
rect 154208 12930 154266 12936
rect 154944 12936 154956 12940
rect 154990 12968 155002 12970
rect 156048 12970 156106 12976
rect 156048 12968 156060 12970
rect 154990 12940 156060 12968
rect 154990 12936 155002 12940
rect 154944 12930 155002 12936
rect 156048 12936 156060 12940
rect 156094 12968 156106 12970
rect 156416 12970 156474 12976
rect 156416 12968 156428 12970
rect 156094 12940 156428 12968
rect 156094 12936 156106 12940
rect 156048 12930 156106 12936
rect 156416 12936 156428 12940
rect 156462 12968 156474 12970
rect 156784 12970 156842 12976
rect 156784 12968 156796 12970
rect 156462 12940 156796 12968
rect 156462 12936 156474 12940
rect 156416 12930 156474 12936
rect 156784 12936 156796 12940
rect 156830 12968 156842 12970
rect 157150 12968 157156 12980
rect 156830 12940 157156 12968
rect 156830 12936 156842 12940
rect 156784 12930 156842 12936
rect 157150 12928 157156 12940
rect 157208 12928 157214 12980
rect 158622 12928 158628 12980
rect 158680 12968 158686 12980
rect 163498 12968 163504 12980
rect 158680 12940 163504 12968
rect 158680 12928 158686 12940
rect 156598 12900 156604 12912
rect 149808 12872 156604 12900
rect 145834 12832 145840 12844
rect 143030 12804 145696 12832
rect 145746 12804 145840 12832
rect 143030 12800 143042 12804
rect 142984 12794 143042 12800
rect 132644 12736 133644 12764
rect 133784 12766 133842 12772
rect 132644 12724 132650 12736
rect 133784 12732 133796 12766
rect 133830 12732 133842 12766
rect 143258 12764 143264 12776
rect 143218 12736 143264 12764
rect 133784 12726 133842 12732
rect 130286 12696 130292 12708
rect 128280 12668 130292 12696
rect 130286 12656 130292 12668
rect 130344 12656 130350 12708
rect 133690 12696 133696 12708
rect 132466 12668 133696 12696
rect 132466 12628 132494 12668
rect 133690 12656 133696 12668
rect 133748 12656 133754 12708
rect 133138 12628 133144 12640
rect 128188 12600 132494 12628
rect 133098 12600 133144 12628
rect 133138 12588 133144 12600
rect 133196 12588 133202 12640
rect 133230 12588 133236 12640
rect 133288 12628 133294 12640
rect 133800 12628 133828 12726
rect 143258 12724 143264 12736
rect 143316 12724 143322 12776
rect 145668 12764 145696 12804
rect 145834 12792 145840 12804
rect 145892 12792 145898 12844
rect 146036 12832 146064 12872
rect 156598 12860 156604 12872
rect 156656 12860 156662 12912
rect 159268 12902 159326 12908
rect 159268 12900 159280 12902
rect 157306 12872 159280 12900
rect 145944 12804 146064 12832
rect 147032 12834 147090 12840
rect 145944 12764 145972 12804
rect 147032 12800 147044 12834
rect 147078 12832 147090 12834
rect 147306 12832 147312 12844
rect 147078 12804 147312 12832
rect 147078 12800 147090 12804
rect 147032 12794 147090 12800
rect 147306 12792 147312 12804
rect 147364 12792 147370 12844
rect 148902 12804 149008 12832
rect 148980 12776 149008 12804
rect 149330 12792 149336 12844
rect 149388 12832 149394 12844
rect 149884 12834 149942 12840
rect 149884 12832 149896 12834
rect 149388 12804 149896 12832
rect 149388 12792 149394 12804
rect 149884 12800 149896 12804
rect 149930 12832 149942 12834
rect 149930 12804 150388 12832
rect 149930 12800 149942 12804
rect 149884 12794 149942 12800
rect 145668 12736 145972 12764
rect 146112 12766 146170 12772
rect 146112 12732 146124 12766
rect 146158 12764 146170 12766
rect 147398 12764 147404 12776
rect 146158 12736 147404 12764
rect 146158 12732 146170 12736
rect 146112 12726 146170 12732
rect 147398 12724 147404 12736
rect 147456 12724 147462 12776
rect 147492 12766 147550 12772
rect 147492 12732 147504 12766
rect 147538 12732 147550 12766
rect 147766 12764 147772 12776
rect 147726 12736 147772 12764
rect 147492 12726 147550 12732
rect 133874 12656 133880 12708
rect 133932 12696 133938 12708
rect 135532 12698 135590 12704
rect 135532 12696 135544 12698
rect 133932 12668 135544 12696
rect 133932 12656 133938 12668
rect 135532 12664 135544 12668
rect 135578 12664 135590 12698
rect 135532 12658 135590 12664
rect 145742 12656 145748 12708
rect 145800 12696 145806 12708
rect 147508 12696 147536 12726
rect 147766 12724 147772 12736
rect 147824 12724 147830 12776
rect 148962 12724 148968 12776
rect 149020 12724 149026 12776
rect 149238 12764 149244 12776
rect 149198 12736 149244 12764
rect 149238 12724 149244 12736
rect 149296 12724 149302 12776
rect 150360 12708 150388 12804
rect 150434 12792 150440 12844
rect 150492 12832 150498 12844
rect 154852 12834 154910 12840
rect 154852 12832 154864 12834
rect 150492 12804 154864 12832
rect 150492 12792 150498 12804
rect 154852 12800 154864 12804
rect 154898 12800 154910 12834
rect 154852 12794 154910 12800
rect 155862 12792 155868 12844
rect 155920 12832 155926 12844
rect 157306 12832 157334 12872
rect 159268 12868 159280 12872
rect 159314 12868 159326 12902
rect 160370 12900 160376 12912
rect 159268 12862 159326 12868
rect 159928 12872 160376 12900
rect 155920 12804 157334 12832
rect 155920 12792 155926 12804
rect 157794 12792 157800 12844
rect 157852 12832 157858 12844
rect 159176 12834 159234 12840
rect 159176 12832 159188 12834
rect 157852 12804 159188 12832
rect 157852 12792 157858 12804
rect 159176 12800 159188 12804
rect 159222 12832 159234 12834
rect 159928 12832 159956 12872
rect 160370 12860 160376 12872
rect 160428 12860 160434 12912
rect 161124 12872 161796 12900
rect 159222 12804 159956 12832
rect 160004 12834 160062 12840
rect 159222 12800 159234 12804
rect 159176 12794 159234 12800
rect 160004 12800 160016 12834
rect 160050 12832 160062 12834
rect 161124 12832 161152 12872
rect 160050 12804 161152 12832
rect 161200 12834 161258 12840
rect 160050 12800 160062 12804
rect 160004 12794 160062 12800
rect 161200 12800 161212 12834
rect 161246 12832 161258 12834
rect 161658 12832 161664 12844
rect 161246 12804 161664 12832
rect 161246 12800 161258 12804
rect 161200 12794 161258 12800
rect 161658 12792 161664 12804
rect 161716 12792 161722 12844
rect 151538 12764 151544 12776
rect 151498 12736 151544 12764
rect 151538 12724 151544 12736
rect 151596 12724 151602 12776
rect 151724 12766 151782 12772
rect 151724 12732 151736 12766
rect 151770 12732 151782 12766
rect 151724 12726 151782 12732
rect 145800 12668 147536 12696
rect 145800 12656 145806 12668
rect 150342 12656 150348 12708
rect 150400 12696 150406 12708
rect 151630 12696 151636 12708
rect 150400 12668 151636 12696
rect 150400 12656 150406 12668
rect 151630 12656 151636 12668
rect 151688 12656 151694 12708
rect 133288 12600 133828 12628
rect 146848 12630 146906 12636
rect 133288 12588 133294 12600
rect 146848 12596 146860 12630
rect 146894 12628 146906 12630
rect 148502 12628 148508 12640
rect 146894 12600 148508 12628
rect 146894 12596 146906 12600
rect 146848 12590 146906 12596
rect 148502 12588 148508 12600
rect 148560 12588 148566 12640
rect 149974 12628 149980 12640
rect 149934 12600 149980 12628
rect 149974 12588 149980 12600
rect 150032 12588 150038 12640
rect 151080 12630 151138 12636
rect 151080 12596 151092 12630
rect 151126 12628 151138 12630
rect 151262 12628 151268 12640
rect 151126 12600 151268 12628
rect 151126 12596 151138 12600
rect 151080 12590 151138 12596
rect 151262 12588 151268 12600
rect 151320 12588 151326 12640
rect 151354 12588 151360 12640
rect 151412 12628 151418 12640
rect 151740 12628 151768 12726
rect 152734 12724 152740 12776
rect 152792 12764 152798 12776
rect 152792 12736 154988 12764
rect 152792 12724 152798 12736
rect 152368 12698 152426 12704
rect 152368 12664 152380 12698
rect 152414 12696 152426 12698
rect 152826 12696 152832 12708
rect 152414 12668 152832 12696
rect 152414 12664 152426 12668
rect 152368 12658 152426 12664
rect 152826 12656 152832 12668
rect 152884 12656 152890 12708
rect 153102 12656 153108 12708
rect 153160 12696 153166 12708
rect 154484 12698 154542 12704
rect 154484 12696 154496 12698
rect 153160 12668 154496 12696
rect 153160 12656 153166 12668
rect 154484 12664 154496 12668
rect 154530 12664 154542 12698
rect 154960 12696 154988 12736
rect 155034 12724 155040 12776
rect 155092 12764 155098 12776
rect 159450 12764 159456 12776
rect 155092 12736 155136 12764
rect 155236 12736 159312 12764
rect 159410 12736 159456 12764
rect 155092 12724 155098 12736
rect 155236 12696 155264 12736
rect 158806 12696 158812 12708
rect 154960 12668 155264 12696
rect 158766 12668 158812 12696
rect 154484 12658 154542 12664
rect 158806 12656 158812 12668
rect 158864 12656 158870 12708
rect 159284 12696 159312 12736
rect 159450 12724 159456 12736
rect 159508 12724 159514 12776
rect 159542 12724 159548 12776
rect 159600 12764 159606 12776
rect 161566 12764 161572 12776
rect 159600 12736 161572 12764
rect 159600 12724 159606 12736
rect 161566 12724 161572 12736
rect 161624 12724 161630 12776
rect 160188 12698 160246 12704
rect 160188 12696 160200 12698
rect 159284 12668 160200 12696
rect 160188 12664 160200 12668
rect 160234 12664 160246 12698
rect 160188 12658 160246 12664
rect 154114 12628 154120 12640
rect 151412 12600 154120 12628
rect 151412 12588 151418 12600
rect 154114 12588 154120 12600
rect 154172 12628 154178 12640
rect 157886 12628 157892 12640
rect 154172 12600 157892 12628
rect 154172 12588 154178 12600
rect 157886 12588 157892 12600
rect 157944 12588 157950 12640
rect 160278 12588 160284 12640
rect 160336 12628 160342 12640
rect 161292 12630 161350 12636
rect 161292 12628 161304 12630
rect 160336 12600 161304 12628
rect 160336 12588 160342 12600
rect 161292 12596 161304 12600
rect 161338 12596 161350 12630
rect 161768 12628 161796 12872
rect 161860 12840 161888 12940
rect 163498 12928 163504 12940
rect 163556 12928 163562 12980
rect 163592 12970 163650 12976
rect 163592 12936 163604 12970
rect 163638 12936 163650 12970
rect 163592 12930 163650 12936
rect 164420 12970 164478 12976
rect 164420 12936 164432 12970
rect 164466 12968 164478 12970
rect 165246 12968 165252 12980
rect 164466 12940 165252 12968
rect 164466 12936 164478 12940
rect 164420 12930 164478 12936
rect 163406 12900 163412 12912
rect 163346 12872 163412 12900
rect 163406 12860 163412 12872
rect 163464 12860 163470 12912
rect 163608 12900 163636 12930
rect 165246 12928 165252 12940
rect 165304 12968 165310 12980
rect 165304 12940 166994 12968
rect 165304 12928 165310 12940
rect 164512 12902 164570 12908
rect 164512 12900 164524 12902
rect 163608 12872 164524 12900
rect 161844 12834 161902 12840
rect 161844 12800 161856 12834
rect 161890 12800 161902 12834
rect 161844 12794 161902 12800
rect 162118 12764 162124 12776
rect 162078 12736 162124 12764
rect 162118 12724 162124 12736
rect 162176 12724 162182 12776
rect 162854 12724 162860 12776
rect 162912 12764 162918 12776
rect 163608 12764 163636 12872
rect 164512 12868 164524 12872
rect 164558 12900 164570 12902
rect 166966 12900 166994 12940
rect 167178 12928 167184 12980
rect 167236 12968 167242 12980
rect 167824 12970 167882 12976
rect 167824 12968 167836 12970
rect 167236 12940 167836 12968
rect 167236 12928 167242 12940
rect 167824 12936 167836 12940
rect 167870 12936 167882 12970
rect 174998 12968 175004 12980
rect 174958 12940 175004 12968
rect 167824 12930 167882 12936
rect 174998 12928 175004 12940
rect 175056 12928 175062 12980
rect 175644 12970 175702 12976
rect 175644 12936 175656 12970
rect 175690 12968 175702 12970
rect 175734 12968 175740 12980
rect 175690 12940 175740 12968
rect 175690 12936 175702 12940
rect 175644 12930 175702 12936
rect 175734 12928 175740 12940
rect 175792 12928 175798 12980
rect 176378 12928 176384 12980
rect 176436 12968 176442 12980
rect 180150 12968 180156 12980
rect 176436 12940 180156 12968
rect 176436 12928 176442 12940
rect 164558 12872 166672 12900
rect 166966 12872 168052 12900
rect 164558 12868 164570 12872
rect 164512 12862 164570 12868
rect 165340 12834 165398 12840
rect 165340 12800 165352 12834
rect 165386 12832 165398 12834
rect 165430 12832 165436 12844
rect 165386 12804 165436 12832
rect 165386 12800 165398 12804
rect 165340 12794 165398 12800
rect 165430 12792 165436 12804
rect 165488 12792 165494 12844
rect 166166 12792 166172 12844
rect 166224 12832 166230 12844
rect 166534 12832 166540 12844
rect 166224 12804 166540 12832
rect 166224 12792 166230 12804
rect 166534 12792 166540 12804
rect 166592 12792 166598 12844
rect 166644 12832 166672 12872
rect 168024 12840 168052 12872
rect 173802 12860 173808 12912
rect 173860 12900 173866 12912
rect 173860 12872 175872 12900
rect 173860 12860 173866 12872
rect 175844 12840 175872 12872
rect 175918 12860 175924 12912
rect 175976 12900 175982 12912
rect 176930 12900 176936 12912
rect 175976 12872 176936 12900
rect 175976 12860 175982 12872
rect 176930 12860 176936 12872
rect 176988 12860 176994 12912
rect 177942 12900 177948 12912
rect 177882 12872 177948 12900
rect 177942 12860 177948 12872
rect 178000 12860 178006 12912
rect 167364 12834 167422 12840
rect 167364 12832 167376 12834
rect 166644 12804 167376 12832
rect 167364 12800 167376 12804
rect 167410 12800 167422 12834
rect 167364 12794 167422 12800
rect 168008 12834 168066 12840
rect 168008 12800 168020 12834
rect 168054 12800 168066 12834
rect 168008 12794 168066 12800
rect 175184 12834 175242 12840
rect 175184 12800 175196 12834
rect 175230 12800 175242 12834
rect 175184 12794 175242 12800
rect 175828 12834 175886 12840
rect 175828 12800 175840 12834
rect 175874 12800 175886 12834
rect 176378 12832 176384 12844
rect 176338 12804 176384 12832
rect 175828 12794 175886 12800
rect 164602 12764 164608 12776
rect 162912 12736 163636 12764
rect 164562 12736 164608 12764
rect 162912 12724 162918 12736
rect 164602 12724 164608 12736
rect 164660 12724 164666 12776
rect 163608 12668 164188 12696
rect 163608 12628 163636 12668
rect 161768 12600 163636 12628
rect 161292 12590 161350 12596
rect 163682 12588 163688 12640
rect 163740 12628 163746 12640
rect 164052 12630 164110 12636
rect 164052 12628 164064 12630
rect 163740 12600 164064 12628
rect 163740 12588 163746 12600
rect 164052 12596 164064 12600
rect 164098 12596 164110 12630
rect 164160 12628 164188 12668
rect 164234 12656 164240 12708
rect 164292 12696 164298 12708
rect 167180 12698 167238 12704
rect 167180 12696 167192 12698
rect 164292 12668 167192 12696
rect 164292 12656 164298 12668
rect 167180 12664 167192 12668
rect 167226 12664 167238 12698
rect 175200 12696 175228 12794
rect 176378 12792 176384 12804
rect 176436 12792 176442 12844
rect 178604 12840 178632 12940
rect 180150 12928 180156 12940
rect 180208 12928 180214 12980
rect 180242 12928 180248 12980
rect 180300 12968 180306 12980
rect 180796 12970 180854 12976
rect 180796 12968 180808 12970
rect 180300 12940 180808 12968
rect 180300 12928 180306 12940
rect 180796 12936 180808 12940
rect 180842 12936 180854 12970
rect 188338 12968 188344 12980
rect 180796 12930 180854 12936
rect 188080 12940 188344 12968
rect 181624 12902 181682 12908
rect 181624 12900 181636 12902
rect 180260 12872 181636 12900
rect 178588 12834 178646 12840
rect 178588 12800 178600 12834
rect 178634 12800 178646 12834
rect 180260 12832 180288 12872
rect 181624 12868 181636 12872
rect 181670 12868 181682 12902
rect 181624 12862 181682 12868
rect 179998 12804 180288 12832
rect 178588 12794 178646 12800
rect 180334 12792 180340 12844
rect 180392 12832 180398 12844
rect 180980 12834 181038 12840
rect 180980 12832 180992 12834
rect 180392 12804 180992 12832
rect 180392 12792 180398 12804
rect 180980 12800 180992 12804
rect 181026 12800 181038 12834
rect 181530 12832 181536 12844
rect 181442 12804 181536 12832
rect 180980 12794 181038 12800
rect 181530 12792 181536 12804
rect 181588 12832 181594 12844
rect 188080 12840 188108 12940
rect 188338 12928 188344 12940
rect 188396 12968 188402 12980
rect 191374 12968 191380 12980
rect 188396 12940 191380 12968
rect 188396 12928 188402 12940
rect 191374 12928 191380 12940
rect 191432 12968 191438 12980
rect 192296 12970 192354 12976
rect 192296 12968 192308 12970
rect 191432 12940 192308 12968
rect 191432 12928 191438 12940
rect 192296 12936 192308 12940
rect 192342 12936 192354 12970
rect 192296 12930 192354 12936
rect 192478 12928 192484 12980
rect 192536 12968 192542 12980
rect 192536 12940 193444 12968
rect 192536 12928 192542 12940
rect 188522 12860 188528 12912
rect 188580 12900 188586 12912
rect 189536 12902 189594 12908
rect 189536 12900 189548 12902
rect 188580 12872 189548 12900
rect 188580 12860 188586 12872
rect 189536 12868 189548 12872
rect 189582 12900 189594 12902
rect 190914 12900 190920 12912
rect 189582 12872 190454 12900
rect 190874 12872 190920 12900
rect 189582 12868 189594 12872
rect 189536 12862 189594 12868
rect 182176 12834 182234 12840
rect 182176 12832 182188 12834
rect 181588 12804 182188 12832
rect 181588 12792 181594 12804
rect 182176 12800 182188 12804
rect 182222 12800 182234 12834
rect 182176 12794 182234 12800
rect 188064 12834 188122 12840
rect 188064 12800 188076 12834
rect 188110 12800 188122 12834
rect 188064 12794 188122 12800
rect 188338 12792 188344 12844
rect 188396 12832 188402 12844
rect 188616 12834 188674 12840
rect 188616 12832 188628 12834
rect 188396 12804 188628 12832
rect 188396 12792 188402 12804
rect 188616 12800 188628 12804
rect 188662 12832 188674 12834
rect 188798 12832 188804 12844
rect 188662 12804 188804 12832
rect 188662 12800 188674 12804
rect 188616 12794 188674 12800
rect 188798 12792 188804 12804
rect 188856 12792 188862 12844
rect 189350 12832 189356 12844
rect 189310 12804 189356 12832
rect 189350 12792 189356 12804
rect 189408 12792 189414 12844
rect 176656 12766 176714 12772
rect 176656 12732 176668 12766
rect 176702 12764 176714 12766
rect 176746 12764 176752 12776
rect 176702 12736 176752 12764
rect 176702 12732 176714 12736
rect 176656 12726 176714 12732
rect 176746 12724 176752 12736
rect 176804 12724 176810 12776
rect 178864 12766 178922 12772
rect 178864 12732 178876 12766
rect 178910 12764 178922 12766
rect 178910 12736 180104 12764
rect 178910 12732 178922 12736
rect 178864 12726 178922 12732
rect 180076 12696 180104 12736
rect 180150 12724 180156 12776
rect 180208 12764 180214 12776
rect 189534 12764 189540 12776
rect 180208 12736 189540 12764
rect 180208 12724 180214 12736
rect 189534 12724 189540 12736
rect 189592 12724 189598 12776
rect 190426 12764 190454 12872
rect 190914 12860 190920 12872
rect 190972 12860 190978 12912
rect 191742 12860 191748 12912
rect 191800 12900 191806 12912
rect 193308 12902 193366 12908
rect 193308 12900 193320 12902
rect 191800 12872 193320 12900
rect 191800 12860 191806 12872
rect 193308 12868 193320 12872
rect 193354 12868 193366 12902
rect 193416 12900 193444 12940
rect 193950 12928 193956 12980
rect 194008 12968 194014 12980
rect 194870 12968 194876 12980
rect 194008 12940 194876 12968
rect 194008 12928 194014 12940
rect 194870 12928 194876 12940
rect 194928 12968 194934 12980
rect 195974 12968 195980 12980
rect 194928 12940 195980 12968
rect 194928 12928 194934 12940
rect 195974 12928 195980 12940
rect 196032 12928 196038 12980
rect 197722 12928 197728 12980
rect 197780 12968 197786 12980
rect 197780 12940 206508 12968
rect 197780 12928 197786 12940
rect 195884 12902 195942 12908
rect 195884 12900 195896 12902
rect 193416 12872 193798 12900
rect 195072 12872 195896 12900
rect 193308 12862 193366 12868
rect 195072 12844 195100 12872
rect 195884 12868 195896 12872
rect 195930 12868 195942 12902
rect 202966 12900 202972 12912
rect 195884 12862 195942 12868
rect 202524 12872 202972 12900
rect 191008 12834 191066 12840
rect 191008 12800 191020 12834
rect 191054 12832 191066 12834
rect 192204 12834 192262 12840
rect 192204 12832 192216 12834
rect 191054 12804 192216 12832
rect 191054 12800 191066 12804
rect 191008 12794 191066 12800
rect 192204 12800 192216 12804
rect 192250 12832 192262 12834
rect 192570 12832 192576 12844
rect 192250 12804 192576 12832
rect 192250 12800 192262 12804
rect 192204 12794 192262 12800
rect 192570 12792 192576 12804
rect 192628 12792 192634 12844
rect 195054 12832 195060 12844
rect 195014 12804 195060 12832
rect 195054 12792 195060 12804
rect 195112 12792 195118 12844
rect 197354 12832 197360 12844
rect 197314 12804 197360 12832
rect 197354 12792 197360 12804
rect 197412 12792 197418 12844
rect 197446 12792 197452 12844
rect 197504 12832 197510 12844
rect 198366 12832 198372 12844
rect 197504 12804 198136 12832
rect 198326 12804 198372 12832
rect 197504 12792 197510 12804
rect 191192 12766 191250 12772
rect 191192 12764 191204 12766
rect 190426 12736 191204 12764
rect 191192 12732 191204 12736
rect 191238 12764 191250 12766
rect 192388 12766 192446 12772
rect 192388 12764 192400 12766
rect 191238 12736 192400 12764
rect 191238 12732 191250 12736
rect 191192 12726 191250 12732
rect 192388 12732 192400 12736
rect 192434 12764 192446 12766
rect 192662 12764 192668 12776
rect 192434 12736 192668 12764
rect 192434 12732 192446 12736
rect 192388 12726 192446 12732
rect 192662 12724 192668 12736
rect 192720 12724 192726 12776
rect 193030 12764 193036 12776
rect 192990 12736 193036 12764
rect 193030 12724 193036 12736
rect 193088 12724 193094 12776
rect 194778 12764 194784 12776
rect 193140 12736 194784 12764
rect 180242 12696 180248 12708
rect 175200 12668 176148 12696
rect 180076 12668 180248 12696
rect 167180 12658 167238 12664
rect 165432 12630 165490 12636
rect 165432 12628 165444 12630
rect 164160 12600 165444 12628
rect 164052 12590 164110 12596
rect 165432 12596 165444 12600
rect 165478 12628 165490 12630
rect 166166 12628 166172 12640
rect 165478 12600 166172 12628
rect 165478 12596 165490 12600
rect 165432 12590 165490 12596
rect 166166 12588 166172 12600
rect 166224 12588 166230 12640
rect 166626 12628 166632 12640
rect 166586 12600 166632 12628
rect 166626 12588 166632 12600
rect 166684 12588 166690 12640
rect 176120 12628 176148 12668
rect 180242 12656 180248 12668
rect 180300 12656 180306 12708
rect 180518 12656 180524 12708
rect 180576 12696 180582 12708
rect 182082 12696 182088 12708
rect 180576 12668 182088 12696
rect 180576 12656 180582 12668
rect 182082 12656 182088 12668
rect 182140 12656 182146 12708
rect 187880 12698 187938 12704
rect 187880 12664 187892 12698
rect 187926 12696 187938 12698
rect 188614 12696 188620 12708
rect 187926 12668 188620 12696
rect 187926 12664 187938 12668
rect 187880 12658 187938 12664
rect 188614 12656 188620 12668
rect 188672 12656 188678 12708
rect 189166 12656 189172 12708
rect 189224 12696 189230 12708
rect 191742 12696 191748 12708
rect 189224 12668 191748 12696
rect 189224 12656 189230 12668
rect 191742 12656 191748 12668
rect 191800 12656 191806 12708
rect 191926 12656 191932 12708
rect 191984 12696 191990 12708
rect 192478 12696 192484 12708
rect 191984 12668 192484 12696
rect 191984 12656 191990 12668
rect 192478 12656 192484 12668
rect 192536 12656 192542 12708
rect 193140 12696 193168 12736
rect 194778 12724 194784 12736
rect 194836 12724 194842 12776
rect 195790 12724 195796 12776
rect 195848 12764 195854 12776
rect 196160 12766 196218 12772
rect 196160 12764 196172 12766
rect 195848 12736 196172 12764
rect 195848 12724 195854 12736
rect 196160 12732 196172 12736
rect 196206 12764 196218 12766
rect 197630 12764 197636 12776
rect 196206 12736 197636 12764
rect 196206 12732 196218 12736
rect 196160 12726 196218 12732
rect 197630 12724 197636 12736
rect 197688 12724 197694 12776
rect 198108 12772 198136 12804
rect 198366 12792 198372 12804
rect 198424 12792 198430 12844
rect 200484 12834 200542 12840
rect 200484 12800 200496 12834
rect 200530 12832 200542 12834
rect 200666 12832 200672 12844
rect 200530 12804 200672 12832
rect 200530 12800 200542 12804
rect 200484 12794 200542 12800
rect 200666 12792 200672 12804
rect 200724 12792 200730 12844
rect 201310 12832 201316 12844
rect 201270 12804 201316 12832
rect 201310 12792 201316 12804
rect 201368 12792 201374 12844
rect 198092 12766 198150 12772
rect 198092 12732 198104 12766
rect 198138 12764 198150 12766
rect 198550 12764 198556 12776
rect 198138 12736 198556 12764
rect 198138 12732 198150 12736
rect 198092 12726 198150 12732
rect 198550 12724 198556 12736
rect 198608 12764 198614 12776
rect 200390 12764 200396 12776
rect 198608 12736 200396 12764
rect 198608 12724 198614 12736
rect 200390 12724 200396 12736
rect 200448 12724 200454 12776
rect 200576 12766 200634 12772
rect 200576 12732 200588 12766
rect 200622 12764 200634 12766
rect 202524 12764 202552 12872
rect 202966 12860 202972 12872
rect 203024 12860 203030 12912
rect 203334 12860 203340 12912
rect 203392 12860 203398 12912
rect 204824 12840 204852 12940
rect 205634 12860 205640 12912
rect 205692 12860 205698 12912
rect 204808 12834 204866 12840
rect 204808 12800 204820 12834
rect 204854 12800 204866 12834
rect 206480 12832 206508 12940
rect 206554 12928 206560 12980
rect 206612 12968 206618 12980
rect 207382 12968 207388 12980
rect 206612 12940 207388 12968
rect 206612 12928 206618 12940
rect 207382 12928 207388 12940
rect 207440 12928 207446 12980
rect 207842 12928 207848 12980
rect 207900 12968 207906 12980
rect 207900 12940 219756 12968
rect 207900 12928 207906 12940
rect 206664 12872 207612 12900
rect 206664 12832 206692 12872
rect 206480 12804 206692 12832
rect 207476 12834 207534 12840
rect 204808 12794 204866 12800
rect 207476 12800 207488 12834
rect 207522 12800 207534 12834
rect 207476 12794 207534 12800
rect 200622 12736 202552 12764
rect 202600 12766 202658 12772
rect 200622 12732 200634 12736
rect 200576 12726 200634 12732
rect 202600 12732 202612 12766
rect 202646 12732 202658 12766
rect 202874 12764 202880 12776
rect 202834 12736 202880 12764
rect 202600 12726 202658 12732
rect 202138 12696 202144 12708
rect 192588 12668 193168 12696
rect 194336 12668 202144 12696
rect 177390 12628 177396 12640
rect 176120 12600 177396 12628
rect 177390 12588 177396 12600
rect 177448 12588 177454 12640
rect 177850 12588 177856 12640
rect 177908 12628 177914 12640
rect 178128 12630 178186 12636
rect 178128 12628 178140 12630
rect 177908 12600 178140 12628
rect 177908 12588 177914 12600
rect 178128 12596 178140 12600
rect 178174 12596 178186 12630
rect 178128 12590 178186 12596
rect 179874 12588 179880 12640
rect 179932 12628 179938 12640
rect 180336 12630 180394 12636
rect 180336 12628 180348 12630
rect 179932 12600 180348 12628
rect 179932 12588 179938 12600
rect 180336 12596 180348 12600
rect 180382 12628 180394 12630
rect 180610 12628 180616 12640
rect 180382 12600 180616 12628
rect 180382 12596 180394 12600
rect 180336 12590 180394 12596
rect 180610 12588 180616 12600
rect 180668 12588 180674 12640
rect 181438 12588 181444 12640
rect 181496 12628 181502 12640
rect 182268 12630 182326 12636
rect 182268 12628 182280 12630
rect 181496 12600 182280 12628
rect 181496 12588 181502 12600
rect 182268 12596 182280 12600
rect 182314 12596 182326 12630
rect 182268 12590 182326 12596
rect 187786 12588 187792 12640
rect 187844 12628 187850 12640
rect 188708 12630 188766 12636
rect 188708 12628 188720 12630
rect 187844 12600 188720 12628
rect 187844 12588 187850 12600
rect 188708 12596 188720 12600
rect 188754 12628 188766 12630
rect 188982 12628 188988 12640
rect 188754 12600 188988 12628
rect 188754 12596 188766 12600
rect 188708 12590 188766 12596
rect 188982 12588 188988 12600
rect 189040 12588 189046 12640
rect 190546 12628 190552 12640
rect 190506 12600 190552 12628
rect 190546 12588 190552 12600
rect 190604 12588 190610 12640
rect 191836 12630 191894 12636
rect 191836 12596 191848 12630
rect 191882 12628 191894 12630
rect 192018 12628 192024 12640
rect 191882 12600 192024 12628
rect 191882 12596 191894 12600
rect 191836 12590 191894 12596
rect 192018 12588 192024 12600
rect 192076 12588 192082 12640
rect 192110 12588 192116 12640
rect 192168 12628 192174 12640
rect 192588 12628 192616 12668
rect 192168 12600 192616 12628
rect 192168 12588 192174 12600
rect 193030 12588 193036 12640
rect 193088 12628 193094 12640
rect 194336 12628 194364 12668
rect 202138 12656 202144 12668
rect 202196 12696 202202 12708
rect 202616 12696 202644 12726
rect 202874 12724 202880 12736
rect 202932 12724 202938 12776
rect 202966 12724 202972 12776
rect 203024 12764 203030 12776
rect 204162 12764 204168 12776
rect 203024 12736 204168 12764
rect 203024 12724 203030 12736
rect 204162 12724 204168 12736
rect 204220 12724 204226 12776
rect 205082 12764 205088 12776
rect 205042 12736 205088 12764
rect 205082 12724 205088 12736
rect 205140 12724 205146 12776
rect 205174 12724 205180 12776
rect 205232 12764 205238 12776
rect 207492 12764 207520 12794
rect 205232 12736 207520 12764
rect 207584 12764 207612 12872
rect 210602 12860 210608 12912
rect 210660 12900 210666 12912
rect 219728 12900 219756 12940
rect 219802 12928 219808 12980
rect 219860 12968 219866 12980
rect 238202 12968 238208 12980
rect 219860 12940 238208 12968
rect 219860 12928 219866 12940
rect 228266 12900 228272 12912
rect 210660 12872 217364 12900
rect 219728 12872 228272 12900
rect 210660 12860 210666 12872
rect 207658 12792 207664 12844
rect 207716 12832 207722 12844
rect 210344 12832 210464 12836
rect 216582 12832 216588 12844
rect 207716 12808 216588 12832
rect 207716 12804 210372 12808
rect 210436 12804 216588 12808
rect 207716 12792 207722 12804
rect 216582 12792 216588 12804
rect 216640 12792 216646 12844
rect 217336 12832 217364 12872
rect 228266 12860 228272 12872
rect 228324 12860 228330 12912
rect 230382 12900 230388 12912
rect 229402 12872 230388 12900
rect 230382 12860 230388 12872
rect 230440 12860 230446 12912
rect 219802 12832 219808 12844
rect 217336 12804 219808 12832
rect 219802 12792 219808 12804
rect 219860 12792 219866 12844
rect 223666 12792 223672 12844
rect 223724 12832 223730 12844
rect 226704 12834 226762 12840
rect 226704 12832 226716 12834
rect 223724 12804 226716 12832
rect 223724 12792 223730 12804
rect 226704 12800 226716 12804
rect 226750 12800 226762 12834
rect 226704 12794 226762 12800
rect 226794 12792 226800 12844
rect 226852 12832 226858 12844
rect 227348 12834 227406 12840
rect 227348 12832 227360 12834
rect 226852 12804 227360 12832
rect 226852 12792 226858 12804
rect 227348 12800 227360 12804
rect 227394 12800 227406 12834
rect 227898 12832 227904 12844
rect 227858 12804 227904 12832
rect 227348 12794 227406 12800
rect 227898 12792 227904 12804
rect 227956 12792 227962 12844
rect 230290 12832 230296 12844
rect 230250 12804 230296 12832
rect 230290 12792 230296 12804
rect 230348 12792 230354 12844
rect 230768 12840 230796 12940
rect 238202 12928 238208 12940
rect 238260 12968 238266 12980
rect 251082 12968 251088 12980
rect 238260 12940 251088 12968
rect 238260 12928 238266 12940
rect 231026 12900 231032 12912
rect 230986 12872 231032 12900
rect 231026 12860 231032 12872
rect 231084 12860 231090 12912
rect 232314 12860 232320 12912
rect 232372 12900 232378 12912
rect 238294 12900 238300 12912
rect 232372 12872 238300 12900
rect 232372 12860 232378 12872
rect 238294 12860 238300 12872
rect 238352 12860 238358 12912
rect 238588 12900 238616 12940
rect 238496 12872 238616 12900
rect 238756 12902 238814 12908
rect 230752 12834 230810 12840
rect 230752 12800 230764 12834
rect 230798 12800 230810 12834
rect 233050 12832 233056 12844
rect 232162 12804 232728 12832
rect 233010 12804 233056 12832
rect 230752 12794 230810 12800
rect 227916 12764 227944 12792
rect 228176 12766 228234 12772
rect 228176 12764 228188 12766
rect 207584 12736 215294 12764
rect 205232 12724 205238 12736
rect 207290 12696 207296 12708
rect 202196 12668 202644 12696
rect 206480 12668 206784 12696
rect 207250 12668 207296 12696
rect 202196 12656 202202 12668
rect 193088 12600 194364 12628
rect 193088 12588 193094 12600
rect 194410 12588 194416 12640
rect 194468 12628 194474 12640
rect 195516 12630 195574 12636
rect 195516 12628 195528 12630
rect 194468 12600 195528 12628
rect 194468 12588 194474 12600
rect 195516 12596 195528 12600
rect 195562 12596 195574 12630
rect 195516 12590 195574 12596
rect 195974 12588 195980 12640
rect 196032 12628 196038 12640
rect 196988 12630 197046 12636
rect 196988 12628 197000 12630
rect 196032 12600 197000 12628
rect 196032 12588 196038 12600
rect 196988 12596 197000 12600
rect 197034 12596 197046 12630
rect 198182 12628 198188 12640
rect 198142 12600 198188 12628
rect 196988 12590 197046 12596
rect 198182 12588 198188 12600
rect 198240 12588 198246 12640
rect 201126 12628 201132 12640
rect 201086 12600 201132 12628
rect 201126 12588 201132 12600
rect 201184 12588 201190 12640
rect 201954 12588 201960 12640
rect 202012 12628 202018 12640
rect 204254 12628 204260 12640
rect 202012 12600 204260 12628
rect 202012 12588 202018 12600
rect 204254 12588 204260 12600
rect 204312 12588 204318 12640
rect 204348 12630 204406 12636
rect 204348 12596 204360 12630
rect 204394 12628 204406 12630
rect 204530 12628 204536 12640
rect 204394 12600 204536 12628
rect 204394 12596 204406 12600
rect 204348 12590 204406 12596
rect 204530 12588 204536 12600
rect 204588 12628 204594 12640
rect 205174 12628 205180 12640
rect 204588 12600 205180 12628
rect 204588 12588 204594 12600
rect 205174 12588 205180 12600
rect 205232 12588 205238 12640
rect 205266 12588 205272 12640
rect 205324 12628 205330 12640
rect 206480 12628 206508 12668
rect 205324 12600 206508 12628
rect 206756 12628 206784 12668
rect 207290 12656 207296 12668
rect 207348 12656 207354 12708
rect 210602 12628 210608 12640
rect 206756 12600 210608 12628
rect 205324 12588 205330 12600
rect 210602 12588 210608 12600
rect 210660 12588 210666 12640
rect 215266 12628 215294 12736
rect 219728 12736 227944 12764
rect 228008 12736 228188 12764
rect 219728 12628 219756 12736
rect 219802 12656 219808 12708
rect 219860 12696 219866 12708
rect 227164 12698 227222 12704
rect 219860 12668 227116 12696
rect 219860 12656 219866 12668
rect 215266 12600 219756 12628
rect 226520 12630 226578 12636
rect 226520 12596 226532 12630
rect 226566 12628 226578 12630
rect 226886 12628 226892 12640
rect 226566 12600 226892 12628
rect 226566 12596 226578 12600
rect 226520 12590 226578 12596
rect 226886 12588 226892 12600
rect 226944 12588 226950 12640
rect 227088 12628 227116 12668
rect 227164 12664 227176 12698
rect 227210 12696 227222 12698
rect 228008 12696 228036 12736
rect 228176 12732 228188 12736
rect 228222 12732 228234 12766
rect 228176 12726 228234 12732
rect 228266 12724 228272 12776
rect 228324 12764 228330 12776
rect 230198 12764 230204 12776
rect 228324 12736 230204 12764
rect 228324 12724 228330 12736
rect 230198 12724 230204 12736
rect 230256 12724 230262 12776
rect 232700 12764 232728 12804
rect 233050 12792 233056 12804
rect 233108 12792 233114 12844
rect 237006 12832 237012 12844
rect 236966 12804 237012 12832
rect 237006 12792 237012 12804
rect 237064 12792 237070 12844
rect 237652 12834 237710 12840
rect 237652 12800 237664 12834
rect 237698 12832 237710 12834
rect 238386 12832 238392 12844
rect 237698 12804 238392 12832
rect 237698 12800 237710 12804
rect 237652 12794 237710 12800
rect 238386 12792 238392 12804
rect 238444 12792 238450 12844
rect 238496 12840 238524 12872
rect 238756 12868 238768 12902
rect 238802 12900 238814 12902
rect 239030 12900 239036 12912
rect 238802 12872 239036 12900
rect 238802 12868 238814 12872
rect 238756 12862 238814 12868
rect 239030 12860 239036 12872
rect 239088 12860 239094 12912
rect 240042 12900 240048 12912
rect 239982 12872 240048 12900
rect 240042 12860 240048 12872
rect 240100 12860 240106 12912
rect 240704 12840 240732 12940
rect 251082 12928 251088 12940
rect 251140 12928 251146 12980
rect 252372 12970 252430 12976
rect 252372 12936 252384 12970
rect 252418 12968 252430 12970
rect 254670 12968 254676 12980
rect 252418 12940 254676 12968
rect 252418 12936 252430 12940
rect 252372 12930 252430 12936
rect 254670 12928 254676 12940
rect 254728 12928 254734 12980
rect 256234 12928 256240 12980
rect 256292 12968 256298 12980
rect 264606 12968 264612 12980
rect 256292 12940 263594 12968
rect 264566 12940 264612 12968
rect 256292 12928 256298 12940
rect 240962 12900 240968 12912
rect 240922 12872 240968 12900
rect 240962 12860 240968 12872
rect 241020 12860 241026 12912
rect 244642 12900 244648 12912
rect 244246 12872 244648 12900
rect 238480 12834 238538 12840
rect 238480 12800 238492 12834
rect 238526 12800 238538 12834
rect 238480 12794 238538 12800
rect 240688 12834 240746 12840
rect 240688 12800 240700 12834
rect 240734 12800 240746 12834
rect 240688 12794 240746 12800
rect 242066 12792 242072 12844
rect 242124 12792 242130 12844
rect 242250 12792 242256 12844
rect 242308 12832 242314 12844
rect 243816 12834 243874 12840
rect 243816 12832 243828 12834
rect 242308 12804 243828 12832
rect 242308 12792 242314 12804
rect 243816 12800 243828 12804
rect 243862 12832 243874 12834
rect 244246 12832 244274 12872
rect 244642 12860 244648 12872
rect 244700 12860 244706 12912
rect 244918 12860 244924 12912
rect 244976 12900 244982 12912
rect 245288 12902 245346 12908
rect 245288 12900 245300 12902
rect 244976 12872 245300 12900
rect 244976 12860 244982 12872
rect 245288 12868 245300 12872
rect 245334 12868 245346 12902
rect 245288 12862 245346 12868
rect 245378 12860 245384 12912
rect 245436 12900 245442 12912
rect 251360 12902 251418 12908
rect 251360 12900 251372 12902
rect 245436 12872 251372 12900
rect 245436 12860 245442 12872
rect 251360 12868 251372 12872
rect 251406 12900 251418 12902
rect 251634 12900 251640 12912
rect 251406 12872 251640 12900
rect 251406 12868 251418 12872
rect 251360 12862 251418 12868
rect 251634 12860 251640 12872
rect 251692 12860 251698 12912
rect 252462 12860 252468 12912
rect 252520 12900 252526 12912
rect 257246 12900 257252 12912
rect 252520 12872 252564 12900
rect 255162 12872 256740 12900
rect 252520 12860 252526 12872
rect 244550 12832 244556 12844
rect 243862 12804 244274 12832
rect 244510 12804 244556 12832
rect 243862 12800 243874 12804
rect 243816 12794 243874 12800
rect 244550 12792 244556 12804
rect 244608 12792 244614 12844
rect 244736 12834 244794 12840
rect 244736 12800 244748 12834
rect 244782 12832 244794 12834
rect 244826 12832 244832 12844
rect 244782 12804 244832 12832
rect 244782 12800 244794 12804
rect 244736 12794 244794 12800
rect 244826 12792 244832 12804
rect 244884 12832 244890 12844
rect 245196 12834 245254 12840
rect 245196 12832 245208 12834
rect 244884 12804 245208 12832
rect 244884 12792 244890 12804
rect 245196 12800 245208 12804
rect 245242 12800 245254 12834
rect 245196 12794 245254 12800
rect 250348 12834 250406 12840
rect 250348 12800 250360 12834
rect 250394 12832 250406 12834
rect 251174 12832 251180 12844
rect 250394 12804 251180 12832
rect 250394 12800 250406 12804
rect 250348 12794 250406 12800
rect 251146 12792 251180 12804
rect 251232 12792 251238 12844
rect 251542 12832 251548 12844
rect 251502 12804 251548 12832
rect 251542 12792 251548 12804
rect 251600 12792 251606 12844
rect 251652 12830 252416 12832
rect 252480 12830 252508 12860
rect 251652 12804 252508 12830
rect 233144 12766 233202 12772
rect 233144 12764 233156 12766
rect 230308 12736 232084 12764
rect 232700 12736 233156 12764
rect 230308 12696 230336 12736
rect 227210 12668 228036 12696
rect 229204 12668 230336 12696
rect 232056 12696 232084 12736
rect 233144 12732 233156 12736
rect 233190 12732 233202 12766
rect 251146 12764 251174 12792
rect 251652 12764 251680 12804
rect 252388 12802 252508 12804
rect 256236 12834 256294 12840
rect 256236 12800 256248 12834
rect 256282 12832 256294 12834
rect 256602 12832 256608 12844
rect 256282 12804 256608 12832
rect 256282 12800 256294 12804
rect 256236 12794 256294 12800
rect 256602 12792 256608 12804
rect 256660 12792 256666 12844
rect 233144 12726 233202 12732
rect 234586 12736 240548 12764
rect 234586 12696 234614 12736
rect 232056 12668 234614 12696
rect 237468 12698 237526 12704
rect 227210 12664 227222 12668
rect 227164 12658 227222 12664
rect 229204 12628 229232 12668
rect 237468 12664 237480 12698
rect 237514 12696 237526 12698
rect 237834 12696 237840 12708
rect 237514 12668 237840 12696
rect 237514 12664 237526 12668
rect 237468 12658 237526 12664
rect 237834 12656 237840 12668
rect 237892 12656 237898 12708
rect 237926 12656 237932 12708
rect 237984 12696 237990 12708
rect 237984 12668 238616 12696
rect 237984 12656 237990 12668
rect 227088 12600 229232 12628
rect 229554 12588 229560 12640
rect 229612 12628 229618 12640
rect 229648 12630 229706 12636
rect 229648 12628 229660 12630
rect 229612 12600 229660 12628
rect 229612 12588 229618 12600
rect 229648 12596 229660 12600
rect 229694 12596 229706 12630
rect 230106 12628 230112 12640
rect 230066 12600 230112 12628
rect 229648 12590 229706 12596
rect 230106 12588 230112 12600
rect 230164 12588 230170 12640
rect 230198 12588 230204 12640
rect 230256 12628 230262 12640
rect 232314 12628 232320 12640
rect 230256 12600 232320 12628
rect 230256 12588 230262 12600
rect 232314 12588 232320 12600
rect 232372 12588 232378 12640
rect 232498 12628 232504 12640
rect 232458 12600 232504 12628
rect 232498 12588 232504 12600
rect 232556 12628 232562 12640
rect 233142 12628 233148 12640
rect 232556 12600 233148 12628
rect 232556 12588 232562 12600
rect 233142 12588 233148 12600
rect 233200 12588 233206 12640
rect 236824 12630 236882 12636
rect 236824 12596 236836 12630
rect 236870 12628 236882 12630
rect 238478 12628 238484 12640
rect 236870 12600 238484 12628
rect 236870 12596 236882 12600
rect 236824 12590 236882 12596
rect 238478 12588 238484 12600
rect 238536 12588 238542 12640
rect 238588 12628 238616 12668
rect 238846 12628 238852 12640
rect 238588 12600 238852 12628
rect 238846 12588 238852 12600
rect 238904 12588 238910 12640
rect 239122 12588 239128 12640
rect 239180 12628 239186 12640
rect 240228 12630 240286 12636
rect 240228 12628 240240 12630
rect 239180 12600 240240 12628
rect 239180 12588 239186 12600
rect 240228 12596 240240 12600
rect 240274 12628 240286 12630
rect 240318 12628 240324 12640
rect 240274 12600 240324 12628
rect 240274 12596 240286 12600
rect 240228 12590 240286 12596
rect 240318 12588 240324 12600
rect 240376 12588 240382 12640
rect 240520 12628 240548 12736
rect 242084 12736 250300 12764
rect 251146 12736 251680 12764
rect 242084 12628 242112 12736
rect 242158 12656 242164 12708
rect 242216 12696 242222 12708
rect 242216 12668 244274 12696
rect 242216 12656 242222 12668
rect 242434 12628 242440 12640
rect 240520 12600 242112 12628
rect 242394 12600 242440 12628
rect 242434 12588 242440 12600
rect 242492 12588 242498 12640
rect 242894 12588 242900 12640
rect 242952 12628 242958 12640
rect 243908 12630 243966 12636
rect 243908 12628 243920 12630
rect 242952 12600 243920 12628
rect 242952 12588 242958 12600
rect 243908 12596 243920 12600
rect 243954 12596 243966 12630
rect 244246 12628 244274 12668
rect 244642 12656 244648 12708
rect 244700 12696 244706 12708
rect 248322 12696 248328 12708
rect 244700 12668 248328 12696
rect 244700 12656 244706 12668
rect 248322 12656 248328 12668
rect 248380 12656 248386 12708
rect 250162 12696 250168 12708
rect 250122 12668 250168 12696
rect 250162 12656 250168 12668
rect 250220 12656 250226 12708
rect 250272 12696 250300 12736
rect 252094 12724 252100 12776
rect 252152 12764 252158 12776
rect 252556 12766 252614 12772
rect 252556 12764 252568 12766
rect 252152 12736 252568 12764
rect 252152 12724 252158 12736
rect 252556 12732 252568 12736
rect 252602 12732 252614 12766
rect 252556 12726 252614 12732
rect 253658 12724 253664 12776
rect 253716 12764 253722 12776
rect 253716 12736 253760 12764
rect 253716 12724 253722 12736
rect 253934 12724 253940 12776
rect 253992 12764 253998 12776
rect 253992 12736 254036 12764
rect 253992 12724 253998 12736
rect 255130 12724 255136 12776
rect 255188 12764 255194 12776
rect 255408 12766 255466 12772
rect 255408 12764 255420 12766
rect 255188 12736 255420 12764
rect 255188 12724 255194 12736
rect 255408 12732 255420 12736
rect 255454 12764 255466 12766
rect 256326 12764 256332 12776
rect 255454 12736 256332 12764
rect 255454 12732 255466 12736
rect 255408 12726 255466 12732
rect 256326 12724 256332 12736
rect 256384 12724 256390 12776
rect 256418 12724 256424 12776
rect 256476 12764 256482 12776
rect 256476 12736 256520 12764
rect 256476 12724 256482 12736
rect 251818 12696 251824 12708
rect 250272 12668 251824 12696
rect 251818 12656 251824 12668
rect 251876 12656 251882 12708
rect 255038 12656 255044 12708
rect 255096 12696 255102 12708
rect 255868 12698 255926 12704
rect 255868 12696 255880 12698
rect 255096 12668 255880 12696
rect 255096 12656 255102 12668
rect 255868 12664 255880 12668
rect 255914 12664 255926 12698
rect 255868 12658 255926 12664
rect 251910 12628 251916 12640
rect 244246 12600 251916 12628
rect 243908 12590 243966 12596
rect 251910 12588 251916 12600
rect 251968 12588 251974 12640
rect 252002 12588 252008 12640
rect 252060 12628 252066 12640
rect 256712 12628 256740 12872
rect 257080 12872 257252 12900
rect 257080 12840 257108 12872
rect 257246 12860 257252 12872
rect 257304 12860 257310 12912
rect 261754 12900 261760 12912
rect 261666 12872 261760 12900
rect 261754 12860 261760 12872
rect 261812 12900 261818 12912
rect 263228 12902 263286 12908
rect 263228 12900 263240 12902
rect 261812 12872 263240 12900
rect 261812 12860 261818 12872
rect 263228 12868 263240 12872
rect 263274 12868 263286 12902
rect 263228 12862 263286 12868
rect 263318 12860 263324 12912
rect 263376 12900 263382 12912
rect 263412 12902 263470 12908
rect 263412 12900 263424 12902
rect 263376 12872 263424 12900
rect 263376 12860 263382 12872
rect 263412 12868 263424 12872
rect 263458 12868 263470 12902
rect 263566 12900 263594 12940
rect 264606 12928 264612 12940
rect 264664 12928 264670 12980
rect 268378 12968 268384 12980
rect 265268 12940 268384 12968
rect 265268 12900 265296 12940
rect 268378 12928 268384 12940
rect 268436 12928 268442 12980
rect 302602 12968 302608 12980
rect 268488 12940 296714 12968
rect 302562 12940 302608 12968
rect 265526 12900 265532 12912
rect 263566 12872 265296 12900
rect 265486 12872 265532 12900
rect 263412 12862 263470 12868
rect 257064 12834 257122 12840
rect 257064 12800 257076 12834
rect 257110 12800 257122 12834
rect 257064 12794 257122 12800
rect 261846 12792 261852 12844
rect 261904 12832 261910 12844
rect 262492 12834 262550 12840
rect 262492 12832 262504 12834
rect 261904 12804 262504 12832
rect 261904 12792 261910 12804
rect 262492 12800 262504 12804
rect 262538 12800 262550 12834
rect 262492 12794 262550 12800
rect 264148 12834 264206 12840
rect 264148 12800 264160 12834
rect 264194 12832 264206 12834
rect 264330 12832 264336 12844
rect 264194 12804 264336 12832
rect 264194 12800 264206 12804
rect 264148 12794 264206 12800
rect 264330 12792 264336 12804
rect 264388 12792 264394 12844
rect 264422 12792 264428 12844
rect 264480 12832 264486 12844
rect 265268 12840 265296 12872
rect 265526 12860 265532 12872
rect 265584 12860 265590 12912
rect 266538 12860 266544 12912
rect 266596 12860 266602 12912
rect 268488 12900 268516 12940
rect 271046 12900 271052 12912
rect 266832 12872 268516 12900
rect 270618 12872 271052 12900
rect 264792 12834 264850 12840
rect 264792 12832 264804 12834
rect 264480 12804 264804 12832
rect 264480 12792 264486 12804
rect 264792 12800 264804 12804
rect 264838 12800 264850 12834
rect 264792 12794 264850 12800
rect 265252 12834 265310 12840
rect 265252 12800 265264 12834
rect 265298 12800 265310 12834
rect 265252 12794 265310 12800
rect 257154 12724 257160 12776
rect 257212 12764 257218 12776
rect 262306 12764 262312 12776
rect 257212 12736 262312 12764
rect 257212 12724 257218 12736
rect 262306 12724 262312 12736
rect 262364 12724 262370 12776
rect 266832 12764 266860 12872
rect 271046 12860 271052 12872
rect 271104 12860 271110 12912
rect 271782 12900 271788 12912
rect 271694 12872 271788 12900
rect 271782 12860 271788 12872
rect 271840 12900 271846 12912
rect 272794 12900 272800 12912
rect 271840 12872 272800 12900
rect 271840 12860 271846 12872
rect 272794 12860 272800 12872
rect 272852 12860 272858 12912
rect 272888 12902 272946 12908
rect 272888 12868 272900 12902
rect 272934 12900 272946 12902
rect 273162 12900 273168 12912
rect 272934 12872 273168 12900
rect 272934 12868 272946 12872
rect 272888 12862 272946 12868
rect 273162 12860 273168 12872
rect 273220 12860 273226 12912
rect 295886 12900 295892 12912
rect 282886 12872 295892 12900
rect 267828 12834 267886 12840
rect 267828 12800 267840 12834
rect 267874 12832 267886 12834
rect 268286 12832 268292 12844
rect 267874 12804 268292 12832
rect 267874 12800 267886 12804
rect 267828 12794 267886 12800
rect 268286 12792 268292 12804
rect 268344 12832 268350 12844
rect 269022 12832 269028 12844
rect 268344 12804 269028 12832
rect 268344 12792 268350 12804
rect 269022 12792 269028 12804
rect 269080 12792 269086 12844
rect 269116 12834 269174 12840
rect 269116 12800 269128 12834
rect 269162 12800 269174 12834
rect 269116 12794 269174 12800
rect 263428 12736 266860 12764
rect 257062 12656 257068 12708
rect 257120 12696 257126 12708
rect 262674 12696 262680 12708
rect 257120 12668 262536 12696
rect 262634 12668 262680 12696
rect 257120 12656 257126 12668
rect 257156 12630 257214 12636
rect 257156 12628 257168 12630
rect 252060 12600 252104 12628
rect 256712 12600 257168 12628
rect 252060 12588 252066 12600
rect 257156 12596 257168 12600
rect 257202 12596 257214 12630
rect 257156 12590 257214 12596
rect 261848 12630 261906 12636
rect 261848 12596 261860 12630
rect 261894 12628 261906 12630
rect 262214 12628 262220 12640
rect 261894 12600 262220 12628
rect 261894 12596 261906 12600
rect 261848 12590 261906 12596
rect 262214 12588 262220 12600
rect 262272 12588 262278 12640
rect 262508 12628 262536 12668
rect 262674 12656 262680 12668
rect 262732 12656 262738 12708
rect 263428 12628 263456 12736
rect 266998 12724 267004 12776
rect 267056 12764 267062 12776
rect 267550 12764 267556 12776
rect 267056 12736 267556 12764
rect 267056 12724 267062 12736
rect 267550 12724 267556 12736
rect 267608 12764 267614 12776
rect 267920 12766 267978 12772
rect 267920 12764 267932 12766
rect 267608 12736 267932 12764
rect 267608 12724 267614 12736
rect 267920 12732 267932 12736
rect 267966 12732 267978 12766
rect 267920 12726 267978 12732
rect 268010 12724 268016 12776
rect 268068 12764 268074 12776
rect 268068 12736 268112 12764
rect 268068 12724 268074 12736
rect 268378 12724 268384 12776
rect 268436 12764 268442 12776
rect 269132 12764 269160 12794
rect 270862 12792 270868 12844
rect 270920 12832 270926 12844
rect 271692 12834 271750 12840
rect 271692 12832 271704 12834
rect 270920 12804 271704 12832
rect 270920 12792 270926 12804
rect 271692 12800 271704 12804
rect 271738 12832 271750 12834
rect 272610 12832 272616 12844
rect 271738 12804 272616 12832
rect 271738 12800 271750 12804
rect 271692 12794 271750 12800
rect 272610 12792 272616 12804
rect 272668 12792 272674 12844
rect 282886 12832 282914 12872
rect 295886 12860 295892 12872
rect 295944 12860 295950 12912
rect 296686 12900 296714 12940
rect 302602 12928 302608 12940
rect 302660 12928 302666 12980
rect 304444 12970 304502 12976
rect 304444 12936 304456 12970
rect 304490 12968 304502 12970
rect 305362 12968 305368 12980
rect 304490 12940 305368 12968
rect 304490 12936 304502 12940
rect 304444 12930 304502 12936
rect 305362 12928 305368 12940
rect 305420 12928 305426 12980
rect 304994 12900 305000 12912
rect 296686 12872 304672 12900
rect 304954 12872 305000 12900
rect 290274 12832 290280 12844
rect 272720 12804 282914 12832
rect 287026 12804 290280 12832
rect 269390 12764 269396 12776
rect 268436 12736 269160 12764
rect 269350 12736 269396 12764
rect 268436 12724 268442 12736
rect 269390 12724 269396 12736
rect 269448 12724 269454 12776
rect 271968 12766 272026 12772
rect 270880 12736 271460 12764
rect 263502 12656 263508 12708
rect 263560 12696 263566 12708
rect 270880 12696 270908 12736
rect 263560 12668 264100 12696
rect 263560 12656 263566 12668
rect 263962 12628 263968 12640
rect 262508 12600 263456 12628
rect 263922 12600 263968 12628
rect 263962 12588 263968 12600
rect 264020 12588 264026 12640
rect 264072 12628 264100 12668
rect 266556 12668 269252 12696
rect 266556 12628 266584 12668
rect 266998 12628 267004 12640
rect 264072 12600 266584 12628
rect 266958 12600 267004 12628
rect 266998 12588 267004 12600
rect 267056 12588 267062 12640
rect 267090 12588 267096 12640
rect 267148 12628 267154 12640
rect 267460 12630 267518 12636
rect 267460 12628 267472 12630
rect 267148 12600 267472 12628
rect 267148 12588 267154 12600
rect 267460 12596 267472 12600
rect 267506 12596 267518 12630
rect 267460 12590 267518 12596
rect 267550 12588 267556 12640
rect 267608 12628 267614 12640
rect 269114 12628 269120 12640
rect 267608 12600 269120 12628
rect 267608 12588 267614 12600
rect 269114 12588 269120 12600
rect 269172 12588 269178 12640
rect 269224 12628 269252 12668
rect 270420 12668 270908 12696
rect 271432 12696 271460 12736
rect 271968 12732 271980 12766
rect 272014 12764 272026 12766
rect 272242 12764 272248 12776
rect 272014 12736 272248 12764
rect 272014 12732 272026 12736
rect 271968 12726 272026 12732
rect 272242 12724 272248 12736
rect 272300 12724 272306 12776
rect 272720 12696 272748 12804
rect 272886 12724 272892 12776
rect 272944 12764 272950 12776
rect 272980 12766 273038 12772
rect 272980 12764 272992 12766
rect 272944 12736 272992 12764
rect 272944 12724 272950 12736
rect 272980 12732 272992 12736
rect 273026 12732 273038 12766
rect 272980 12726 273038 12732
rect 273072 12766 273130 12772
rect 273072 12732 273084 12766
rect 273118 12732 273130 12766
rect 273072 12726 273130 12732
rect 271432 12668 272748 12696
rect 270420 12628 270448 12668
rect 272794 12656 272800 12708
rect 272852 12696 272858 12708
rect 273088 12696 273116 12726
rect 273162 12724 273168 12776
rect 273220 12764 273226 12776
rect 287026 12764 287054 12804
rect 290274 12792 290280 12804
rect 290332 12792 290338 12844
rect 302786 12832 302792 12844
rect 302746 12804 302792 12832
rect 302786 12792 302792 12804
rect 302844 12792 302850 12844
rect 304644 12840 304672 12872
rect 304994 12860 305000 12872
rect 305052 12900 305058 12912
rect 305454 12900 305460 12912
rect 305052 12872 305460 12900
rect 305052 12860 305058 12872
rect 305454 12860 305460 12872
rect 305512 12860 305518 12912
rect 304628 12834 304686 12840
rect 304628 12800 304640 12834
rect 304674 12800 304686 12834
rect 304628 12794 304686 12800
rect 273220 12736 287054 12764
rect 273220 12724 273226 12736
rect 272852 12668 273116 12696
rect 272852 12656 272858 12668
rect 270862 12628 270868 12640
rect 269224 12600 270448 12628
rect 270822 12600 270868 12628
rect 270862 12588 270868 12600
rect 270920 12588 270926 12640
rect 271138 12588 271144 12640
rect 271196 12628 271202 12640
rect 271324 12630 271382 12636
rect 271324 12628 271336 12630
rect 271196 12600 271336 12628
rect 271196 12588 271202 12600
rect 271324 12596 271336 12600
rect 271370 12596 271382 12630
rect 272518 12628 272524 12640
rect 272478 12600 272524 12628
rect 271324 12590 271382 12596
rect 272518 12588 272524 12600
rect 272576 12588 272582 12640
rect 272610 12588 272616 12640
rect 272668 12628 272674 12640
rect 281074 12628 281080 12640
rect 272668 12600 281080 12628
rect 272668 12588 272674 12600
rect 281074 12588 281080 12600
rect 281132 12588 281138 12640
rect 1104 12538 305808 12560
rect 1104 12486 39048 12538
rect 39100 12486 39112 12538
rect 39164 12486 39176 12538
rect 39228 12486 39240 12538
rect 39292 12486 39304 12538
rect 39356 12486 115246 12538
rect 115298 12486 115310 12538
rect 115362 12486 115374 12538
rect 115426 12486 115438 12538
rect 115490 12486 115502 12538
rect 115554 12486 191444 12538
rect 191496 12486 191508 12538
rect 191560 12486 191572 12538
rect 191624 12486 191636 12538
rect 191688 12486 191700 12538
rect 191752 12486 267642 12538
rect 267694 12486 267706 12538
rect 267758 12486 267770 12538
rect 267822 12486 267834 12538
rect 267886 12486 267898 12538
rect 267950 12486 305808 12538
rect 1104 12464 305808 12486
rect 26970 12384 26976 12436
rect 27028 12424 27034 12436
rect 28074 12424 28080 12436
rect 27028 12396 28080 12424
rect 27028 12384 27034 12396
rect 28074 12384 28080 12396
rect 28132 12424 28138 12436
rect 28132 12396 28488 12424
rect 28132 12384 28138 12396
rect 14274 12316 14280 12368
rect 14332 12356 14338 12368
rect 28460 12356 28488 12396
rect 28810 12384 28816 12436
rect 28868 12424 28874 12436
rect 31296 12426 31354 12432
rect 31296 12424 31308 12426
rect 28868 12396 31308 12424
rect 28868 12384 28874 12396
rect 31296 12392 31308 12396
rect 31342 12392 31354 12426
rect 31296 12386 31354 12392
rect 32582 12384 32588 12436
rect 32640 12424 32646 12436
rect 33964 12426 34022 12432
rect 32640 12396 33088 12424
rect 32640 12384 32646 12396
rect 33060 12356 33088 12396
rect 33964 12392 33976 12426
rect 34010 12424 34022 12426
rect 34514 12424 34520 12436
rect 34010 12396 34520 12424
rect 34010 12392 34022 12396
rect 33964 12386 34022 12392
rect 34514 12384 34520 12396
rect 34572 12384 34578 12436
rect 34792 12426 34850 12432
rect 34792 12392 34804 12426
rect 34838 12424 34850 12426
rect 35986 12424 35992 12436
rect 34838 12396 35992 12424
rect 34838 12392 34850 12396
rect 34792 12386 34850 12392
rect 35986 12384 35992 12396
rect 36044 12384 36050 12436
rect 37184 12426 37242 12432
rect 37184 12392 37196 12426
rect 37230 12392 37242 12426
rect 37184 12386 37242 12392
rect 34882 12356 34888 12368
rect 14332 12328 28396 12356
rect 28460 12328 28948 12356
rect 33060 12328 34888 12356
rect 14332 12316 14338 12328
rect 26878 12288 26884 12300
rect 16960 12260 26884 12288
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 16960 12084 16988 12260
rect 26878 12248 26884 12260
rect 26936 12248 26942 12300
rect 27708 12290 27766 12296
rect 27708 12256 27720 12290
rect 27754 12288 27766 12290
rect 28074 12288 28080 12300
rect 27754 12260 28080 12288
rect 27754 12256 27766 12260
rect 27708 12250 27766 12256
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 28368 12288 28396 12328
rect 28718 12288 28724 12300
rect 28368 12260 28724 12288
rect 28718 12248 28724 12260
rect 28776 12248 28782 12300
rect 28920 12296 28948 12328
rect 34882 12316 34888 12328
rect 34940 12356 34946 12368
rect 37200 12356 37228 12386
rect 37826 12384 37832 12436
rect 37884 12424 37890 12436
rect 38472 12426 38530 12432
rect 38472 12424 38484 12426
rect 37884 12396 38484 12424
rect 37884 12384 37890 12396
rect 38472 12392 38484 12396
rect 38518 12392 38530 12426
rect 38472 12386 38530 12392
rect 38930 12384 38936 12436
rect 38988 12424 38994 12436
rect 39208 12426 39266 12432
rect 39208 12424 39220 12426
rect 38988 12396 39220 12424
rect 38988 12384 38994 12396
rect 39208 12392 39220 12396
rect 39254 12392 39266 12426
rect 39208 12386 39266 12392
rect 39390 12384 39396 12436
rect 39448 12424 39454 12436
rect 40954 12424 40960 12436
rect 39448 12396 40960 12424
rect 39448 12384 39454 12396
rect 40954 12384 40960 12396
rect 41012 12384 41018 12436
rect 43162 12424 43168 12436
rect 41524 12396 43024 12424
rect 43122 12396 43168 12424
rect 41524 12356 41552 12396
rect 34940 12328 37228 12356
rect 37292 12328 41552 12356
rect 42996 12356 43024 12396
rect 43162 12384 43168 12396
rect 43220 12384 43226 12436
rect 43806 12424 43812 12436
rect 43766 12396 43812 12424
rect 43806 12384 43812 12396
rect 43864 12384 43870 12436
rect 54018 12384 54024 12436
rect 54076 12424 54082 12436
rect 54112 12426 54170 12432
rect 54112 12424 54124 12426
rect 54076 12396 54124 12424
rect 54076 12384 54082 12396
rect 54112 12392 54124 12396
rect 54158 12392 54170 12426
rect 54112 12386 54170 12392
rect 54664 12426 54722 12432
rect 54664 12392 54676 12426
rect 54710 12424 54722 12426
rect 55490 12424 55496 12436
rect 54710 12396 55496 12424
rect 54710 12392 54722 12396
rect 54664 12386 54722 12392
rect 55490 12384 55496 12396
rect 55548 12384 55554 12436
rect 56686 12384 56692 12436
rect 56744 12424 56750 12436
rect 57332 12426 57390 12432
rect 57332 12424 57344 12426
rect 56744 12396 57344 12424
rect 56744 12384 56750 12396
rect 57332 12392 57344 12396
rect 57378 12392 57390 12426
rect 57974 12424 57980 12436
rect 57934 12396 57980 12424
rect 57332 12386 57390 12392
rect 57974 12384 57980 12396
rect 58032 12384 58038 12436
rect 75086 12384 75092 12436
rect 75144 12424 75150 12436
rect 75180 12426 75238 12432
rect 75180 12424 75192 12426
rect 75144 12396 75192 12424
rect 75144 12384 75150 12396
rect 75180 12392 75192 12396
rect 75226 12392 75238 12426
rect 79318 12424 79324 12436
rect 75180 12386 75238 12392
rect 75288 12396 78536 12424
rect 79278 12396 79324 12424
rect 43714 12356 43720 12368
rect 42996 12328 43720 12356
rect 34940 12316 34946 12328
rect 28904 12290 28962 12296
rect 28904 12256 28916 12290
rect 28950 12288 28962 12290
rect 28994 12288 29000 12300
rect 28950 12260 29000 12288
rect 28950 12256 28962 12260
rect 28904 12250 28962 12256
rect 28994 12248 29000 12260
rect 29052 12248 29058 12300
rect 29546 12288 29552 12300
rect 29458 12260 29552 12288
rect 29546 12248 29552 12260
rect 29604 12288 29610 12300
rect 31756 12290 31814 12296
rect 31756 12288 31768 12290
rect 29604 12260 31768 12288
rect 29604 12248 29610 12260
rect 31756 12256 31768 12260
rect 31802 12288 31814 12290
rect 31802 12260 35572 12288
rect 31802 12256 31814 12260
rect 31756 12250 31814 12256
rect 17034 12180 17040 12232
rect 17092 12220 17098 12232
rect 17092 12192 22094 12220
rect 17092 12180 17098 12192
rect 22066 12152 22094 12192
rect 27080 12192 27384 12220
rect 27080 12152 27108 12192
rect 22066 12124 27108 12152
rect 27356 12152 27384 12192
rect 27430 12180 27436 12232
rect 27488 12220 27494 12232
rect 28628 12222 28686 12228
rect 28628 12220 28640 12222
rect 27488 12192 27532 12220
rect 28000 12192 28640 12220
rect 27488 12180 27494 12192
rect 28000 12152 28028 12192
rect 28628 12188 28640 12192
rect 28674 12220 28686 12222
rect 29362 12220 29368 12232
rect 28674 12192 29368 12220
rect 28674 12188 28686 12192
rect 28628 12182 28686 12188
rect 29362 12180 29368 12192
rect 29420 12180 29426 12232
rect 34146 12220 34152 12232
rect 34106 12192 34152 12220
rect 34146 12180 34152 12192
rect 34204 12180 34210 12232
rect 34698 12220 34704 12232
rect 34610 12192 34704 12220
rect 34698 12180 34704 12192
rect 34756 12220 34762 12232
rect 35342 12220 35348 12232
rect 34756 12192 35348 12220
rect 34756 12180 34762 12192
rect 35342 12180 35348 12192
rect 35400 12180 35406 12232
rect 29454 12152 29460 12164
rect 27356 12124 28028 12152
rect 28276 12124 29460 12152
rect 27062 12084 27068 12096
rect 4856 12056 16988 12084
rect 27022 12056 27068 12084
rect 4856 12044 4862 12056
rect 27062 12044 27068 12056
rect 27120 12044 27126 12096
rect 27154 12044 27160 12096
rect 27212 12084 27218 12096
rect 27524 12086 27582 12092
rect 27524 12084 27536 12086
rect 27212 12056 27536 12084
rect 27212 12044 27218 12056
rect 27524 12052 27536 12056
rect 27570 12084 27582 12086
rect 27982 12084 27988 12096
rect 27570 12056 27988 12084
rect 27570 12052 27582 12056
rect 27524 12046 27582 12052
rect 27982 12044 27988 12056
rect 28040 12044 28046 12096
rect 28276 12092 28304 12124
rect 29454 12112 29460 12124
rect 29512 12112 29518 12164
rect 29822 12152 29828 12164
rect 29782 12124 29828 12152
rect 29822 12112 29828 12124
rect 29880 12112 29886 12164
rect 31202 12152 31208 12164
rect 31050 12124 31208 12152
rect 31202 12112 31208 12124
rect 31260 12112 31266 12164
rect 32030 12152 32036 12164
rect 31990 12124 32036 12152
rect 32030 12112 32036 12124
rect 32088 12112 32094 12164
rect 35436 12154 35494 12160
rect 35436 12152 35448 12154
rect 33258 12124 35448 12152
rect 35436 12120 35448 12124
rect 35482 12120 35494 12154
rect 35544 12152 35572 12260
rect 36356 12222 36414 12228
rect 36356 12188 36368 12222
rect 36402 12220 36414 12222
rect 37092 12222 37150 12228
rect 37092 12220 37104 12222
rect 36402 12192 37104 12220
rect 36402 12188 36414 12192
rect 36356 12182 36414 12188
rect 37092 12188 37104 12192
rect 37138 12220 37150 12222
rect 37292 12220 37320 12328
rect 43714 12316 43720 12328
rect 43772 12316 43778 12368
rect 75288 12356 75316 12396
rect 53668 12328 75316 12356
rect 40864 12290 40922 12296
rect 40864 12256 40876 12290
rect 40910 12288 40922 12290
rect 40954 12288 40960 12300
rect 40910 12260 40960 12288
rect 40910 12256 40922 12260
rect 40864 12250 40922 12256
rect 40954 12248 40960 12260
rect 41012 12248 41018 12300
rect 52364 12290 52422 12296
rect 52364 12288 52376 12290
rect 41432 12260 52376 12288
rect 37138 12192 37320 12220
rect 37138 12188 37150 12192
rect 37092 12182 37150 12188
rect 38010 12180 38016 12232
rect 38068 12220 38074 12232
rect 38656 12222 38714 12228
rect 38656 12220 38668 12222
rect 38068 12192 38668 12220
rect 38068 12180 38074 12192
rect 38656 12188 38668 12192
rect 38702 12188 38714 12222
rect 38656 12182 38714 12188
rect 39116 12222 39174 12228
rect 39116 12188 39128 12222
rect 39162 12220 39174 12222
rect 40310 12220 40316 12232
rect 39162 12192 40316 12220
rect 39162 12188 39174 12192
rect 39116 12182 39174 12188
rect 40310 12180 40316 12192
rect 40368 12180 40374 12232
rect 40586 12220 40592 12232
rect 40546 12192 40592 12220
rect 40586 12180 40592 12192
rect 40644 12180 40650 12232
rect 41432 12228 41460 12260
rect 52364 12256 52376 12260
rect 52410 12288 52422 12290
rect 53668 12288 53696 12328
rect 76006 12316 76012 12368
rect 76064 12356 76070 12368
rect 77202 12356 77208 12368
rect 76064 12328 77208 12356
rect 76064 12316 76070 12328
rect 52410 12260 53696 12288
rect 52410 12256 52422 12260
rect 52364 12250 52422 12256
rect 53834 12248 53840 12300
rect 53892 12248 53898 12300
rect 55676 12290 55734 12296
rect 55676 12288 55688 12290
rect 55186 12260 55688 12288
rect 41416 12222 41474 12228
rect 41416 12188 41428 12222
rect 41462 12188 41474 12222
rect 43714 12220 43720 12232
rect 43674 12192 43720 12220
rect 41416 12182 41474 12188
rect 41432 12152 41460 12182
rect 43714 12180 43720 12192
rect 43772 12220 43778 12232
rect 53852 12220 53880 12248
rect 54572 12222 54630 12228
rect 54572 12220 54584 12222
rect 43772 12192 48314 12220
rect 53852 12192 54584 12220
rect 43772 12180 43778 12192
rect 35544 12124 41460 12152
rect 35436 12114 35494 12120
rect 41598 12112 41604 12164
rect 41656 12152 41662 12164
rect 41692 12154 41750 12160
rect 41692 12152 41704 12154
rect 41656 12124 41704 12152
rect 41656 12112 41662 12124
rect 41692 12120 41704 12124
rect 41738 12120 41750 12154
rect 41692 12114 41750 12120
rect 41782 12112 41788 12164
rect 41840 12152 41846 12164
rect 41840 12124 42182 12152
rect 41840 12112 41846 12124
rect 28260 12086 28318 12092
rect 28260 12052 28272 12086
rect 28306 12052 28318 12086
rect 28260 12046 28318 12052
rect 28902 12044 28908 12096
rect 28960 12084 28966 12096
rect 31110 12084 31116 12096
rect 28960 12056 31116 12084
rect 28960 12044 28966 12056
rect 31110 12044 31116 12056
rect 31168 12044 31174 12096
rect 32306 12044 32312 12096
rect 32364 12084 32370 12096
rect 32950 12084 32956 12096
rect 32364 12056 32956 12084
rect 32364 12044 32370 12056
rect 32950 12044 32956 12056
rect 33008 12084 33014 12096
rect 33504 12086 33562 12092
rect 33504 12084 33516 12086
rect 33008 12056 33516 12084
rect 33008 12044 33014 12056
rect 33504 12052 33516 12056
rect 33550 12052 33562 12086
rect 36446 12084 36452 12096
rect 36406 12056 36452 12084
rect 33504 12046 33562 12052
rect 36446 12044 36452 12056
rect 36504 12044 36510 12096
rect 40220 12086 40278 12092
rect 40220 12052 40232 12086
rect 40266 12084 40278 12086
rect 40494 12084 40500 12096
rect 40266 12056 40500 12084
rect 40266 12052 40278 12056
rect 40220 12046 40278 12052
rect 40494 12044 40500 12056
rect 40552 12044 40558 12096
rect 40678 12084 40684 12096
rect 40638 12056 40684 12084
rect 40678 12044 40684 12056
rect 40736 12044 40742 12096
rect 48286 12084 48314 12192
rect 54572 12188 54584 12192
rect 54618 12220 54630 12222
rect 55186 12220 55214 12260
rect 55676 12256 55688 12260
rect 55722 12256 55734 12290
rect 55676 12250 55734 12256
rect 56410 12248 56416 12300
rect 56468 12288 56474 12300
rect 56688 12290 56746 12296
rect 56688 12288 56700 12290
rect 56468 12260 56700 12288
rect 56468 12248 56474 12260
rect 56688 12256 56700 12260
rect 56734 12256 56746 12290
rect 56688 12250 56746 12256
rect 74810 12248 74816 12300
rect 74868 12288 74874 12300
rect 76760 12296 76788 12328
rect 77202 12316 77208 12328
rect 77260 12316 77266 12368
rect 77480 12358 77538 12364
rect 77480 12324 77492 12358
rect 77526 12356 77538 12358
rect 78398 12356 78404 12368
rect 77526 12328 78404 12356
rect 77526 12324 77538 12328
rect 77480 12318 77538 12324
rect 78398 12316 78404 12328
rect 78456 12316 78462 12368
rect 76744 12290 76802 12296
rect 74868 12260 76696 12288
rect 74868 12248 74874 12260
rect 54618 12192 55214 12220
rect 54618 12188 54630 12192
rect 54572 12182 54630 12188
rect 55306 12180 55312 12232
rect 55364 12220 55370 12232
rect 56502 12220 56508 12232
rect 55364 12192 56508 12220
rect 55364 12180 55370 12192
rect 56502 12180 56508 12192
rect 56560 12220 56566 12232
rect 76668 12228 76696 12260
rect 76744 12256 76756 12290
rect 76790 12256 76802 12290
rect 76744 12250 76802 12256
rect 76926 12248 76932 12300
rect 76984 12288 76990 12300
rect 78122 12288 78128 12300
rect 76984 12260 78128 12288
rect 76984 12248 76990 12260
rect 78122 12248 78128 12260
rect 78180 12248 78186 12300
rect 56596 12222 56654 12228
rect 56596 12220 56608 12222
rect 56560 12192 56608 12220
rect 56560 12180 56566 12192
rect 56596 12188 56608 12192
rect 56642 12220 56654 12222
rect 57516 12222 57574 12228
rect 57516 12220 57528 12222
rect 56642 12192 57528 12220
rect 56642 12188 56654 12192
rect 56596 12182 56654 12188
rect 57516 12188 57528 12192
rect 57562 12188 57574 12222
rect 57516 12182 57574 12188
rect 58160 12222 58218 12228
rect 58160 12188 58172 12222
rect 58206 12188 58218 12222
rect 58160 12182 58218 12188
rect 75364 12222 75422 12228
rect 75364 12188 75376 12222
rect 75410 12220 75422 12222
rect 76652 12222 76710 12228
rect 75410 12192 76604 12220
rect 75410 12188 75422 12192
rect 75364 12182 75422 12188
rect 52638 12152 52644 12164
rect 52598 12124 52644 12152
rect 52638 12112 52644 12124
rect 52696 12112 52702 12164
rect 53098 12112 53104 12164
rect 53156 12112 53162 12164
rect 55492 12154 55550 12160
rect 53944 12124 55214 12152
rect 53944 12084 53972 12124
rect 48286 12056 53972 12084
rect 55186 12084 55214 12124
rect 55492 12120 55504 12154
rect 55538 12152 55550 12154
rect 58176 12152 58204 12182
rect 55538 12124 56088 12152
rect 55538 12120 55550 12124
rect 55492 12114 55550 12120
rect 56060 12096 56088 12124
rect 56152 12124 58204 12152
rect 76576 12152 76604 12192
rect 76652 12188 76664 12222
rect 76698 12220 76710 12222
rect 77938 12220 77944 12232
rect 76698 12192 77944 12220
rect 76698 12188 76710 12192
rect 76652 12182 76710 12188
rect 77938 12180 77944 12192
rect 77996 12180 78002 12232
rect 78508 12152 78536 12396
rect 79318 12384 79324 12396
rect 79376 12384 79382 12436
rect 80240 12426 80298 12432
rect 80240 12392 80252 12426
rect 80286 12424 80298 12426
rect 80514 12424 80520 12436
rect 80286 12396 80520 12424
rect 80286 12392 80298 12396
rect 80240 12386 80298 12392
rect 80514 12384 80520 12396
rect 80572 12384 80578 12436
rect 85482 12384 85488 12436
rect 85540 12424 85546 12436
rect 85576 12426 85634 12432
rect 85576 12424 85588 12426
rect 85540 12396 85588 12424
rect 85540 12384 85546 12396
rect 85576 12392 85588 12396
rect 85622 12392 85634 12426
rect 86402 12424 86408 12436
rect 86362 12396 86408 12424
rect 85576 12386 85634 12392
rect 86402 12384 86408 12396
rect 86460 12384 86466 12436
rect 87874 12384 87880 12436
rect 87932 12424 87938 12436
rect 88888 12426 88946 12432
rect 88888 12424 88900 12426
rect 87932 12396 88900 12424
rect 87932 12384 87938 12396
rect 88888 12392 88900 12396
rect 88934 12392 88946 12426
rect 90174 12424 90180 12436
rect 90134 12396 90180 12424
rect 88888 12386 88946 12392
rect 90174 12384 90180 12396
rect 90232 12384 90238 12436
rect 99100 12426 99158 12432
rect 99100 12392 99112 12426
rect 99146 12424 99158 12426
rect 99466 12424 99472 12436
rect 99146 12396 99472 12424
rect 99146 12392 99158 12396
rect 99100 12386 99158 12392
rect 99466 12384 99472 12396
rect 99524 12384 99530 12436
rect 99836 12426 99894 12432
rect 99836 12392 99848 12426
rect 99882 12424 99894 12426
rect 99926 12424 99932 12436
rect 99882 12396 99932 12424
rect 99882 12392 99894 12396
rect 99836 12386 99894 12392
rect 99926 12384 99932 12396
rect 99984 12384 99990 12436
rect 103884 12426 103942 12432
rect 103884 12392 103896 12426
rect 103930 12424 103942 12426
rect 104986 12424 104992 12436
rect 103930 12396 104992 12424
rect 103930 12392 103942 12396
rect 103884 12386 103942 12392
rect 104986 12384 104992 12396
rect 105044 12384 105050 12436
rect 105170 12424 105176 12436
rect 105130 12396 105176 12424
rect 105170 12384 105176 12396
rect 105228 12384 105234 12436
rect 112530 12384 112536 12436
rect 112588 12424 112594 12436
rect 113084 12426 113142 12432
rect 113084 12424 113096 12426
rect 112588 12396 113096 12424
rect 112588 12384 112594 12396
rect 113084 12392 113096 12396
rect 113130 12392 113142 12426
rect 113084 12386 113142 12392
rect 113728 12426 113786 12432
rect 113728 12392 113740 12426
rect 113774 12424 113786 12426
rect 115014 12424 115020 12436
rect 113774 12396 115020 12424
rect 113774 12392 113786 12396
rect 113728 12386 113786 12392
rect 115014 12384 115020 12396
rect 115072 12384 115078 12436
rect 116946 12384 116952 12436
rect 117004 12424 117010 12436
rect 118420 12426 118478 12432
rect 118420 12424 118432 12426
rect 117004 12396 118432 12424
rect 117004 12384 117010 12396
rect 118420 12392 118432 12396
rect 118466 12392 118478 12426
rect 118420 12386 118478 12392
rect 127712 12426 127770 12432
rect 127712 12392 127724 12426
rect 127758 12424 127770 12426
rect 127802 12424 127808 12436
rect 127758 12396 127808 12424
rect 127758 12392 127770 12396
rect 127712 12386 127770 12392
rect 127802 12384 127808 12396
rect 127860 12384 127866 12436
rect 129090 12384 129096 12436
rect 129148 12424 129154 12436
rect 130840 12426 130898 12432
rect 130840 12424 130852 12426
rect 129148 12396 130852 12424
rect 129148 12384 129154 12396
rect 130840 12392 130852 12396
rect 130886 12424 130898 12426
rect 130930 12424 130936 12436
rect 130886 12396 130936 12424
rect 130886 12392 130898 12396
rect 130840 12386 130898 12392
rect 130930 12384 130936 12396
rect 130988 12384 130994 12436
rect 132402 12384 132408 12436
rect 132460 12424 132466 12436
rect 132680 12426 132738 12432
rect 132680 12424 132692 12426
rect 132460 12396 132692 12424
rect 132460 12384 132466 12396
rect 132680 12392 132692 12396
rect 132726 12392 132738 12426
rect 132680 12386 132738 12392
rect 147308 12426 147366 12432
rect 147308 12392 147320 12426
rect 147354 12424 147366 12426
rect 147766 12424 147772 12436
rect 147354 12396 147772 12424
rect 147354 12392 147366 12396
rect 147308 12386 147366 12392
rect 147766 12384 147772 12396
rect 147824 12384 147830 12436
rect 152458 12384 152464 12436
rect 152516 12424 152522 12436
rect 152552 12426 152610 12432
rect 152552 12424 152564 12426
rect 152516 12396 152564 12424
rect 152516 12384 152522 12396
rect 152552 12392 152564 12396
rect 152598 12392 152610 12426
rect 152552 12386 152610 12392
rect 152844 12396 153424 12424
rect 86126 12356 86132 12368
rect 80164 12328 86132 12356
rect 78582 12180 78588 12232
rect 78640 12220 78646 12232
rect 80164 12228 80192 12328
rect 86126 12316 86132 12328
rect 86184 12316 86190 12368
rect 87414 12316 87420 12368
rect 87472 12356 87478 12368
rect 89440 12358 89498 12364
rect 89440 12356 89452 12358
rect 87472 12328 89452 12356
rect 87472 12316 87478 12328
rect 89440 12324 89452 12328
rect 89486 12324 89498 12358
rect 89440 12318 89498 12324
rect 94516 12328 113174 12356
rect 81434 12248 81440 12300
rect 81492 12288 81498 12300
rect 84472 12290 84530 12296
rect 84472 12288 84484 12290
rect 81492 12260 84484 12288
rect 81492 12248 81498 12260
rect 84472 12256 84484 12260
rect 84518 12256 84530 12290
rect 84654 12288 84660 12300
rect 84614 12260 84660 12288
rect 84472 12250 84530 12256
rect 84654 12248 84660 12260
rect 84712 12248 84718 12300
rect 85758 12288 85764 12300
rect 85040 12260 85764 12288
rect 79228 12222 79286 12228
rect 79228 12220 79240 12222
rect 78640 12192 79240 12220
rect 78640 12180 78646 12192
rect 79228 12188 79240 12192
rect 79274 12220 79286 12222
rect 80148 12222 80206 12228
rect 80148 12220 80160 12222
rect 79274 12192 80160 12220
rect 79274 12188 79286 12192
rect 79228 12182 79286 12188
rect 80148 12188 80160 12192
rect 80194 12188 80206 12222
rect 80148 12182 80206 12188
rect 83826 12180 83832 12232
rect 83884 12220 83890 12232
rect 84380 12222 84438 12228
rect 84380 12220 84392 12222
rect 83884 12192 84392 12220
rect 83884 12180 83890 12192
rect 84380 12188 84392 12192
rect 84426 12220 84438 12222
rect 85040 12220 85068 12260
rect 85758 12248 85764 12260
rect 85816 12248 85822 12300
rect 86310 12248 86316 12300
rect 86368 12288 86374 12300
rect 87048 12290 87106 12296
rect 87048 12288 87060 12290
rect 86368 12260 87060 12288
rect 86368 12248 86374 12260
rect 87048 12256 87060 12260
rect 87094 12288 87106 12290
rect 88150 12288 88156 12300
rect 87094 12260 88156 12288
rect 87094 12256 87106 12260
rect 87048 12250 87106 12256
rect 88150 12248 88156 12260
rect 88208 12248 88214 12300
rect 89162 12288 89168 12300
rect 88904 12260 89168 12288
rect 85482 12220 85488 12232
rect 84426 12192 85068 12220
rect 85442 12192 85488 12220
rect 84426 12188 84438 12192
rect 84380 12182 84438 12188
rect 85482 12180 85488 12192
rect 85540 12180 85546 12232
rect 86034 12180 86040 12232
rect 86092 12220 86098 12232
rect 86864 12222 86922 12228
rect 86864 12220 86876 12222
rect 86092 12192 86876 12220
rect 86092 12180 86098 12192
rect 86864 12188 86876 12192
rect 86910 12188 86922 12222
rect 86864 12182 86922 12188
rect 87968 12222 88026 12228
rect 87968 12188 87980 12222
rect 88014 12220 88026 12222
rect 88242 12220 88248 12232
rect 88014 12192 88248 12220
rect 88014 12188 88026 12192
rect 87968 12182 88026 12188
rect 88242 12180 88248 12192
rect 88300 12180 88306 12232
rect 88796 12222 88854 12228
rect 88904 12222 88932 12260
rect 89162 12248 89168 12260
rect 89220 12288 89226 12300
rect 89220 12260 90128 12288
rect 89220 12248 89226 12260
rect 88796 12188 88808 12222
rect 88842 12194 88932 12222
rect 88842 12188 88854 12194
rect 88796 12182 88854 12188
rect 88978 12180 88984 12232
rect 89036 12220 89042 12232
rect 90100 12228 90128 12260
rect 89624 12222 89682 12228
rect 89624 12220 89636 12222
rect 89036 12192 89636 12220
rect 89036 12180 89042 12192
rect 89624 12188 89636 12192
rect 89670 12188 89682 12222
rect 89624 12182 89682 12188
rect 90084 12222 90142 12228
rect 90084 12188 90096 12222
rect 90130 12220 90142 12222
rect 92014 12220 92020 12232
rect 90130 12192 92020 12220
rect 90130 12188 90142 12192
rect 90084 12182 90142 12188
rect 92014 12180 92020 12192
rect 92072 12180 92078 12232
rect 94516 12152 94544 12328
rect 99098 12248 99104 12300
rect 99156 12288 99162 12300
rect 100940 12290 100998 12296
rect 100940 12288 100952 12290
rect 99156 12260 100952 12288
rect 99156 12248 99162 12260
rect 100940 12256 100952 12260
rect 100986 12288 100998 12290
rect 102042 12288 102048 12300
rect 100986 12260 102048 12288
rect 100986 12256 100998 12260
rect 100940 12250 100998 12256
rect 102042 12248 102048 12260
rect 102100 12288 102106 12300
rect 103148 12290 103206 12296
rect 103148 12288 103160 12290
rect 102100 12260 103160 12288
rect 102100 12248 102106 12260
rect 103148 12256 103160 12260
rect 103194 12288 103206 12290
rect 103238 12288 103244 12300
rect 103194 12260 103244 12288
rect 103194 12256 103206 12260
rect 103148 12250 103206 12256
rect 103238 12248 103244 12260
rect 103296 12248 103302 12300
rect 103330 12248 103336 12300
rect 103388 12288 103394 12300
rect 104528 12290 104586 12296
rect 104528 12288 104540 12290
rect 103388 12260 104540 12288
rect 103388 12248 103394 12260
rect 104528 12256 104540 12260
rect 104574 12256 104586 12290
rect 113146 12288 113174 12328
rect 115750 12316 115756 12368
rect 115808 12356 115814 12368
rect 141970 12356 141976 12368
rect 115808 12328 117820 12356
rect 115808 12316 115814 12328
rect 117792 12296 117820 12328
rect 130396 12328 141976 12356
rect 114372 12290 114430 12296
rect 114372 12288 114384 12290
rect 113146 12260 114384 12288
rect 104528 12250 104586 12256
rect 114372 12256 114384 12260
rect 114418 12288 114430 12290
rect 117776 12290 117834 12296
rect 114418 12260 116808 12288
rect 114418 12256 114430 12260
rect 114372 12250 114430 12256
rect 97534 12180 97540 12232
rect 97592 12220 97598 12232
rect 99284 12222 99342 12228
rect 99284 12220 99296 12222
rect 97592 12192 99296 12220
rect 97592 12180 97598 12192
rect 99284 12188 99296 12192
rect 99330 12188 99342 12222
rect 99284 12182 99342 12188
rect 99744 12222 99802 12228
rect 99744 12188 99756 12222
rect 99790 12220 99802 12222
rect 102964 12222 103022 12228
rect 99790 12192 102180 12220
rect 99790 12188 99802 12192
rect 99744 12182 99802 12188
rect 102152 12164 102180 12192
rect 102964 12188 102976 12222
rect 103010 12220 103022 12222
rect 103698 12220 103704 12232
rect 103010 12192 103704 12220
rect 103010 12188 103022 12192
rect 102964 12182 103022 12188
rect 103698 12180 103704 12192
rect 103756 12180 103762 12232
rect 103792 12222 103850 12228
rect 103792 12188 103804 12222
rect 103838 12220 103850 12222
rect 104436 12222 104494 12228
rect 104436 12220 104448 12222
rect 103838 12192 104448 12220
rect 103838 12188 103850 12192
rect 103792 12182 103850 12188
rect 104436 12188 104448 12192
rect 104482 12220 104494 12222
rect 105080 12222 105138 12228
rect 105080 12220 105092 12222
rect 104482 12192 105092 12220
rect 104482 12188 104494 12192
rect 104436 12182 104494 12188
rect 105080 12188 105092 12192
rect 105126 12188 105138 12222
rect 105080 12182 105138 12188
rect 100754 12152 100760 12164
rect 76576 12124 77892 12152
rect 78508 12124 88840 12152
rect 55858 12084 55864 12096
rect 55186 12056 55864 12084
rect 55858 12044 55864 12056
rect 55916 12044 55922 12096
rect 56042 12084 56048 12096
rect 56002 12056 56048 12084
rect 56042 12044 56048 12056
rect 56100 12044 56106 12096
rect 56152 12092 56180 12124
rect 56136 12086 56194 12092
rect 56136 12052 56148 12086
rect 56182 12052 56194 12086
rect 56136 12046 56194 12052
rect 56504 12086 56562 12092
rect 56504 12052 56516 12086
rect 56550 12084 56562 12086
rect 57330 12084 57336 12096
rect 56550 12056 57336 12084
rect 56550 12052 56562 12056
rect 56504 12046 56562 12052
rect 57330 12044 57336 12056
rect 57388 12044 57394 12096
rect 76282 12084 76288 12096
rect 76242 12056 76288 12084
rect 76282 12044 76288 12056
rect 76340 12044 76346 12096
rect 77864 12092 77892 12124
rect 77848 12086 77906 12092
rect 77848 12052 77860 12086
rect 77894 12084 77906 12086
rect 80238 12084 80244 12096
rect 77894 12056 80244 12084
rect 77894 12052 77906 12056
rect 77848 12046 77906 12052
rect 80238 12044 80244 12056
rect 80296 12044 80302 12096
rect 84010 12084 84016 12096
rect 83970 12056 84016 12084
rect 84010 12044 84016 12056
rect 84068 12044 84074 12096
rect 84654 12044 84660 12096
rect 84712 12084 84718 12096
rect 86310 12084 86316 12096
rect 84712 12056 86316 12084
rect 84712 12044 84718 12056
rect 86310 12044 86316 12056
rect 86368 12044 86374 12096
rect 86772 12086 86830 12092
rect 86772 12052 86784 12086
rect 86818 12084 86830 12086
rect 87506 12084 87512 12096
rect 86818 12056 87512 12084
rect 86818 12052 86830 12056
rect 86772 12046 86830 12052
rect 87506 12044 87512 12056
rect 87564 12044 87570 12096
rect 87600 12086 87658 12092
rect 87600 12052 87612 12086
rect 87646 12084 87658 12086
rect 87782 12084 87788 12096
rect 87646 12056 87788 12084
rect 87646 12052 87658 12056
rect 87600 12046 87658 12052
rect 87782 12044 87788 12056
rect 87840 12044 87846 12096
rect 87966 12044 87972 12096
rect 88024 12084 88030 12096
rect 88060 12086 88118 12092
rect 88060 12084 88072 12086
rect 88024 12056 88072 12084
rect 88024 12044 88030 12056
rect 88060 12052 88072 12056
rect 88106 12084 88118 12086
rect 88702 12084 88708 12096
rect 88106 12056 88708 12084
rect 88106 12052 88118 12056
rect 88060 12046 88118 12052
rect 88702 12044 88708 12056
rect 88760 12044 88766 12096
rect 88812 12084 88840 12124
rect 89686 12124 94544 12152
rect 100714 12124 100760 12152
rect 89686 12084 89714 12124
rect 100754 12112 100760 12124
rect 100812 12112 100818 12164
rect 100848 12154 100906 12160
rect 100848 12120 100860 12154
rect 100894 12152 100906 12154
rect 101030 12152 101036 12164
rect 100894 12124 101036 12152
rect 100894 12120 100906 12124
rect 100848 12114 100906 12120
rect 101030 12112 101036 12124
rect 101088 12112 101094 12164
rect 101950 12152 101956 12164
rect 101910 12124 101956 12152
rect 101950 12112 101956 12124
rect 102008 12112 102014 12164
rect 102134 12112 102140 12164
rect 102192 12152 102198 12164
rect 103808 12152 103836 12182
rect 111886 12180 111892 12232
rect 111944 12220 111950 12232
rect 113268 12222 113326 12228
rect 113268 12220 113280 12222
rect 111944 12192 113280 12220
rect 111944 12180 111950 12192
rect 113268 12188 113280 12192
rect 113314 12188 113326 12222
rect 113268 12182 113326 12188
rect 113912 12222 113970 12228
rect 113912 12188 113924 12222
rect 113958 12220 113970 12222
rect 114278 12220 114284 12232
rect 113958 12192 114284 12220
rect 113958 12188 113970 12192
rect 113912 12182 113970 12188
rect 114278 12180 114284 12192
rect 114336 12180 114342 12232
rect 116780 12220 116808 12260
rect 117776 12256 117788 12290
rect 117822 12288 117834 12290
rect 118878 12288 118884 12300
rect 117822 12260 118884 12288
rect 117822 12256 117834 12260
rect 117776 12250 117834 12256
rect 118878 12248 118884 12260
rect 118936 12248 118942 12300
rect 130396 12288 130424 12328
rect 141970 12316 141976 12328
rect 142028 12316 142034 12368
rect 147582 12316 147588 12368
rect 147640 12356 147646 12368
rect 148412 12358 148470 12364
rect 148412 12356 148424 12358
rect 147640 12328 148424 12356
rect 147640 12316 147646 12328
rect 148412 12324 148424 12328
rect 148458 12324 148470 12358
rect 148412 12318 148470 12324
rect 151630 12316 151636 12368
rect 151688 12356 151694 12368
rect 152734 12356 152740 12368
rect 151688 12328 152740 12356
rect 151688 12316 151694 12328
rect 129108 12260 130424 12288
rect 117592 12222 117650 12228
rect 116780 12192 117268 12220
rect 102192 12124 103836 12152
rect 102192 12112 102198 12124
rect 113818 12112 113824 12164
rect 113876 12152 113882 12164
rect 114648 12154 114706 12160
rect 114648 12152 114660 12154
rect 113876 12124 114660 12152
rect 113876 12112 113882 12124
rect 114648 12120 114660 12124
rect 114694 12120 114706 12154
rect 114648 12114 114706 12120
rect 114756 12124 115138 12152
rect 100386 12084 100392 12096
rect 88812 12056 89714 12084
rect 100346 12056 100392 12084
rect 100386 12044 100392 12056
rect 100444 12044 100450 12096
rect 101968 12084 101996 12112
rect 102318 12084 102324 12096
rect 101968 12056 102324 12084
rect 102318 12044 102324 12056
rect 102376 12044 102382 12096
rect 102594 12084 102600 12096
rect 102554 12056 102600 12084
rect 102594 12044 102600 12056
rect 102652 12044 102658 12096
rect 103054 12084 103060 12096
rect 103014 12056 103060 12084
rect 103054 12044 103060 12056
rect 103112 12044 103118 12096
rect 113910 12044 113916 12096
rect 113968 12084 113974 12096
rect 114756 12084 114784 12124
rect 113968 12056 114784 12084
rect 113968 12044 113974 12056
rect 115658 12044 115664 12096
rect 115716 12084 115722 12096
rect 116120 12086 116178 12092
rect 116120 12084 116132 12086
rect 115716 12056 116132 12084
rect 115716 12044 115722 12056
rect 116120 12052 116132 12056
rect 116166 12052 116178 12086
rect 116120 12046 116178 12052
rect 116394 12044 116400 12096
rect 116452 12084 116458 12096
rect 117132 12086 117190 12092
rect 117132 12084 117144 12086
rect 116452 12056 117144 12084
rect 116452 12044 116458 12056
rect 117132 12052 117144 12056
rect 117178 12052 117190 12086
rect 117240 12084 117268 12192
rect 117592 12188 117604 12222
rect 117638 12220 117650 12222
rect 118050 12220 118056 12232
rect 117638 12192 118056 12220
rect 117638 12188 117650 12192
rect 117592 12182 117650 12188
rect 118050 12180 118056 12192
rect 118108 12180 118114 12232
rect 118326 12220 118332 12232
rect 118286 12192 118332 12220
rect 118326 12180 118332 12192
rect 118384 12180 118390 12232
rect 126146 12180 126152 12232
rect 126204 12220 126210 12232
rect 127896 12222 127954 12228
rect 127896 12220 127908 12222
rect 126204 12192 127908 12220
rect 126204 12180 126210 12192
rect 127896 12188 127908 12192
rect 127942 12188 127954 12222
rect 128630 12220 128636 12232
rect 128590 12192 128636 12220
rect 127896 12182 127954 12188
rect 128630 12180 128636 12192
rect 128688 12180 128694 12232
rect 129108 12228 129136 12260
rect 131022 12248 131028 12300
rect 131080 12288 131086 12300
rect 131852 12290 131910 12296
rect 131852 12288 131864 12290
rect 131080 12260 131864 12288
rect 131080 12248 131086 12260
rect 131852 12256 131864 12260
rect 131898 12288 131910 12290
rect 133230 12288 133236 12300
rect 131898 12260 133236 12288
rect 131898 12256 131910 12260
rect 131852 12250 131910 12256
rect 133230 12248 133236 12260
rect 133288 12248 133294 12300
rect 149054 12248 149060 12300
rect 149112 12288 149118 12300
rect 152092 12290 152150 12296
rect 152092 12288 152104 12290
rect 149112 12260 152104 12288
rect 149112 12248 149118 12260
rect 152092 12256 152104 12260
rect 152138 12256 152150 12290
rect 152092 12250 152150 12256
rect 152184 12290 152242 12296
rect 152184 12256 152196 12290
rect 152230 12256 152242 12290
rect 152184 12250 152242 12256
rect 129092 12222 129150 12228
rect 129092 12188 129104 12222
rect 129138 12188 129150 12222
rect 129092 12182 129150 12188
rect 117500 12154 117558 12160
rect 117500 12120 117512 12154
rect 117546 12152 117558 12154
rect 118234 12152 118240 12164
rect 117546 12124 118240 12152
rect 117546 12120 117558 12124
rect 117500 12114 117558 12120
rect 118234 12112 118240 12124
rect 118292 12112 118298 12164
rect 129108 12152 129136 12182
rect 130470 12180 130476 12232
rect 130528 12180 130534 12232
rect 131668 12222 131726 12228
rect 131668 12188 131680 12222
rect 131714 12220 131726 12222
rect 132402 12220 132408 12232
rect 131714 12192 132408 12220
rect 131714 12188 131726 12192
rect 131668 12182 131726 12188
rect 132402 12180 132408 12192
rect 132460 12180 132466 12232
rect 132586 12220 132592 12232
rect 132546 12192 132592 12220
rect 132586 12180 132592 12192
rect 132644 12180 132650 12232
rect 137738 12220 137744 12232
rect 137698 12192 137744 12220
rect 137738 12180 137744 12192
rect 137796 12180 137802 12232
rect 147492 12222 147550 12228
rect 147492 12188 147504 12222
rect 147538 12220 147550 12222
rect 148042 12220 148048 12232
rect 147538 12192 148048 12220
rect 147538 12188 147550 12192
rect 147492 12182 147550 12188
rect 148042 12180 148048 12192
rect 148100 12180 148106 12232
rect 148320 12222 148378 12228
rect 148320 12188 148332 12222
rect 148366 12220 148378 12222
rect 149330 12220 149336 12232
rect 148366 12192 149336 12220
rect 148366 12188 148378 12192
rect 148320 12182 148378 12188
rect 149330 12180 149336 12192
rect 149388 12180 149394 12232
rect 149422 12180 149428 12232
rect 149480 12220 149486 12232
rect 149480 12192 149524 12220
rect 149480 12180 149486 12192
rect 151354 12180 151360 12232
rect 151412 12220 151418 12232
rect 152200 12220 152228 12250
rect 152476 12228 152504 12328
rect 152734 12316 152740 12328
rect 152792 12316 152798 12368
rect 151412 12192 152228 12220
rect 152460 12222 152518 12228
rect 151412 12180 151418 12192
rect 152460 12188 152472 12222
rect 152506 12188 152518 12222
rect 152460 12182 152518 12188
rect 122806 12124 129136 12152
rect 129368 12154 129426 12160
rect 122806 12084 122834 12124
rect 129368 12120 129380 12154
rect 129414 12120 129426 12154
rect 132494 12152 132500 12164
rect 129368 12114 129426 12120
rect 131316 12124 132500 12152
rect 117240 12056 122834 12084
rect 128448 12086 128506 12092
rect 117132 12046 117190 12052
rect 128448 12052 128460 12086
rect 128494 12084 128506 12086
rect 129384 12084 129412 12114
rect 131316 12092 131344 12124
rect 132494 12112 132500 12124
rect 132552 12112 132558 12164
rect 138014 12152 138020 12164
rect 137974 12124 138020 12152
rect 138014 12112 138020 12124
rect 138072 12152 138078 12164
rect 145836 12154 145894 12160
rect 145836 12152 145848 12154
rect 138072 12124 145848 12152
rect 138072 12112 138078 12124
rect 145836 12120 145848 12124
rect 145882 12120 145894 12154
rect 145836 12114 145894 12120
rect 146204 12154 146262 12160
rect 146204 12120 146216 12154
rect 146250 12152 146262 12154
rect 152844 12152 152872 12396
rect 153288 12358 153346 12364
rect 153288 12324 153300 12358
rect 153334 12324 153346 12358
rect 153396 12356 153424 12396
rect 153746 12384 153752 12436
rect 153804 12424 153810 12436
rect 154116 12426 154174 12432
rect 154116 12424 154128 12426
rect 153804 12396 154128 12424
rect 153804 12384 153810 12396
rect 154116 12392 154128 12396
rect 154162 12392 154174 12426
rect 154116 12386 154174 12392
rect 157242 12384 157248 12436
rect 157300 12424 157306 12436
rect 160922 12424 160928 12436
rect 157300 12396 160928 12424
rect 157300 12384 157306 12396
rect 160922 12384 160928 12396
rect 160980 12384 160986 12436
rect 161566 12384 161572 12436
rect 161624 12424 161630 12436
rect 165340 12426 165398 12432
rect 161624 12396 164924 12424
rect 161624 12384 161630 12396
rect 155034 12356 155040 12368
rect 153396 12328 155040 12356
rect 153288 12318 153346 12324
rect 153304 12220 153332 12318
rect 155034 12316 155040 12328
rect 155092 12316 155098 12368
rect 158898 12316 158904 12368
rect 158956 12356 158962 12368
rect 160004 12358 160062 12364
rect 160004 12356 160016 12358
rect 158956 12328 160016 12356
rect 158956 12316 158962 12328
rect 160004 12324 160016 12328
rect 160050 12324 160062 12358
rect 164896 12356 164924 12396
rect 165340 12392 165352 12426
rect 165386 12424 165398 12426
rect 166442 12424 166448 12436
rect 165386 12396 166448 12424
rect 165386 12392 165398 12396
rect 165340 12386 165398 12392
rect 166442 12384 166448 12396
rect 166500 12384 166506 12436
rect 175920 12426 175978 12432
rect 175920 12392 175932 12426
rect 175966 12424 175978 12426
rect 176470 12424 176476 12436
rect 175966 12396 176476 12424
rect 175966 12392 175978 12396
rect 175920 12386 175978 12392
rect 176470 12384 176476 12396
rect 176528 12384 176534 12436
rect 179506 12384 179512 12436
rect 179564 12424 179570 12436
rect 181348 12426 181406 12432
rect 181348 12424 181360 12426
rect 179564 12396 181360 12424
rect 179564 12384 179570 12396
rect 181348 12392 181360 12396
rect 181394 12392 181406 12426
rect 181348 12386 181406 12392
rect 188524 12426 188582 12432
rect 188524 12392 188536 12426
rect 188570 12424 188582 12426
rect 189166 12424 189172 12436
rect 188570 12396 189172 12424
rect 188570 12392 188582 12396
rect 188524 12386 188582 12392
rect 189166 12384 189172 12396
rect 189224 12384 189230 12436
rect 189626 12384 189632 12436
rect 189684 12424 189690 12436
rect 190180 12426 190238 12432
rect 190180 12424 190192 12426
rect 189684 12396 190192 12424
rect 189684 12384 189690 12396
rect 190180 12392 190192 12396
rect 190226 12392 190238 12426
rect 190180 12386 190238 12392
rect 190822 12384 190828 12436
rect 190880 12424 190886 12436
rect 194042 12424 194048 12436
rect 190880 12396 194048 12424
rect 190880 12384 190886 12396
rect 194042 12384 194048 12396
rect 194100 12384 194106 12436
rect 201680 12426 201738 12432
rect 194152 12396 197584 12424
rect 165430 12356 165436 12368
rect 164896 12328 165436 12356
rect 160004 12318 160062 12324
rect 165430 12316 165436 12328
rect 165488 12316 165494 12368
rect 166074 12356 166080 12368
rect 166034 12328 166080 12356
rect 166074 12316 166080 12328
rect 166132 12316 166138 12368
rect 177758 12356 177764 12368
rect 177040 12328 177764 12356
rect 153932 12290 153990 12296
rect 153932 12256 153944 12290
rect 153978 12288 153990 12290
rect 154114 12288 154120 12300
rect 153978 12260 154120 12288
rect 153978 12256 153990 12260
rect 153932 12250 153990 12256
rect 154114 12248 154120 12260
rect 154172 12248 154178 12300
rect 160370 12248 160376 12300
rect 160428 12288 160434 12300
rect 161292 12290 161350 12296
rect 161292 12288 161304 12290
rect 160428 12260 161304 12288
rect 160428 12248 160434 12260
rect 161292 12256 161304 12260
rect 161338 12256 161350 12290
rect 161292 12250 161350 12256
rect 161474 12248 161480 12300
rect 161532 12288 161538 12300
rect 162486 12288 162492 12300
rect 161532 12260 161576 12288
rect 162446 12260 162492 12288
rect 161532 12248 161538 12260
rect 162486 12248 162492 12260
rect 162544 12248 162550 12300
rect 162670 12288 162676 12300
rect 162630 12260 162676 12288
rect 162670 12248 162676 12260
rect 162728 12248 162734 12300
rect 163590 12288 163596 12300
rect 163550 12260 163596 12288
rect 163590 12248 163596 12260
rect 163648 12248 163654 12300
rect 177040 12296 177068 12328
rect 177758 12316 177764 12328
rect 177816 12316 177822 12368
rect 180886 12356 180892 12368
rect 180846 12328 180892 12356
rect 180886 12316 180892 12328
rect 180944 12316 180950 12368
rect 192570 12356 192576 12368
rect 185596 12328 190500 12356
rect 192530 12328 192576 12356
rect 177024 12290 177082 12296
rect 177024 12256 177036 12290
rect 177070 12256 177082 12290
rect 177024 12250 177082 12256
rect 177114 12248 177120 12300
rect 177172 12288 177178 12300
rect 185596 12288 185624 12328
rect 177172 12260 177216 12288
rect 179156 12260 185624 12288
rect 177172 12248 177178 12260
rect 154300 12222 154358 12228
rect 154300 12220 154312 12222
rect 153304 12192 154312 12220
rect 154300 12188 154312 12192
rect 154346 12188 154358 12222
rect 154300 12182 154358 12188
rect 158806 12180 158812 12232
rect 158864 12220 158870 12232
rect 160188 12222 160246 12228
rect 160188 12220 160200 12222
rect 158864 12192 160200 12220
rect 158864 12180 158870 12192
rect 160188 12188 160200 12192
rect 160234 12188 160246 12222
rect 160188 12182 160246 12188
rect 161200 12222 161258 12228
rect 161200 12188 161212 12222
rect 161246 12220 161258 12222
rect 161750 12220 161756 12232
rect 161246 12192 161756 12220
rect 161246 12188 161258 12192
rect 161200 12182 161258 12188
rect 161750 12180 161756 12192
rect 161808 12220 161814 12232
rect 162504 12220 162532 12248
rect 179156 12232 179184 12260
rect 187970 12248 187976 12300
rect 188028 12288 188034 12300
rect 188028 12260 190408 12288
rect 188028 12248 188034 12260
rect 161808 12192 162532 12220
rect 176104 12222 176162 12228
rect 161808 12180 161814 12192
rect 176104 12188 176116 12222
rect 176150 12220 176162 12222
rect 176932 12222 176990 12228
rect 176932 12220 176944 12222
rect 176150 12192 176944 12220
rect 176150 12188 176162 12192
rect 176104 12182 176162 12188
rect 176932 12188 176944 12192
rect 176978 12220 176990 12222
rect 177850 12220 177856 12232
rect 176978 12192 177856 12220
rect 176978 12188 176990 12192
rect 176932 12182 176990 12188
rect 177850 12180 177856 12192
rect 177908 12180 177914 12232
rect 179138 12220 179144 12232
rect 179098 12192 179144 12220
rect 179138 12180 179144 12192
rect 179196 12180 179202 12232
rect 180702 12180 180708 12232
rect 180760 12220 180766 12232
rect 181532 12222 181590 12228
rect 181532 12220 181544 12222
rect 180760 12192 181544 12220
rect 180760 12180 180766 12192
rect 181532 12188 181544 12192
rect 181578 12188 181590 12222
rect 181532 12182 181590 12188
rect 188708 12222 188766 12228
rect 188708 12188 188720 12222
rect 188754 12188 188766 12222
rect 189534 12220 189540 12232
rect 189494 12192 189540 12220
rect 188708 12182 188766 12188
rect 146250 12124 147674 12152
rect 146250 12120 146262 12124
rect 146204 12114 146262 12120
rect 128494 12056 129412 12084
rect 131300 12086 131358 12092
rect 128494 12052 128506 12056
rect 128448 12046 128506 12052
rect 131300 12052 131312 12086
rect 131346 12052 131358 12086
rect 131300 12046 131358 12052
rect 131574 12044 131580 12096
rect 131632 12084 131638 12096
rect 131760 12086 131818 12092
rect 131760 12084 131772 12086
rect 131632 12056 131772 12084
rect 131632 12044 131638 12056
rect 131760 12052 131772 12056
rect 131806 12052 131818 12086
rect 147646 12084 147674 12124
rect 149440 12124 152872 12152
rect 153656 12154 153714 12160
rect 149440 12084 149468 12124
rect 153656 12120 153668 12154
rect 153702 12152 153714 12154
rect 155862 12152 155868 12164
rect 153702 12124 155868 12152
rect 153702 12120 153714 12124
rect 153656 12114 153714 12120
rect 155862 12112 155868 12124
rect 155920 12112 155926 12164
rect 156414 12112 156420 12164
rect 156472 12152 156478 12164
rect 162578 12152 162584 12164
rect 156472 12124 162584 12152
rect 156472 12112 156478 12124
rect 162578 12112 162584 12124
rect 162636 12112 162642 12164
rect 162670 12112 162676 12164
rect 162728 12152 162734 12164
rect 163868 12154 163926 12160
rect 163868 12152 163880 12154
rect 162728 12124 163880 12152
rect 162728 12112 162734 12124
rect 163868 12120 163880 12124
rect 163914 12120 163926 12154
rect 163868 12114 163926 12120
rect 164326 12112 164332 12164
rect 164384 12112 164390 12164
rect 165890 12152 165896 12164
rect 165850 12124 165896 12152
rect 165890 12112 165896 12124
rect 165948 12112 165954 12164
rect 166534 12112 166540 12164
rect 166592 12152 166598 12164
rect 177944 12154 178002 12160
rect 177944 12152 177956 12154
rect 166592 12124 177956 12152
rect 166592 12112 166598 12124
rect 177944 12120 177956 12124
rect 177990 12152 178002 12154
rect 179414 12152 179420 12164
rect 177990 12124 179276 12152
rect 179374 12124 179420 12152
rect 177990 12120 178002 12124
rect 177944 12114 178002 12120
rect 147646 12056 149468 12084
rect 131760 12046 131818 12052
rect 149514 12044 149520 12096
rect 149572 12084 149578 12096
rect 150712 12086 150770 12092
rect 150712 12084 150724 12086
rect 149572 12056 150724 12084
rect 149572 12044 149578 12056
rect 150712 12052 150724 12056
rect 150758 12052 150770 12086
rect 151630 12084 151636 12096
rect 151590 12056 151636 12084
rect 150712 12046 150770 12052
rect 151630 12044 151636 12056
rect 151688 12044 151694 12096
rect 151722 12044 151728 12096
rect 151780 12084 151786 12096
rect 152000 12086 152058 12092
rect 152000 12084 152012 12086
rect 151780 12056 152012 12084
rect 151780 12044 151786 12056
rect 152000 12052 152012 12056
rect 152046 12052 152058 12086
rect 152000 12046 152058 12052
rect 152182 12044 152188 12096
rect 152240 12084 152246 12096
rect 152550 12084 152556 12096
rect 152240 12056 152556 12084
rect 152240 12044 152246 12056
rect 152550 12044 152556 12056
rect 152608 12084 152614 12096
rect 153748 12086 153806 12092
rect 153748 12084 153760 12086
rect 152608 12056 153760 12084
rect 152608 12044 152614 12056
rect 153748 12052 153760 12056
rect 153794 12052 153806 12086
rect 153748 12046 153806 12052
rect 160832 12086 160890 12092
rect 160832 12052 160844 12086
rect 160878 12084 160890 12086
rect 161106 12084 161112 12096
rect 160878 12056 161112 12084
rect 160878 12052 160890 12056
rect 160832 12046 160890 12052
rect 161106 12044 161112 12056
rect 161164 12044 161170 12096
rect 162028 12086 162086 12092
rect 162028 12052 162040 12086
rect 162074 12084 162086 12086
rect 162210 12084 162216 12096
rect 162074 12056 162216 12084
rect 162074 12052 162086 12056
rect 162028 12046 162086 12052
rect 162210 12044 162216 12056
rect 162268 12044 162274 12096
rect 162396 12086 162454 12092
rect 162396 12052 162408 12086
rect 162442 12084 162454 12086
rect 162854 12084 162860 12096
rect 162442 12056 162860 12084
rect 162442 12052 162454 12056
rect 162396 12046 162454 12052
rect 162854 12044 162860 12056
rect 162912 12044 162918 12096
rect 176564 12086 176622 12092
rect 176564 12052 176576 12086
rect 176610 12084 176622 12086
rect 176654 12084 176660 12096
rect 176610 12056 176660 12084
rect 176610 12052 176622 12056
rect 176564 12046 176622 12052
rect 176654 12044 176660 12056
rect 176712 12044 176718 12096
rect 178034 12084 178040 12096
rect 177994 12056 178040 12084
rect 178034 12044 178040 12056
rect 178092 12044 178098 12096
rect 179248 12084 179276 12124
rect 179414 12112 179420 12124
rect 179472 12112 179478 12164
rect 181438 12152 181444 12164
rect 180642 12124 181444 12152
rect 181438 12112 181444 12124
rect 181496 12112 181502 12164
rect 188724 12152 188752 12182
rect 189534 12180 189540 12192
rect 189592 12180 189598 12232
rect 190380 12228 190408 12260
rect 190364 12222 190422 12228
rect 190364 12188 190376 12222
rect 190410 12188 190422 12222
rect 190472 12220 190500 12328
rect 192570 12316 192576 12328
rect 192628 12316 192634 12368
rect 190824 12290 190882 12296
rect 190824 12256 190836 12290
rect 190870 12288 190882 12290
rect 191834 12288 191840 12300
rect 190870 12260 191840 12288
rect 190870 12256 190882 12260
rect 190824 12250 190882 12256
rect 190840 12220 190868 12250
rect 191834 12248 191840 12260
rect 191892 12248 191898 12300
rect 192662 12248 192668 12300
rect 192720 12288 192726 12300
rect 193676 12290 193734 12296
rect 193676 12288 193688 12290
rect 192720 12260 193688 12288
rect 192720 12248 192726 12260
rect 193676 12256 193688 12260
rect 193722 12288 193734 12290
rect 194152 12288 194180 12396
rect 197446 12356 197452 12368
rect 196452 12328 197452 12356
rect 193722 12260 194180 12288
rect 194428 12260 196020 12288
rect 193722 12256 193734 12260
rect 193676 12250 193734 12256
rect 194428 12232 194456 12260
rect 194410 12220 194416 12232
rect 190472 12192 190868 12220
rect 192404 12192 193812 12220
rect 194370 12192 194416 12220
rect 190364 12182 190422 12188
rect 190822 12152 190828 12164
rect 188724 12124 190828 12152
rect 190822 12112 190828 12124
rect 190880 12112 190886 12164
rect 191098 12152 191104 12164
rect 191058 12124 191104 12152
rect 191098 12112 191104 12124
rect 191156 12112 191162 12164
rect 191190 12112 191196 12164
rect 191248 12152 191254 12164
rect 191248 12124 191590 12152
rect 191248 12112 191254 12124
rect 180150 12084 180156 12096
rect 179248 12056 180156 12084
rect 180150 12044 180156 12056
rect 180208 12044 180214 12096
rect 189628 12086 189686 12092
rect 189628 12052 189640 12086
rect 189674 12084 189686 12086
rect 192404 12084 192432 12192
rect 193398 12152 193404 12164
rect 193358 12124 193404 12152
rect 193398 12112 193404 12124
rect 193456 12112 193462 12164
rect 193030 12084 193036 12096
rect 189674 12056 192432 12084
rect 192990 12056 193036 12084
rect 189674 12052 189686 12056
rect 189628 12046 189686 12052
rect 193030 12044 193036 12056
rect 193088 12044 193094 12096
rect 193492 12086 193550 12092
rect 193492 12052 193504 12086
rect 193538 12084 193550 12086
rect 193674 12084 193680 12096
rect 193538 12056 193680 12084
rect 193538 12052 193550 12056
rect 193492 12046 193550 12052
rect 193674 12044 193680 12056
rect 193732 12044 193738 12096
rect 193784 12084 193812 12192
rect 194410 12180 194416 12192
rect 194468 12180 194474 12232
rect 194686 12152 194692 12164
rect 194646 12124 194692 12152
rect 194686 12112 194692 12124
rect 194744 12112 194750 12164
rect 195992 12152 196020 12260
rect 196452 12228 196480 12328
rect 197446 12316 197452 12328
rect 197504 12316 197510 12368
rect 197556 12296 197584 12396
rect 201680 12392 201692 12426
rect 201726 12424 201738 12426
rect 202414 12424 202420 12436
rect 201726 12396 202420 12424
rect 201726 12392 201738 12396
rect 201680 12386 201738 12392
rect 202414 12384 202420 12396
rect 202472 12384 202478 12436
rect 205634 12424 205640 12436
rect 203628 12396 205640 12424
rect 201128 12358 201186 12364
rect 201128 12324 201140 12358
rect 201174 12356 201186 12358
rect 203628 12356 203656 12396
rect 205634 12384 205640 12396
rect 205692 12384 205698 12436
rect 206464 12426 206522 12432
rect 206464 12392 206476 12426
rect 206510 12424 206522 12426
rect 207658 12424 207664 12436
rect 206510 12396 207664 12424
rect 206510 12392 206522 12396
rect 206464 12386 206522 12392
rect 207658 12384 207664 12396
rect 207716 12384 207722 12436
rect 227796 12426 227854 12432
rect 227796 12392 227808 12426
rect 227842 12424 227854 12426
rect 230106 12424 230112 12436
rect 227842 12396 230112 12424
rect 227842 12392 227854 12396
rect 227796 12386 227854 12392
rect 230106 12384 230112 12396
rect 230164 12384 230170 12436
rect 231854 12384 231860 12436
rect 231912 12424 231918 12436
rect 232224 12426 232282 12432
rect 232224 12424 232236 12426
rect 231912 12396 232236 12424
rect 231912 12384 231918 12396
rect 232224 12392 232236 12396
rect 232270 12392 232282 12426
rect 232224 12386 232282 12392
rect 239030 12384 239036 12436
rect 239088 12424 239094 12436
rect 239952 12426 240010 12432
rect 239952 12424 239964 12426
rect 239088 12396 239964 12424
rect 239088 12384 239094 12396
rect 239952 12392 239964 12396
rect 239998 12392 240010 12426
rect 239952 12386 240010 12392
rect 240134 12384 240140 12436
rect 240192 12424 240198 12436
rect 243540 12426 243598 12432
rect 240192 12396 241192 12424
rect 240192 12384 240198 12396
rect 201174 12328 203656 12356
rect 201174 12324 201186 12328
rect 201128 12318 201186 12324
rect 228818 12316 228824 12368
rect 228876 12356 228882 12368
rect 229740 12358 229798 12364
rect 229740 12356 229752 12358
rect 228876 12328 229752 12356
rect 228876 12316 228882 12328
rect 229740 12324 229752 12328
rect 229786 12324 229798 12358
rect 229740 12318 229798 12324
rect 231118 12316 231124 12368
rect 231176 12356 231182 12368
rect 232498 12356 232504 12368
rect 231176 12328 232504 12356
rect 231176 12316 231182 12328
rect 232498 12316 232504 12328
rect 232556 12316 232562 12368
rect 238756 12358 238814 12364
rect 238756 12324 238768 12358
rect 238802 12356 238814 12358
rect 241164 12356 241192 12396
rect 242360 12396 243124 12424
rect 242250 12356 242256 12368
rect 238802 12328 239720 12356
rect 238802 12324 238814 12328
rect 238756 12318 238814 12324
rect 197540 12290 197598 12296
rect 196544 12260 196848 12288
rect 196436 12222 196494 12228
rect 196436 12188 196448 12222
rect 196482 12188 196494 12222
rect 196436 12182 196494 12188
rect 196544 12152 196572 12260
rect 196712 12222 196770 12228
rect 196712 12220 196724 12222
rect 194796 12124 195178 12152
rect 195992 12124 196572 12152
rect 196636 12192 196724 12220
rect 194796 12084 194824 12124
rect 193784 12056 194824 12084
rect 194962 12044 194968 12096
rect 195020 12084 195026 12096
rect 196636 12084 196664 12192
rect 196712 12188 196724 12192
rect 196758 12188 196770 12222
rect 196712 12182 196770 12188
rect 196820 12152 196848 12260
rect 197540 12256 197552 12290
rect 197586 12256 197598 12290
rect 197540 12250 197598 12256
rect 200482 12248 200488 12300
rect 200540 12288 200546 12300
rect 200540 12260 201908 12288
rect 200540 12248 200546 12260
rect 197446 12220 197452 12232
rect 197358 12192 197452 12220
rect 197446 12180 197452 12192
rect 197504 12220 197510 12232
rect 198366 12220 198372 12232
rect 197504 12192 198372 12220
rect 197504 12180 197510 12192
rect 198366 12180 198372 12192
rect 198424 12180 198430 12232
rect 200574 12180 200580 12232
rect 200632 12220 200638 12232
rect 201034 12220 201040 12232
rect 200632 12192 201040 12220
rect 200632 12180 200638 12192
rect 201034 12180 201040 12192
rect 201092 12180 201098 12232
rect 201880 12228 201908 12260
rect 202046 12248 202052 12300
rect 202104 12288 202110 12300
rect 203518 12288 203524 12300
rect 202104 12260 203524 12288
rect 202104 12248 202110 12260
rect 203518 12248 203524 12260
rect 203576 12248 203582 12300
rect 204716 12290 204774 12296
rect 204716 12256 204728 12290
rect 204762 12288 204774 12290
rect 231580 12290 231638 12296
rect 204762 12260 209774 12288
rect 204762 12256 204774 12260
rect 204716 12250 204774 12256
rect 201864 12222 201922 12228
rect 201864 12188 201876 12222
rect 201910 12188 201922 12222
rect 201864 12182 201922 12188
rect 203244 12222 203302 12228
rect 203244 12188 203256 12222
rect 203290 12220 203302 12222
rect 204530 12220 204536 12232
rect 203290 12192 204536 12220
rect 203290 12188 203302 12192
rect 203244 12182 203302 12188
rect 204530 12180 204536 12192
rect 204588 12180 204594 12232
rect 204732 12152 204760 12250
rect 209746 12220 209774 12260
rect 227548 12260 231440 12288
rect 227548 12228 227576 12260
rect 227532 12222 227590 12228
rect 227532 12220 227544 12222
rect 209746 12192 227544 12220
rect 227532 12188 227544 12192
rect 227578 12188 227590 12222
rect 229922 12220 229928 12232
rect 229834 12192 229928 12220
rect 227532 12182 227590 12188
rect 229922 12180 229928 12192
rect 229980 12220 229986 12232
rect 231302 12220 231308 12232
rect 229980 12192 231308 12220
rect 229980 12180 229986 12192
rect 231302 12180 231308 12192
rect 231360 12180 231366 12232
rect 204990 12152 204996 12164
rect 196820 12124 204760 12152
rect 204950 12124 204996 12152
rect 204990 12112 204996 12124
rect 205048 12112 205054 12164
rect 230842 12152 230848 12164
rect 205100 12124 205482 12152
rect 229034 12124 230848 12152
rect 196802 12084 196808 12096
rect 195020 12056 196664 12084
rect 196762 12056 196808 12084
rect 195020 12044 195026 12056
rect 196802 12044 196808 12056
rect 196860 12044 196866 12096
rect 196986 12084 196992 12096
rect 196946 12056 196992 12084
rect 196986 12044 196992 12056
rect 197044 12044 197050 12096
rect 197354 12084 197360 12096
rect 197314 12056 197360 12084
rect 197354 12044 197360 12056
rect 197412 12044 197418 12096
rect 202876 12086 202934 12092
rect 202876 12052 202888 12086
rect 202922 12084 202934 12086
rect 203058 12084 203064 12096
rect 202922 12056 203064 12084
rect 202922 12052 202934 12056
rect 202876 12046 202934 12052
rect 203058 12044 203064 12056
rect 203116 12044 203122 12096
rect 203336 12086 203394 12092
rect 203336 12052 203348 12086
rect 203382 12084 203394 12086
rect 203426 12084 203432 12096
rect 203382 12056 203432 12084
rect 203382 12052 203394 12056
rect 203336 12046 203394 12052
rect 203426 12044 203432 12056
rect 203484 12044 203490 12096
rect 204254 12044 204260 12096
rect 204312 12084 204318 12096
rect 205100 12084 205128 12124
rect 230842 12112 230848 12124
rect 230900 12112 230906 12164
rect 231118 12112 231124 12164
rect 231176 12152 231182 12164
rect 231412 12152 231440 12260
rect 231580 12256 231592 12290
rect 231626 12288 231638 12290
rect 231670 12288 231676 12300
rect 231626 12260 231676 12288
rect 231626 12256 231638 12260
rect 231580 12250 231638 12256
rect 231670 12248 231676 12260
rect 231728 12248 231734 12300
rect 238846 12248 238852 12300
rect 238904 12288 238910 12300
rect 239306 12288 239312 12300
rect 238904 12260 239312 12288
rect 238904 12248 238910 12260
rect 239306 12248 239312 12260
rect 239364 12248 239370 12300
rect 232130 12220 232136 12232
rect 232042 12192 232136 12220
rect 232130 12180 232136 12192
rect 232188 12220 232194 12232
rect 233050 12220 233056 12232
rect 232188 12192 233056 12220
rect 232188 12180 232194 12192
rect 233050 12180 233056 12192
rect 233108 12180 233114 12232
rect 238018 12220 238024 12232
rect 237978 12192 238024 12220
rect 238018 12180 238024 12192
rect 238076 12180 238082 12232
rect 238386 12180 238392 12232
rect 238444 12220 238450 12232
rect 239122 12220 239128 12232
rect 238444 12192 239128 12220
rect 238444 12180 238450 12192
rect 239122 12180 239128 12192
rect 239180 12180 239186 12232
rect 239216 12222 239274 12228
rect 239216 12188 239228 12222
rect 239262 12220 239274 12222
rect 239490 12220 239496 12232
rect 239262 12192 239496 12220
rect 239262 12188 239274 12192
rect 239216 12182 239274 12188
rect 239490 12180 239496 12192
rect 239548 12180 239554 12232
rect 239692 12220 239720 12328
rect 239968 12328 241008 12356
rect 241164 12328 242256 12356
rect 239968 12300 239996 12328
rect 239950 12248 239956 12300
rect 240008 12248 240014 12300
rect 240980 12288 241008 12328
rect 242250 12316 242256 12328
rect 242308 12316 242314 12368
rect 242360 12364 242388 12396
rect 242344 12358 242402 12364
rect 242344 12324 242356 12358
rect 242390 12324 242402 12358
rect 242986 12356 242992 12368
rect 242344 12318 242402 12324
rect 242728 12328 242992 12356
rect 241424 12290 241482 12296
rect 241424 12288 241436 12290
rect 240980 12260 241436 12288
rect 241424 12256 241436 12260
rect 241470 12288 241482 12290
rect 241470 12260 242296 12288
rect 241470 12256 241482 12260
rect 241424 12250 241482 12256
rect 242268 12236 242296 12260
rect 242434 12248 242440 12300
rect 242492 12288 242498 12300
rect 242728 12288 242756 12328
rect 242986 12316 242992 12328
rect 243044 12316 243050 12368
rect 242804 12290 242862 12296
rect 242804 12288 242816 12290
rect 242492 12260 242816 12288
rect 242492 12248 242498 12260
rect 242804 12256 242816 12260
rect 242850 12256 242862 12290
rect 242804 12250 242862 12256
rect 242894 12248 242900 12300
rect 242952 12288 242958 12300
rect 242952 12260 243044 12288
rect 242952 12248 242958 12260
rect 240136 12222 240194 12228
rect 240136 12220 240148 12222
rect 239692 12192 240148 12220
rect 240136 12188 240148 12192
rect 240182 12188 240194 12222
rect 240136 12182 240194 12188
rect 241240 12222 241298 12228
rect 241240 12188 241252 12222
rect 241286 12220 241298 12222
rect 242158 12220 242164 12232
rect 241286 12192 242164 12220
rect 241286 12188 241298 12192
rect 241240 12182 241298 12188
rect 242158 12180 242164 12192
rect 242216 12180 242222 12232
rect 242268 12220 242388 12236
rect 242268 12216 242848 12220
rect 242912 12216 242940 12248
rect 242268 12208 242940 12216
rect 242360 12192 242940 12208
rect 243096 12220 243124 12396
rect 243540 12392 243552 12426
rect 243586 12424 243598 12426
rect 243630 12424 243636 12436
rect 243586 12396 243636 12424
rect 243586 12392 243598 12396
rect 243540 12386 243598 12392
rect 243630 12384 243636 12396
rect 243688 12384 243694 12436
rect 244182 12424 244188 12436
rect 244142 12396 244188 12424
rect 244182 12384 244188 12396
rect 244240 12384 244246 12436
rect 251084 12426 251142 12432
rect 251084 12392 251096 12426
rect 251130 12424 251142 12426
rect 251358 12424 251364 12436
rect 251130 12396 251364 12424
rect 251130 12392 251142 12396
rect 251084 12386 251142 12392
rect 251358 12384 251364 12396
rect 251416 12384 251422 12436
rect 251910 12384 251916 12436
rect 251968 12424 251974 12436
rect 251968 12396 256280 12424
rect 251968 12384 251974 12396
rect 251450 12316 251456 12368
rect 251508 12356 251514 12368
rect 252094 12356 252100 12368
rect 251508 12328 252100 12356
rect 251508 12316 251514 12328
rect 252094 12316 252100 12328
rect 252152 12316 252158 12368
rect 254302 12356 254308 12368
rect 254214 12328 254308 12356
rect 254302 12316 254308 12328
rect 254360 12356 254366 12368
rect 255222 12356 255228 12368
rect 254360 12328 255228 12356
rect 254360 12316 254366 12328
rect 255222 12316 255228 12328
rect 255280 12316 255286 12368
rect 243170 12248 243176 12300
rect 243228 12288 243234 12300
rect 243228 12260 244412 12288
rect 243228 12248 243234 12260
rect 244384 12228 244412 12260
rect 248322 12248 248328 12300
rect 248380 12288 248386 12300
rect 249242 12288 249248 12300
rect 248380 12260 249248 12288
rect 248380 12248 248386 12260
rect 249242 12248 249248 12260
rect 249300 12248 249306 12300
rect 252556 12290 252614 12296
rect 252556 12288 252568 12290
rect 251146 12260 252568 12288
rect 243724 12222 243782 12228
rect 243724 12220 243736 12222
rect 243096 12192 243736 12220
rect 242820 12188 242940 12192
rect 243724 12188 243736 12192
rect 243770 12188 243782 12222
rect 243724 12182 243782 12188
rect 244368 12222 244426 12228
rect 244368 12188 244380 12222
rect 244414 12188 244426 12222
rect 251146 12220 251174 12260
rect 252556 12256 252568 12260
rect 252602 12288 252614 12290
rect 255316 12290 255374 12296
rect 252602 12260 255268 12288
rect 252602 12256 252614 12260
rect 252556 12250 252614 12256
rect 244368 12182 244426 12188
rect 248386 12192 251174 12220
rect 248386 12152 248414 12192
rect 251266 12180 251272 12232
rect 251324 12220 251330 12232
rect 251910 12220 251916 12232
rect 251324 12192 251368 12220
rect 251870 12192 251916 12220
rect 251324 12180 251330 12192
rect 251910 12180 251916 12192
rect 251968 12180 251974 12232
rect 255130 12220 255136 12232
rect 255090 12192 255136 12220
rect 255130 12180 255136 12192
rect 255188 12180 255194 12232
rect 249058 12152 249064 12164
rect 231176 12124 231348 12152
rect 231412 12124 248414 12152
rect 249018 12124 249064 12152
rect 231176 12112 231182 12124
rect 204312 12056 205128 12084
rect 204312 12044 204318 12056
rect 228818 12044 228824 12096
rect 228876 12084 228882 12096
rect 229280 12086 229338 12092
rect 229280 12084 229292 12086
rect 228876 12056 229292 12084
rect 228876 12044 228882 12056
rect 229280 12052 229292 12056
rect 229326 12052 229338 12086
rect 229280 12046 229338 12052
rect 230936 12086 230994 12092
rect 230936 12052 230948 12086
rect 230982 12084 230994 12086
rect 231210 12084 231216 12096
rect 230982 12056 231216 12084
rect 230982 12052 230994 12056
rect 230936 12046 230994 12052
rect 231210 12044 231216 12056
rect 231268 12044 231274 12096
rect 231320 12092 231348 12124
rect 249058 12112 249064 12124
rect 249116 12112 249122 12164
rect 249242 12112 249248 12164
rect 249300 12152 249306 12164
rect 251928 12152 251956 12180
rect 249300 12124 251956 12152
rect 252832 12154 252890 12160
rect 249300 12112 249306 12124
rect 252832 12120 252844 12154
rect 252878 12152 252890 12154
rect 253106 12152 253112 12164
rect 252878 12124 253112 12152
rect 252878 12120 252890 12124
rect 252832 12114 252890 12120
rect 253106 12112 253112 12124
rect 253164 12112 253170 12164
rect 255240 12152 255268 12260
rect 255316 12256 255328 12290
rect 255362 12288 255374 12290
rect 255590 12288 255596 12300
rect 255362 12260 255596 12288
rect 255362 12256 255374 12260
rect 255316 12250 255374 12256
rect 255590 12248 255596 12260
rect 255648 12248 255654 12300
rect 256252 12288 256280 12396
rect 256510 12384 256516 12436
rect 256568 12424 256574 12436
rect 256880 12426 256938 12432
rect 256880 12424 256892 12426
rect 256568 12396 256892 12424
rect 256568 12384 256574 12396
rect 256880 12392 256892 12396
rect 256926 12392 256938 12426
rect 262490 12424 262496 12436
rect 262450 12396 262496 12424
rect 256880 12386 256938 12392
rect 262490 12384 262496 12396
rect 262548 12384 262554 12436
rect 264608 12426 264666 12432
rect 264608 12392 264620 12426
rect 264654 12424 264666 12426
rect 265526 12424 265532 12436
rect 264654 12396 265532 12424
rect 264654 12392 264666 12396
rect 264608 12386 264666 12392
rect 265526 12384 265532 12396
rect 265584 12384 265590 12436
rect 268010 12424 268016 12436
rect 265912 12396 268016 12424
rect 256328 12358 256386 12364
rect 256328 12324 256340 12358
rect 256374 12356 256386 12358
rect 256970 12356 256976 12368
rect 256374 12328 256976 12356
rect 256374 12324 256386 12328
rect 256328 12318 256386 12324
rect 256970 12316 256976 12328
rect 257028 12316 257034 12368
rect 264056 12358 264114 12364
rect 264056 12324 264068 12358
rect 264102 12356 264114 12358
rect 264974 12356 264980 12368
rect 264102 12328 264980 12356
rect 264102 12324 264114 12328
rect 264056 12318 264114 12324
rect 264974 12316 264980 12328
rect 265032 12316 265038 12368
rect 265912 12356 265940 12396
rect 268010 12384 268016 12396
rect 268068 12384 268074 12436
rect 268378 12384 268384 12436
rect 268436 12424 268442 12436
rect 271046 12424 271052 12436
rect 268436 12396 270080 12424
rect 271006 12396 271052 12424
rect 268436 12384 268442 12396
rect 265084 12328 265940 12356
rect 270052 12356 270080 12396
rect 271046 12384 271052 12396
rect 271104 12384 271110 12436
rect 305454 12424 305460 12436
rect 305414 12396 305460 12424
rect 305454 12384 305460 12396
rect 305512 12384 305518 12436
rect 271692 12358 271750 12364
rect 271692 12356 271704 12358
rect 270052 12328 271704 12356
rect 261846 12288 261852 12300
rect 256252 12260 261852 12288
rect 261846 12248 261852 12260
rect 261904 12248 261910 12300
rect 262398 12248 262404 12300
rect 262456 12288 262462 12300
rect 262456 12260 264008 12288
rect 262456 12248 262462 12260
rect 256234 12220 256240 12232
rect 256194 12192 256240 12220
rect 256234 12180 256240 12192
rect 256292 12180 256298 12232
rect 256326 12180 256332 12232
rect 256384 12220 256390 12232
rect 257064 12222 257122 12228
rect 257064 12220 257076 12222
rect 256384 12192 257076 12220
rect 256384 12180 256390 12192
rect 257064 12188 257076 12192
rect 257110 12188 257122 12222
rect 257064 12182 257122 12188
rect 262676 12222 262734 12228
rect 262676 12188 262688 12222
rect 262722 12220 262734 12222
rect 263042 12220 263048 12232
rect 262722 12192 263048 12220
rect 262722 12188 262734 12192
rect 262676 12182 262734 12188
rect 263042 12180 263048 12192
rect 263100 12180 263106 12232
rect 263980 12228 264008 12260
rect 264146 12248 264152 12300
rect 264204 12288 264210 12300
rect 265084 12288 265112 12328
rect 264204 12260 265112 12288
rect 264204 12248 264210 12260
rect 265158 12248 265164 12300
rect 265216 12288 265222 12300
rect 265216 12260 265388 12288
rect 265216 12248 265222 12260
rect 263964 12222 264022 12228
rect 263964 12188 263976 12222
rect 264010 12220 264022 12222
rect 264330 12220 264336 12232
rect 264010 12192 264336 12220
rect 264010 12188 264022 12192
rect 263964 12182 264022 12188
rect 264330 12180 264336 12192
rect 264388 12180 264394 12232
rect 264792 12222 264850 12228
rect 264792 12188 264804 12222
rect 264838 12220 264850 12222
rect 265360 12220 265388 12260
rect 265618 12248 265624 12300
rect 265676 12288 265682 12300
rect 265912 12296 265940 12328
rect 271692 12324 271704 12328
rect 271738 12324 271750 12358
rect 271692 12318 271750 12324
rect 265712 12290 265770 12296
rect 265712 12288 265724 12290
rect 265676 12260 265724 12288
rect 265676 12248 265682 12260
rect 265712 12256 265724 12260
rect 265758 12256 265770 12290
rect 265712 12250 265770 12256
rect 265896 12290 265954 12296
rect 265896 12256 265908 12290
rect 265942 12256 265954 12290
rect 268748 12290 268806 12296
rect 268748 12288 268760 12290
rect 265896 12250 265954 12256
rect 266556 12260 268760 12288
rect 266556 12228 266584 12260
rect 268748 12256 268760 12260
rect 268794 12288 268806 12290
rect 269114 12288 269120 12300
rect 268794 12260 269120 12288
rect 268794 12256 268806 12260
rect 268748 12250 268806 12256
rect 269114 12248 269120 12260
rect 269172 12248 269178 12300
rect 269666 12248 269672 12300
rect 269724 12288 269730 12300
rect 271138 12288 271144 12300
rect 269724 12260 271144 12288
rect 269724 12248 269730 12260
rect 271138 12248 271144 12260
rect 271196 12248 271202 12300
rect 272242 12288 272248 12300
rect 272202 12260 272248 12288
rect 272242 12248 272248 12260
rect 272300 12288 272306 12300
rect 272794 12288 272800 12300
rect 272300 12260 272800 12288
rect 272300 12248 272306 12260
rect 272794 12248 272800 12260
rect 272852 12248 272858 12300
rect 266540 12222 266598 12228
rect 266540 12220 266552 12222
rect 264838 12192 265296 12220
rect 265360 12192 266552 12220
rect 264838 12188 264850 12192
rect 264792 12182 264850 12188
rect 265158 12152 265164 12164
rect 254058 12124 255084 12152
rect 255240 12124 256464 12152
rect 255056 12096 255084 12124
rect 231304 12086 231362 12092
rect 231304 12052 231316 12086
rect 231350 12052 231362 12086
rect 231304 12046 231362 12052
rect 231394 12044 231400 12096
rect 231452 12084 231458 12096
rect 231762 12084 231768 12096
rect 231452 12056 231768 12084
rect 231452 12044 231458 12056
rect 231762 12044 231768 12056
rect 231820 12044 231826 12096
rect 233050 12044 233056 12096
rect 233108 12084 233114 12096
rect 238204 12086 238262 12092
rect 238204 12084 238216 12086
rect 233108 12056 238216 12084
rect 233108 12044 233114 12056
rect 238204 12052 238216 12056
rect 238250 12052 238262 12086
rect 240870 12084 240876 12096
rect 240830 12056 240876 12084
rect 238204 12046 238262 12052
rect 240870 12044 240876 12056
rect 240928 12044 240934 12096
rect 241332 12086 241390 12092
rect 241332 12052 241344 12086
rect 241378 12084 241390 12086
rect 241514 12084 241520 12096
rect 241378 12056 241520 12084
rect 241378 12052 241390 12056
rect 241332 12046 241390 12052
rect 241514 12044 241520 12056
rect 241572 12084 241578 12096
rect 242526 12084 242532 12096
rect 241572 12056 242532 12084
rect 241572 12044 241578 12056
rect 242526 12044 242532 12056
rect 242584 12044 242590 12096
rect 242712 12086 242770 12092
rect 242712 12052 242724 12086
rect 242758 12084 242770 12086
rect 244090 12084 244096 12096
rect 242758 12056 244096 12084
rect 242758 12052 242770 12056
rect 242712 12046 242770 12052
rect 244090 12044 244096 12056
rect 244148 12044 244154 12096
rect 254394 12044 254400 12096
rect 254452 12084 254458 12096
rect 254764 12086 254822 12092
rect 254764 12084 254776 12086
rect 254452 12056 254776 12084
rect 254452 12044 254458 12056
rect 254764 12052 254776 12056
rect 254810 12052 254822 12086
rect 254764 12046 254822 12052
rect 255038 12044 255044 12096
rect 255096 12044 255102 12096
rect 255222 12044 255228 12096
rect 255280 12084 255286 12096
rect 256326 12084 256332 12096
rect 255280 12056 256332 12084
rect 255280 12044 255286 12056
rect 256326 12044 256332 12056
rect 256384 12044 256390 12096
rect 256436 12084 256464 12124
rect 263566 12124 265164 12152
rect 263566 12084 263594 12124
rect 265158 12112 265164 12124
rect 265216 12112 265222 12164
rect 265268 12092 265296 12192
rect 266540 12188 266552 12192
rect 266586 12188 266598 12222
rect 266540 12182 266598 12188
rect 268102 12180 268108 12232
rect 268160 12220 268166 12232
rect 268654 12220 268660 12232
rect 268160 12192 268660 12220
rect 268160 12180 268166 12192
rect 268654 12180 268660 12192
rect 268712 12180 268718 12232
rect 270956 12222 271014 12228
rect 270956 12220 270968 12222
rect 270328 12192 270968 12220
rect 265620 12154 265678 12160
rect 265620 12120 265632 12154
rect 265666 12152 265678 12154
rect 266814 12152 266820 12164
rect 265666 12124 266676 12152
rect 266774 12124 266820 12152
rect 265666 12120 265678 12124
rect 265620 12114 265678 12120
rect 256436 12056 263594 12084
rect 265252 12086 265310 12092
rect 265252 12052 265264 12086
rect 265298 12052 265310 12086
rect 266648 12084 266676 12124
rect 266814 12112 266820 12124
rect 266872 12112 266878 12164
rect 267274 12112 267280 12164
rect 267332 12112 267338 12164
rect 268194 12112 268200 12164
rect 268252 12152 268258 12164
rect 269024 12154 269082 12160
rect 269024 12152 269036 12154
rect 268252 12124 269036 12152
rect 268252 12112 268258 12124
rect 269024 12120 269036 12124
rect 269070 12120 269082 12154
rect 269024 12114 269082 12120
rect 269482 12112 269488 12164
rect 269540 12112 269546 12164
rect 266998 12084 267004 12096
rect 266648 12056 267004 12084
rect 265252 12046 265310 12052
rect 266998 12044 267004 12056
rect 267056 12044 267062 12096
rect 268288 12086 268346 12092
rect 268288 12052 268300 12086
rect 268334 12084 268346 12086
rect 268470 12084 268476 12096
rect 268334 12056 268476 12084
rect 268334 12052 268346 12056
rect 268288 12046 268346 12052
rect 268470 12044 268476 12056
rect 268528 12044 268534 12096
rect 268654 12044 268660 12096
rect 268712 12084 268718 12096
rect 270328 12084 270356 12192
rect 270956 12188 270968 12192
rect 271002 12220 271014 12222
rect 271322 12220 271328 12232
rect 271002 12192 271328 12220
rect 271002 12188 271014 12192
rect 270956 12182 271014 12188
rect 271322 12180 271328 12192
rect 271380 12180 271386 12232
rect 272060 12222 272118 12228
rect 272060 12188 272072 12222
rect 272106 12220 272118 12222
rect 272886 12220 272892 12232
rect 272106 12192 272892 12220
rect 272106 12188 272118 12192
rect 272060 12182 272118 12188
rect 272886 12180 272892 12192
rect 272944 12180 272950 12232
rect 270512 12124 272196 12152
rect 268712 12056 270356 12084
rect 268712 12044 268718 12056
rect 270402 12044 270408 12096
rect 270460 12084 270466 12096
rect 270512 12092 270540 12124
rect 272168 12092 272196 12124
rect 270496 12086 270554 12092
rect 270496 12084 270508 12086
rect 270460 12056 270508 12084
rect 270460 12044 270466 12056
rect 270496 12052 270508 12056
rect 270542 12052 270554 12086
rect 270496 12046 270554 12052
rect 272152 12086 272210 12092
rect 272152 12052 272164 12086
rect 272198 12084 272210 12086
rect 284754 12084 284760 12096
rect 272198 12056 284760 12084
rect 272198 12052 272210 12056
rect 272152 12046 272210 12052
rect 284754 12044 284760 12056
rect 284812 12044 284818 12096
rect 1104 11994 305808 12016
rect 1104 11942 77148 11994
rect 77200 11942 77212 11994
rect 77264 11942 77276 11994
rect 77328 11942 77340 11994
rect 77392 11942 77404 11994
rect 77456 11942 153346 11994
rect 153398 11942 153410 11994
rect 153462 11942 153474 11994
rect 153526 11942 153538 11994
rect 153590 11942 153602 11994
rect 153654 11942 229544 11994
rect 229596 11942 229608 11994
rect 229660 11942 229672 11994
rect 229724 11942 229736 11994
rect 229788 11942 229800 11994
rect 229852 11942 305808 11994
rect 1104 11920 305808 11942
rect 27800 11882 27858 11888
rect 27800 11848 27812 11882
rect 27846 11880 27858 11882
rect 29086 11880 29092 11892
rect 27846 11852 29092 11880
rect 27846 11848 27858 11852
rect 27800 11842 27858 11848
rect 29086 11840 29092 11852
rect 29144 11840 29150 11892
rect 29454 11840 29460 11892
rect 29512 11880 29518 11892
rect 30926 11880 30932 11892
rect 29512 11852 30932 11880
rect 29512 11840 29518 11852
rect 30926 11840 30932 11852
rect 30984 11840 30990 11892
rect 32214 11840 32220 11892
rect 32272 11880 32278 11892
rect 32584 11882 32642 11888
rect 32584 11880 32596 11882
rect 32272 11852 32596 11880
rect 32272 11840 32278 11852
rect 32584 11848 32596 11852
rect 32630 11848 32642 11882
rect 33778 11880 33784 11892
rect 33738 11852 33784 11880
rect 32584 11842 32642 11848
rect 33778 11840 33784 11852
rect 33836 11840 33842 11892
rect 34422 11880 34428 11892
rect 34382 11852 34428 11880
rect 34422 11840 34428 11852
rect 34480 11840 34486 11892
rect 34976 11882 35034 11888
rect 34976 11848 34988 11882
rect 35022 11848 35034 11882
rect 38378 11880 38384 11892
rect 38338 11852 38384 11880
rect 34976 11842 35034 11848
rect 27706 11772 27712 11824
rect 27764 11812 27770 11824
rect 27764 11784 28120 11812
rect 27764 11772 27770 11784
rect 27984 11746 28042 11752
rect 27984 11712 27996 11746
rect 28030 11712 28042 11746
rect 27984 11706 28042 11712
rect 28000 11608 28028 11706
rect 28092 11676 28120 11784
rect 28718 11772 28724 11824
rect 28776 11812 28782 11824
rect 28812 11814 28870 11820
rect 28812 11812 28824 11814
rect 28776 11784 28824 11812
rect 28776 11772 28782 11784
rect 28812 11780 28824 11784
rect 28858 11780 28870 11814
rect 28812 11774 28870 11780
rect 28994 11772 29000 11824
rect 29052 11812 29058 11824
rect 30006 11812 30012 11824
rect 29052 11784 30012 11812
rect 29052 11772 29058 11784
rect 28902 11676 28908 11688
rect 28092 11648 28908 11676
rect 28902 11636 28908 11648
rect 28960 11636 28966 11688
rect 29104 11684 29132 11784
rect 30006 11772 30012 11784
rect 30064 11772 30070 11824
rect 32030 11772 32036 11824
rect 32088 11812 32094 11824
rect 34992 11812 35020 11842
rect 38378 11840 38384 11852
rect 38436 11840 38442 11892
rect 39024 11882 39082 11888
rect 39024 11848 39036 11882
rect 39070 11880 39082 11882
rect 39574 11880 39580 11892
rect 39070 11852 39580 11880
rect 39070 11848 39082 11852
rect 39024 11842 39082 11848
rect 39574 11840 39580 11852
rect 39632 11840 39638 11892
rect 39668 11882 39726 11888
rect 39668 11848 39680 11882
rect 39714 11848 39726 11882
rect 39668 11842 39726 11848
rect 32088 11784 35020 11812
rect 32088 11772 32094 11784
rect 29546 11704 29552 11756
rect 29604 11744 29610 11756
rect 29640 11746 29698 11752
rect 29640 11744 29652 11746
rect 29604 11716 29652 11744
rect 29604 11704 29610 11716
rect 29640 11712 29652 11716
rect 29686 11712 29698 11746
rect 32398 11744 32404 11756
rect 31050 11716 32404 11744
rect 29640 11706 29698 11712
rect 32398 11704 32404 11716
rect 32456 11704 32462 11756
rect 32492 11746 32550 11752
rect 32492 11712 32504 11746
rect 32538 11744 32550 11746
rect 33688 11746 33746 11752
rect 32538 11716 32812 11744
rect 32538 11712 32550 11716
rect 32492 11706 32550 11712
rect 29088 11678 29146 11684
rect 29088 11644 29100 11678
rect 29134 11644 29146 11678
rect 29914 11676 29920 11688
rect 29874 11648 29920 11676
rect 29088 11638 29146 11644
rect 29914 11636 29920 11648
rect 29972 11636 29978 11688
rect 32508 11676 32536 11706
rect 30944 11648 32536 11676
rect 28000 11580 29776 11608
rect 28442 11540 28448 11552
rect 28402 11512 28448 11540
rect 28442 11500 28448 11512
rect 28500 11500 28506 11552
rect 29748 11540 29776 11580
rect 30944 11540 30972 11648
rect 32582 11636 32588 11688
rect 32640 11676 32646 11688
rect 32676 11678 32734 11684
rect 32676 11676 32688 11678
rect 32640 11648 32688 11676
rect 32640 11636 32646 11648
rect 32676 11644 32688 11648
rect 32722 11644 32734 11678
rect 32784 11676 32812 11716
rect 33688 11712 33700 11746
rect 33734 11744 33746 11746
rect 34332 11746 34390 11752
rect 34332 11744 34344 11746
rect 33734 11716 34344 11744
rect 33734 11712 33746 11716
rect 33688 11706 33746 11712
rect 34332 11712 34344 11716
rect 34378 11744 34390 11746
rect 34698 11744 34704 11756
rect 34378 11716 34704 11744
rect 34378 11712 34390 11716
rect 34332 11706 34390 11712
rect 34698 11704 34704 11716
rect 34756 11704 34762 11756
rect 35160 11746 35218 11752
rect 35160 11712 35172 11746
rect 35206 11712 35218 11746
rect 35160 11706 35218 11712
rect 38564 11746 38622 11752
rect 38564 11712 38576 11746
rect 38610 11712 38622 11746
rect 38564 11706 38622 11712
rect 39208 11746 39266 11752
rect 39208 11712 39220 11746
rect 39254 11744 39266 11746
rect 39684 11744 39712 11842
rect 39942 11840 39948 11892
rect 40000 11880 40006 11892
rect 40128 11882 40186 11888
rect 40128 11880 40140 11882
rect 40000 11852 40140 11880
rect 40000 11840 40006 11852
rect 40128 11848 40140 11852
rect 40174 11848 40186 11882
rect 40128 11842 40186 11848
rect 41140 11882 41198 11888
rect 41140 11848 41152 11882
rect 41186 11880 41198 11882
rect 41414 11880 41420 11892
rect 41186 11852 41420 11880
rect 41186 11848 41198 11852
rect 41140 11842 41198 11848
rect 41414 11840 41420 11852
rect 41472 11840 41478 11892
rect 41692 11882 41750 11888
rect 41692 11848 41704 11882
rect 41738 11880 41750 11882
rect 42886 11880 42892 11892
rect 41738 11852 42892 11880
rect 41738 11848 41750 11852
rect 41692 11842 41750 11848
rect 42886 11840 42892 11852
rect 42944 11840 42950 11892
rect 52638 11840 52644 11892
rect 52696 11880 52702 11892
rect 52824 11882 52882 11888
rect 52824 11880 52836 11882
rect 52696 11852 52836 11880
rect 52696 11840 52702 11852
rect 52824 11848 52836 11852
rect 52870 11848 52882 11882
rect 53650 11880 53656 11892
rect 53610 11852 53656 11880
rect 52824 11842 52882 11848
rect 53650 11840 53656 11852
rect 53708 11840 53714 11892
rect 54386 11880 54392 11892
rect 54346 11852 54392 11880
rect 54386 11840 54392 11852
rect 54444 11840 54450 11892
rect 55306 11880 55312 11892
rect 55266 11852 55312 11880
rect 55306 11840 55312 11852
rect 55364 11840 55370 11892
rect 56504 11882 56562 11888
rect 56504 11848 56516 11882
rect 56550 11880 56562 11882
rect 56594 11880 56600 11892
rect 56550 11852 56600 11880
rect 56550 11848 56562 11852
rect 56504 11842 56562 11848
rect 56594 11840 56600 11852
rect 56652 11840 56658 11892
rect 57148 11882 57206 11888
rect 57148 11848 57160 11882
rect 57194 11880 57206 11882
rect 58618 11880 58624 11892
rect 57194 11852 58624 11880
rect 57194 11848 57206 11852
rect 57148 11842 57206 11848
rect 58618 11840 58624 11852
rect 58676 11840 58682 11892
rect 75454 11840 75460 11892
rect 75512 11880 75518 11892
rect 75548 11882 75606 11888
rect 75548 11880 75560 11882
rect 75512 11852 75560 11880
rect 75512 11840 75518 11852
rect 75548 11848 75560 11852
rect 75594 11848 75606 11882
rect 75548 11842 75606 11848
rect 75638 11840 75644 11892
rect 75696 11880 75702 11892
rect 76008 11882 76066 11888
rect 76008 11880 76020 11882
rect 75696 11852 76020 11880
rect 75696 11840 75702 11852
rect 76008 11848 76020 11852
rect 76054 11848 76066 11882
rect 76008 11842 76066 11848
rect 76466 11840 76472 11892
rect 76524 11880 76530 11892
rect 76928 11882 76986 11888
rect 76928 11880 76940 11882
rect 76524 11852 76940 11880
rect 76524 11840 76530 11852
rect 76928 11848 76940 11852
rect 76974 11848 76986 11882
rect 77846 11880 77852 11892
rect 77806 11852 77852 11880
rect 76928 11842 76986 11848
rect 77846 11840 77852 11852
rect 77904 11840 77910 11892
rect 78490 11880 78496 11892
rect 78450 11852 78496 11880
rect 78490 11840 78496 11852
rect 78548 11840 78554 11892
rect 84286 11840 84292 11892
rect 84344 11880 84350 11892
rect 84380 11882 84438 11888
rect 84380 11880 84392 11882
rect 84344 11852 84392 11880
rect 84344 11840 84350 11852
rect 84380 11848 84392 11852
rect 84426 11848 84438 11882
rect 86034 11880 86040 11892
rect 84380 11842 84438 11848
rect 85040 11852 86040 11880
rect 40036 11814 40094 11820
rect 40036 11780 40048 11814
rect 40082 11812 40094 11814
rect 40678 11812 40684 11824
rect 40082 11784 40684 11812
rect 40082 11780 40094 11784
rect 40036 11774 40094 11780
rect 39254 11716 39712 11744
rect 39254 11712 39266 11716
rect 39208 11706 39266 11712
rect 34054 11676 34060 11688
rect 32784 11648 34060 11676
rect 32676 11638 32734 11644
rect 34054 11636 34060 11648
rect 34112 11636 34118 11688
rect 31110 11568 31116 11620
rect 31168 11608 31174 11620
rect 35176 11608 35204 11706
rect 38580 11676 38608 11706
rect 40052 11676 40080 11774
rect 40678 11772 40684 11784
rect 40736 11812 40742 11824
rect 41230 11812 41236 11824
rect 40736 11784 41236 11812
rect 40736 11772 40742 11784
rect 41230 11772 41236 11784
rect 41288 11772 41294 11824
rect 53742 11772 53748 11824
rect 53800 11812 53806 11824
rect 53800 11784 56456 11812
rect 53800 11772 53806 11784
rect 40310 11704 40316 11756
rect 40368 11744 40374 11756
rect 41048 11746 41106 11752
rect 41048 11744 41060 11746
rect 40368 11716 41060 11744
rect 40368 11704 40374 11716
rect 41048 11712 41060 11716
rect 41094 11744 41106 11746
rect 41876 11746 41934 11752
rect 41094 11716 41414 11744
rect 41094 11712 41106 11716
rect 41048 11706 41106 11712
rect 41386 11688 41414 11716
rect 41876 11712 41888 11746
rect 41922 11744 41934 11746
rect 42794 11744 42800 11756
rect 41922 11716 42800 11744
rect 41922 11712 41934 11716
rect 41876 11706 41934 11712
rect 42794 11704 42800 11716
rect 42852 11704 42858 11756
rect 42888 11746 42946 11752
rect 42888 11712 42900 11746
rect 42934 11744 42946 11746
rect 42978 11744 42984 11756
rect 42934 11716 42984 11744
rect 42934 11712 42946 11716
rect 42888 11706 42946 11712
rect 42978 11704 42984 11716
rect 43036 11744 43042 11756
rect 53006 11744 53012 11756
rect 43036 11716 43484 11744
rect 52966 11716 53012 11744
rect 43036 11704 43042 11716
rect 38580 11648 40080 11676
rect 40220 11678 40278 11684
rect 40220 11644 40232 11678
rect 40266 11676 40278 11678
rect 40954 11676 40960 11688
rect 40266 11648 40960 11676
rect 40266 11644 40278 11648
rect 40220 11638 40278 11644
rect 40954 11636 40960 11648
rect 41012 11636 41018 11688
rect 41386 11648 41420 11688
rect 41414 11636 41420 11648
rect 41472 11676 41478 11688
rect 43072 11678 43130 11684
rect 43072 11676 43084 11678
rect 41472 11648 43084 11676
rect 41472 11636 41478 11648
rect 43072 11644 43084 11648
rect 43118 11644 43130 11678
rect 43072 11638 43130 11644
rect 43456 11616 43484 11716
rect 53006 11704 53012 11716
rect 53064 11704 53070 11756
rect 54312 11752 54340 11784
rect 56428 11752 56456 11784
rect 57422 11772 57428 11824
rect 57480 11812 57486 11824
rect 84930 11812 84936 11824
rect 57480 11784 84936 11812
rect 57480 11772 57486 11784
rect 84930 11772 84936 11784
rect 84988 11772 84994 11824
rect 53836 11746 53894 11752
rect 53836 11712 53848 11746
rect 53882 11712 53894 11746
rect 53836 11706 53894 11712
rect 54296 11746 54354 11752
rect 54296 11712 54308 11746
rect 54342 11712 54354 11746
rect 54296 11706 54354 11712
rect 56412 11746 56470 11752
rect 56412 11712 56424 11746
rect 56458 11744 56470 11746
rect 57056 11746 57114 11752
rect 57056 11744 57068 11746
rect 56458 11716 57068 11744
rect 56458 11712 56470 11716
rect 56412 11706 56470 11712
rect 57056 11712 57068 11716
rect 57102 11712 57114 11746
rect 57056 11706 57114 11712
rect 53852 11676 53880 11706
rect 54662 11676 54668 11688
rect 53852 11648 54668 11676
rect 54662 11636 54668 11648
rect 54720 11676 54726 11688
rect 55400 11678 55458 11684
rect 55400 11676 55412 11678
rect 54720 11648 55412 11676
rect 54720 11636 54726 11648
rect 55400 11644 55412 11648
rect 55446 11644 55458 11678
rect 55582 11676 55588 11688
rect 55542 11648 55588 11676
rect 55400 11638 55458 11644
rect 55582 11636 55588 11648
rect 55640 11636 55646 11688
rect 55858 11636 55864 11688
rect 55916 11676 55922 11688
rect 57440 11676 57468 11772
rect 75916 11746 75974 11752
rect 75916 11712 75928 11746
rect 75962 11744 75974 11746
rect 76006 11744 76012 11756
rect 75962 11716 76012 11744
rect 75962 11712 75974 11716
rect 75916 11706 75974 11712
rect 76006 11704 76012 11716
rect 76064 11704 76070 11756
rect 76282 11704 76288 11756
rect 76340 11744 76346 11756
rect 77112 11746 77170 11752
rect 77112 11744 77124 11746
rect 76340 11716 77124 11744
rect 76340 11704 76346 11716
rect 77112 11712 77124 11716
rect 77158 11712 77170 11746
rect 77112 11706 77170 11712
rect 77756 11746 77814 11752
rect 77756 11712 77768 11746
rect 77802 11744 77814 11746
rect 78582 11744 78588 11756
rect 77802 11716 78588 11744
rect 77802 11712 77814 11716
rect 77756 11706 77814 11712
rect 78582 11704 78588 11716
rect 78640 11704 78646 11756
rect 78676 11746 78734 11752
rect 78676 11712 78688 11746
rect 78722 11744 78734 11746
rect 81434 11744 81440 11756
rect 78722 11716 81440 11744
rect 78722 11712 78734 11716
rect 78676 11706 78734 11712
rect 81434 11704 81440 11716
rect 81492 11704 81498 11756
rect 84564 11746 84622 11752
rect 84564 11712 84576 11746
rect 84610 11744 84622 11746
rect 85040 11744 85068 11852
rect 86034 11840 86040 11852
rect 86092 11840 86098 11892
rect 86126 11840 86132 11892
rect 86184 11880 86190 11892
rect 87140 11882 87198 11888
rect 87140 11880 87152 11882
rect 86184 11852 87152 11880
rect 86184 11840 86190 11852
rect 87140 11848 87152 11852
rect 87186 11848 87198 11882
rect 87874 11880 87880 11892
rect 87834 11852 87880 11880
rect 87140 11842 87198 11848
rect 87874 11840 87880 11852
rect 87932 11840 87938 11892
rect 88888 11882 88946 11888
rect 88888 11848 88900 11882
rect 88934 11880 88946 11882
rect 89530 11880 89536 11892
rect 88934 11852 89536 11880
rect 88934 11848 88946 11852
rect 88888 11842 88946 11848
rect 89530 11840 89536 11852
rect 89588 11840 89594 11892
rect 99650 11840 99656 11892
rect 99708 11880 99714 11892
rect 100204 11882 100262 11888
rect 100204 11880 100216 11882
rect 99708 11852 100216 11880
rect 99708 11840 99714 11852
rect 100204 11848 100216 11852
rect 100250 11848 100262 11882
rect 100938 11880 100944 11892
rect 100898 11852 100944 11880
rect 100204 11842 100262 11848
rect 100938 11840 100944 11852
rect 100996 11840 101002 11892
rect 101860 11882 101918 11888
rect 101860 11848 101872 11882
rect 101906 11880 101918 11882
rect 103054 11880 103060 11892
rect 101906 11852 103060 11880
rect 101906 11848 101918 11852
rect 101860 11842 101918 11848
rect 103054 11840 103060 11852
rect 103112 11840 103118 11892
rect 103514 11840 103520 11892
rect 103572 11880 103578 11892
rect 113818 11880 113824 11892
rect 103572 11852 113174 11880
rect 113778 11852 113824 11880
rect 103572 11840 103578 11852
rect 85298 11772 85304 11824
rect 85356 11812 85362 11824
rect 113146 11812 113174 11852
rect 113818 11840 113824 11852
rect 113876 11840 113882 11892
rect 114278 11840 114284 11892
rect 114336 11880 114342 11892
rect 115016 11882 115074 11888
rect 115016 11880 115028 11882
rect 114336 11852 115028 11880
rect 114336 11840 114342 11852
rect 115016 11848 115028 11852
rect 115062 11880 115074 11882
rect 115658 11880 115664 11892
rect 115062 11852 115664 11880
rect 115062 11848 115074 11852
rect 115016 11842 115074 11848
rect 115658 11840 115664 11852
rect 115716 11840 115722 11892
rect 116212 11882 116270 11888
rect 116212 11848 116224 11882
rect 116258 11880 116270 11882
rect 116762 11880 116768 11892
rect 116258 11852 116768 11880
rect 116258 11848 116270 11852
rect 116212 11842 116270 11848
rect 116762 11840 116768 11852
rect 116820 11840 116826 11892
rect 116948 11882 117006 11888
rect 116948 11848 116960 11882
rect 116994 11880 117006 11882
rect 117314 11880 117320 11892
rect 116994 11852 117320 11880
rect 116994 11848 117006 11852
rect 116948 11842 117006 11848
rect 117314 11840 117320 11852
rect 117372 11840 117378 11892
rect 117592 11882 117650 11888
rect 117592 11848 117604 11882
rect 117638 11880 117650 11882
rect 118786 11880 118792 11892
rect 117638 11852 118792 11880
rect 117638 11848 117650 11852
rect 117592 11842 117650 11848
rect 118786 11840 118792 11852
rect 118844 11840 118850 11892
rect 129366 11880 129372 11892
rect 129326 11852 129372 11880
rect 129366 11840 129372 11852
rect 129424 11840 129430 11892
rect 130286 11840 130292 11892
rect 130344 11880 130350 11892
rect 130472 11882 130530 11888
rect 130472 11880 130484 11882
rect 130344 11852 130484 11880
rect 130344 11840 130350 11852
rect 130472 11848 130484 11852
rect 130518 11848 130530 11882
rect 130930 11880 130936 11892
rect 130890 11852 130936 11880
rect 130472 11842 130530 11848
rect 130930 11840 130936 11852
rect 130988 11840 130994 11892
rect 131114 11840 131120 11892
rect 131172 11880 131178 11892
rect 132404 11882 132462 11888
rect 132404 11880 132416 11882
rect 131172 11852 132416 11880
rect 131172 11840 131178 11852
rect 132404 11848 132416 11852
rect 132450 11848 132462 11882
rect 132404 11842 132462 11848
rect 137738 11840 137744 11892
rect 137796 11880 137802 11892
rect 151078 11880 151084 11892
rect 137796 11852 150940 11880
rect 151038 11852 151084 11880
rect 137796 11840 137802 11852
rect 114554 11812 114560 11824
rect 85356 11784 108252 11812
rect 113146 11784 114560 11812
rect 85356 11772 85362 11784
rect 84610 11716 85068 11744
rect 85208 11746 85266 11752
rect 84610 11712 84622 11716
rect 84564 11706 84622 11712
rect 85208 11712 85220 11746
rect 85254 11712 85266 11746
rect 85208 11706 85266 11712
rect 55916 11648 57468 11676
rect 55916 11636 55922 11648
rect 74994 11636 75000 11688
rect 75052 11676 75058 11688
rect 76192 11678 76250 11684
rect 76192 11676 76204 11678
rect 75052 11648 76204 11676
rect 75052 11636 75058 11648
rect 76192 11644 76204 11648
rect 76238 11676 76250 11678
rect 76926 11676 76932 11688
rect 76238 11648 76932 11676
rect 76238 11644 76250 11648
rect 76192 11638 76250 11644
rect 76926 11636 76932 11648
rect 76984 11636 76990 11688
rect 84010 11636 84016 11688
rect 84068 11676 84074 11688
rect 85224 11676 85252 11706
rect 85758 11704 85764 11756
rect 85816 11744 85822 11756
rect 86128 11746 86186 11752
rect 86128 11744 86140 11746
rect 85816 11716 86140 11744
rect 85816 11704 85822 11716
rect 86128 11712 86140 11716
rect 86174 11712 86186 11746
rect 86128 11706 86186 11712
rect 86954 11704 86960 11756
rect 87012 11744 87018 11756
rect 87784 11746 87842 11752
rect 87012 11716 87056 11744
rect 87012 11704 87018 11716
rect 87784 11712 87796 11746
rect 87830 11744 87842 11746
rect 88796 11746 88854 11752
rect 87830 11716 87920 11744
rect 87830 11712 87842 11716
rect 87784 11706 87842 11712
rect 86310 11676 86316 11688
rect 84068 11648 85252 11676
rect 86270 11648 86316 11676
rect 84068 11636 84074 11648
rect 86310 11636 86316 11648
rect 86368 11636 86374 11688
rect 87892 11676 87920 11716
rect 88796 11712 88808 11746
rect 88842 11744 88854 11746
rect 89162 11744 89168 11756
rect 88842 11716 89168 11744
rect 88842 11712 88854 11716
rect 88796 11706 88854 11712
rect 89162 11704 89168 11716
rect 89220 11704 89226 11756
rect 100386 11744 100392 11756
rect 100346 11716 100392 11744
rect 100386 11704 100392 11716
rect 100444 11704 100450 11756
rect 100848 11746 100906 11752
rect 100848 11712 100860 11746
rect 100894 11744 100906 11746
rect 102134 11744 102140 11756
rect 100894 11716 102140 11744
rect 100894 11712 100906 11716
rect 100848 11706 100906 11712
rect 102134 11704 102140 11716
rect 102192 11704 102198 11756
rect 103148 11746 103206 11752
rect 103148 11712 103160 11746
rect 103194 11744 103206 11746
rect 103606 11744 103612 11756
rect 103194 11716 103612 11744
rect 103194 11712 103206 11716
rect 103148 11706 103206 11712
rect 103606 11704 103612 11716
rect 103664 11704 103670 11756
rect 90450 11676 90456 11688
rect 86420 11648 86954 11676
rect 87892 11648 90456 11676
rect 31168 11580 35204 11608
rect 43440 11610 43498 11616
rect 31168 11568 31174 11580
rect 43440 11576 43452 11610
rect 43486 11608 43498 11610
rect 56042 11608 56048 11620
rect 43486 11580 56048 11608
rect 43486 11576 43498 11580
rect 43440 11570 43498 11576
rect 56042 11568 56048 11580
rect 56100 11608 56106 11620
rect 86420 11608 86448 11648
rect 56100 11580 86448 11608
rect 86926 11608 86954 11648
rect 90450 11636 90456 11648
rect 90508 11636 90514 11688
rect 100754 11636 100760 11688
rect 100812 11676 100818 11688
rect 101952 11678 102010 11684
rect 101952 11676 101964 11678
rect 100812 11648 101964 11676
rect 100812 11636 100818 11648
rect 101952 11644 101964 11648
rect 101998 11644 102010 11678
rect 101952 11638 102010 11644
rect 102042 11636 102048 11688
rect 102100 11676 102106 11688
rect 102100 11648 102144 11676
rect 102100 11636 102106 11648
rect 102318 11636 102324 11688
rect 102376 11676 102382 11688
rect 103514 11676 103520 11688
rect 102376 11648 103520 11676
rect 102376 11636 102382 11648
rect 103514 11636 103520 11648
rect 103572 11636 103578 11688
rect 108224 11676 108252 11784
rect 114554 11772 114560 11784
rect 114612 11772 114618 11824
rect 138014 11812 138020 11824
rect 114940 11784 138020 11812
rect 114002 11744 114008 11756
rect 113962 11716 114008 11744
rect 114002 11704 114008 11716
rect 114060 11704 114066 11756
rect 114940 11676 114968 11784
rect 138014 11772 138020 11784
rect 138072 11772 138078 11824
rect 149974 11812 149980 11824
rect 149822 11784 149980 11812
rect 149974 11772 149980 11784
rect 150032 11772 150038 11824
rect 150912 11812 150940 11852
rect 151078 11840 151084 11852
rect 151136 11840 151142 11892
rect 151998 11880 152004 11892
rect 151958 11852 152004 11880
rect 151998 11840 152004 11852
rect 152056 11840 152062 11892
rect 152736 11882 152794 11888
rect 152736 11848 152748 11882
rect 152782 11880 152794 11882
rect 154206 11880 154212 11892
rect 152782 11852 154212 11880
rect 152782 11848 152794 11852
rect 152736 11842 152794 11848
rect 154206 11840 154212 11852
rect 154264 11840 154270 11892
rect 157306 11852 161980 11880
rect 157306 11812 157334 11852
rect 150912 11784 157334 11812
rect 115014 11704 115020 11756
rect 115072 11744 115078 11756
rect 115108 11746 115166 11752
rect 115108 11744 115120 11746
rect 115072 11716 115120 11744
rect 115072 11704 115078 11716
rect 115108 11712 115120 11716
rect 115154 11712 115166 11746
rect 116394 11744 116400 11756
rect 116354 11716 116400 11744
rect 115108 11706 115166 11712
rect 116394 11704 116400 11716
rect 116452 11704 116458 11756
rect 116856 11746 116914 11752
rect 116856 11712 116868 11746
rect 116902 11744 116914 11746
rect 117500 11746 117558 11752
rect 117500 11744 117512 11746
rect 116902 11716 117512 11744
rect 116902 11712 116914 11716
rect 116856 11706 116914 11712
rect 117500 11712 117512 11716
rect 117546 11744 117558 11746
rect 118326 11744 118332 11756
rect 117546 11716 118332 11744
rect 117546 11712 117558 11716
rect 117500 11706 117558 11712
rect 108224 11648 114968 11676
rect 115292 11678 115350 11684
rect 115292 11644 115304 11678
rect 115338 11676 115350 11678
rect 115658 11676 115664 11688
rect 115338 11648 115664 11676
rect 115338 11644 115350 11648
rect 115292 11638 115350 11644
rect 115658 11636 115664 11648
rect 115716 11636 115722 11688
rect 115750 11636 115756 11688
rect 115808 11676 115814 11688
rect 116872 11676 116900 11706
rect 118326 11704 118332 11716
rect 118384 11704 118390 11756
rect 128354 11704 128360 11756
rect 128412 11744 128418 11756
rect 129276 11746 129334 11752
rect 129276 11744 129288 11746
rect 128412 11716 129288 11744
rect 128412 11704 128418 11716
rect 129276 11712 129288 11716
rect 129322 11744 129334 11746
rect 130286 11744 130292 11756
rect 129322 11716 130292 11744
rect 129322 11712 129334 11716
rect 129276 11706 129334 11712
rect 130286 11704 130292 11716
rect 130344 11704 130350 11756
rect 130840 11746 130898 11752
rect 130840 11712 130852 11746
rect 130886 11744 130898 11746
rect 131574 11744 131580 11756
rect 130886 11716 131580 11744
rect 130886 11712 130898 11716
rect 130840 11706 130898 11712
rect 131574 11704 131580 11716
rect 131632 11704 131638 11756
rect 131668 11746 131726 11752
rect 131668 11712 131680 11746
rect 131714 11712 131726 11746
rect 131668 11706 131726 11712
rect 115808 11648 116900 11676
rect 115808 11636 115814 11648
rect 129734 11636 129740 11688
rect 129792 11676 129798 11688
rect 131022 11676 131028 11688
rect 129792 11648 131028 11676
rect 129792 11636 129798 11648
rect 131022 11636 131028 11648
rect 131080 11636 131086 11688
rect 131684 11676 131712 11706
rect 132494 11704 132500 11756
rect 132552 11744 132558 11756
rect 132588 11746 132646 11752
rect 132588 11744 132600 11746
rect 132552 11716 132600 11744
rect 132552 11704 132558 11716
rect 132588 11712 132600 11716
rect 132634 11712 132646 11746
rect 132588 11706 132646 11712
rect 147674 11704 147680 11756
rect 147732 11744 147738 11756
rect 147768 11746 147826 11752
rect 147768 11744 147780 11746
rect 147732 11716 147780 11744
rect 147732 11704 147738 11716
rect 147768 11712 147780 11716
rect 147814 11712 147826 11746
rect 151262 11744 151268 11756
rect 151222 11716 151268 11744
rect 147768 11706 147826 11712
rect 151262 11704 151268 11716
rect 151320 11704 151326 11756
rect 152182 11744 152188 11756
rect 152142 11716 152188 11744
rect 152182 11704 152188 11716
rect 152240 11704 152246 11756
rect 152644 11746 152702 11752
rect 152644 11712 152656 11746
rect 152690 11744 152702 11746
rect 152734 11744 152740 11756
rect 152690 11716 152740 11744
rect 152690 11712 152702 11716
rect 152644 11706 152702 11712
rect 152734 11704 152740 11716
rect 152792 11704 152798 11756
rect 161106 11744 161112 11756
rect 161066 11716 161112 11744
rect 161106 11704 161112 11716
rect 161164 11704 161170 11756
rect 161750 11744 161756 11756
rect 161710 11716 161756 11744
rect 161750 11704 161756 11716
rect 161808 11704 161814 11756
rect 137738 11676 137744 11688
rect 131684 11648 137744 11676
rect 137738 11636 137744 11648
rect 137796 11636 137802 11688
rect 148318 11676 148324 11688
rect 148278 11648 148324 11676
rect 148318 11636 148324 11648
rect 148376 11636 148382 11688
rect 148594 11676 148600 11688
rect 148554 11648 148600 11676
rect 148594 11636 148600 11648
rect 148652 11636 148658 11688
rect 143258 11608 143264 11620
rect 86926 11580 143264 11608
rect 56100 11568 56106 11580
rect 143258 11568 143264 11580
rect 143316 11568 143322 11620
rect 146018 11568 146024 11620
rect 146076 11608 146082 11620
rect 147584 11610 147642 11616
rect 147584 11608 147596 11610
rect 146076 11580 147596 11608
rect 146076 11568 146082 11580
rect 147584 11576 147596 11580
rect 147630 11576 147642 11610
rect 147584 11570 147642 11576
rect 160924 11610 160982 11616
rect 160924 11576 160936 11610
rect 160970 11608 160982 11610
rect 161198 11608 161204 11620
rect 160970 11580 161204 11608
rect 160970 11576 160982 11580
rect 160924 11570 160982 11576
rect 161198 11568 161204 11580
rect 161256 11568 161262 11620
rect 161290 11568 161296 11620
rect 161348 11608 161354 11620
rect 161568 11610 161626 11616
rect 161568 11608 161580 11610
rect 161348 11580 161580 11608
rect 161348 11568 161354 11580
rect 161568 11576 161580 11580
rect 161614 11576 161626 11610
rect 161952 11608 161980 11852
rect 162026 11840 162032 11892
rect 162084 11880 162090 11892
rect 162304 11882 162362 11888
rect 162304 11880 162316 11882
rect 162084 11852 162316 11880
rect 162084 11840 162090 11852
rect 162304 11848 162316 11852
rect 162350 11848 162362 11882
rect 162304 11842 162362 11848
rect 162762 11840 162768 11892
rect 162820 11880 162826 11892
rect 162948 11882 163006 11888
rect 162948 11880 162960 11882
rect 162820 11852 162960 11880
rect 162820 11840 162826 11852
rect 162948 11848 162960 11852
rect 162994 11848 163006 11882
rect 162948 11842 163006 11848
rect 163500 11882 163558 11888
rect 163500 11848 163512 11882
rect 163546 11880 163558 11882
rect 163774 11880 163780 11892
rect 163546 11852 163780 11880
rect 163546 11848 163558 11852
rect 163500 11842 163558 11848
rect 163774 11840 163780 11852
rect 163832 11840 163838 11892
rect 164236 11882 164294 11888
rect 164236 11848 164248 11882
rect 164282 11880 164294 11882
rect 164326 11880 164332 11892
rect 164282 11852 164332 11880
rect 164282 11848 164294 11852
rect 164236 11842 164294 11848
rect 164326 11840 164332 11852
rect 164384 11840 164390 11892
rect 164878 11880 164884 11892
rect 164838 11852 164884 11880
rect 164878 11840 164884 11852
rect 164936 11840 164942 11892
rect 176472 11882 176530 11888
rect 176472 11848 176484 11882
rect 176518 11880 176530 11882
rect 176746 11880 176752 11892
rect 176518 11852 176752 11880
rect 176518 11848 176530 11852
rect 176472 11842 176530 11848
rect 176746 11840 176752 11852
rect 176804 11840 176810 11892
rect 177390 11840 177396 11892
rect 177448 11880 177454 11892
rect 177576 11882 177634 11888
rect 177576 11880 177588 11882
rect 177448 11852 177588 11880
rect 177448 11840 177454 11852
rect 177576 11848 177588 11852
rect 177622 11848 177634 11882
rect 177576 11842 177634 11848
rect 177850 11840 177856 11892
rect 177908 11880 177914 11892
rect 178036 11882 178094 11888
rect 178036 11880 178048 11882
rect 177908 11852 178048 11880
rect 177908 11840 177914 11852
rect 178036 11848 178048 11852
rect 178082 11848 178094 11882
rect 178036 11842 178094 11848
rect 179140 11882 179198 11888
rect 179140 11848 179152 11882
rect 179186 11880 179198 11882
rect 179874 11880 179880 11892
rect 179186 11852 179880 11880
rect 179186 11848 179198 11852
rect 179140 11842 179198 11848
rect 179874 11840 179880 11852
rect 179932 11840 179938 11892
rect 179966 11840 179972 11892
rect 180024 11880 180030 11892
rect 180060 11882 180118 11888
rect 180060 11880 180072 11882
rect 180024 11852 180072 11880
rect 180024 11840 180030 11852
rect 180060 11848 180072 11852
rect 180106 11848 180118 11882
rect 180060 11842 180118 11848
rect 180150 11840 180156 11892
rect 180208 11880 180214 11892
rect 188338 11880 188344 11892
rect 180208 11852 188344 11880
rect 180208 11840 180214 11852
rect 188338 11840 188344 11852
rect 188396 11840 188402 11892
rect 190824 11882 190882 11888
rect 190824 11848 190836 11882
rect 190870 11880 190882 11882
rect 191742 11880 191748 11892
rect 190870 11852 191748 11880
rect 190870 11848 190882 11852
rect 190824 11842 190882 11848
rect 191742 11840 191748 11852
rect 191800 11840 191806 11892
rect 191834 11840 191840 11892
rect 191892 11880 191898 11892
rect 194410 11880 194416 11892
rect 191892 11852 194416 11880
rect 191892 11840 191898 11852
rect 162578 11772 162584 11824
rect 162636 11812 162642 11824
rect 189534 11812 189540 11824
rect 162636 11784 189540 11812
rect 162636 11772 162642 11784
rect 189534 11772 189540 11784
rect 189592 11772 189598 11824
rect 193858 11812 193864 11824
rect 193338 11784 193864 11812
rect 193858 11772 193864 11784
rect 193916 11772 193922 11824
rect 162212 11746 162270 11752
rect 162212 11712 162224 11746
rect 162258 11744 162270 11746
rect 162856 11746 162914 11752
rect 162856 11744 162868 11746
rect 162258 11716 162868 11744
rect 162258 11712 162270 11716
rect 162212 11706 162270 11712
rect 162856 11712 162868 11716
rect 162902 11712 162914 11746
rect 163682 11744 163688 11756
rect 163642 11716 163688 11744
rect 162856 11706 162914 11712
rect 162872 11676 162900 11706
rect 163682 11704 163688 11716
rect 163740 11704 163746 11756
rect 164144 11746 164202 11752
rect 164144 11712 164156 11746
rect 164190 11744 164202 11746
rect 164788 11746 164846 11752
rect 164788 11744 164800 11746
rect 164190 11716 164800 11744
rect 164190 11712 164202 11716
rect 164144 11706 164202 11712
rect 164788 11712 164800 11716
rect 164834 11744 164846 11746
rect 166626 11744 166632 11756
rect 164834 11716 166632 11744
rect 164834 11712 164846 11716
rect 164788 11706 164846 11712
rect 163498 11676 163504 11688
rect 162872 11648 163504 11676
rect 163498 11636 163504 11648
rect 163556 11676 163562 11688
rect 164160 11676 164188 11706
rect 166626 11704 166632 11716
rect 166684 11704 166690 11756
rect 176654 11744 176660 11756
rect 176614 11716 176660 11744
rect 176654 11704 176660 11716
rect 176712 11704 176718 11756
rect 177944 11746 178002 11752
rect 177944 11712 177956 11746
rect 177990 11744 178002 11746
rect 179232 11746 179290 11752
rect 179232 11744 179244 11746
rect 177990 11716 179244 11744
rect 177990 11712 178002 11716
rect 177944 11706 178002 11712
rect 179232 11712 179244 11716
rect 179278 11744 179290 11746
rect 179874 11744 179880 11756
rect 179278 11716 179880 11744
rect 179278 11712 179290 11716
rect 179232 11706 179290 11712
rect 179874 11704 179880 11716
rect 179932 11704 179938 11756
rect 179968 11746 180026 11752
rect 179968 11712 179980 11746
rect 180014 11712 180026 11746
rect 179968 11706 180026 11712
rect 163556 11648 164188 11676
rect 163556 11636 163562 11648
rect 177114 11636 177120 11688
rect 177172 11676 177178 11688
rect 178128 11678 178186 11684
rect 178128 11676 178140 11678
rect 177172 11648 178140 11676
rect 177172 11636 177178 11648
rect 178128 11644 178140 11648
rect 178174 11676 178186 11678
rect 179324 11678 179382 11684
rect 179324 11676 179336 11678
rect 178174 11648 179336 11676
rect 178174 11644 178186 11648
rect 178128 11638 178186 11644
rect 165890 11608 165896 11620
rect 161952 11580 165896 11608
rect 161568 11570 161626 11576
rect 165890 11568 165896 11580
rect 165948 11568 165954 11620
rect 31386 11540 31392 11552
rect 29748 11512 30972 11540
rect 31346 11512 31392 11540
rect 31386 11500 31392 11512
rect 31444 11500 31450 11552
rect 32124 11542 32182 11548
rect 32124 11508 32136 11542
rect 32170 11540 32182 11542
rect 32950 11540 32956 11552
rect 32170 11512 32956 11540
rect 32170 11508 32182 11512
rect 32124 11502 32182 11508
rect 32950 11500 32956 11512
rect 33008 11500 33014 11552
rect 54940 11542 54998 11548
rect 54940 11508 54952 11542
rect 54986 11540 54998 11542
rect 55490 11540 55496 11552
rect 54986 11512 55496 11540
rect 54986 11508 54998 11512
rect 54940 11502 54998 11508
rect 55490 11500 55496 11512
rect 55548 11500 55554 11552
rect 84838 11500 84844 11552
rect 84896 11540 84902 11552
rect 85024 11542 85082 11548
rect 85024 11540 85036 11542
rect 84896 11512 85036 11540
rect 84896 11500 84902 11512
rect 85024 11508 85036 11512
rect 85070 11508 85082 11542
rect 85024 11502 85082 11508
rect 85668 11542 85726 11548
rect 85668 11508 85680 11542
rect 85714 11540 85726 11542
rect 86402 11540 86408 11552
rect 85714 11512 86408 11540
rect 85714 11508 85726 11512
rect 85668 11502 85726 11508
rect 86402 11500 86408 11512
rect 86460 11500 86466 11552
rect 101492 11542 101550 11548
rect 101492 11508 101504 11542
rect 101538 11540 101550 11542
rect 101858 11540 101864 11552
rect 101538 11512 101864 11540
rect 101538 11508 101550 11512
rect 101492 11502 101550 11508
rect 101858 11500 101864 11512
rect 101916 11500 101922 11552
rect 102964 11542 103022 11548
rect 102964 11508 102976 11542
rect 103010 11540 103022 11542
rect 104066 11540 104072 11552
rect 103010 11512 104072 11540
rect 103010 11508 103022 11512
rect 102964 11502 103022 11508
rect 104066 11500 104072 11512
rect 104124 11500 104130 11552
rect 114002 11500 114008 11552
rect 114060 11540 114066 11552
rect 114648 11542 114706 11548
rect 114648 11540 114660 11542
rect 114060 11512 114660 11540
rect 114060 11500 114066 11512
rect 114648 11508 114660 11512
rect 114694 11508 114706 11542
rect 131850 11540 131856 11552
rect 131810 11512 131856 11540
rect 114648 11502 114706 11508
rect 131850 11500 131856 11512
rect 131908 11500 131914 11552
rect 147306 11500 147312 11552
rect 147364 11540 147370 11552
rect 150068 11542 150126 11548
rect 150068 11540 150080 11542
rect 147364 11512 150080 11540
rect 147364 11500 147370 11512
rect 150068 11508 150080 11512
rect 150114 11540 150126 11542
rect 151722 11540 151728 11552
rect 150114 11512 151728 11540
rect 150114 11508 150126 11512
rect 150068 11502 150126 11508
rect 151722 11500 151728 11512
rect 151780 11500 151786 11552
rect 178696 11540 178724 11648
rect 179324 11644 179336 11648
rect 179370 11644 179382 11678
rect 179984 11676 180012 11706
rect 180058 11704 180064 11756
rect 180116 11744 180122 11756
rect 180610 11744 180616 11756
rect 180116 11716 180616 11744
rect 180116 11704 180122 11716
rect 180610 11704 180616 11716
rect 180668 11704 180674 11756
rect 180794 11676 180800 11688
rect 179984 11648 180800 11676
rect 179324 11638 179382 11644
rect 180794 11636 180800 11648
rect 180852 11676 180858 11688
rect 181530 11676 181536 11688
rect 180852 11648 181536 11676
rect 180852 11636 180858 11648
rect 181530 11636 181536 11648
rect 181588 11636 181594 11688
rect 189552 11676 189580 11772
rect 189626 11704 189632 11756
rect 189684 11744 189690 11756
rect 190088 11746 190146 11752
rect 189684 11716 189728 11744
rect 189684 11704 189690 11716
rect 190088 11712 190100 11746
rect 190134 11744 190146 11746
rect 190732 11746 190790 11752
rect 190732 11744 190744 11746
rect 190134 11716 190744 11744
rect 190134 11712 190146 11716
rect 190088 11706 190146 11712
rect 190732 11712 190744 11716
rect 190778 11744 190790 11746
rect 190822 11744 190828 11756
rect 190778 11716 190828 11744
rect 190778 11712 190790 11716
rect 190732 11706 190790 11712
rect 190104 11676 190132 11706
rect 190822 11704 190828 11716
rect 190880 11704 190886 11756
rect 191834 11744 191840 11756
rect 191794 11716 191840 11744
rect 191834 11704 191840 11716
rect 191892 11704 191898 11756
rect 194060 11752 194088 11852
rect 194410 11840 194416 11852
rect 194468 11840 194474 11892
rect 194686 11840 194692 11892
rect 194744 11880 194750 11892
rect 196252 11882 196310 11888
rect 196252 11880 196264 11882
rect 194744 11852 196264 11880
rect 194744 11840 194750 11852
rect 196252 11848 196264 11852
rect 196298 11848 196310 11882
rect 202874 11880 202880 11892
rect 202834 11852 202880 11880
rect 196252 11842 196310 11848
rect 202874 11840 202880 11852
rect 202932 11840 202938 11892
rect 204072 11882 204130 11888
rect 204072 11848 204084 11882
rect 204118 11880 204130 11882
rect 204530 11880 204536 11892
rect 204118 11852 204536 11880
rect 204118 11848 204130 11852
rect 204072 11842 204130 11848
rect 204530 11840 204536 11852
rect 204588 11840 204594 11892
rect 205176 11882 205234 11888
rect 205176 11848 205188 11882
rect 205222 11880 205234 11882
rect 206554 11880 206560 11892
rect 205222 11852 206560 11880
rect 205222 11848 205234 11852
rect 205176 11842 205234 11848
rect 206554 11840 206560 11852
rect 206612 11840 206618 11892
rect 227806 11840 227812 11892
rect 227864 11880 227870 11892
rect 228268 11882 228326 11888
rect 228268 11880 228280 11882
rect 227864 11852 228280 11880
rect 227864 11840 227870 11852
rect 228268 11848 228280 11852
rect 228314 11880 228326 11882
rect 228818 11880 228824 11892
rect 228314 11852 228824 11880
rect 228314 11848 228326 11852
rect 228268 11842 228326 11848
rect 228818 11840 228824 11852
rect 228876 11880 228882 11892
rect 229464 11882 229522 11888
rect 228876 11852 229094 11880
rect 228876 11840 228882 11852
rect 196802 11812 196808 11824
rect 195546 11784 196808 11812
rect 196802 11772 196808 11784
rect 196860 11772 196866 11824
rect 202324 11814 202382 11820
rect 202324 11780 202336 11814
rect 202370 11812 202382 11814
rect 203150 11812 203156 11824
rect 202370 11784 203156 11812
rect 202370 11780 202382 11784
rect 202324 11774 202382 11780
rect 203150 11772 203156 11784
rect 203208 11772 203214 11824
rect 203980 11814 204038 11820
rect 203980 11780 203992 11814
rect 204026 11812 204038 11814
rect 205268 11814 205326 11820
rect 205268 11812 205280 11814
rect 204026 11784 205280 11812
rect 204026 11780 204038 11784
rect 203980 11774 204038 11780
rect 205268 11780 205280 11784
rect 205314 11812 205326 11814
rect 205542 11812 205548 11824
rect 205314 11784 205548 11812
rect 205314 11780 205326 11784
rect 205268 11774 205326 11780
rect 205542 11772 205548 11784
rect 205600 11772 205606 11824
rect 227714 11772 227720 11824
rect 227772 11812 227778 11824
rect 228360 11814 228418 11820
rect 228360 11812 228372 11814
rect 227772 11784 228372 11812
rect 227772 11772 227778 11784
rect 228360 11780 228372 11784
rect 228406 11780 228418 11814
rect 229066 11812 229094 11852
rect 229464 11848 229476 11882
rect 229510 11880 229522 11882
rect 229922 11880 229928 11892
rect 229510 11852 229928 11880
rect 229510 11848 229522 11852
rect 229464 11842 229522 11848
rect 229922 11840 229928 11852
rect 229980 11840 229986 11892
rect 230382 11880 230388 11892
rect 230342 11852 230388 11880
rect 230382 11840 230388 11852
rect 230440 11840 230446 11892
rect 231026 11840 231032 11892
rect 231084 11880 231090 11892
rect 231580 11882 231638 11888
rect 231580 11880 231592 11882
rect 231084 11852 231592 11880
rect 231084 11840 231090 11852
rect 231580 11848 231592 11852
rect 231626 11848 231638 11882
rect 231580 11842 231638 11848
rect 231670 11840 231676 11892
rect 231728 11880 231734 11892
rect 238756 11882 238814 11888
rect 238756 11880 238768 11882
rect 231728 11852 238768 11880
rect 231728 11840 231734 11852
rect 238756 11848 238768 11852
rect 238802 11848 238814 11882
rect 240318 11880 240324 11892
rect 240278 11852 240324 11880
rect 238756 11842 238814 11848
rect 240318 11840 240324 11852
rect 240376 11840 240382 11892
rect 241054 11880 241060 11892
rect 241014 11852 241060 11880
rect 241054 11840 241060 11852
rect 241112 11840 241118 11892
rect 241790 11880 241796 11892
rect 241750 11852 241796 11880
rect 241790 11840 241796 11852
rect 241848 11840 241854 11892
rect 251820 11882 251878 11888
rect 251820 11848 251832 11882
rect 251866 11880 251878 11882
rect 252922 11880 252928 11892
rect 251866 11852 252928 11880
rect 251866 11848 251878 11852
rect 251820 11842 251878 11848
rect 252922 11840 252928 11852
rect 252980 11840 252986 11892
rect 254120 11882 254178 11888
rect 254120 11848 254132 11882
rect 254166 11880 254178 11882
rect 254670 11880 254676 11892
rect 254166 11852 254676 11880
rect 254166 11848 254178 11852
rect 254120 11842 254178 11848
rect 254670 11840 254676 11852
rect 254728 11840 254734 11892
rect 254762 11840 254768 11892
rect 254820 11880 254826 11892
rect 254948 11882 255006 11888
rect 254948 11880 254960 11882
rect 254820 11852 254960 11880
rect 254820 11840 254826 11852
rect 254948 11848 254960 11852
rect 254994 11848 255006 11882
rect 254948 11842 255006 11848
rect 255038 11840 255044 11892
rect 255096 11880 255102 11892
rect 255592 11882 255650 11888
rect 255592 11880 255604 11882
rect 255096 11852 255604 11880
rect 255096 11840 255102 11852
rect 255592 11848 255604 11852
rect 255638 11848 255650 11882
rect 255592 11842 255650 11848
rect 264976 11882 265034 11888
rect 264976 11848 264988 11882
rect 265022 11880 265034 11882
rect 266814 11880 266820 11892
rect 265022 11852 266820 11880
rect 265022 11848 265034 11852
rect 264976 11842 265034 11848
rect 266814 11840 266820 11852
rect 266872 11840 266878 11892
rect 267368 11882 267426 11888
rect 267368 11848 267380 11882
rect 267414 11880 267426 11882
rect 268196 11882 268254 11888
rect 267414 11852 267734 11880
rect 267414 11848 267426 11852
rect 267368 11842 267426 11848
rect 229556 11814 229614 11820
rect 229556 11812 229568 11814
rect 229066 11784 229568 11812
rect 228360 11774 228418 11780
rect 229556 11780 229568 11784
rect 229602 11780 229614 11814
rect 229556 11774 229614 11780
rect 194044 11746 194102 11752
rect 194044 11712 194056 11746
rect 194090 11712 194102 11746
rect 194044 11706 194102 11712
rect 196436 11746 196494 11752
rect 196436 11712 196448 11746
rect 196482 11744 196494 11746
rect 197906 11744 197912 11756
rect 196482 11716 197912 11744
rect 196482 11712 196494 11716
rect 196436 11706 196494 11712
rect 197906 11704 197912 11716
rect 197964 11704 197970 11756
rect 201034 11704 201040 11756
rect 201092 11744 201098 11756
rect 202232 11746 202290 11752
rect 202232 11744 202244 11746
rect 201092 11716 202244 11744
rect 201092 11704 201098 11716
rect 202232 11712 202244 11716
rect 202278 11712 202290 11746
rect 203058 11744 203064 11756
rect 203018 11716 203064 11744
rect 202232 11706 202290 11712
rect 203058 11704 203064 11716
rect 203116 11704 203122 11756
rect 206370 11744 206376 11756
rect 203168 11716 206376 11744
rect 192110 11676 192116 11688
rect 189552 11648 190132 11676
rect 192070 11648 192116 11676
rect 192110 11636 192116 11648
rect 192168 11636 192174 11688
rect 194318 11676 194324 11688
rect 194278 11648 194324 11676
rect 194318 11636 194324 11648
rect 194376 11636 194382 11688
rect 194410 11636 194416 11688
rect 194468 11676 194474 11688
rect 195792 11678 195850 11684
rect 194468 11648 195376 11676
rect 194468 11636 194474 11648
rect 178772 11610 178830 11616
rect 178772 11576 178784 11610
rect 178818 11608 178830 11610
rect 180334 11608 180340 11620
rect 178818 11580 180340 11608
rect 178818 11576 178830 11580
rect 178772 11570 178830 11576
rect 180334 11568 180340 11580
rect 180392 11568 180398 11620
rect 190180 11610 190238 11616
rect 190180 11576 190192 11610
rect 190226 11608 190238 11610
rect 195348 11608 195376 11648
rect 195792 11644 195804 11678
rect 195838 11676 195850 11678
rect 197354 11676 197360 11688
rect 195838 11648 197360 11676
rect 195838 11644 195850 11648
rect 195792 11638 195850 11644
rect 197354 11636 197360 11648
rect 197412 11676 197418 11688
rect 201310 11676 201316 11688
rect 197412 11648 201316 11676
rect 197412 11636 197418 11648
rect 201310 11636 201316 11648
rect 201368 11636 201374 11688
rect 202874 11636 202880 11688
rect 202932 11676 202938 11688
rect 203168 11676 203196 11716
rect 206370 11704 206376 11716
rect 206428 11704 206434 11756
rect 228376 11744 228404 11774
rect 230842 11772 230848 11824
rect 230900 11812 230906 11824
rect 238664 11814 238722 11820
rect 230900 11784 231072 11812
rect 230900 11772 230906 11784
rect 229370 11744 229376 11756
rect 228376 11716 229376 11744
rect 229370 11704 229376 11716
rect 229428 11704 229434 11756
rect 231044 11752 231072 11784
rect 238664 11780 238676 11814
rect 238710 11812 238722 11814
rect 240134 11812 240140 11824
rect 238710 11784 240140 11812
rect 238710 11780 238722 11784
rect 238664 11774 238722 11780
rect 240134 11772 240140 11784
rect 240192 11772 240198 11824
rect 241514 11812 241520 11824
rect 240244 11784 241520 11812
rect 230292 11746 230350 11752
rect 230292 11712 230304 11746
rect 230338 11744 230350 11746
rect 230936 11746 230994 11752
rect 230936 11744 230948 11746
rect 230338 11716 230948 11744
rect 230338 11712 230350 11716
rect 230292 11706 230350 11712
rect 230936 11712 230948 11716
rect 230982 11712 230994 11746
rect 230936 11706 230994 11712
rect 231028 11746 231086 11752
rect 231028 11712 231040 11746
rect 231074 11712 231086 11746
rect 231028 11706 231086 11712
rect 202932 11648 203196 11676
rect 202932 11636 202938 11648
rect 203518 11636 203524 11688
rect 203576 11676 203582 11688
rect 204256 11678 204314 11684
rect 204256 11676 204268 11678
rect 203576 11648 204268 11676
rect 203576 11636 203582 11648
rect 204256 11644 204268 11648
rect 204302 11676 204314 11678
rect 205452 11678 205510 11684
rect 205452 11676 205464 11678
rect 204302 11648 205464 11676
rect 204302 11644 204314 11648
rect 204256 11638 204314 11644
rect 205452 11644 205464 11648
rect 205498 11676 205510 11678
rect 207842 11676 207848 11688
rect 205498 11648 207848 11676
rect 205498 11644 205510 11648
rect 205452 11638 205510 11644
rect 207842 11636 207848 11648
rect 207900 11636 207906 11688
rect 227254 11636 227260 11688
rect 227312 11676 227318 11688
rect 228452 11678 228510 11684
rect 228452 11676 228464 11678
rect 227312 11648 228464 11676
rect 227312 11636 227318 11648
rect 228452 11644 228464 11648
rect 228498 11676 228510 11678
rect 229740 11678 229798 11684
rect 229740 11676 229752 11678
rect 228498 11648 229752 11676
rect 228498 11644 228510 11648
rect 228452 11638 228510 11644
rect 229740 11644 229752 11648
rect 229786 11676 229798 11678
rect 229786 11648 230888 11676
rect 229786 11644 229798 11648
rect 229740 11638 229798 11644
rect 197446 11608 197452 11620
rect 190226 11580 191972 11608
rect 195348 11580 197452 11608
rect 190226 11576 190238 11580
rect 190180 11570 190238 11576
rect 180518 11540 180524 11552
rect 178696 11512 180524 11540
rect 180518 11500 180524 11512
rect 180576 11500 180582 11552
rect 189442 11540 189448 11552
rect 189402 11512 189448 11540
rect 189442 11500 189448 11512
rect 189500 11500 189506 11552
rect 191944 11540 191972 11580
rect 197446 11568 197452 11580
rect 197504 11568 197510 11620
rect 203426 11568 203432 11620
rect 203484 11608 203490 11620
rect 204898 11608 204904 11620
rect 203484 11580 204904 11608
rect 203484 11568 203490 11580
rect 204898 11568 204904 11580
rect 204956 11568 204962 11620
rect 227900 11610 227958 11616
rect 227900 11576 227912 11610
rect 227946 11608 227958 11610
rect 230290 11608 230296 11620
rect 227946 11580 230296 11608
rect 227946 11576 227958 11580
rect 227900 11570 227958 11576
rect 230290 11568 230296 11580
rect 230348 11568 230354 11620
rect 193306 11540 193312 11552
rect 191944 11512 193312 11540
rect 193306 11500 193312 11512
rect 193364 11500 193370 11552
rect 193490 11500 193496 11552
rect 193548 11540 193554 11552
rect 193584 11542 193642 11548
rect 193584 11540 193596 11542
rect 193548 11512 193596 11540
rect 193548 11500 193554 11512
rect 193584 11508 193596 11512
rect 193630 11540 193642 11542
rect 195790 11540 195796 11552
rect 193630 11512 195796 11540
rect 193630 11508 193642 11512
rect 193584 11502 193642 11508
rect 195790 11500 195796 11512
rect 195848 11500 195854 11552
rect 195882 11500 195888 11552
rect 195940 11540 195946 11552
rect 196986 11540 196992 11552
rect 195940 11512 196992 11540
rect 195940 11500 195946 11512
rect 196986 11500 196992 11512
rect 197044 11500 197050 11552
rect 201494 11500 201500 11552
rect 201552 11540 201558 11552
rect 203612 11542 203670 11548
rect 203612 11540 203624 11542
rect 201552 11512 203624 11540
rect 201552 11500 201558 11512
rect 203612 11508 203624 11512
rect 203658 11508 203670 11542
rect 204806 11540 204812 11552
rect 204766 11512 204812 11540
rect 203612 11502 203670 11508
rect 204806 11500 204812 11512
rect 204864 11500 204870 11552
rect 229096 11542 229154 11548
rect 229096 11508 229108 11542
rect 229142 11540 229154 11542
rect 229370 11540 229376 11552
rect 229142 11512 229376 11540
rect 229142 11508 229154 11512
rect 229096 11502 229154 11508
rect 229370 11500 229376 11512
rect 229428 11500 229434 11552
rect 230860 11540 230888 11648
rect 230952 11608 230980 11706
rect 231210 11704 231216 11756
rect 231268 11744 231274 11756
rect 240244 11752 240272 11784
rect 241514 11772 241520 11784
rect 241572 11772 241578 11824
rect 244826 11812 244832 11824
rect 242636 11784 244832 11812
rect 231764 11746 231822 11752
rect 231764 11744 231776 11746
rect 231268 11716 231776 11744
rect 231268 11704 231274 11716
rect 231764 11712 231776 11716
rect 231810 11712 231822 11746
rect 231764 11706 231822 11712
rect 240228 11746 240286 11752
rect 240228 11712 240240 11746
rect 240274 11712 240286 11746
rect 241240 11746 241298 11752
rect 241240 11744 241252 11746
rect 240228 11706 240286 11712
rect 240612 11716 241252 11744
rect 239306 11636 239312 11688
rect 239364 11676 239370 11688
rect 239950 11676 239956 11688
rect 239364 11648 239956 11676
rect 239364 11636 239370 11648
rect 239950 11636 239956 11648
rect 240008 11676 240014 11688
rect 240412 11678 240470 11684
rect 240412 11676 240424 11678
rect 240008 11648 240424 11676
rect 240008 11636 240014 11648
rect 240412 11644 240424 11648
rect 240458 11644 240470 11678
rect 240412 11638 240470 11644
rect 232130 11608 232136 11620
rect 230952 11580 232136 11608
rect 232130 11568 232136 11580
rect 232188 11568 232194 11620
rect 239860 11610 239918 11616
rect 239860 11576 239872 11610
rect 239906 11608 239918 11610
rect 240612 11608 240640 11716
rect 241240 11712 241252 11716
rect 241286 11712 241298 11746
rect 241240 11706 241298 11712
rect 241700 11746 241758 11752
rect 241700 11712 241712 11746
rect 241746 11712 241758 11746
rect 242526 11744 242532 11756
rect 242486 11716 242532 11744
rect 241700 11706 241758 11712
rect 241716 11676 241744 11706
rect 242526 11704 242532 11716
rect 242584 11704 242590 11756
rect 241974 11676 241980 11688
rect 241716 11648 241980 11676
rect 241974 11636 241980 11648
rect 242032 11676 242038 11688
rect 242636 11676 242664 11784
rect 244826 11772 244832 11784
rect 244884 11772 244890 11824
rect 254028 11814 254086 11820
rect 254028 11780 254040 11814
rect 254074 11812 254086 11814
rect 254302 11812 254308 11824
rect 254074 11784 254308 11812
rect 254074 11780 254086 11784
rect 254028 11774 254086 11780
rect 254302 11772 254308 11784
rect 254360 11772 254366 11824
rect 264424 11814 264482 11820
rect 264424 11780 264436 11814
rect 264470 11812 264482 11814
rect 267706 11812 267734 11852
rect 268196 11848 268208 11882
rect 268242 11880 268254 11882
rect 270678 11880 270684 11892
rect 268242 11852 270684 11880
rect 268242 11848 268254 11852
rect 268196 11842 268254 11848
rect 270678 11840 270684 11852
rect 270736 11840 270742 11892
rect 270770 11840 270776 11892
rect 270828 11880 270834 11892
rect 271416 11882 271474 11888
rect 271416 11880 271428 11882
rect 270828 11852 271428 11880
rect 270828 11840 270834 11852
rect 271416 11848 271428 11852
rect 271462 11848 271474 11882
rect 271416 11842 271474 11848
rect 268286 11812 268292 11824
rect 264470 11784 266386 11812
rect 267706 11784 268292 11812
rect 264470 11780 264482 11784
rect 264424 11774 264482 11780
rect 268286 11772 268292 11784
rect 268344 11772 268350 11824
rect 269850 11772 269856 11824
rect 269908 11772 269914 11824
rect 252002 11744 252008 11756
rect 251962 11716 252008 11744
rect 252002 11704 252008 11716
rect 252060 11704 252066 11756
rect 252372 11746 252430 11752
rect 252372 11712 252384 11746
rect 252418 11744 252430 11746
rect 252738 11744 252744 11756
rect 252418 11716 252744 11744
rect 252418 11712 252430 11716
rect 252372 11706 252430 11712
rect 252738 11704 252744 11716
rect 252796 11704 252802 11756
rect 253014 11704 253020 11756
rect 253072 11744 253078 11756
rect 254856 11746 254914 11752
rect 254856 11744 254868 11746
rect 253072 11716 254868 11744
rect 253072 11704 253078 11716
rect 254856 11712 254868 11716
rect 254902 11744 254914 11746
rect 255500 11746 255558 11752
rect 255500 11744 255512 11746
rect 254902 11716 255512 11744
rect 254902 11712 254914 11716
rect 254856 11706 254914 11712
rect 255500 11712 255512 11716
rect 255546 11744 255558 11746
rect 256234 11744 256240 11756
rect 255546 11716 256240 11744
rect 255546 11712 255558 11716
rect 255500 11706 255558 11712
rect 256234 11704 256240 11716
rect 256292 11744 256298 11756
rect 257246 11744 257252 11756
rect 256292 11716 257252 11744
rect 256292 11704 256298 11716
rect 257246 11704 257252 11716
rect 257304 11704 257310 11756
rect 264330 11744 264336 11756
rect 264290 11716 264336 11744
rect 264330 11704 264336 11716
rect 264388 11704 264394 11756
rect 265158 11744 265164 11756
rect 265118 11716 265164 11744
rect 265158 11704 265164 11716
rect 265216 11704 265222 11756
rect 265250 11704 265256 11756
rect 265308 11744 265314 11756
rect 265620 11746 265678 11752
rect 265620 11744 265632 11746
rect 265308 11716 265632 11744
rect 265308 11704 265314 11716
rect 265620 11712 265632 11716
rect 265666 11712 265678 11746
rect 268470 11744 268476 11756
rect 265620 11706 265678 11712
rect 268304 11716 268476 11744
rect 242032 11648 242664 11676
rect 242032 11636 242038 11648
rect 242710 11636 242716 11688
rect 242768 11676 242774 11688
rect 244550 11676 244556 11688
rect 242768 11648 244556 11676
rect 242768 11636 242774 11648
rect 244550 11636 244556 11648
rect 244608 11636 244614 11688
rect 252094 11636 252100 11688
rect 252152 11676 252158 11688
rect 254212 11678 254270 11684
rect 254212 11676 254224 11678
rect 252152 11648 254224 11676
rect 252152 11636 252158 11648
rect 254212 11644 254224 11648
rect 254258 11676 254270 11678
rect 255590 11676 255596 11688
rect 254258 11648 255596 11676
rect 254258 11644 254270 11648
rect 254212 11638 254270 11644
rect 255590 11636 255596 11648
rect 255648 11676 255654 11688
rect 256418 11676 256424 11688
rect 255648 11648 256424 11676
rect 255648 11636 255654 11648
rect 256418 11636 256424 11648
rect 256476 11636 256482 11688
rect 263962 11636 263968 11688
rect 264020 11676 264026 11688
rect 268304 11684 268332 11716
rect 268470 11704 268476 11716
rect 268528 11704 268534 11756
rect 269114 11744 269120 11756
rect 269074 11716 269120 11744
rect 269114 11704 269120 11716
rect 269172 11704 269178 11756
rect 271322 11744 271328 11756
rect 271282 11716 271328 11744
rect 271322 11704 271328 11716
rect 271380 11704 271386 11756
rect 265896 11678 265954 11684
rect 265896 11676 265908 11678
rect 264020 11648 265908 11676
rect 264020 11636 264026 11648
rect 265896 11644 265908 11648
rect 265942 11644 265954 11678
rect 265896 11638 265954 11644
rect 268288 11678 268346 11684
rect 268288 11644 268300 11678
rect 268334 11644 268346 11678
rect 268288 11638 268346 11644
rect 268380 11678 268438 11684
rect 268380 11644 268392 11678
rect 268426 11644 268438 11678
rect 268380 11638 268438 11644
rect 239906 11580 240640 11608
rect 240704 11580 248414 11608
rect 239906 11576 239918 11580
rect 239860 11570 239918 11576
rect 231670 11540 231676 11552
rect 230860 11512 231676 11540
rect 231670 11500 231676 11512
rect 231728 11500 231734 11552
rect 239398 11500 239404 11552
rect 239456 11540 239462 11552
rect 240704 11540 240732 11580
rect 239456 11512 240732 11540
rect 239456 11500 239462 11512
rect 241238 11500 241244 11552
rect 241296 11540 241302 11552
rect 242344 11542 242402 11548
rect 242344 11540 242356 11542
rect 241296 11512 242356 11540
rect 241296 11500 241302 11512
rect 242344 11508 242356 11512
rect 242390 11508 242402 11542
rect 248386 11540 248414 11580
rect 251634 11568 251640 11620
rect 251692 11608 251698 11620
rect 252924 11610 252982 11616
rect 252924 11608 252936 11610
rect 251692 11580 252936 11608
rect 251692 11568 251698 11580
rect 252924 11576 252936 11580
rect 252970 11608 252982 11610
rect 252970 11580 260834 11608
rect 252970 11576 252982 11580
rect 252924 11570 252982 11576
rect 249058 11540 249064 11552
rect 248386 11512 249064 11540
rect 242344 11502 242402 11508
rect 249058 11500 249064 11512
rect 249116 11500 249122 11552
rect 253290 11500 253296 11552
rect 253348 11540 253354 11552
rect 253660 11542 253718 11548
rect 253660 11540 253672 11542
rect 253348 11512 253672 11540
rect 253348 11500 253354 11512
rect 253660 11508 253672 11512
rect 253706 11508 253718 11542
rect 260806 11540 260834 11580
rect 268010 11568 268016 11620
rect 268068 11608 268074 11620
rect 268396 11608 268424 11638
rect 268068 11580 268424 11608
rect 268068 11568 268074 11580
rect 261754 11540 261760 11552
rect 260806 11512 261760 11540
rect 253660 11502 253718 11508
rect 261754 11500 261760 11512
rect 261812 11500 261818 11552
rect 262674 11500 262680 11552
rect 262732 11540 262738 11552
rect 266262 11540 266268 11552
rect 262732 11512 266268 11540
rect 262732 11500 262738 11512
rect 266262 11500 266268 11512
rect 266320 11500 266326 11552
rect 266354 11500 266360 11552
rect 266412 11540 266418 11552
rect 267828 11542 267886 11548
rect 267828 11540 267840 11542
rect 266412 11512 267840 11540
rect 266412 11500 266418 11512
rect 267828 11508 267840 11512
rect 267874 11508 267886 11542
rect 268488 11540 268516 11704
rect 269390 11676 269396 11688
rect 269350 11648 269396 11676
rect 269390 11636 269396 11648
rect 269448 11636 269454 11688
rect 269942 11636 269948 11688
rect 270000 11676 270006 11688
rect 270864 11678 270922 11684
rect 270864 11676 270876 11678
rect 270000 11648 270876 11676
rect 270000 11636 270006 11648
rect 270864 11644 270876 11648
rect 270910 11676 270922 11678
rect 273162 11676 273168 11688
rect 270910 11648 273168 11676
rect 270910 11644 270922 11648
rect 270864 11638 270922 11644
rect 273162 11636 273168 11648
rect 273220 11636 273226 11688
rect 275094 11540 275100 11552
rect 268488 11512 275100 11540
rect 267828 11502 267886 11508
rect 275094 11500 275100 11512
rect 275152 11500 275158 11552
rect 1104 11450 305808 11472
rect 1104 11398 39048 11450
rect 39100 11398 39112 11450
rect 39164 11398 39176 11450
rect 39228 11398 39240 11450
rect 39292 11398 39304 11450
rect 39356 11398 115246 11450
rect 115298 11398 115310 11450
rect 115362 11398 115374 11450
rect 115426 11398 115438 11450
rect 115490 11398 115502 11450
rect 115554 11398 191444 11450
rect 191496 11398 191508 11450
rect 191560 11398 191572 11450
rect 191624 11398 191636 11450
rect 191688 11398 191700 11450
rect 191752 11398 267642 11450
rect 267694 11398 267706 11450
rect 267758 11398 267770 11450
rect 267822 11398 267834 11450
rect 267886 11398 267898 11450
rect 267950 11398 305808 11450
rect 1104 11376 305808 11398
rect 28812 11338 28870 11344
rect 28812 11304 28824 11338
rect 28858 11336 28870 11338
rect 29914 11336 29920 11348
rect 28858 11308 29920 11336
rect 28858 11304 28870 11308
rect 28812 11298 28870 11304
rect 29914 11296 29920 11308
rect 29972 11296 29978 11348
rect 30006 11296 30012 11348
rect 30064 11336 30070 11348
rect 30064 11308 31754 11336
rect 30064 11296 30070 11308
rect 28902 11228 28908 11280
rect 28960 11268 28966 11280
rect 31726 11268 31754 11308
rect 32398 11296 32404 11348
rect 32456 11336 32462 11348
rect 33318 11336 33324 11348
rect 32456 11308 33324 11336
rect 32456 11296 32462 11308
rect 33318 11296 33324 11308
rect 33376 11296 33382 11348
rect 33594 11336 33600 11348
rect 33554 11308 33600 11336
rect 33594 11296 33600 11308
rect 33652 11296 33658 11348
rect 40312 11338 40370 11344
rect 40312 11304 40324 11338
rect 40358 11336 40370 11338
rect 40402 11336 40408 11348
rect 40358 11308 40408 11336
rect 40358 11304 40370 11308
rect 40312 11298 40370 11304
rect 40402 11296 40408 11308
rect 40460 11296 40466 11348
rect 41046 11336 41052 11348
rect 41006 11308 41052 11336
rect 41046 11296 41052 11308
rect 41104 11296 41110 11348
rect 41598 11336 41604 11348
rect 41558 11308 41604 11336
rect 41598 11296 41604 11308
rect 41656 11296 41662 11348
rect 55030 11296 55036 11348
rect 55088 11336 55094 11348
rect 55308 11338 55366 11344
rect 55308 11336 55320 11338
rect 55088 11308 55320 11336
rect 55088 11296 55094 11308
rect 55308 11304 55320 11308
rect 55354 11304 55366 11338
rect 55308 11298 55366 11304
rect 56228 11338 56286 11344
rect 56228 11304 56240 11338
rect 56274 11336 56286 11338
rect 57698 11336 57704 11348
rect 56274 11308 57704 11336
rect 56274 11304 56286 11308
rect 56228 11298 56286 11304
rect 57698 11296 57704 11308
rect 57756 11296 57762 11348
rect 76374 11296 76380 11348
rect 76432 11336 76438 11348
rect 76468 11338 76526 11344
rect 76468 11336 76480 11338
rect 76432 11308 76480 11336
rect 76432 11296 76438 11308
rect 76468 11304 76480 11308
rect 76514 11304 76526 11338
rect 76468 11298 76526 11304
rect 78216 11338 78274 11344
rect 78216 11304 78228 11338
rect 78262 11336 78274 11338
rect 78766 11336 78772 11348
rect 78262 11308 78772 11336
rect 78262 11304 78274 11308
rect 78216 11298 78274 11304
rect 78766 11296 78772 11308
rect 78824 11296 78830 11348
rect 84470 11296 84476 11348
rect 84528 11336 84534 11348
rect 86220 11338 86278 11344
rect 86220 11336 86232 11338
rect 84528 11308 86232 11336
rect 84528 11296 84534 11308
rect 86220 11304 86232 11308
rect 86266 11304 86278 11338
rect 86220 11298 86278 11304
rect 86956 11338 87014 11344
rect 86956 11304 86968 11338
rect 87002 11336 87014 11338
rect 87138 11336 87144 11348
rect 87002 11308 87144 11336
rect 87002 11304 87014 11308
rect 86956 11298 87014 11304
rect 87138 11296 87144 11308
rect 87196 11296 87202 11348
rect 88244 11338 88302 11344
rect 88244 11304 88256 11338
rect 88290 11336 88302 11338
rect 89070 11336 89076 11348
rect 88290 11308 89076 11336
rect 88290 11304 88302 11308
rect 88244 11298 88302 11304
rect 89070 11296 89076 11308
rect 89128 11296 89134 11348
rect 102870 11336 102876 11348
rect 102830 11308 102876 11336
rect 102870 11296 102876 11308
rect 102928 11296 102934 11348
rect 115106 11296 115112 11348
rect 115164 11336 115170 11348
rect 116028 11338 116086 11344
rect 116028 11336 116040 11338
rect 115164 11308 116040 11336
rect 115164 11296 115170 11308
rect 116028 11304 116040 11308
rect 116074 11304 116086 11338
rect 116028 11298 116086 11304
rect 117132 11338 117190 11344
rect 117132 11304 117144 11338
rect 117178 11336 117190 11338
rect 117682 11336 117688 11348
rect 117178 11308 117688 11336
rect 117178 11304 117190 11308
rect 117132 11298 117190 11304
rect 117682 11296 117688 11308
rect 117740 11296 117746 11348
rect 130378 11296 130384 11348
rect 130436 11336 130442 11348
rect 130472 11338 130530 11344
rect 130472 11336 130484 11338
rect 130436 11308 130484 11336
rect 130436 11296 130442 11308
rect 130472 11304 130484 11308
rect 130518 11304 130530 11338
rect 131206 11336 131212 11348
rect 131166 11308 131212 11336
rect 130472 11298 130530 11304
rect 131206 11296 131212 11308
rect 131264 11296 131270 11348
rect 131760 11338 131818 11344
rect 131760 11304 131772 11338
rect 131806 11336 131818 11338
rect 132862 11336 132868 11348
rect 131806 11308 132868 11336
rect 131806 11304 131818 11308
rect 131760 11298 131818 11304
rect 132862 11296 132868 11308
rect 132920 11296 132926 11348
rect 148042 11336 148048 11348
rect 148002 11308 148048 11336
rect 148042 11296 148048 11308
rect 148100 11296 148106 11348
rect 150802 11336 150808 11348
rect 150762 11308 150808 11336
rect 150802 11296 150808 11308
rect 150860 11296 150866 11348
rect 157242 11296 157248 11348
rect 157300 11336 157306 11348
rect 157336 11338 157394 11344
rect 157336 11336 157348 11338
rect 157300 11308 157348 11336
rect 157300 11296 157306 11308
rect 157336 11304 157348 11308
rect 157382 11304 157394 11338
rect 157336 11298 157394 11304
rect 162028 11338 162086 11344
rect 162028 11304 162040 11338
rect 162074 11336 162086 11338
rect 162118 11336 162124 11348
rect 162074 11308 162124 11336
rect 162074 11304 162086 11308
rect 162028 11298 162086 11304
rect 162118 11296 162124 11308
rect 162176 11296 162182 11348
rect 162670 11336 162676 11348
rect 162630 11308 162676 11336
rect 162670 11296 162676 11308
rect 162728 11296 162734 11348
rect 163406 11296 163412 11348
rect 163464 11336 163470 11348
rect 163592 11338 163650 11344
rect 163592 11336 163604 11338
rect 163464 11308 163604 11336
rect 163464 11296 163470 11308
rect 163592 11304 163604 11308
rect 163638 11304 163650 11338
rect 163592 11298 163650 11304
rect 165890 11296 165896 11348
rect 165948 11336 165954 11348
rect 239398 11336 239404 11348
rect 165948 11308 239404 11336
rect 165948 11296 165954 11308
rect 239398 11296 239404 11308
rect 239456 11296 239462 11348
rect 239766 11296 239772 11348
rect 239824 11336 239830 11348
rect 239952 11338 240010 11344
rect 239952 11336 239964 11338
rect 239824 11308 239964 11336
rect 239824 11296 239830 11308
rect 239952 11304 239964 11308
rect 239998 11304 240010 11338
rect 239952 11298 240010 11304
rect 240042 11296 240048 11348
rect 240100 11336 240106 11348
rect 240872 11338 240930 11344
rect 240872 11336 240884 11338
rect 240100 11308 240884 11336
rect 240100 11296 240106 11308
rect 240872 11304 240884 11308
rect 240918 11304 240930 11338
rect 240872 11298 240930 11304
rect 240962 11296 240968 11348
rect 241020 11336 241026 11348
rect 241424 11338 241482 11344
rect 241424 11336 241436 11338
rect 241020 11308 241436 11336
rect 241020 11296 241026 11308
rect 241424 11304 241436 11308
rect 241470 11304 241482 11338
rect 241424 11298 241482 11304
rect 242066 11296 242072 11348
rect 242124 11336 242130 11348
rect 242160 11338 242218 11344
rect 242160 11336 242172 11338
rect 242124 11308 242172 11336
rect 242124 11296 242130 11308
rect 242160 11304 242172 11308
rect 242206 11304 242218 11338
rect 242160 11298 242218 11304
rect 252462 11296 252468 11348
rect 252520 11336 252526 11348
rect 252556 11338 252614 11344
rect 252556 11336 252568 11338
rect 252520 11308 252568 11336
rect 252520 11296 252526 11308
rect 252556 11304 252568 11308
rect 252602 11304 252614 11338
rect 253106 11336 253112 11348
rect 253066 11308 253112 11336
rect 252556 11298 252614 11304
rect 253106 11296 253112 11308
rect 253164 11296 253170 11348
rect 253752 11338 253810 11344
rect 253752 11304 253764 11338
rect 253798 11336 253810 11338
rect 254026 11336 254032 11348
rect 253798 11308 254032 11336
rect 253798 11304 253810 11308
rect 253752 11298 253810 11304
rect 254026 11296 254032 11308
rect 254084 11296 254090 11348
rect 265434 11296 265440 11348
rect 265492 11336 265498 11348
rect 265528 11338 265586 11344
rect 265528 11336 265540 11338
rect 265492 11308 265540 11336
rect 265492 11296 265498 11308
rect 265528 11304 265540 11308
rect 265574 11304 265586 11338
rect 265528 11298 265586 11304
rect 266262 11296 266268 11348
rect 266320 11336 266326 11348
rect 268012 11338 268070 11344
rect 266320 11308 267964 11336
rect 266320 11296 266326 11308
rect 36446 11268 36452 11280
rect 28960 11240 29776 11268
rect 31726 11240 36452 11268
rect 28960 11228 28966 11240
rect 27062 11160 27068 11212
rect 27120 11200 27126 11212
rect 29454 11200 29460 11212
rect 27120 11172 29460 11200
rect 27120 11160 27126 11172
rect 29454 11160 29460 11172
rect 29512 11160 29518 11212
rect 29546 11160 29552 11212
rect 29604 11200 29610 11212
rect 29640 11202 29698 11208
rect 29640 11200 29652 11202
rect 29604 11172 29652 11200
rect 29604 11160 29610 11172
rect 29640 11168 29652 11172
rect 29686 11168 29698 11202
rect 29748 11200 29776 11240
rect 36446 11228 36452 11240
rect 36504 11228 36510 11280
rect 41322 11228 41328 11280
rect 41380 11268 41386 11280
rect 42244 11270 42302 11276
rect 42244 11268 42256 11270
rect 41380 11240 42256 11268
rect 41380 11228 41386 11240
rect 42244 11236 42256 11240
rect 42290 11236 42302 11270
rect 42244 11230 42302 11236
rect 86770 11228 86776 11280
rect 86828 11268 86834 11280
rect 87600 11270 87658 11276
rect 87600 11268 87612 11270
rect 86828 11240 87612 11268
rect 86828 11228 86834 11240
rect 87600 11236 87612 11240
rect 87646 11236 87658 11270
rect 87600 11230 87658 11236
rect 102226 11228 102232 11280
rect 102284 11268 102290 11280
rect 103516 11270 103574 11276
rect 103516 11268 103528 11270
rect 102284 11240 103528 11268
rect 102284 11228 102290 11240
rect 103516 11236 103528 11240
rect 103562 11236 103574 11270
rect 103516 11230 103574 11236
rect 114186 11228 114192 11280
rect 114244 11268 114250 11280
rect 115384 11270 115442 11276
rect 115384 11268 115396 11270
rect 114244 11240 115396 11268
rect 114244 11228 114250 11240
rect 115384 11236 115396 11240
rect 115430 11236 115442 11270
rect 115384 11230 115442 11236
rect 147398 11228 147404 11280
rect 147456 11268 147462 11280
rect 149884 11270 149942 11276
rect 147456 11240 148732 11268
rect 147456 11228 147462 11240
rect 31386 11200 31392 11212
rect 29748 11172 31392 11200
rect 29640 11162 29698 11168
rect 31386 11160 31392 11172
rect 31444 11160 31450 11212
rect 32306 11200 32312 11212
rect 32266 11172 32312 11200
rect 32306 11160 32312 11172
rect 32364 11160 32370 11212
rect 32492 11202 32550 11208
rect 32492 11168 32504 11202
rect 32538 11200 32550 11202
rect 32582 11200 32588 11212
rect 32538 11172 32588 11200
rect 32538 11168 32550 11172
rect 32492 11162 32550 11168
rect 27614 11092 27620 11144
rect 27672 11132 27678 11144
rect 28996 11134 29054 11140
rect 28996 11132 29008 11134
rect 27672 11104 29008 11132
rect 27672 11092 27678 11104
rect 28996 11100 29008 11104
rect 29042 11100 29054 11134
rect 32214 11132 32220 11144
rect 32174 11104 32220 11132
rect 28996 11094 29054 11100
rect 32214 11092 32220 11104
rect 32272 11092 32278 11144
rect 27982 11024 27988 11076
rect 28040 11064 28046 11076
rect 29914 11064 29920 11076
rect 28040 11036 29776 11064
rect 29874 11036 29920 11064
rect 28040 11024 28046 11036
rect 29748 10996 29776 11036
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 31662 11064 31668 11076
rect 31142 11036 31668 11064
rect 31662 11024 31668 11036
rect 31720 11024 31726 11076
rect 31754 11024 31760 11076
rect 31812 11064 31818 11076
rect 32508 11064 32536 11162
rect 32582 11160 32588 11172
rect 32640 11160 32646 11212
rect 45002 11200 45008 11212
rect 41800 11172 45008 11200
rect 33504 11134 33562 11140
rect 33504 11100 33516 11134
rect 33550 11132 33562 11134
rect 34698 11132 34704 11144
rect 33550 11104 34704 11132
rect 33550 11100 33562 11104
rect 33504 11094 33562 11100
rect 34698 11092 34704 11104
rect 34756 11092 34762 11144
rect 40494 11132 40500 11144
rect 40454 11104 40500 11132
rect 40494 11092 40500 11104
rect 40552 11092 40558 11144
rect 40956 11134 41014 11140
rect 40956 11100 40968 11134
rect 41002 11132 41014 11134
rect 41414 11132 41420 11144
rect 41002 11104 41420 11132
rect 41002 11100 41014 11104
rect 40956 11094 41014 11100
rect 41414 11092 41420 11104
rect 41472 11092 41478 11144
rect 41800 11140 41828 11172
rect 45002 11160 45008 11172
rect 45060 11160 45066 11212
rect 85482 11160 85488 11212
rect 85540 11200 85546 11212
rect 89162 11200 89168 11212
rect 85540 11172 89168 11200
rect 85540 11160 85546 11172
rect 41784 11134 41842 11140
rect 41784 11100 41796 11134
rect 41830 11100 41842 11134
rect 42426 11132 42432 11144
rect 42386 11104 42432 11132
rect 41784 11094 41842 11100
rect 42426 11092 42432 11104
rect 42484 11092 42490 11144
rect 55490 11132 55496 11144
rect 55450 11104 55496 11132
rect 55490 11092 55496 11104
rect 55548 11092 55554 11144
rect 56412 11134 56470 11140
rect 56412 11100 56424 11134
rect 56458 11132 56470 11134
rect 57238 11132 57244 11144
rect 56458 11104 57244 11132
rect 56458 11100 56470 11104
rect 56412 11094 56470 11100
rect 57238 11092 57244 11104
rect 57296 11092 57302 11144
rect 74718 11092 74724 11144
rect 74776 11132 74782 11144
rect 76652 11134 76710 11140
rect 76652 11132 76664 11134
rect 74776 11104 76664 11132
rect 74776 11092 74782 11104
rect 76652 11100 76664 11104
rect 76698 11100 76710 11134
rect 78398 11132 78404 11144
rect 78358 11104 78404 11132
rect 76652 11094 76710 11100
rect 78398 11092 78404 11104
rect 78456 11092 78462 11144
rect 86402 11132 86408 11144
rect 86362 11104 86408 11132
rect 86402 11092 86408 11104
rect 86460 11092 86466 11144
rect 86880 11140 86908 11172
rect 89162 11160 89168 11172
rect 89220 11160 89226 11212
rect 102042 11160 102048 11212
rect 102100 11200 102106 11212
rect 102320 11202 102378 11208
rect 102320 11200 102332 11202
rect 102100 11172 102332 11200
rect 102100 11160 102106 11172
rect 102320 11168 102332 11172
rect 102366 11168 102378 11202
rect 102320 11162 102378 11168
rect 102594 11160 102600 11212
rect 102652 11200 102658 11212
rect 102652 11172 103514 11200
rect 102652 11160 102658 11172
rect 86864 11134 86922 11140
rect 86864 11100 86876 11134
rect 86910 11100 86922 11134
rect 87782 11132 87788 11144
rect 87742 11104 87788 11132
rect 86864 11094 86922 11100
rect 87782 11092 87788 11104
rect 87840 11092 87846 11144
rect 88426 11132 88432 11144
rect 88386 11104 88432 11132
rect 88426 11092 88432 11104
rect 88484 11092 88490 11144
rect 102136 11134 102194 11140
rect 102136 11100 102148 11134
rect 102182 11132 102194 11134
rect 102410 11132 102416 11144
rect 102182 11104 102416 11132
rect 102182 11100 102194 11104
rect 102136 11094 102194 11100
rect 102410 11092 102416 11104
rect 102468 11092 102474 11144
rect 103054 11132 103060 11144
rect 103014 11104 103060 11132
rect 103054 11092 103060 11104
rect 103112 11092 103118 11144
rect 103486 11132 103514 11172
rect 130286 11160 130292 11212
rect 130344 11200 130350 11212
rect 132586 11200 132592 11212
rect 130344 11172 132592 11200
rect 130344 11160 130350 11172
rect 103700 11134 103758 11140
rect 103700 11132 103712 11134
rect 103486 11104 103712 11132
rect 103700 11100 103712 11104
rect 103746 11100 103758 11134
rect 103700 11094 103758 11100
rect 114738 11092 114744 11144
rect 114796 11132 114802 11144
rect 115292 11134 115350 11140
rect 115292 11132 115304 11134
rect 114796 11104 115304 11132
rect 114796 11092 114802 11104
rect 115292 11100 115304 11104
rect 115338 11132 115350 11134
rect 115750 11132 115756 11144
rect 115338 11104 115756 11132
rect 115338 11100 115350 11104
rect 115292 11094 115350 11100
rect 115750 11092 115756 11104
rect 115808 11092 115814 11144
rect 115842 11092 115848 11144
rect 115900 11132 115906 11144
rect 116212 11134 116270 11140
rect 116212 11132 116224 11134
rect 115900 11104 116224 11132
rect 115900 11092 115906 11104
rect 116212 11100 116224 11104
rect 116258 11100 116270 11134
rect 116212 11094 116270 11100
rect 117316 11134 117374 11140
rect 117316 11100 117328 11134
rect 117362 11132 117374 11134
rect 119706 11132 119712 11144
rect 117362 11104 119712 11132
rect 117362 11100 117374 11104
rect 117316 11094 117374 11100
rect 119706 11092 119712 11104
rect 119764 11092 119770 11144
rect 130656 11134 130714 11140
rect 130656 11100 130668 11134
rect 130702 11132 130714 11134
rect 130930 11132 130936 11144
rect 130702 11104 130936 11132
rect 130702 11100 130714 11104
rect 130656 11094 130714 11100
rect 130930 11092 130936 11104
rect 130988 11092 130994 11144
rect 131132 11140 131160 11172
rect 132586 11160 132592 11172
rect 132644 11160 132650 11212
rect 143258 11160 143264 11212
rect 143316 11200 143322 11212
rect 143316 11172 145880 11200
rect 143316 11160 143322 11172
rect 131116 11134 131174 11140
rect 131116 11100 131128 11134
rect 131162 11100 131174 11134
rect 131116 11094 131174 11100
rect 131944 11134 132002 11140
rect 131944 11100 131956 11134
rect 131990 11132 132002 11134
rect 133138 11132 133144 11144
rect 131990 11104 133144 11132
rect 131990 11100 132002 11104
rect 131944 11094 132002 11100
rect 133138 11092 133144 11104
rect 133196 11092 133202 11144
rect 142062 11132 142068 11144
rect 141974 11104 142068 11132
rect 142062 11092 142068 11104
rect 142120 11132 142126 11144
rect 145742 11132 145748 11144
rect 142120 11104 145748 11132
rect 142120 11092 142126 11104
rect 145742 11092 145748 11104
rect 145800 11092 145806 11144
rect 145852 11132 145880 11172
rect 147490 11160 147496 11212
rect 147548 11200 147554 11212
rect 148704 11208 148732 11240
rect 149884 11236 149896 11270
rect 149930 11268 149942 11270
rect 156414 11268 156420 11280
rect 149930 11240 156420 11268
rect 149930 11236 149942 11240
rect 149884 11230 149942 11236
rect 156414 11228 156420 11240
rect 156472 11228 156478 11280
rect 165430 11228 165436 11280
rect 165488 11268 165494 11280
rect 252738 11268 252744 11280
rect 165488 11240 192156 11268
rect 165488 11228 165494 11240
rect 148504 11202 148562 11208
rect 148504 11200 148516 11202
rect 147548 11172 148516 11200
rect 147548 11160 147554 11172
rect 148504 11168 148516 11172
rect 148550 11168 148562 11202
rect 148504 11162 148562 11168
rect 148688 11202 148746 11208
rect 148688 11168 148700 11202
rect 148734 11200 148746 11202
rect 151354 11200 151360 11212
rect 148734 11172 151360 11200
rect 148734 11168 148746 11172
rect 148688 11162 148746 11168
rect 151354 11160 151360 11172
rect 151412 11160 151418 11212
rect 165338 11200 165344 11212
rect 162872 11172 165344 11200
rect 150988 11134 151046 11140
rect 145852 11104 149560 11132
rect 31812 11036 32536 11064
rect 31812 11024 31818 11036
rect 81618 11024 81624 11076
rect 81676 11064 81682 11076
rect 87874 11064 87880 11076
rect 81676 11036 87880 11064
rect 81676 11024 81682 11036
rect 87874 11024 87880 11036
rect 87932 11024 87938 11076
rect 102428 11064 102456 11092
rect 113726 11064 113732 11076
rect 102428 11036 113732 11064
rect 113726 11024 113732 11036
rect 113784 11024 113790 11076
rect 140408 11066 140466 11072
rect 140408 11032 140420 11066
rect 140454 11064 140466 11066
rect 140682 11064 140688 11076
rect 140454 11036 140688 11064
rect 140454 11032 140466 11036
rect 140408 11026 140466 11032
rect 140682 11024 140688 11036
rect 140740 11064 140746 11076
rect 149532 11064 149560 11104
rect 150988 11100 151000 11134
rect 151034 11132 151046 11134
rect 153102 11132 153108 11144
rect 151034 11104 153108 11132
rect 151034 11100 151046 11104
rect 150988 11094 151046 11100
rect 153102 11092 153108 11104
rect 153160 11092 153166 11144
rect 162210 11132 162216 11144
rect 162170 11104 162216 11132
rect 162210 11092 162216 11104
rect 162268 11092 162274 11144
rect 162872 11140 162900 11172
rect 165338 11160 165344 11172
rect 165396 11160 165402 11212
rect 177576 11202 177634 11208
rect 177576 11168 177588 11202
rect 177622 11200 177634 11202
rect 177666 11200 177672 11212
rect 177622 11172 177672 11200
rect 177622 11168 177634 11172
rect 177576 11162 177634 11168
rect 177666 11160 177672 11172
rect 177724 11160 177730 11212
rect 177942 11160 177948 11212
rect 178000 11200 178006 11212
rect 178220 11202 178278 11208
rect 178220 11200 178232 11202
rect 178000 11172 178232 11200
rect 178000 11160 178006 11172
rect 178220 11168 178232 11172
rect 178266 11168 178278 11202
rect 180794 11200 180800 11212
rect 178220 11162 178278 11168
rect 178604 11172 180800 11200
rect 162856 11134 162914 11140
rect 162856 11100 162868 11134
rect 162902 11100 162914 11134
rect 163498 11132 163504 11144
rect 163458 11104 163504 11132
rect 162856 11094 162914 11100
rect 163498 11092 163504 11104
rect 163556 11092 163562 11144
rect 177484 11134 177542 11140
rect 177484 11100 177496 11134
rect 177530 11132 177542 11134
rect 178034 11132 178040 11144
rect 177530 11104 178040 11132
rect 177530 11100 177542 11104
rect 177484 11094 177542 11100
rect 178034 11092 178040 11104
rect 178092 11132 178098 11144
rect 178128 11134 178186 11140
rect 178128 11132 178140 11134
rect 178092 11104 178140 11132
rect 178092 11092 178098 11104
rect 178128 11100 178140 11104
rect 178174 11132 178186 11134
rect 178604 11132 178632 11172
rect 180794 11160 180800 11172
rect 180852 11160 180858 11212
rect 190272 11202 190330 11208
rect 190272 11168 190284 11202
rect 190318 11200 190330 11202
rect 191190 11200 191196 11212
rect 190318 11172 191196 11200
rect 190318 11168 190330 11172
rect 190272 11162 190330 11168
rect 191190 11160 191196 11172
rect 191248 11160 191254 11212
rect 191834 11160 191840 11212
rect 191892 11200 191898 11212
rect 192020 11202 192078 11208
rect 192020 11200 192032 11202
rect 191892 11172 192032 11200
rect 191892 11160 191898 11172
rect 192020 11168 192032 11172
rect 192066 11168 192078 11202
rect 192128 11200 192156 11240
rect 193324 11240 252744 11268
rect 193324 11200 193352 11240
rect 252738 11228 252744 11240
rect 252796 11228 252802 11280
rect 253198 11228 253204 11280
rect 253256 11268 253262 11280
rect 254396 11270 254454 11276
rect 254396 11268 254408 11270
rect 253256 11240 254408 11268
rect 253256 11228 253262 11240
rect 254396 11236 254408 11240
rect 254442 11236 254454 11270
rect 254396 11230 254454 11236
rect 265158 11228 265164 11280
rect 265216 11268 265222 11280
rect 266816 11270 266874 11276
rect 266816 11268 266828 11270
rect 265216 11240 266828 11268
rect 265216 11228 265222 11240
rect 266816 11236 266828 11240
rect 266862 11236 266874 11270
rect 267936 11268 267964 11308
rect 268012 11304 268024 11338
rect 268058 11336 268070 11338
rect 269298 11336 269304 11348
rect 268058 11308 269304 11336
rect 268058 11304 268070 11308
rect 268012 11298 268070 11304
rect 269298 11296 269304 11308
rect 269356 11296 269362 11348
rect 267936 11240 269436 11268
rect 266816 11230 266874 11236
rect 192128 11172 193352 11200
rect 192020 11162 192078 11168
rect 193490 11160 193496 11212
rect 193548 11200 193554 11212
rect 193768 11202 193826 11208
rect 193768 11200 193780 11202
rect 193548 11172 193780 11200
rect 193548 11160 193554 11172
rect 193768 11168 193780 11172
rect 193814 11200 193826 11202
rect 194410 11200 194416 11212
rect 193814 11172 194416 11200
rect 193814 11168 193826 11172
rect 193768 11162 193826 11168
rect 194410 11160 194416 11172
rect 194468 11160 194474 11212
rect 194594 11160 194600 11212
rect 194652 11200 194658 11212
rect 194964 11202 195022 11208
rect 194964 11200 194976 11202
rect 194652 11172 194976 11200
rect 194652 11160 194658 11172
rect 194964 11168 194976 11172
rect 195010 11168 195022 11202
rect 196434 11200 196440 11212
rect 194964 11162 195022 11168
rect 195440 11172 196440 11200
rect 178174 11104 178632 11132
rect 179140 11134 179198 11140
rect 178174 11100 178186 11104
rect 178128 11094 178186 11100
rect 179140 11100 179152 11134
rect 179186 11132 179198 11134
rect 180426 11132 180432 11144
rect 179186 11104 180432 11132
rect 179186 11100 179198 11104
rect 179140 11094 179198 11100
rect 180426 11092 180432 11104
rect 180484 11092 180490 11144
rect 188982 11092 188988 11144
rect 189040 11132 189046 11144
rect 190180 11134 190238 11140
rect 190180 11132 190192 11134
rect 189040 11104 190192 11132
rect 189040 11092 189046 11104
rect 190180 11100 190192 11104
rect 190226 11132 190238 11134
rect 190638 11132 190644 11144
rect 190226 11104 190644 11132
rect 190226 11100 190238 11104
rect 190180 11094 190238 11100
rect 190638 11092 190644 11104
rect 190696 11092 190702 11144
rect 190822 11132 190828 11144
rect 190782 11104 190828 11132
rect 190822 11092 190828 11104
rect 190880 11092 190886 11144
rect 190916 11134 190974 11140
rect 190916 11100 190928 11134
rect 190962 11132 190974 11134
rect 191926 11132 191932 11144
rect 190962 11104 191932 11132
rect 190962 11100 190974 11104
rect 190916 11094 190974 11100
rect 191926 11092 191932 11104
rect 191984 11092 191990 11144
rect 194780 11134 194838 11140
rect 194780 11100 194792 11134
rect 194826 11132 194838 11134
rect 194870 11132 194876 11144
rect 194826 11104 194876 11132
rect 194826 11100 194838 11104
rect 194780 11094 194838 11100
rect 194870 11092 194876 11104
rect 194928 11092 194934 11144
rect 195440 11132 195468 11172
rect 196434 11160 196440 11172
rect 196492 11160 196498 11212
rect 201034 11160 201040 11212
rect 201092 11200 201098 11212
rect 202876 11202 202934 11208
rect 201092 11172 202828 11200
rect 201092 11160 201098 11172
rect 195790 11132 195796 11144
rect 195164 11104 195468 11132
rect 195750 11104 195796 11132
rect 149608 11066 149666 11072
rect 149608 11064 149620 11066
rect 140740 11036 149468 11064
rect 149532 11036 149620 11064
rect 140740 11024 140746 11036
rect 31388 10998 31446 11004
rect 31388 10996 31400 10998
rect 29748 10968 31400 10996
rect 31388 10964 31400 10968
rect 31434 10964 31446 10998
rect 31846 10996 31852 11008
rect 31806 10968 31852 10996
rect 31388 10958 31446 10964
rect 31846 10956 31852 10968
rect 31904 10956 31910 11008
rect 148412 10998 148470 11004
rect 148412 10964 148424 10998
rect 148458 10996 148470 10998
rect 149054 10996 149060 11008
rect 148458 10968 149060 10996
rect 148458 10964 148470 10968
rect 148412 10958 148470 10964
rect 149054 10956 149060 10968
rect 149112 10956 149118 11008
rect 149440 10996 149468 11036
rect 149608 11032 149620 11036
rect 149654 11032 149666 11066
rect 156048 11066 156106 11072
rect 156048 11064 156060 11066
rect 149608 11026 149666 11032
rect 149716 11036 156060 11064
rect 149514 10996 149520 11008
rect 149440 10968 149520 10996
rect 149514 10956 149520 10968
rect 149572 10996 149578 11008
rect 149716 10996 149744 11036
rect 156048 11032 156060 11036
rect 156094 11064 156106 11066
rect 156138 11064 156144 11076
rect 156094 11036 156144 11064
rect 156094 11032 156106 11036
rect 156048 11026 156106 11032
rect 156138 11024 156144 11036
rect 156196 11024 156202 11076
rect 179414 11064 179420 11076
rect 178972 11036 179420 11064
rect 178972 11004 179000 11036
rect 179414 11024 179420 11036
rect 179472 11024 179478 11076
rect 189442 11024 189448 11076
rect 189500 11064 189506 11076
rect 192296 11066 192354 11072
rect 192296 11064 192308 11066
rect 189500 11036 192308 11064
rect 189500 11024 189506 11036
rect 192296 11032 192308 11036
rect 192342 11032 192354 11066
rect 192296 11026 192354 11032
rect 193306 11024 193312 11076
rect 193364 11024 193370 11076
rect 195164 11064 195192 11104
rect 195790 11092 195796 11104
rect 195848 11092 195854 11144
rect 202324 11134 202382 11140
rect 202324 11100 202336 11134
rect 202370 11132 202382 11134
rect 202690 11132 202696 11144
rect 202370 11104 202696 11132
rect 202370 11100 202382 11104
rect 202324 11094 202382 11100
rect 202690 11092 202696 11104
rect 202748 11092 202754 11144
rect 202800 11140 202828 11172
rect 202876 11168 202888 11202
rect 202922 11200 202934 11202
rect 203334 11200 203340 11212
rect 202922 11172 203340 11200
rect 202922 11168 202934 11172
rect 202876 11162 202934 11168
rect 203334 11160 203340 11172
rect 203392 11160 203398 11212
rect 204990 11200 204996 11212
rect 203536 11172 204996 11200
rect 202784 11134 202842 11140
rect 202784 11100 202796 11134
rect 202830 11132 202842 11134
rect 203428 11134 203486 11140
rect 203428 11132 203440 11134
rect 202830 11104 203440 11132
rect 202830 11100 202842 11104
rect 202784 11094 202842 11100
rect 203428 11100 203440 11104
rect 203474 11100 203486 11134
rect 203428 11094 203486 11100
rect 194888 11036 195192 11064
rect 149572 10968 149744 10996
rect 178956 10998 179014 11004
rect 149572 10956 149578 10968
rect 178956 10964 178968 10998
rect 179002 10964 179014 10998
rect 194410 10996 194416 11008
rect 194370 10968 194416 10996
rect 178956 10958 179014 10964
rect 194410 10956 194416 10968
rect 194468 10956 194474 11008
rect 194888 11004 194916 11036
rect 195238 11024 195244 11076
rect 195296 11064 195302 11076
rect 203536 11064 203564 11172
rect 204990 11160 204996 11172
rect 205048 11160 205054 11212
rect 238018 11160 238024 11212
rect 238076 11200 238082 11212
rect 242710 11200 242716 11212
rect 238076 11172 242716 11200
rect 238076 11160 238082 11172
rect 242710 11160 242716 11172
rect 242768 11160 242774 11212
rect 264976 11202 265034 11208
rect 264976 11168 264988 11202
rect 265022 11200 265034 11202
rect 267274 11200 267280 11212
rect 265022 11172 267280 11200
rect 265022 11168 265034 11172
rect 264976 11162 265034 11168
rect 267274 11160 267280 11172
rect 267332 11160 267338 11212
rect 267460 11202 267518 11208
rect 267460 11168 267472 11202
rect 267506 11200 267518 11202
rect 268010 11200 268016 11212
rect 267506 11172 268016 11200
rect 267506 11168 267518 11172
rect 267460 11162 267518 11168
rect 268010 11160 268016 11172
rect 268068 11160 268074 11212
rect 268470 11200 268476 11212
rect 268120 11172 268476 11200
rect 195296 11036 195652 11064
rect 195296 11024 195302 11036
rect 195624 11004 195652 11036
rect 202156 11036 203564 11064
rect 203628 11104 204852 11132
rect 202156 11004 202184 11036
rect 194872 10998 194930 11004
rect 194872 10964 194884 10998
rect 194918 10964 194930 10998
rect 194872 10958 194930 10964
rect 195608 10998 195666 11004
rect 195608 10964 195620 10998
rect 195654 10964 195666 10998
rect 195608 10958 195666 10964
rect 202140 10998 202198 11004
rect 202140 10964 202152 10998
rect 202186 10964 202198 10998
rect 202140 10958 202198 10964
rect 203520 10998 203578 11004
rect 203520 10964 203532 10998
rect 203566 10996 203578 10998
rect 203628 10996 203656 11104
rect 204070 11024 204076 11076
rect 204128 11064 204134 11076
rect 204824 11064 204852 11104
rect 204898 11092 204904 11144
rect 204956 11132 204962 11144
rect 229370 11132 229376 11144
rect 204956 11104 205000 11132
rect 229330 11104 229376 11132
rect 204956 11092 204962 11104
rect 229370 11092 229376 11104
rect 229428 11092 229434 11144
rect 239860 11134 239918 11140
rect 239860 11100 239872 11134
rect 239906 11132 239918 11134
rect 240780 11134 240838 11140
rect 240780 11132 240792 11134
rect 239906 11104 240792 11132
rect 239906 11100 239918 11104
rect 239860 11094 239918 11100
rect 240780 11100 240792 11104
rect 240826 11100 240838 11134
rect 240780 11094 240838 11100
rect 205450 11064 205456 11076
rect 204128 11036 204760 11064
rect 204824 11036 205456 11064
rect 204128 11024 204134 11036
rect 204732 11004 204760 11036
rect 205450 11024 205456 11036
rect 205508 11024 205514 11076
rect 230750 11064 230756 11076
rect 229204 11036 230756 11064
rect 229204 11004 229232 11036
rect 230750 11024 230756 11036
rect 230808 11024 230814 11076
rect 240796 11064 240824 11094
rect 240870 11092 240876 11144
rect 240928 11132 240934 11144
rect 241608 11134 241666 11140
rect 241608 11132 241620 11134
rect 240928 11104 241620 11132
rect 240928 11092 240934 11104
rect 241608 11100 241620 11104
rect 241654 11100 241666 11134
rect 241608 11094 241666 11100
rect 241974 11092 241980 11144
rect 242032 11132 242038 11144
rect 242068 11134 242126 11140
rect 242068 11132 242080 11134
rect 242032 11104 242080 11132
rect 242032 11092 242038 11104
rect 242068 11100 242080 11104
rect 242114 11100 242126 11134
rect 242068 11094 242126 11100
rect 251542 11092 251548 11144
rect 251600 11132 251606 11144
rect 252464 11134 252522 11140
rect 252464 11132 252476 11134
rect 251600 11104 252476 11132
rect 251600 11092 251606 11104
rect 252464 11100 252476 11104
rect 252510 11132 252522 11134
rect 253014 11132 253020 11144
rect 252510 11104 253020 11132
rect 252510 11100 252522 11104
rect 252464 11094 252522 11100
rect 253014 11092 253020 11104
rect 253072 11092 253078 11144
rect 253290 11132 253296 11144
rect 253250 11104 253296 11132
rect 253290 11092 253296 11104
rect 253348 11092 253354 11144
rect 253936 11134 253994 11140
rect 253936 11100 253948 11134
rect 253982 11132 253994 11134
rect 254394 11132 254400 11144
rect 253982 11104 254400 11132
rect 253982 11100 253994 11104
rect 253936 11094 253994 11100
rect 254394 11092 254400 11104
rect 254452 11092 254458 11144
rect 254580 11134 254638 11140
rect 254580 11100 254592 11134
rect 254626 11132 254638 11134
rect 254670 11132 254676 11144
rect 254626 11104 254676 11132
rect 254626 11100 254638 11104
rect 254580 11094 254638 11100
rect 254670 11092 254676 11104
rect 254728 11092 254734 11144
rect 264330 11092 264336 11144
rect 264388 11132 264394 11144
rect 264882 11132 264888 11144
rect 264388 11104 264888 11132
rect 264388 11092 264394 11104
rect 264882 11092 264888 11104
rect 264940 11092 264946 11144
rect 265618 11092 265624 11144
rect 265676 11132 265682 11144
rect 265712 11134 265770 11140
rect 265712 11132 265724 11134
rect 265676 11104 265724 11132
rect 265676 11092 265682 11104
rect 265712 11100 265724 11104
rect 265758 11100 265770 11134
rect 265712 11094 265770 11100
rect 267184 11134 267242 11140
rect 267184 11100 267196 11134
rect 267230 11132 267242 11134
rect 268120 11132 268148 11172
rect 268470 11160 268476 11172
rect 268528 11160 268534 11212
rect 268564 11202 268622 11208
rect 268564 11168 268576 11202
rect 268610 11200 268622 11202
rect 268930 11200 268936 11212
rect 268610 11172 268936 11200
rect 268610 11168 268622 11172
rect 268564 11162 268622 11168
rect 268930 11160 268936 11172
rect 268988 11160 268994 11212
rect 269408 11208 269436 11240
rect 269392 11202 269450 11208
rect 269392 11168 269404 11202
rect 269438 11200 269450 11202
rect 270588 11202 270646 11208
rect 270588 11200 270600 11202
rect 269438 11172 270600 11200
rect 269438 11168 269450 11172
rect 269392 11162 269450 11168
rect 270588 11168 270600 11172
rect 270634 11200 270646 11202
rect 272242 11200 272248 11212
rect 270634 11172 272248 11200
rect 270634 11168 270646 11172
rect 270588 11162 270646 11168
rect 272242 11160 272248 11172
rect 272300 11160 272306 11212
rect 267230 11104 268148 11132
rect 268196 11134 268254 11140
rect 267230 11100 267242 11104
rect 267184 11094 267242 11100
rect 268196 11100 268208 11134
rect 268242 11132 268254 11134
rect 269666 11132 269672 11144
rect 268242 11104 269672 11132
rect 268242 11100 268254 11104
rect 268196 11094 268254 11100
rect 269666 11092 269672 11104
rect 269724 11092 269730 11144
rect 270402 11132 270408 11144
rect 270362 11104 270408 11132
rect 270402 11092 270408 11104
rect 270460 11092 270466 11144
rect 270496 11134 270554 11140
rect 270496 11100 270508 11134
rect 270542 11132 270554 11134
rect 270862 11132 270868 11144
rect 270542 11104 270868 11132
rect 270542 11100 270554 11104
rect 270496 11094 270554 11100
rect 270862 11092 270868 11104
rect 270920 11092 270926 11144
rect 241992 11064 242020 11092
rect 240796 11036 242020 11064
rect 267276 11066 267334 11072
rect 267276 11032 267288 11066
rect 267322 11064 267334 11066
rect 268286 11064 268292 11076
rect 267322 11036 268292 11064
rect 267322 11032 267334 11036
rect 267276 11026 267334 11032
rect 268286 11024 268292 11036
rect 268344 11024 268350 11076
rect 268930 11024 268936 11076
rect 268988 11064 268994 11076
rect 269208 11066 269266 11072
rect 269208 11064 269220 11066
rect 268988 11036 269220 11064
rect 268988 11024 268994 11036
rect 269208 11032 269220 11036
rect 269254 11032 269266 11066
rect 269208 11026 269266 11032
rect 269300 11066 269358 11072
rect 269300 11032 269312 11066
rect 269346 11064 269358 11066
rect 269942 11064 269948 11076
rect 269346 11036 269948 11064
rect 269346 11032 269358 11036
rect 269300 11026 269358 11032
rect 269942 11024 269948 11036
rect 270000 11024 270006 11076
rect 203566 10968 203656 10996
rect 204716 10998 204774 11004
rect 203566 10964 203578 10968
rect 203520 10958 203578 10964
rect 204716 10964 204728 10998
rect 204762 10964 204774 10998
rect 204716 10958 204774 10964
rect 229188 10998 229246 11004
rect 229188 10964 229200 10998
rect 229234 10964 229246 10998
rect 268838 10996 268844 11008
rect 268798 10968 268844 10996
rect 229188 10958 229246 10964
rect 268838 10956 268844 10968
rect 268896 10956 268902 11008
rect 270034 10996 270040 11008
rect 269994 10968 270040 10996
rect 270034 10956 270040 10968
rect 270092 10956 270098 11008
rect 1104 10906 305808 10928
rect 1104 10854 77148 10906
rect 77200 10854 77212 10906
rect 77264 10854 77276 10906
rect 77328 10854 77340 10906
rect 77392 10854 77404 10906
rect 77456 10854 153346 10906
rect 153398 10854 153410 10906
rect 153462 10854 153474 10906
rect 153526 10854 153538 10906
rect 153590 10854 153602 10906
rect 153654 10854 229544 10906
rect 229596 10854 229608 10906
rect 229660 10854 229672 10906
rect 229724 10854 229736 10906
rect 229788 10854 229800 10906
rect 229852 10854 305808 10906
rect 1104 10832 305808 10854
rect 29640 10794 29698 10800
rect 29640 10760 29652 10794
rect 29686 10792 29698 10794
rect 29822 10792 29828 10804
rect 29686 10764 29828 10792
rect 29686 10760 29698 10764
rect 29640 10754 29698 10760
rect 29822 10752 29828 10764
rect 29880 10752 29886 10804
rect 30466 10752 30472 10804
rect 30524 10792 30530 10804
rect 30652 10794 30710 10800
rect 30652 10792 30664 10794
rect 30524 10764 30664 10792
rect 30524 10752 30530 10764
rect 30652 10760 30664 10764
rect 30698 10760 30710 10794
rect 30652 10754 30710 10760
rect 30742 10752 30748 10804
rect 30800 10792 30806 10804
rect 32124 10794 32182 10800
rect 32124 10792 32136 10794
rect 30800 10764 30844 10792
rect 30944 10764 32136 10792
rect 30800 10752 30806 10764
rect 29730 10684 29736 10736
rect 29788 10724 29794 10736
rect 29788 10696 30144 10724
rect 29788 10684 29794 10696
rect 28442 10616 28448 10668
rect 28500 10656 28506 10668
rect 29824 10658 29882 10664
rect 29824 10656 29836 10658
rect 28500 10628 29836 10656
rect 28500 10616 28506 10628
rect 29824 10624 29836 10628
rect 29870 10624 29882 10658
rect 30116 10656 30144 10696
rect 30190 10684 30196 10736
rect 30248 10724 30254 10736
rect 30944 10724 30972 10764
rect 32124 10760 32136 10764
rect 32170 10760 32182 10794
rect 32124 10754 32182 10760
rect 32674 10752 32680 10804
rect 32732 10792 32738 10804
rect 32768 10794 32826 10800
rect 32768 10792 32780 10794
rect 32732 10764 32780 10792
rect 32732 10752 32738 10764
rect 32768 10760 32780 10764
rect 32814 10760 32826 10794
rect 32768 10754 32826 10760
rect 33042 10752 33048 10804
rect 33100 10792 33106 10804
rect 33412 10794 33470 10800
rect 33412 10792 33424 10794
rect 33100 10764 33424 10792
rect 33100 10752 33106 10764
rect 33412 10760 33424 10764
rect 33458 10760 33470 10794
rect 101674 10792 101680 10804
rect 101634 10764 101680 10792
rect 33412 10754 33470 10760
rect 101674 10752 101680 10764
rect 101732 10752 101738 10804
rect 130470 10792 130476 10804
rect 130430 10764 130476 10792
rect 130470 10752 130476 10764
rect 130528 10752 130534 10804
rect 141970 10792 141976 10804
rect 141930 10764 141976 10792
rect 141970 10752 141976 10764
rect 142028 10752 142034 10804
rect 148594 10752 148600 10804
rect 148652 10792 148658 10804
rect 148872 10794 148930 10800
rect 148872 10792 148884 10794
rect 148652 10764 148884 10792
rect 148652 10752 148658 10764
rect 148872 10760 148884 10764
rect 148918 10760 148930 10794
rect 148872 10754 148930 10760
rect 148962 10752 148968 10804
rect 149020 10792 149026 10804
rect 150712 10794 150770 10800
rect 150712 10792 150724 10794
rect 149020 10764 150724 10792
rect 149020 10752 149026 10764
rect 150712 10760 150724 10764
rect 150758 10760 150770 10794
rect 150712 10754 150770 10760
rect 191098 10752 191104 10804
rect 191156 10792 191162 10804
rect 191836 10794 191894 10800
rect 191836 10792 191848 10794
rect 191156 10764 191848 10792
rect 191156 10752 191162 10764
rect 191836 10760 191848 10764
rect 191882 10760 191894 10794
rect 191836 10754 191894 10760
rect 192128 10764 193812 10792
rect 31754 10724 31760 10736
rect 30248 10696 30972 10724
rect 31036 10696 31760 10724
rect 30248 10684 30254 10696
rect 31036 10656 31064 10696
rect 31754 10684 31760 10696
rect 31812 10684 31818 10736
rect 31846 10684 31852 10736
rect 31904 10724 31910 10736
rect 140682 10724 140688 10736
rect 31904 10696 33640 10724
rect 140642 10696 140688 10724
rect 31904 10684 31910 10696
rect 32308 10658 32366 10664
rect 32308 10656 32320 10658
rect 30116 10628 31064 10656
rect 31726 10628 32320 10656
rect 29824 10618 29882 10624
rect 30852 10596 30880 10628
rect 30836 10590 30894 10596
rect 30836 10556 30848 10590
rect 30882 10556 30894 10590
rect 30836 10550 30894 10556
rect 30284 10522 30342 10528
rect 30284 10488 30296 10522
rect 30330 10520 30342 10522
rect 31726 10520 31754 10628
rect 32308 10624 32320 10628
rect 32354 10624 32366 10658
rect 32950 10656 32956 10668
rect 32910 10628 32956 10656
rect 32308 10618 32366 10624
rect 32950 10616 32956 10628
rect 33008 10616 33014 10668
rect 33612 10664 33640 10696
rect 140682 10684 140688 10696
rect 140740 10684 140746 10736
rect 151630 10724 151636 10736
rect 149072 10696 151636 10724
rect 33596 10658 33654 10664
rect 33596 10624 33608 10658
rect 33642 10624 33654 10658
rect 101858 10656 101864 10668
rect 101818 10628 101864 10656
rect 33596 10618 33654 10624
rect 101858 10616 101864 10628
rect 101916 10616 101922 10668
rect 130286 10616 130292 10668
rect 130344 10656 130350 10668
rect 149072 10664 149100 10696
rect 151630 10684 151636 10696
rect 151688 10684 151694 10736
rect 156138 10724 156144 10736
rect 156098 10696 156144 10724
rect 156138 10684 156144 10696
rect 156196 10684 156202 10736
rect 192128 10724 192156 10764
rect 187252 10696 192156 10724
rect 130380 10658 130438 10664
rect 130380 10656 130392 10658
rect 130344 10628 130392 10656
rect 130344 10616 130350 10628
rect 130380 10624 130392 10628
rect 130426 10624 130438 10658
rect 130380 10618 130438 10624
rect 149056 10658 149114 10664
rect 149056 10624 149068 10658
rect 149102 10624 149114 10658
rect 149056 10618 149114 10624
rect 150342 10616 150348 10668
rect 150400 10656 150406 10668
rect 187252 10664 187280 10696
rect 192202 10684 192208 10736
rect 192260 10724 192266 10736
rect 192260 10696 192708 10724
rect 192260 10684 192266 10696
rect 150620 10658 150678 10664
rect 150620 10656 150632 10658
rect 150400 10628 150632 10656
rect 150400 10616 150406 10628
rect 150620 10624 150632 10628
rect 150666 10624 150678 10658
rect 150620 10618 150678 10624
rect 187236 10658 187294 10664
rect 187236 10624 187248 10658
rect 187282 10624 187294 10658
rect 187236 10618 187294 10624
rect 190546 10616 190552 10668
rect 190604 10656 190610 10668
rect 191284 10658 191342 10664
rect 191284 10656 191296 10658
rect 190604 10628 191296 10656
rect 190604 10616 190610 10628
rect 191284 10624 191296 10628
rect 191330 10624 191342 10658
rect 191284 10618 191342 10624
rect 192020 10658 192078 10664
rect 192020 10624 192032 10658
rect 192066 10656 192078 10658
rect 192294 10656 192300 10668
rect 192066 10628 192300 10656
rect 192066 10624 192078 10628
rect 192020 10618 192078 10624
rect 192294 10616 192300 10628
rect 192352 10616 192358 10668
rect 192680 10664 192708 10696
rect 193214 10684 193220 10736
rect 193272 10724 193278 10736
rect 193492 10726 193550 10732
rect 193492 10724 193504 10726
rect 193272 10696 193504 10724
rect 193272 10684 193278 10696
rect 193492 10692 193504 10696
rect 193538 10692 193550 10726
rect 193784 10724 193812 10764
rect 193858 10752 193864 10804
rect 193916 10792 193922 10804
rect 194228 10794 194286 10800
rect 194228 10792 194240 10794
rect 193916 10764 194240 10792
rect 193916 10752 193922 10764
rect 194228 10760 194240 10764
rect 194274 10760 194286 10794
rect 194228 10754 194286 10760
rect 202876 10794 202934 10800
rect 202876 10760 202888 10794
rect 202922 10792 202934 10794
rect 205082 10792 205088 10804
rect 202922 10764 205088 10792
rect 202922 10760 202934 10764
rect 202876 10754 202934 10760
rect 205082 10752 205088 10764
rect 205140 10752 205146 10804
rect 253660 10794 253718 10800
rect 253660 10760 253672 10794
rect 253706 10792 253718 10794
rect 255222 10792 255228 10804
rect 253706 10764 255228 10792
rect 253706 10760 253718 10764
rect 253660 10754 253718 10760
rect 255222 10752 255228 10764
rect 255280 10752 255286 10804
rect 266538 10792 266544 10804
rect 266498 10764 266544 10792
rect 266538 10752 266544 10764
rect 266596 10752 266602 10804
rect 267736 10794 267794 10800
rect 267736 10760 267748 10794
rect 267782 10792 267794 10794
rect 268194 10792 268200 10804
rect 267782 10764 268200 10792
rect 267782 10760 267794 10764
rect 267736 10754 267794 10760
rect 268194 10752 268200 10764
rect 268252 10752 268258 10804
rect 268380 10794 268438 10800
rect 268380 10760 268392 10794
rect 268426 10792 268438 10794
rect 269390 10792 269396 10804
rect 268426 10764 269396 10792
rect 268426 10760 268438 10764
rect 268380 10754 268438 10760
rect 269390 10752 269396 10764
rect 269448 10752 269454 10804
rect 195054 10724 195060 10736
rect 193784 10696 195060 10724
rect 193492 10686 193550 10692
rect 195054 10684 195060 10696
rect 195112 10684 195118 10736
rect 264882 10684 264888 10736
rect 264940 10724 264946 10736
rect 270034 10724 270040 10736
rect 264940 10696 266492 10724
rect 264940 10684 264946 10696
rect 192664 10658 192722 10664
rect 192664 10624 192676 10658
rect 192710 10624 192722 10658
rect 194134 10656 194140 10668
rect 194094 10628 194140 10656
rect 192664 10618 192722 10624
rect 194134 10616 194140 10628
rect 194192 10656 194198 10668
rect 194962 10656 194968 10668
rect 194192 10628 194968 10656
rect 194192 10616 194198 10628
rect 194962 10616 194968 10628
rect 195020 10616 195026 10668
rect 203060 10658 203118 10664
rect 203060 10624 203072 10658
rect 203106 10656 203118 10658
rect 204806 10656 204812 10668
rect 203106 10628 204812 10656
rect 203106 10624 203118 10628
rect 203060 10618 203118 10624
rect 204806 10616 204812 10628
rect 204864 10616 204870 10668
rect 253844 10658 253902 10664
rect 253844 10624 253856 10658
rect 253890 10656 253902 10658
rect 254946 10656 254952 10668
rect 253890 10628 254952 10656
rect 253890 10624 253902 10628
rect 253844 10618 253902 10624
rect 254946 10616 254952 10628
rect 255004 10616 255010 10668
rect 265988 10658 266046 10664
rect 265988 10624 266000 10658
rect 266034 10656 266046 10658
rect 266354 10656 266360 10668
rect 266034 10628 266360 10656
rect 266034 10624 266046 10628
rect 265988 10618 266046 10624
rect 266354 10616 266360 10628
rect 266412 10616 266418 10668
rect 266464 10664 266492 10696
rect 267936 10696 270040 10724
rect 267936 10664 267964 10696
rect 270034 10684 270040 10696
rect 270092 10684 270098 10736
rect 266448 10658 266506 10664
rect 266448 10624 266460 10658
rect 266494 10656 266506 10658
rect 267092 10658 267150 10664
rect 267092 10656 267104 10658
rect 266494 10628 267104 10656
rect 266494 10624 266506 10628
rect 266448 10618 266506 10624
rect 267092 10624 267104 10628
rect 267138 10624 267150 10658
rect 267092 10618 267150 10624
rect 267920 10658 267978 10664
rect 267920 10624 267932 10658
rect 267966 10624 267978 10658
rect 267920 10618 267978 10624
rect 268564 10658 268622 10664
rect 268564 10624 268576 10658
rect 268610 10624 268622 10658
rect 268564 10618 268622 10624
rect 187510 10588 187516 10600
rect 187470 10560 187516 10588
rect 187510 10548 187516 10560
rect 187568 10548 187574 10600
rect 201034 10588 201040 10600
rect 192864 10560 201040 10588
rect 30330 10492 31754 10520
rect 191100 10522 191158 10528
rect 30330 10488 30342 10492
rect 30284 10482 30342 10488
rect 191100 10488 191112 10522
rect 191146 10520 191158 10522
rect 192110 10520 192116 10532
rect 191146 10492 192116 10520
rect 191146 10488 191158 10492
rect 191100 10482 191158 10488
rect 192110 10480 192116 10492
rect 192168 10480 192174 10532
rect 192864 10528 192892 10560
rect 201034 10548 201040 10560
rect 201092 10548 201098 10600
rect 268580 10588 268608 10618
rect 269022 10616 269028 10668
rect 269080 10656 269086 10668
rect 269116 10658 269174 10664
rect 269116 10656 269128 10658
rect 269080 10628 269128 10656
rect 269080 10616 269086 10628
rect 269116 10624 269128 10628
rect 269162 10624 269174 10658
rect 269116 10618 269174 10624
rect 269208 10658 269266 10664
rect 269208 10624 269220 10658
rect 269254 10656 269266 10658
rect 270310 10656 270316 10668
rect 269254 10628 270316 10656
rect 269254 10624 269266 10628
rect 269208 10618 269266 10624
rect 270310 10616 270316 10628
rect 270368 10616 270374 10668
rect 272518 10588 272524 10600
rect 268580 10560 272524 10588
rect 272518 10548 272524 10560
rect 272576 10548 272582 10600
rect 192848 10522 192906 10528
rect 192848 10488 192860 10522
rect 192894 10488 192906 10522
rect 192848 10482 192906 10488
rect 193676 10522 193734 10528
rect 193676 10488 193688 10522
rect 193722 10520 193734 10522
rect 267184 10522 267242 10528
rect 193722 10492 196848 10520
rect 193722 10488 193734 10492
rect 193676 10482 193734 10488
rect 157612 10454 157670 10460
rect 157612 10420 157624 10454
rect 157658 10452 157670 10454
rect 179138 10452 179144 10464
rect 157658 10424 179144 10452
rect 157658 10420 157670 10424
rect 157612 10414 157670 10420
rect 179138 10412 179144 10424
rect 179196 10412 179202 10464
rect 196820 10452 196848 10492
rect 267184 10488 267196 10522
rect 267230 10520 267242 10522
rect 268746 10520 268752 10532
rect 267230 10492 268752 10520
rect 267230 10488 267242 10492
rect 267184 10482 267242 10488
rect 268746 10480 268752 10492
rect 268804 10480 268810 10532
rect 203518 10452 203524 10464
rect 196820 10424 203524 10452
rect 203518 10412 203524 10424
rect 203576 10412 203582 10464
rect 265804 10454 265862 10460
rect 265804 10420 265816 10454
rect 265850 10452 265862 10454
rect 269574 10452 269580 10464
rect 265850 10424 269580 10452
rect 265850 10420 265862 10424
rect 265804 10414 265862 10420
rect 269574 10412 269580 10424
rect 269632 10412 269638 10464
rect 1104 10362 305808 10384
rect 1104 10310 39048 10362
rect 39100 10310 39112 10362
rect 39164 10310 39176 10362
rect 39228 10310 39240 10362
rect 39292 10310 39304 10362
rect 39356 10310 115246 10362
rect 115298 10310 115310 10362
rect 115362 10310 115374 10362
rect 115426 10310 115438 10362
rect 115490 10310 115502 10362
rect 115554 10310 191444 10362
rect 191496 10310 191508 10362
rect 191560 10310 191572 10362
rect 191624 10310 191636 10362
rect 191688 10310 191700 10362
rect 191752 10310 267642 10362
rect 267694 10310 267706 10362
rect 267758 10310 267770 10362
rect 267822 10310 267834 10362
rect 267886 10310 267898 10362
rect 267950 10310 305808 10362
rect 1104 10288 305808 10310
rect 30098 10208 30104 10260
rect 30156 10248 30162 10260
rect 30928 10250 30986 10256
rect 30928 10248 30940 10250
rect 30156 10220 30940 10248
rect 30156 10208 30162 10220
rect 30928 10216 30940 10220
rect 30974 10216 30986 10250
rect 31662 10248 31668 10260
rect 31622 10220 31668 10248
rect 30928 10210 30986 10216
rect 31662 10208 31668 10220
rect 31720 10208 31726 10260
rect 32122 10208 32128 10260
rect 32180 10248 32186 10260
rect 32860 10250 32918 10256
rect 32860 10248 32872 10250
rect 32180 10220 32872 10248
rect 32180 10208 32186 10220
rect 32860 10216 32872 10220
rect 32906 10216 32918 10250
rect 32860 10210 32918 10216
rect 33318 10208 33324 10260
rect 33376 10248 33382 10260
rect 33596 10250 33654 10256
rect 33596 10248 33608 10250
rect 33376 10220 33608 10248
rect 33376 10208 33382 10220
rect 33596 10216 33608 10220
rect 33642 10216 33654 10250
rect 33596 10210 33654 10216
rect 191282 10208 191288 10260
rect 191340 10248 191346 10260
rect 191836 10250 191894 10256
rect 191836 10248 191848 10250
rect 191340 10220 191848 10248
rect 191340 10208 191346 10220
rect 191836 10216 191848 10220
rect 191882 10216 191894 10250
rect 191836 10210 191894 10216
rect 192478 10208 192484 10260
rect 192536 10248 192542 10260
rect 193124 10250 193182 10256
rect 193124 10248 193136 10250
rect 192536 10220 193136 10248
rect 192536 10208 192542 10220
rect 193124 10216 193136 10220
rect 193170 10216 193182 10250
rect 193124 10210 193182 10216
rect 266906 10208 266912 10260
rect 266964 10248 266970 10260
rect 267736 10250 267794 10256
rect 267736 10248 267748 10250
rect 266964 10220 267748 10248
rect 266964 10208 266970 10220
rect 267736 10216 267748 10220
rect 267782 10216 267794 10250
rect 267736 10210 267794 10216
rect 268562 10208 268568 10260
rect 268620 10248 268626 10260
rect 269024 10250 269082 10256
rect 269024 10248 269036 10250
rect 268620 10220 269036 10248
rect 268620 10208 268626 10220
rect 269024 10216 269036 10220
rect 269070 10216 269082 10250
rect 269024 10210 269082 10216
rect 27522 10140 27528 10192
rect 27580 10180 27586 10192
rect 30284 10182 30342 10188
rect 30284 10180 30296 10182
rect 27580 10152 30296 10180
rect 27580 10140 27586 10152
rect 30284 10148 30296 10152
rect 30330 10148 30342 10182
rect 30284 10142 30342 10148
rect 31570 10140 31576 10192
rect 31628 10180 31634 10192
rect 32308 10182 32366 10188
rect 32308 10180 32320 10182
rect 31628 10152 32320 10180
rect 31628 10140 31634 10152
rect 32308 10148 32320 10152
rect 32354 10148 32366 10182
rect 32308 10142 32366 10148
rect 267092 10182 267150 10188
rect 267092 10148 267104 10182
rect 267138 10180 267150 10182
rect 268378 10180 268384 10192
rect 267138 10152 267734 10180
rect 267138 10148 267150 10152
rect 267092 10142 267150 10148
rect 267706 10124 267734 10152
rect 267844 10152 268384 10180
rect 157796 10114 157854 10120
rect 157796 10080 157808 10114
rect 157842 10112 157854 10114
rect 163590 10112 163596 10124
rect 157842 10084 163596 10112
rect 157842 10080 157854 10084
rect 157796 10074 157854 10080
rect 163590 10072 163596 10084
rect 163648 10072 163654 10124
rect 195882 10112 195888 10124
rect 192680 10084 195888 10112
rect 29454 10004 29460 10056
rect 29512 10044 29518 10056
rect 30468 10046 30526 10052
rect 30468 10044 30480 10046
rect 29512 10016 30480 10044
rect 29512 10004 29518 10016
rect 30468 10012 30480 10016
rect 30514 10012 30526 10046
rect 30468 10006 30526 10012
rect 30926 10004 30932 10056
rect 30984 10044 30990 10056
rect 31112 10046 31170 10052
rect 31112 10044 31124 10046
rect 30984 10016 31124 10044
rect 30984 10004 30990 10016
rect 31112 10012 31124 10016
rect 31158 10012 31170 10046
rect 31112 10006 31170 10012
rect 31572 10046 31630 10052
rect 31572 10012 31584 10046
rect 31618 10044 31630 10046
rect 32216 10046 32274 10052
rect 32216 10044 32228 10046
rect 31618 10016 32228 10044
rect 31618 10012 31630 10016
rect 31572 10006 31630 10012
rect 32216 10012 32228 10016
rect 32262 10012 32274 10046
rect 32216 10006 32274 10012
rect 33044 10046 33102 10052
rect 33044 10012 33056 10046
rect 33090 10044 33102 10046
rect 33410 10044 33416 10056
rect 33090 10016 33416 10044
rect 33090 10012 33102 10016
rect 33044 10006 33102 10012
rect 32232 9976 32260 10006
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 33504 10046 33562 10052
rect 33504 10012 33516 10046
rect 33550 10044 33562 10046
rect 33686 10044 33692 10056
rect 33550 10016 33692 10044
rect 33550 10012 33562 10016
rect 33504 10006 33562 10012
rect 33520 9976 33548 10006
rect 33686 10004 33692 10016
rect 33744 10004 33750 10056
rect 140408 10046 140466 10052
rect 140408 10012 140420 10046
rect 140454 10044 140466 10046
rect 140682 10044 140688 10056
rect 140454 10016 140688 10044
rect 140454 10012 140466 10016
rect 140408 10006 140466 10012
rect 140682 10004 140688 10016
rect 140740 10004 140746 10056
rect 156048 10046 156106 10052
rect 156048 10012 156060 10046
rect 156094 10044 156106 10046
rect 156138 10044 156144 10056
rect 156094 10016 156144 10044
rect 156094 10012 156106 10016
rect 156048 10006 156106 10012
rect 156138 10004 156144 10016
rect 156196 10004 156202 10056
rect 192020 10046 192078 10052
rect 192020 10012 192032 10046
rect 192066 10044 192078 10046
rect 192570 10044 192576 10056
rect 192066 10016 192576 10044
rect 192066 10012 192078 10016
rect 192020 10006 192078 10012
rect 192570 10004 192576 10016
rect 192628 10004 192634 10056
rect 192680 10052 192708 10084
rect 195882 10072 195888 10084
rect 195940 10072 195946 10124
rect 267706 10084 267740 10124
rect 267734 10072 267740 10084
rect 267792 10072 267798 10124
rect 192664 10046 192722 10052
rect 192664 10012 192676 10046
rect 192710 10012 192722 10046
rect 192664 10006 192722 10012
rect 193308 10046 193366 10052
rect 193308 10012 193320 10046
rect 193354 10044 193366 10046
rect 194410 10044 194416 10056
rect 193354 10016 194416 10044
rect 193354 10012 193366 10016
rect 193308 10006 193366 10012
rect 194410 10004 194416 10016
rect 194468 10004 194474 10056
rect 267276 10046 267334 10052
rect 267276 10012 267288 10046
rect 267322 10044 267334 10046
rect 267844 10044 267872 10152
rect 268378 10140 268384 10152
rect 268436 10140 268442 10192
rect 268472 10182 268530 10188
rect 268472 10148 268484 10182
rect 268518 10180 268530 10182
rect 269482 10180 269488 10192
rect 268518 10152 269488 10180
rect 268518 10148 268530 10152
rect 268472 10142 268530 10148
rect 269482 10140 269488 10152
rect 269540 10140 269546 10192
rect 268838 10112 268844 10124
rect 267936 10084 268844 10112
rect 267936 10052 267964 10084
rect 268838 10072 268844 10084
rect 268896 10072 268902 10124
rect 267322 10016 267872 10044
rect 267920 10046 267978 10052
rect 267322 10012 267334 10016
rect 267276 10006 267334 10012
rect 267920 10012 267932 10046
rect 267966 10012 267978 10046
rect 267920 10006 267978 10012
rect 268102 10004 268108 10056
rect 268160 10044 268166 10056
rect 268380 10046 268438 10052
rect 268380 10044 268392 10046
rect 268160 10016 268392 10044
rect 268160 10004 268166 10016
rect 268380 10012 268392 10016
rect 268426 10044 268438 10046
rect 269022 10044 269028 10056
rect 268426 10016 269028 10044
rect 268426 10012 268438 10016
rect 268380 10006 268438 10012
rect 269022 10004 269028 10016
rect 269080 10004 269086 10056
rect 269206 10044 269212 10056
rect 269166 10016 269212 10044
rect 269206 10004 269212 10016
rect 269264 10004 269270 10056
rect 304442 10044 304448 10056
rect 304402 10016 304448 10044
rect 304442 10004 304448 10016
rect 304500 10004 304506 10056
rect 32232 9948 33548 9976
rect 252738 9936 252744 9988
rect 252796 9976 252802 9988
rect 304812 9978 304870 9984
rect 304812 9976 304824 9978
rect 252796 9948 304824 9976
rect 252796 9936 252802 9948
rect 304812 9944 304824 9948
rect 304858 9944 304870 9978
rect 304812 9938 304870 9944
rect 117406 9868 117412 9920
rect 117464 9908 117470 9920
rect 141696 9910 141754 9916
rect 141696 9908 141708 9910
rect 117464 9880 141708 9908
rect 117464 9868 117470 9880
rect 141696 9876 141708 9880
rect 141742 9876 141754 9910
rect 141696 9870 141754 9876
rect 192480 9910 192538 9916
rect 192480 9876 192492 9910
rect 192526 9908 192538 9910
rect 194318 9908 194324 9920
rect 192526 9880 194324 9908
rect 192526 9876 192538 9880
rect 192480 9870 192538 9876
rect 194318 9868 194324 9880
rect 194376 9868 194382 9920
rect 267734 9868 267740 9920
rect 267792 9908 267798 9920
rect 270954 9908 270960 9920
rect 267792 9880 270960 9908
rect 267792 9868 267798 9880
rect 270954 9868 270960 9880
rect 271012 9868 271018 9920
rect 1104 9818 305808 9840
rect 1104 9766 77148 9818
rect 77200 9766 77212 9818
rect 77264 9766 77276 9818
rect 77328 9766 77340 9818
rect 77392 9766 77404 9818
rect 77456 9766 153346 9818
rect 153398 9766 153410 9818
rect 153462 9766 153474 9818
rect 153526 9766 153538 9818
rect 153590 9766 153602 9818
rect 153654 9766 229544 9818
rect 229596 9766 229608 9818
rect 229660 9766 229672 9818
rect 229724 9766 229736 9818
rect 229788 9766 229800 9818
rect 229852 9766 305808 9818
rect 1104 9744 305808 9766
rect 31202 9596 31208 9648
rect 31260 9636 31266 9648
rect 32860 9638 32918 9644
rect 32860 9636 32872 9638
rect 31260 9608 32872 9636
rect 31260 9596 31266 9608
rect 32860 9604 32872 9608
rect 32906 9604 32918 9638
rect 140682 9636 140688 9648
rect 140642 9608 140688 9636
rect 32860 9598 32918 9604
rect 140682 9596 140688 9608
rect 140740 9596 140746 9648
rect 156138 9636 156144 9648
rect 156098 9608 156144 9636
rect 156138 9596 156144 9608
rect 156196 9596 156202 9648
rect 157888 9638 157946 9644
rect 157888 9604 157900 9638
rect 157934 9636 157946 9638
rect 158622 9636 158628 9648
rect 157934 9608 158628 9636
rect 157934 9604 157946 9608
rect 157888 9598 157946 9604
rect 158622 9596 158628 9608
rect 158680 9596 158686 9648
rect 190638 9596 190644 9648
rect 190696 9636 190702 9648
rect 193032 9638 193090 9644
rect 190696 9608 192984 9636
rect 190696 9596 190702 9608
rect 27338 9528 27344 9580
rect 27396 9568 27402 9580
rect 31296 9570 31354 9576
rect 31296 9568 31308 9570
rect 27396 9540 31308 9568
rect 27396 9528 27402 9540
rect 31296 9536 31308 9540
rect 31342 9536 31354 9570
rect 31296 9530 31354 9536
rect 32124 9570 32182 9576
rect 32124 9536 32136 9570
rect 32170 9568 32182 9570
rect 32768 9570 32826 9576
rect 32768 9568 32780 9570
rect 32170 9540 32780 9568
rect 32170 9536 32182 9540
rect 32124 9530 32182 9536
rect 32768 9536 32780 9540
rect 32814 9568 32826 9570
rect 33686 9568 33692 9580
rect 32814 9540 33692 9568
rect 32814 9536 32826 9540
rect 32768 9530 32826 9536
rect 33686 9528 33692 9540
rect 33744 9528 33750 9580
rect 192956 9576 192984 9608
rect 193032 9604 193044 9638
rect 193078 9636 193090 9638
rect 193306 9636 193312 9648
rect 193078 9608 193312 9636
rect 193078 9604 193090 9608
rect 193032 9598 193090 9604
rect 193306 9596 193312 9608
rect 193364 9596 193370 9648
rect 267920 9638 267978 9644
rect 267920 9604 267932 9638
rect 267966 9636 267978 9638
rect 269850 9636 269856 9648
rect 267966 9608 269856 9636
rect 267966 9604 267978 9608
rect 267920 9598 267978 9604
rect 269850 9596 269856 9608
rect 269908 9596 269914 9648
rect 192480 9570 192538 9576
rect 192480 9536 192492 9570
rect 192526 9536 192538 9570
rect 192480 9530 192538 9536
rect 192940 9570 192998 9576
rect 192940 9536 192952 9570
rect 192986 9568 192998 9570
rect 194134 9568 194140 9580
rect 192986 9540 194140 9568
rect 192986 9536 192998 9540
rect 192940 9530 192998 9536
rect 30558 9460 30564 9512
rect 30616 9500 30622 9512
rect 32216 9502 32274 9508
rect 32216 9500 32228 9502
rect 30616 9472 32228 9500
rect 30616 9460 30622 9472
rect 32216 9468 32228 9472
rect 32262 9468 32274 9502
rect 192496 9500 192524 9530
rect 194134 9528 194140 9540
rect 194192 9528 194198 9580
rect 267828 9570 267886 9576
rect 267828 9536 267840 9570
rect 267874 9568 267886 9570
rect 268102 9568 268108 9580
rect 267874 9540 268108 9568
rect 267874 9536 267886 9540
rect 267828 9530 267886 9536
rect 268102 9528 268108 9540
rect 268160 9528 268166 9580
rect 195974 9500 195980 9512
rect 192496 9472 195980 9500
rect 32216 9462 32274 9468
rect 195974 9460 195980 9472
rect 196032 9460 196038 9512
rect 29914 9392 29920 9444
rect 29972 9432 29978 9444
rect 31112 9434 31170 9440
rect 31112 9432 31124 9434
rect 29972 9404 31124 9432
rect 29972 9392 29978 9404
rect 31112 9400 31124 9404
rect 31158 9400 31170 9434
rect 31112 9394 31170 9400
rect 192296 9434 192354 9440
rect 192296 9400 192308 9434
rect 192342 9432 192354 9434
rect 194502 9432 194508 9444
rect 192342 9404 194508 9432
rect 192342 9400 192354 9404
rect 192296 9394 192354 9400
rect 194502 9392 194508 9404
rect 194560 9392 194566 9444
rect 104250 9324 104256 9376
rect 104308 9364 104314 9376
rect 141972 9366 142030 9372
rect 141972 9364 141984 9366
rect 104308 9336 141984 9364
rect 104308 9324 104314 9336
rect 141972 9332 141984 9336
rect 142018 9364 142030 9366
rect 148318 9364 148324 9376
rect 142018 9336 148324 9364
rect 142018 9332 142030 9336
rect 141972 9326 142030 9332
rect 148318 9324 148324 9336
rect 148376 9324 148382 9376
rect 1104 9274 305808 9296
rect 1104 9222 39048 9274
rect 39100 9222 39112 9274
rect 39164 9222 39176 9274
rect 39228 9222 39240 9274
rect 39292 9222 39304 9274
rect 39356 9222 115246 9274
rect 115298 9222 115310 9274
rect 115362 9222 115374 9274
rect 115426 9222 115438 9274
rect 115490 9222 115502 9274
rect 115554 9222 191444 9274
rect 191496 9222 191508 9274
rect 191560 9222 191572 9274
rect 191624 9222 191636 9274
rect 191688 9222 191700 9274
rect 191752 9222 267642 9274
rect 267694 9222 267706 9274
rect 267758 9222 267770 9274
rect 267822 9222 267834 9274
rect 267886 9222 267898 9274
rect 267950 9222 305808 9274
rect 1104 9200 305808 9222
rect 1104 8730 305808 8752
rect 1104 8678 77148 8730
rect 77200 8678 77212 8730
rect 77264 8678 77276 8730
rect 77328 8678 77340 8730
rect 77392 8678 77404 8730
rect 77456 8678 153346 8730
rect 153398 8678 153410 8730
rect 153462 8678 153474 8730
rect 153526 8678 153538 8730
rect 153590 8678 153602 8730
rect 153654 8678 229544 8730
rect 229596 8678 229608 8730
rect 229660 8678 229672 8730
rect 229724 8678 229736 8730
rect 229788 8678 229800 8730
rect 229852 8678 305808 8730
rect 1104 8656 305808 8678
rect 1580 8482 1638 8488
rect 1580 8448 1592 8482
rect 1626 8480 1638 8482
rect 1626 8452 1992 8480
rect 1626 8448 1638 8452
rect 1580 8442 1638 8448
rect 1394 8344 1400 8356
rect 1354 8316 1400 8344
rect 1394 8304 1400 8316
rect 1452 8304 1458 8356
rect 1964 8352 1992 8452
rect 1948 8346 2006 8352
rect 1948 8312 1960 8346
rect 1994 8344 2006 8346
rect 2316 8346 2374 8352
rect 2316 8344 2328 8346
rect 1994 8316 2328 8344
rect 1994 8312 2006 8316
rect 1948 8306 2006 8312
rect 2316 8312 2328 8316
rect 2362 8344 2374 8346
rect 2684 8346 2742 8352
rect 2684 8344 2696 8346
rect 2362 8316 2696 8344
rect 2362 8312 2374 8316
rect 2316 8306 2374 8312
rect 2684 8312 2696 8316
rect 2730 8344 2742 8346
rect 3052 8346 3110 8352
rect 3052 8344 3064 8346
rect 2730 8316 3064 8344
rect 2730 8312 2742 8316
rect 2684 8306 2742 8312
rect 3052 8312 3064 8316
rect 3098 8344 3110 8346
rect 187510 8344 187516 8356
rect 3098 8316 187516 8344
rect 3098 8312 3110 8316
rect 3052 8306 3110 8312
rect 187510 8304 187516 8316
rect 187568 8304 187574 8356
rect 1104 8186 305808 8208
rect 1104 8134 39048 8186
rect 39100 8134 39112 8186
rect 39164 8134 39176 8186
rect 39228 8134 39240 8186
rect 39292 8134 39304 8186
rect 39356 8134 115246 8186
rect 115298 8134 115310 8186
rect 115362 8134 115374 8186
rect 115426 8134 115438 8186
rect 115490 8134 115502 8186
rect 115554 8134 191444 8186
rect 191496 8134 191508 8186
rect 191560 8134 191572 8186
rect 191624 8134 191636 8186
rect 191688 8134 191700 8186
rect 191752 8134 267642 8186
rect 267694 8134 267706 8186
rect 267758 8134 267770 8186
rect 267822 8134 267834 8186
rect 267886 8134 267898 8186
rect 267950 8134 305808 8186
rect 1104 8112 305808 8134
rect 1104 7642 305808 7664
rect 1104 7590 77148 7642
rect 77200 7590 77212 7642
rect 77264 7590 77276 7642
rect 77328 7590 77340 7642
rect 77392 7590 77404 7642
rect 77456 7590 153346 7642
rect 153398 7590 153410 7642
rect 153462 7590 153474 7642
rect 153526 7590 153538 7642
rect 153590 7590 153602 7642
rect 153654 7590 229544 7642
rect 229596 7590 229608 7642
rect 229660 7590 229672 7642
rect 229724 7590 229736 7642
rect 229788 7590 229800 7642
rect 229852 7590 305808 7642
rect 1104 7568 305808 7590
rect 1104 7098 305808 7120
rect 1104 7046 39048 7098
rect 39100 7046 39112 7098
rect 39164 7046 39176 7098
rect 39228 7046 39240 7098
rect 39292 7046 39304 7098
rect 39356 7046 115246 7098
rect 115298 7046 115310 7098
rect 115362 7046 115374 7098
rect 115426 7046 115438 7098
rect 115490 7046 115502 7098
rect 115554 7046 191444 7098
rect 191496 7046 191508 7098
rect 191560 7046 191572 7098
rect 191624 7046 191636 7098
rect 191688 7046 191700 7098
rect 191752 7046 267642 7098
rect 267694 7046 267706 7098
rect 267758 7046 267770 7098
rect 267822 7046 267834 7098
rect 267886 7046 267898 7098
rect 267950 7046 305808 7098
rect 1104 7024 305808 7046
rect 1104 6554 305808 6576
rect 1104 6502 77148 6554
rect 77200 6502 77212 6554
rect 77264 6502 77276 6554
rect 77328 6502 77340 6554
rect 77392 6502 77404 6554
rect 77456 6502 153346 6554
rect 153398 6502 153410 6554
rect 153462 6502 153474 6554
rect 153526 6502 153538 6554
rect 153590 6502 153602 6554
rect 153654 6502 229544 6554
rect 229596 6502 229608 6554
rect 229660 6502 229672 6554
rect 229724 6502 229736 6554
rect 229788 6502 229800 6554
rect 229852 6502 305808 6554
rect 1104 6480 305808 6502
rect 303982 6304 303988 6316
rect 303942 6276 303988 6304
rect 303982 6264 303988 6276
rect 304040 6264 304046 6316
rect 249058 6196 249064 6248
rect 249116 6236 249122 6248
rect 304260 6238 304318 6244
rect 304260 6236 304272 6238
rect 249116 6208 304272 6236
rect 249116 6196 249122 6208
rect 304260 6204 304272 6208
rect 304306 6204 304318 6238
rect 304260 6198 304318 6204
rect 1104 6010 305808 6032
rect 1104 5958 39048 6010
rect 39100 5958 39112 6010
rect 39164 5958 39176 6010
rect 39228 5958 39240 6010
rect 39292 5958 39304 6010
rect 39356 5958 115246 6010
rect 115298 5958 115310 6010
rect 115362 5958 115374 6010
rect 115426 5958 115438 6010
rect 115490 5958 115502 6010
rect 115554 5958 191444 6010
rect 191496 5958 191508 6010
rect 191560 5958 191572 6010
rect 191624 5958 191636 6010
rect 191688 5958 191700 6010
rect 191752 5958 267642 6010
rect 267694 5958 267706 6010
rect 267758 5958 267770 6010
rect 267822 5958 267834 6010
rect 267886 5958 267898 6010
rect 267950 5958 305808 6010
rect 1104 5936 305808 5958
rect 1104 5466 305808 5488
rect 1104 5414 77148 5466
rect 77200 5414 77212 5466
rect 77264 5414 77276 5466
rect 77328 5414 77340 5466
rect 77392 5414 77404 5466
rect 77456 5414 153346 5466
rect 153398 5414 153410 5466
rect 153462 5414 153474 5466
rect 153526 5414 153538 5466
rect 153590 5414 153602 5466
rect 153654 5414 229544 5466
rect 229596 5414 229608 5466
rect 229660 5414 229672 5466
rect 229724 5414 229736 5466
rect 229788 5414 229800 5466
rect 229852 5414 305808 5466
rect 1104 5392 305808 5414
rect 1104 4922 305808 4944
rect 1104 4870 39048 4922
rect 39100 4870 39112 4922
rect 39164 4870 39176 4922
rect 39228 4870 39240 4922
rect 39292 4870 39304 4922
rect 39356 4870 115246 4922
rect 115298 4870 115310 4922
rect 115362 4870 115374 4922
rect 115426 4870 115438 4922
rect 115490 4870 115502 4922
rect 115554 4870 191444 4922
rect 191496 4870 191508 4922
rect 191560 4870 191572 4922
rect 191624 4870 191636 4922
rect 191688 4870 191700 4922
rect 191752 4870 267642 4922
rect 267694 4870 267706 4922
rect 267758 4870 267770 4922
rect 267822 4870 267834 4922
rect 267886 4870 267898 4922
rect 267950 4870 305808 4922
rect 1104 4848 305808 4870
rect 1104 4378 305808 4400
rect 1104 4326 77148 4378
rect 77200 4326 77212 4378
rect 77264 4326 77276 4378
rect 77328 4326 77340 4378
rect 77392 4326 77404 4378
rect 77456 4326 153346 4378
rect 153398 4326 153410 4378
rect 153462 4326 153474 4378
rect 153526 4326 153538 4378
rect 153590 4326 153602 4378
rect 153654 4326 229544 4378
rect 229596 4326 229608 4378
rect 229660 4326 229672 4378
rect 229724 4326 229736 4378
rect 229788 4326 229800 4378
rect 229852 4326 305808 4378
rect 1104 4304 305808 4326
rect 1104 3834 305808 3856
rect 1104 3782 39048 3834
rect 39100 3782 39112 3834
rect 39164 3782 39176 3834
rect 39228 3782 39240 3834
rect 39292 3782 39304 3834
rect 39356 3782 115246 3834
rect 115298 3782 115310 3834
rect 115362 3782 115374 3834
rect 115426 3782 115438 3834
rect 115490 3782 115502 3834
rect 115554 3782 191444 3834
rect 191496 3782 191508 3834
rect 191560 3782 191572 3834
rect 191624 3782 191636 3834
rect 191688 3782 191700 3834
rect 191752 3782 267642 3834
rect 267694 3782 267706 3834
rect 267758 3782 267770 3834
rect 267822 3782 267834 3834
rect 267886 3782 267898 3834
rect 267950 3782 305808 3834
rect 1104 3760 305808 3782
rect 1104 3290 305808 3312
rect 1104 3238 77148 3290
rect 77200 3238 77212 3290
rect 77264 3238 77276 3290
rect 77328 3238 77340 3290
rect 77392 3238 77404 3290
rect 77456 3238 153346 3290
rect 153398 3238 153410 3290
rect 153462 3238 153474 3290
rect 153526 3238 153538 3290
rect 153590 3238 153602 3290
rect 153654 3238 229544 3290
rect 229596 3238 229608 3290
rect 229660 3238 229672 3290
rect 229724 3238 229736 3290
rect 229788 3238 229800 3290
rect 229852 3238 305808 3290
rect 1104 3216 305808 3238
rect 1104 2746 305808 2768
rect 1104 2694 39048 2746
rect 39100 2694 39112 2746
rect 39164 2694 39176 2746
rect 39228 2694 39240 2746
rect 39292 2694 39304 2746
rect 39356 2694 115246 2746
rect 115298 2694 115310 2746
rect 115362 2694 115374 2746
rect 115426 2694 115438 2746
rect 115490 2694 115502 2746
rect 115554 2694 191444 2746
rect 191496 2694 191508 2746
rect 191560 2694 191572 2746
rect 191624 2694 191636 2746
rect 191688 2694 191700 2746
rect 191752 2694 267642 2746
rect 267694 2694 267706 2746
rect 267758 2694 267770 2746
rect 267822 2694 267834 2746
rect 267886 2694 267898 2746
rect 267950 2694 305808 2746
rect 1104 2672 305808 2694
rect 149422 2592 149428 2644
rect 149480 2632 149486 2644
rect 302234 2632 302240 2644
rect 149480 2604 302240 2632
rect 149480 2592 149486 2604
rect 302234 2592 302240 2604
rect 302292 2592 302298 2644
rect 1104 2202 305808 2224
rect 1104 2150 77148 2202
rect 77200 2150 77212 2202
rect 77264 2150 77276 2202
rect 77328 2150 77340 2202
rect 77392 2150 77404 2202
rect 77456 2150 153346 2202
rect 153398 2150 153410 2202
rect 153462 2150 153474 2202
rect 153526 2150 153538 2202
rect 153590 2150 153602 2202
rect 153654 2150 229544 2202
rect 229596 2150 229608 2202
rect 229660 2150 229672 2202
rect 229724 2150 229736 2202
rect 229788 2150 229800 2202
rect 229852 2150 305808 2202
rect 1104 2128 305808 2150
<< via1 >>
rect 29000 13744 29052 13796
rect 32956 13744 33008 13796
rect 46204 13744 46256 13796
rect 63408 13744 63460 13796
rect 69296 13744 69348 13796
rect 75368 13744 75420 13796
rect 76012 13744 76064 13796
rect 90640 13744 90692 13796
rect 102416 13744 102468 13796
rect 113824 13744 113876 13796
rect 125508 13744 125560 13796
rect 131856 13744 131908 13796
rect 161664 13744 161716 13796
rect 166080 13744 166132 13796
rect 167368 13744 167420 13796
rect 174176 13744 174228 13796
rect 177764 13744 177816 13796
rect 181904 13744 181956 13796
rect 189908 13812 189960 13864
rect 189356 13744 189408 13796
rect 193220 13744 193272 13796
rect 195980 13744 196032 13796
rect 302792 13744 302844 13796
rect 27160 13676 27212 13728
rect 36544 13676 36596 13728
rect 42524 13676 42576 13728
rect 47860 13676 47912 13728
rect 51632 13676 51684 13728
rect 54116 13676 54168 13728
rect 66168 13676 66220 13728
rect 72424 13676 72476 13728
rect 73896 13676 73948 13728
rect 76380 13676 76432 13728
rect 83096 13676 83148 13728
rect 86408 13676 86460 13728
rect 91836 13676 91888 13728
rect 101956 13676 102008 13728
rect 114652 13676 114704 13728
rect 127440 13676 127492 13728
rect 127532 13676 127584 13728
rect 129740 13676 129792 13728
rect 133604 13676 133656 13728
rect 136824 13676 136876 13728
rect 148140 13676 148192 13728
rect 150440 13676 150492 13728
rect 157156 13676 157208 13728
rect 301412 13676 301464 13728
rect 39048 13574 39100 13626
rect 39112 13574 39164 13626
rect 39176 13574 39228 13626
rect 39240 13574 39292 13626
rect 39304 13574 39356 13626
rect 115246 13574 115298 13626
rect 115310 13574 115362 13626
rect 115374 13574 115426 13626
rect 115438 13574 115490 13626
rect 115502 13574 115554 13626
rect 191444 13574 191496 13626
rect 191508 13574 191560 13626
rect 191572 13574 191624 13626
rect 191636 13574 191688 13626
rect 191700 13574 191752 13626
rect 267642 13574 267694 13626
rect 267706 13574 267758 13626
rect 267770 13574 267822 13626
rect 267834 13574 267886 13626
rect 267898 13574 267950 13626
rect 1584 13514 1636 13524
rect 1584 13480 1592 13514
rect 1592 13480 1626 13514
rect 1626 13480 1636 13514
rect 1584 13472 1636 13480
rect 4620 13514 4672 13524
rect 4620 13480 4628 13514
rect 4628 13480 4662 13514
rect 4662 13480 4672 13514
rect 4620 13472 4672 13480
rect 7656 13514 7708 13524
rect 7656 13480 7664 13514
rect 7664 13480 7698 13514
rect 7698 13480 7708 13514
rect 7656 13472 7708 13480
rect 10784 13514 10836 13524
rect 10784 13480 10792 13514
rect 10792 13480 10826 13514
rect 10826 13480 10836 13514
rect 10784 13472 10836 13480
rect 13820 13472 13872 13524
rect 16856 13514 16908 13524
rect 16856 13480 16864 13514
rect 16864 13480 16898 13514
rect 16898 13480 16908 13514
rect 16856 13472 16908 13480
rect 19984 13514 20036 13524
rect 19984 13480 19992 13514
rect 19992 13480 20026 13514
rect 20026 13480 20036 13514
rect 19984 13472 20036 13480
rect 23020 13514 23072 13524
rect 23020 13480 23028 13514
rect 23028 13480 23062 13514
rect 23062 13480 23072 13514
rect 23020 13472 23072 13480
rect 27620 13472 27672 13524
rect 27712 13472 27764 13524
rect 30472 13472 30524 13524
rect 36544 13472 36596 13524
rect 46204 13472 46256 13524
rect 47584 13514 47636 13524
rect 47584 13480 47592 13514
rect 47592 13480 47626 13514
rect 47626 13480 47636 13514
rect 47584 13472 47636 13480
rect 50528 13472 50580 13524
rect 53012 13472 53064 13524
rect 55588 13472 55640 13524
rect 57888 13472 57940 13524
rect 61752 13472 61804 13524
rect 63408 13472 63460 13524
rect 142896 13514 142948 13524
rect 27160 13404 27212 13456
rect 44180 13404 44232 13456
rect 4804 13310 4856 13320
rect 4804 13276 4812 13310
rect 4812 13276 4846 13310
rect 4846 13276 4856 13310
rect 4804 13268 4856 13276
rect 14280 13310 14332 13320
rect 14280 13276 14288 13310
rect 14288 13276 14322 13310
rect 14322 13276 14332 13310
rect 14280 13268 14332 13276
rect 17040 13310 17092 13320
rect 17040 13276 17048 13310
rect 17048 13276 17082 13310
rect 17082 13276 17092 13310
rect 17040 13268 17092 13276
rect 20168 13310 20220 13320
rect 20168 13276 20176 13310
rect 20176 13276 20210 13310
rect 20210 13276 20220 13310
rect 20168 13268 20220 13276
rect 23204 13310 23256 13320
rect 23204 13276 23212 13310
rect 23212 13276 23246 13310
rect 23246 13276 23256 13310
rect 23204 13268 23256 13276
rect 26976 13336 27028 13388
rect 29828 13310 29880 13320
rect 29828 13276 29836 13310
rect 29836 13276 29870 13310
rect 29870 13276 29880 13310
rect 29828 13268 29880 13276
rect 32404 13310 32456 13320
rect 32404 13276 32412 13310
rect 32412 13276 32446 13310
rect 32446 13276 32456 13310
rect 32404 13268 32456 13276
rect 33784 13268 33836 13320
rect 44364 13404 44416 13456
rect 45560 13378 45612 13388
rect 45560 13344 45568 13378
rect 45568 13344 45602 13378
rect 45602 13344 45612 13378
rect 51632 13378 51684 13388
rect 45560 13336 45612 13344
rect 51632 13344 51640 13378
rect 51640 13344 51674 13378
rect 51674 13344 51684 13378
rect 51632 13336 51684 13344
rect 59820 13404 59872 13456
rect 63040 13446 63092 13456
rect 63040 13412 63048 13446
rect 63048 13412 63082 13446
rect 63082 13412 63092 13446
rect 63040 13404 63092 13412
rect 75368 13446 75420 13456
rect 72700 13378 72752 13388
rect 27528 13242 27580 13252
rect 27252 13132 27304 13184
rect 27528 13208 27536 13242
rect 27536 13208 27570 13242
rect 27570 13208 27580 13242
rect 27528 13200 27580 13208
rect 27712 13132 27764 13184
rect 30196 13200 30248 13252
rect 32680 13242 32732 13252
rect 30472 13132 30524 13184
rect 32680 13208 32688 13242
rect 32688 13208 32722 13242
rect 32722 13208 32732 13242
rect 32680 13200 32732 13208
rect 34520 13200 34572 13252
rect 35992 13200 36044 13252
rect 33600 13132 33652 13184
rect 34152 13174 34204 13184
rect 34152 13140 34160 13174
rect 34160 13140 34194 13174
rect 34194 13140 34204 13174
rect 34152 13132 34204 13140
rect 34336 13132 34388 13184
rect 37464 13132 37516 13184
rect 38936 13268 38988 13320
rect 37832 13242 37884 13252
rect 37832 13208 37840 13242
rect 37840 13208 37874 13242
rect 37874 13208 37884 13242
rect 37832 13200 37884 13208
rect 42524 13310 42576 13320
rect 39304 13174 39356 13184
rect 39304 13140 39312 13174
rect 39312 13140 39346 13174
rect 39346 13140 39356 13174
rect 39304 13132 39356 13140
rect 39948 13132 40000 13184
rect 42524 13276 42532 13310
rect 42532 13276 42566 13310
rect 42566 13276 42576 13310
rect 42524 13268 42576 13276
rect 44272 13268 44324 13320
rect 51356 13310 51408 13320
rect 40408 13242 40460 13252
rect 40408 13208 40416 13242
rect 40416 13208 40450 13242
rect 40450 13208 40460 13242
rect 40408 13200 40460 13208
rect 41420 13200 41472 13252
rect 42892 13200 42944 13252
rect 43260 13200 43312 13252
rect 42432 13132 42484 13184
rect 45008 13174 45060 13184
rect 45008 13140 45016 13174
rect 45016 13140 45050 13174
rect 45050 13140 45060 13174
rect 45008 13132 45060 13140
rect 45376 13174 45428 13184
rect 45376 13140 45384 13174
rect 45384 13140 45418 13174
rect 45418 13140 45428 13174
rect 45376 13132 45428 13140
rect 51356 13276 51364 13310
rect 51364 13276 51398 13310
rect 51398 13276 51408 13310
rect 51356 13268 51408 13276
rect 47860 13200 47912 13252
rect 54392 13268 54444 13320
rect 54760 13268 54812 13320
rect 55588 13310 55640 13320
rect 55588 13276 55596 13310
rect 55596 13276 55630 13310
rect 55630 13276 55640 13310
rect 55588 13268 55640 13276
rect 57888 13310 57940 13320
rect 57888 13276 57896 13310
rect 57896 13276 57930 13310
rect 57930 13276 57940 13310
rect 57888 13268 57940 13276
rect 60648 13310 60700 13320
rect 60648 13276 60656 13310
rect 60656 13276 60690 13310
rect 60690 13276 60700 13310
rect 60648 13268 60700 13276
rect 53288 13242 53340 13252
rect 53288 13208 53296 13242
rect 53296 13208 53330 13242
rect 53330 13208 53340 13242
rect 53288 13200 53340 13208
rect 55864 13242 55916 13252
rect 54668 13132 54720 13184
rect 55864 13208 55872 13242
rect 55872 13208 55906 13242
rect 55906 13208 55916 13242
rect 55864 13200 55916 13208
rect 56600 13200 56652 13252
rect 57336 13174 57388 13184
rect 57336 13140 57344 13174
rect 57344 13140 57378 13174
rect 57378 13140 57388 13174
rect 57336 13132 57388 13140
rect 57704 13200 57756 13252
rect 58624 13200 58676 13252
rect 61476 13200 61528 13252
rect 59636 13174 59688 13184
rect 59636 13140 59644 13174
rect 59644 13140 59678 13174
rect 59678 13140 59688 13174
rect 66168 13310 66220 13320
rect 66168 13276 66176 13310
rect 66176 13276 66210 13310
rect 66210 13276 66220 13310
rect 66168 13268 66220 13276
rect 69296 13310 69348 13320
rect 69296 13276 69304 13310
rect 69304 13276 69338 13310
rect 69338 13276 69348 13310
rect 69296 13268 69348 13276
rect 72700 13344 72708 13378
rect 72708 13344 72742 13378
rect 72742 13344 72752 13378
rect 72700 13336 72752 13344
rect 75368 13412 75376 13446
rect 75376 13412 75410 13446
rect 75410 13412 75420 13446
rect 75368 13404 75420 13412
rect 75644 13404 75696 13456
rect 80244 13378 80296 13388
rect 80244 13344 80252 13378
rect 80252 13344 80286 13378
rect 80286 13344 80296 13378
rect 80244 13336 80296 13344
rect 81624 13378 81676 13388
rect 81624 13344 81632 13378
rect 81632 13344 81666 13378
rect 81666 13344 81676 13378
rect 93860 13404 93912 13456
rect 81624 13336 81676 13344
rect 61752 13200 61804 13252
rect 59636 13132 59688 13140
rect 61660 13132 61712 13184
rect 65892 13132 65944 13184
rect 65984 13174 66036 13184
rect 65984 13140 65992 13174
rect 65992 13140 66026 13174
rect 66026 13140 66036 13174
rect 69112 13174 69164 13184
rect 65984 13132 66036 13140
rect 69112 13140 69120 13174
rect 69120 13140 69154 13174
rect 69154 13140 69164 13174
rect 69112 13132 69164 13140
rect 72332 13132 72384 13184
rect 72424 13174 72476 13184
rect 72424 13140 72432 13174
rect 72432 13140 72466 13174
rect 72466 13140 72476 13174
rect 73896 13242 73948 13252
rect 73896 13208 73904 13242
rect 73904 13208 73938 13242
rect 73938 13208 73948 13242
rect 73896 13200 73948 13208
rect 75184 13200 75236 13252
rect 78404 13268 78456 13320
rect 81440 13268 81492 13320
rect 83096 13310 83148 13320
rect 76472 13242 76524 13252
rect 76472 13208 76480 13242
rect 76480 13208 76514 13242
rect 76514 13208 76524 13242
rect 76472 13200 76524 13208
rect 78772 13242 78824 13252
rect 72424 13132 72476 13140
rect 77944 13174 77996 13184
rect 77944 13140 77952 13174
rect 77952 13140 77986 13174
rect 77986 13140 77996 13174
rect 78772 13208 78780 13242
rect 78780 13208 78814 13242
rect 78814 13208 78824 13242
rect 78772 13200 78824 13208
rect 79324 13200 79376 13252
rect 80060 13200 80112 13252
rect 83096 13276 83104 13310
rect 83104 13276 83138 13310
rect 83138 13276 83148 13310
rect 83096 13268 83148 13276
rect 83924 13310 83976 13320
rect 83924 13276 83932 13310
rect 83932 13276 83966 13310
rect 83966 13276 83976 13310
rect 83924 13268 83976 13276
rect 77944 13132 77996 13140
rect 80796 13132 80848 13184
rect 81440 13174 81492 13184
rect 81440 13140 81448 13174
rect 81448 13140 81482 13174
rect 81482 13140 81492 13174
rect 81440 13132 81492 13140
rect 83832 13200 83884 13252
rect 84476 13200 84528 13252
rect 85488 13200 85540 13252
rect 82912 13174 82964 13184
rect 82912 13140 82920 13174
rect 82920 13140 82954 13174
rect 82954 13140 82964 13174
rect 82912 13132 82964 13140
rect 83924 13132 83976 13184
rect 86040 13132 86092 13184
rect 87880 13268 87932 13320
rect 86776 13242 86828 13252
rect 86776 13208 86784 13242
rect 86784 13208 86818 13242
rect 86818 13208 86828 13242
rect 86776 13200 86828 13208
rect 88248 13174 88300 13184
rect 88248 13140 88256 13174
rect 88256 13140 88290 13174
rect 88290 13140 88300 13174
rect 88248 13132 88300 13140
rect 89076 13242 89128 13252
rect 89076 13208 89084 13242
rect 89084 13208 89118 13242
rect 89118 13208 89128 13242
rect 89076 13200 89128 13208
rect 89536 13200 89588 13252
rect 91652 13200 91704 13252
rect 91836 13242 91888 13252
rect 91836 13208 91844 13242
rect 91844 13208 91878 13242
rect 91878 13208 91888 13242
rect 91836 13200 91888 13208
rect 92020 13242 92072 13252
rect 92020 13208 92028 13242
rect 92028 13208 92062 13242
rect 92062 13208 92072 13242
rect 92020 13200 92072 13208
rect 90548 13174 90600 13184
rect 90548 13140 90556 13174
rect 90556 13140 90590 13174
rect 90590 13140 90600 13174
rect 99104 13336 99156 13388
rect 100760 13404 100812 13456
rect 109040 13404 109092 13456
rect 111708 13404 111760 13456
rect 118884 13404 118936 13456
rect 121276 13446 121328 13456
rect 118240 13336 118292 13388
rect 121276 13412 121284 13446
rect 121284 13412 121318 13446
rect 121318 13412 121328 13446
rect 121276 13404 121328 13412
rect 124128 13446 124180 13456
rect 124128 13412 124136 13446
rect 124136 13412 124170 13446
rect 124170 13412 124180 13446
rect 124128 13404 124180 13412
rect 127532 13404 127584 13456
rect 136640 13446 136692 13456
rect 136640 13412 136648 13446
rect 136648 13412 136682 13446
rect 136682 13412 136692 13446
rect 136640 13404 136692 13412
rect 139584 13404 139636 13456
rect 142896 13480 142904 13514
rect 142904 13480 142938 13514
rect 142938 13480 142948 13514
rect 142896 13472 142948 13480
rect 145748 13472 145800 13524
rect 148140 13472 148192 13524
rect 150808 13472 150860 13524
rect 96712 13174 96764 13184
rect 90548 13132 90600 13140
rect 96712 13140 96720 13174
rect 96720 13140 96754 13174
rect 96754 13140 96764 13174
rect 96712 13132 96764 13140
rect 97540 13174 97592 13184
rect 97540 13140 97548 13174
rect 97548 13140 97582 13174
rect 97582 13140 97592 13174
rect 97540 13132 97592 13140
rect 98000 13200 98052 13252
rect 99196 13200 99248 13252
rect 101404 13268 101456 13320
rect 99656 13242 99708 13252
rect 99656 13208 99664 13242
rect 99664 13208 99698 13242
rect 99698 13208 99708 13242
rect 99656 13200 99708 13208
rect 100944 13200 100996 13252
rect 101036 13132 101088 13184
rect 103336 13268 103388 13320
rect 104256 13310 104308 13320
rect 102232 13242 102284 13252
rect 102232 13208 102240 13242
rect 102240 13208 102274 13242
rect 102274 13208 102284 13242
rect 102232 13200 102284 13208
rect 104256 13276 104264 13310
rect 104264 13276 104298 13310
rect 104298 13276 104308 13310
rect 104256 13268 104308 13276
rect 109592 13310 109644 13320
rect 109592 13276 109600 13310
rect 109600 13276 109634 13310
rect 109634 13276 109644 13310
rect 109592 13268 109644 13276
rect 111432 13310 111484 13320
rect 111432 13276 111440 13310
rect 111440 13276 111474 13310
rect 111474 13276 111484 13310
rect 111432 13268 111484 13276
rect 114836 13310 114888 13320
rect 114836 13276 114844 13310
rect 114844 13276 114878 13310
rect 114878 13276 114888 13310
rect 114836 13268 114888 13276
rect 117412 13310 117464 13320
rect 117412 13276 117420 13310
rect 117420 13276 117454 13310
rect 117454 13276 117464 13310
rect 117412 13268 117464 13276
rect 118792 13268 118844 13320
rect 130292 13378 130344 13388
rect 130292 13344 130300 13378
rect 130300 13344 130334 13378
rect 130334 13344 130344 13378
rect 130292 13336 130344 13344
rect 142068 13336 142120 13388
rect 104072 13200 104124 13252
rect 104992 13200 105044 13252
rect 112536 13242 112588 13252
rect 112536 13208 112544 13242
rect 112544 13208 112578 13242
rect 112578 13208 112588 13242
rect 112536 13200 112588 13208
rect 114192 13200 114244 13252
rect 115112 13242 115164 13252
rect 115112 13208 115120 13242
rect 115120 13208 115154 13242
rect 115154 13208 115164 13242
rect 115112 13200 115164 13208
rect 116952 13200 117004 13252
rect 117688 13242 117740 13252
rect 117688 13208 117696 13242
rect 117696 13208 117730 13242
rect 117730 13208 117740 13242
rect 117688 13200 117740 13208
rect 103704 13174 103756 13184
rect 103704 13140 103712 13174
rect 103712 13140 103746 13174
rect 103746 13140 103756 13174
rect 103704 13132 103756 13140
rect 104440 13132 104492 13184
rect 104624 13132 104676 13184
rect 109592 13132 109644 13184
rect 114560 13132 114612 13184
rect 114928 13132 114980 13184
rect 115756 13132 115808 13184
rect 118056 13132 118108 13184
rect 127532 13310 127584 13320
rect 127532 13276 127540 13310
rect 127540 13276 127574 13310
rect 127574 13276 127584 13310
rect 127532 13268 127584 13276
rect 129372 13268 129424 13320
rect 136824 13310 136876 13320
rect 136824 13276 136832 13310
rect 136832 13276 136866 13310
rect 136866 13276 136876 13310
rect 136824 13268 136876 13276
rect 143080 13310 143132 13320
rect 125508 13242 125560 13252
rect 125508 13208 125516 13242
rect 125516 13208 125550 13242
rect 125550 13208 125560 13242
rect 125508 13200 125560 13208
rect 127808 13242 127860 13252
rect 127808 13208 127816 13242
rect 127816 13208 127850 13242
rect 127850 13208 127860 13242
rect 127808 13200 127860 13208
rect 119712 13174 119764 13184
rect 119712 13140 119720 13174
rect 119720 13140 119754 13174
rect 119754 13140 119764 13174
rect 119712 13132 119764 13140
rect 126152 13174 126204 13184
rect 126152 13140 126160 13174
rect 126160 13140 126194 13174
rect 126194 13140 126204 13174
rect 126152 13132 126204 13140
rect 126520 13174 126572 13184
rect 126520 13140 126528 13174
rect 126528 13140 126562 13174
rect 126562 13140 126572 13174
rect 126520 13132 126572 13140
rect 128084 13132 128136 13184
rect 131212 13200 131264 13252
rect 132868 13242 132920 13252
rect 132868 13208 132876 13242
rect 132876 13208 132910 13242
rect 132910 13208 132920 13242
rect 132868 13200 132920 13208
rect 133328 13200 133380 13252
rect 143080 13276 143088 13310
rect 143088 13276 143122 13310
rect 143122 13276 143132 13310
rect 143080 13268 143132 13276
rect 145748 13310 145800 13320
rect 145748 13276 145756 13310
rect 145756 13276 145790 13310
rect 145790 13276 145800 13310
rect 145748 13268 145800 13276
rect 157248 13472 157300 13524
rect 157984 13472 158036 13524
rect 159456 13472 159508 13524
rect 161572 13472 161624 13524
rect 162676 13472 162728 13524
rect 163504 13472 163556 13524
rect 176384 13472 176436 13524
rect 182732 13514 182784 13524
rect 154948 13404 155000 13456
rect 166448 13404 166500 13456
rect 170404 13446 170456 13456
rect 160928 13378 160980 13388
rect 160928 13344 160936 13378
rect 160936 13344 160970 13378
rect 160970 13344 160980 13378
rect 160928 13336 160980 13344
rect 165252 13336 165304 13388
rect 129188 13132 129240 13184
rect 131580 13132 131632 13184
rect 133696 13132 133748 13184
rect 134156 13132 134208 13184
rect 145932 13200 145984 13252
rect 146024 13242 146076 13252
rect 146024 13208 146032 13242
rect 146032 13208 146066 13242
rect 146066 13208 146076 13242
rect 146024 13200 146076 13208
rect 147588 13200 147640 13252
rect 145840 13132 145892 13184
rect 147496 13174 147548 13184
rect 147496 13140 147504 13174
rect 147504 13140 147538 13174
rect 147538 13140 147548 13174
rect 147496 13132 147548 13140
rect 155224 13268 155276 13320
rect 155868 13268 155920 13320
rect 156420 13310 156472 13320
rect 156420 13276 156428 13310
rect 156428 13276 156462 13310
rect 156462 13276 156472 13310
rect 156420 13268 156472 13276
rect 157800 13310 157852 13320
rect 157800 13276 157808 13310
rect 157808 13276 157842 13310
rect 157842 13276 157852 13310
rect 157800 13268 157852 13276
rect 158628 13310 158680 13320
rect 158628 13276 158636 13310
rect 158636 13276 158670 13310
rect 158670 13276 158680 13310
rect 158628 13268 158680 13276
rect 162676 13268 162728 13320
rect 163504 13310 163556 13320
rect 149244 13132 149296 13184
rect 150440 13200 150492 13252
rect 151084 13200 151136 13252
rect 152464 13200 152516 13252
rect 153752 13242 153804 13252
rect 152648 13174 152700 13184
rect 152648 13140 152656 13174
rect 152656 13140 152690 13174
rect 152690 13140 152700 13174
rect 153752 13208 153760 13242
rect 153760 13208 153794 13242
rect 153794 13208 153804 13242
rect 153752 13200 153804 13208
rect 154212 13200 154264 13252
rect 156604 13200 156656 13252
rect 158904 13242 158956 13252
rect 155224 13174 155276 13184
rect 152648 13132 152700 13140
rect 155224 13140 155232 13174
rect 155232 13140 155266 13174
rect 155266 13140 155276 13174
rect 155224 13132 155276 13140
rect 158904 13208 158912 13242
rect 158912 13208 158946 13242
rect 158946 13208 158956 13242
rect 158904 13200 158956 13208
rect 161204 13242 161256 13252
rect 159548 13132 159600 13184
rect 160376 13174 160428 13184
rect 160376 13140 160384 13174
rect 160384 13140 160418 13174
rect 160418 13140 160428 13174
rect 160376 13132 160428 13140
rect 161204 13208 161212 13242
rect 161212 13208 161246 13242
rect 161246 13208 161256 13242
rect 161204 13200 161256 13208
rect 162768 13200 162820 13252
rect 162032 13132 162084 13184
rect 162492 13132 162544 13184
rect 163504 13276 163512 13310
rect 163512 13276 163546 13310
rect 163546 13276 163556 13310
rect 163504 13268 163556 13276
rect 164884 13268 164936 13320
rect 170404 13412 170412 13446
rect 170412 13412 170446 13446
rect 170446 13412 170456 13446
rect 170404 13404 170456 13412
rect 173072 13446 173124 13456
rect 173072 13412 173080 13446
rect 173080 13412 173114 13446
rect 173114 13412 173124 13446
rect 173072 13404 173124 13412
rect 173808 13446 173860 13456
rect 173808 13412 173816 13446
rect 173816 13412 173850 13446
rect 173850 13412 173860 13446
rect 173808 13404 173860 13412
rect 175924 13404 175976 13456
rect 176016 13404 176068 13456
rect 177764 13404 177816 13456
rect 180432 13404 180484 13456
rect 163780 13242 163832 13252
rect 163780 13208 163788 13242
rect 163788 13208 163822 13242
rect 163822 13208 163832 13242
rect 163780 13200 163832 13208
rect 164608 13132 164660 13184
rect 165160 13200 165212 13252
rect 167368 13242 167420 13252
rect 167368 13208 167376 13242
rect 167376 13208 167410 13242
rect 167410 13208 167420 13242
rect 167368 13200 167420 13208
rect 174176 13310 174228 13320
rect 174176 13276 174184 13310
rect 174184 13276 174218 13310
rect 174218 13276 174228 13310
rect 174176 13268 174228 13276
rect 165252 13174 165304 13184
rect 165252 13140 165260 13174
rect 165260 13140 165294 13174
rect 165294 13140 165304 13174
rect 165252 13132 165304 13140
rect 165344 13132 165396 13184
rect 166448 13174 166500 13184
rect 166448 13140 166456 13174
rect 166456 13140 166490 13174
rect 166490 13140 166500 13174
rect 166448 13132 166500 13140
rect 175832 13268 175884 13320
rect 181904 13336 181956 13388
rect 182088 13378 182140 13388
rect 182088 13344 182096 13378
rect 182096 13344 182130 13378
rect 182130 13344 182140 13378
rect 182732 13480 182740 13514
rect 182740 13480 182774 13514
rect 182774 13480 182784 13514
rect 182732 13472 182784 13480
rect 185768 13514 185820 13524
rect 185768 13480 185776 13514
rect 185776 13480 185810 13514
rect 185810 13480 185820 13514
rect 185768 13472 185820 13480
rect 189356 13472 189408 13524
rect 188804 13404 188856 13456
rect 189540 13404 189592 13456
rect 190920 13472 190972 13524
rect 193496 13472 193548 13524
rect 188528 13378 188580 13388
rect 182088 13336 182140 13344
rect 176384 13310 176436 13320
rect 176384 13276 176392 13310
rect 176392 13276 176426 13310
rect 176426 13276 176436 13310
rect 176384 13268 176436 13276
rect 180616 13268 180668 13320
rect 188528 13344 188536 13378
rect 188536 13344 188570 13378
rect 188570 13344 188580 13378
rect 188528 13336 188580 13344
rect 191840 13404 191892 13456
rect 207112 13472 207164 13524
rect 210332 13514 210384 13524
rect 189908 13336 189960 13388
rect 201960 13404 202012 13456
rect 203432 13404 203484 13456
rect 206008 13404 206060 13456
rect 207756 13404 207808 13456
rect 197636 13336 197688 13388
rect 202052 13336 202104 13388
rect 189540 13310 189592 13320
rect 175740 13200 175792 13252
rect 177672 13200 177724 13252
rect 175004 13132 175056 13184
rect 179972 13200 180024 13252
rect 180892 13200 180944 13252
rect 180708 13174 180760 13184
rect 180708 13140 180716 13174
rect 180716 13140 180750 13174
rect 180750 13140 180760 13174
rect 180708 13132 180760 13140
rect 189540 13276 189548 13310
rect 189548 13276 189582 13310
rect 189582 13276 189592 13310
rect 189540 13268 189592 13276
rect 187792 13132 187844 13184
rect 187976 13174 188028 13184
rect 187976 13140 187984 13174
rect 187984 13140 188018 13174
rect 188018 13140 188028 13174
rect 187976 13132 188028 13140
rect 188344 13174 188396 13184
rect 188344 13140 188352 13174
rect 188352 13140 188386 13174
rect 188386 13140 188396 13174
rect 188344 13132 188396 13140
rect 189540 13132 189592 13184
rect 191380 13132 191432 13184
rect 192392 13200 192444 13252
rect 193404 13200 193456 13252
rect 193956 13200 194008 13252
rect 201500 13268 201552 13320
rect 202144 13310 202196 13320
rect 202144 13276 202152 13310
rect 202152 13276 202186 13310
rect 202186 13276 202196 13310
rect 202144 13268 202196 13276
rect 194600 13200 194652 13252
rect 194784 13200 194836 13252
rect 196440 13242 196492 13252
rect 196440 13208 196448 13242
rect 196448 13208 196482 13242
rect 196482 13208 196492 13242
rect 196440 13200 196492 13208
rect 197360 13200 197412 13252
rect 202420 13242 202472 13252
rect 197728 13132 197780 13184
rect 197912 13132 197964 13184
rect 198556 13174 198608 13184
rect 198556 13140 198564 13174
rect 198564 13140 198598 13174
rect 198598 13140 198608 13174
rect 198556 13132 198608 13140
rect 200488 13174 200540 13184
rect 200488 13140 200496 13174
rect 200496 13140 200530 13174
rect 200530 13140 200540 13174
rect 200488 13132 200540 13140
rect 200856 13174 200908 13184
rect 200856 13140 200864 13174
rect 200864 13140 200898 13174
rect 200898 13140 200908 13174
rect 200856 13132 200908 13140
rect 201316 13132 201368 13184
rect 202420 13208 202428 13242
rect 202428 13208 202462 13242
rect 202462 13208 202472 13242
rect 202420 13200 202472 13208
rect 203156 13200 203208 13252
rect 204260 13200 204312 13252
rect 205456 13200 205508 13252
rect 205640 13132 205692 13184
rect 205732 13132 205784 13184
rect 207204 13268 207256 13320
rect 206376 13200 206428 13252
rect 207572 13200 207624 13252
rect 210332 13480 210340 13514
rect 210340 13480 210374 13514
rect 210374 13480 210384 13514
rect 210332 13472 210384 13480
rect 213368 13514 213420 13524
rect 213368 13480 213376 13514
rect 213376 13480 213410 13514
rect 213410 13480 213420 13514
rect 213368 13472 213420 13480
rect 208032 13404 208084 13456
rect 213276 13404 213328 13456
rect 268936 13472 268988 13524
rect 269580 13472 269632 13524
rect 271788 13472 271840 13524
rect 274916 13514 274968 13524
rect 274916 13480 274924 13514
rect 274924 13480 274958 13514
rect 274958 13480 274968 13514
rect 274916 13472 274968 13480
rect 277860 13514 277912 13524
rect 277860 13480 277868 13514
rect 277868 13480 277902 13514
rect 277902 13480 277912 13514
rect 277860 13472 277912 13480
rect 280896 13514 280948 13524
rect 280896 13480 280904 13514
rect 280904 13480 280938 13514
rect 280938 13480 280948 13514
rect 280896 13472 280948 13480
rect 284300 13472 284352 13524
rect 287060 13472 287112 13524
rect 290096 13514 290148 13524
rect 290096 13480 290104 13514
rect 290104 13480 290138 13514
rect 290138 13480 290148 13514
rect 290096 13472 290148 13480
rect 293224 13514 293276 13524
rect 293224 13480 293232 13514
rect 293232 13480 293266 13514
rect 293266 13480 293276 13514
rect 293224 13472 293276 13480
rect 296260 13514 296312 13524
rect 296260 13480 296268 13514
rect 296268 13480 296302 13514
rect 296302 13480 296312 13514
rect 296260 13472 296312 13480
rect 299296 13514 299348 13524
rect 299296 13480 299304 13514
rect 299304 13480 299338 13514
rect 299338 13480 299348 13514
rect 299296 13472 299348 13480
rect 301412 13514 301464 13524
rect 301412 13480 301420 13514
rect 301420 13480 301454 13514
rect 301454 13480 301464 13514
rect 301412 13472 301464 13480
rect 216404 13446 216456 13456
rect 216404 13412 216412 13446
rect 216412 13412 216446 13446
rect 216446 13412 216456 13446
rect 216404 13404 216456 13412
rect 219440 13404 219492 13456
rect 207940 13268 207992 13320
rect 213552 13310 213604 13320
rect 213552 13276 213560 13310
rect 213560 13276 213594 13310
rect 213594 13276 213604 13310
rect 213552 13268 213604 13276
rect 216588 13310 216640 13320
rect 216588 13276 216596 13310
rect 216596 13276 216630 13310
rect 216630 13276 216640 13310
rect 224132 13404 224184 13456
rect 224040 13336 224092 13388
rect 226432 13404 226484 13456
rect 226616 13446 226668 13456
rect 226616 13412 226624 13446
rect 226624 13412 226658 13446
rect 226658 13412 226668 13446
rect 226616 13404 226668 13412
rect 226892 13404 226944 13456
rect 227904 13404 227956 13456
rect 229192 13404 229244 13456
rect 224408 13336 224460 13388
rect 227076 13378 227128 13388
rect 227076 13344 227084 13378
rect 227084 13344 227118 13378
rect 227118 13344 227128 13378
rect 227076 13336 227128 13344
rect 227168 13378 227220 13388
rect 227168 13344 227176 13378
rect 227176 13344 227210 13378
rect 227210 13344 227220 13378
rect 227168 13336 227220 13344
rect 216588 13268 216640 13276
rect 224224 13200 224276 13252
rect 207388 13132 207440 13184
rect 213552 13132 213604 13184
rect 222752 13174 222804 13184
rect 222752 13140 222760 13174
rect 222760 13140 222794 13174
rect 222794 13140 222804 13174
rect 222752 13132 222804 13140
rect 223672 13174 223724 13184
rect 223672 13140 223680 13174
rect 223680 13140 223714 13174
rect 223714 13140 223724 13174
rect 223672 13132 223724 13140
rect 224040 13174 224092 13184
rect 224040 13140 224048 13174
rect 224048 13140 224082 13174
rect 224082 13140 224092 13174
rect 224040 13132 224092 13140
rect 224132 13174 224184 13184
rect 224132 13140 224140 13174
rect 224140 13140 224174 13174
rect 224174 13140 224184 13174
rect 224408 13200 224460 13252
rect 227720 13268 227772 13320
rect 231952 13336 232004 13388
rect 230388 13268 230440 13320
rect 231860 13268 231912 13320
rect 232044 13268 232096 13320
rect 233148 13336 233200 13388
rect 233332 13336 233384 13388
rect 233056 13310 233108 13320
rect 233056 13276 233064 13310
rect 233064 13276 233098 13310
rect 233098 13276 233108 13310
rect 233056 13268 233108 13276
rect 228088 13200 228140 13252
rect 230756 13242 230808 13252
rect 230756 13208 230764 13242
rect 230764 13208 230798 13242
rect 230798 13208 230808 13242
rect 230756 13200 230808 13208
rect 237932 13336 237984 13388
rect 238116 13336 238168 13388
rect 239496 13404 239548 13456
rect 244648 13404 244700 13456
rect 245384 13404 245436 13456
rect 247132 13446 247184 13456
rect 247132 13412 247140 13446
rect 247140 13412 247174 13446
rect 247174 13412 247184 13446
rect 247132 13404 247184 13412
rect 251088 13404 251140 13456
rect 252468 13404 252520 13456
rect 254952 13404 255004 13456
rect 259460 13446 259512 13456
rect 259460 13412 259468 13446
rect 259468 13412 259502 13446
rect 259502 13412 259512 13446
rect 259460 13404 259512 13412
rect 263508 13404 263560 13456
rect 265532 13404 265584 13456
rect 270408 13404 270460 13456
rect 244096 13336 244148 13388
rect 238208 13310 238260 13320
rect 238208 13276 238216 13310
rect 238216 13276 238250 13310
rect 238250 13276 238260 13310
rect 238208 13268 238260 13276
rect 239772 13268 239824 13320
rect 250996 13336 251048 13388
rect 251088 13310 251140 13320
rect 251088 13276 251096 13310
rect 251096 13276 251130 13310
rect 251130 13276 251140 13310
rect 251088 13268 251140 13276
rect 224132 13132 224184 13140
rect 225420 13132 225472 13184
rect 225696 13174 225748 13184
rect 225696 13140 225704 13174
rect 225704 13140 225738 13174
rect 225738 13140 225748 13174
rect 225696 13132 225748 13140
rect 227076 13132 227128 13184
rect 227628 13132 227680 13184
rect 227904 13132 227956 13184
rect 232136 13132 232188 13184
rect 233240 13132 233292 13184
rect 234896 13174 234948 13184
rect 234896 13140 234904 13174
rect 234904 13140 234938 13174
rect 234938 13140 234948 13174
rect 234896 13132 234948 13140
rect 237012 13132 237064 13184
rect 238484 13242 238536 13252
rect 238484 13208 238492 13242
rect 238492 13208 238526 13242
rect 238526 13208 238536 13242
rect 241060 13242 241112 13252
rect 238484 13200 238536 13208
rect 241060 13208 241068 13242
rect 241068 13208 241102 13242
rect 241102 13208 241112 13242
rect 241060 13200 241112 13208
rect 241796 13200 241848 13252
rect 243636 13242 243688 13252
rect 242532 13174 242584 13184
rect 242532 13140 242540 13174
rect 242540 13140 242574 13174
rect 242574 13140 242584 13174
rect 242532 13132 242584 13140
rect 243636 13208 243644 13242
rect 243644 13208 243678 13242
rect 243678 13208 243688 13242
rect 243636 13200 243688 13208
rect 244924 13200 244976 13252
rect 251180 13132 251232 13184
rect 251364 13242 251416 13252
rect 251364 13208 251372 13242
rect 251372 13208 251406 13242
rect 251406 13208 251416 13242
rect 251364 13200 251416 13208
rect 252376 13200 252428 13252
rect 256240 13310 256292 13320
rect 253020 13200 253072 13252
rect 254952 13200 255004 13252
rect 253480 13132 253532 13184
rect 256240 13276 256248 13310
rect 256248 13276 256282 13310
rect 256282 13276 256292 13310
rect 256240 13268 256292 13276
rect 255320 13200 255372 13252
rect 256976 13200 257028 13252
rect 256332 13132 256384 13184
rect 264152 13336 264204 13388
rect 272984 13404 273036 13456
rect 268936 13268 268988 13320
rect 273168 13336 273220 13388
rect 273260 13268 273312 13320
rect 275100 13310 275152 13320
rect 275100 13276 275108 13310
rect 275108 13276 275142 13310
rect 275142 13276 275152 13310
rect 275100 13268 275152 13276
rect 261852 13242 261904 13252
rect 261852 13208 261860 13242
rect 261860 13208 261894 13242
rect 261894 13208 261904 13242
rect 261852 13200 261904 13208
rect 263416 13200 263468 13252
rect 263508 13200 263560 13252
rect 264428 13200 264480 13252
rect 264612 13200 264664 13252
rect 264980 13200 265032 13252
rect 257988 13174 258040 13184
rect 257988 13140 257996 13174
rect 257996 13140 258030 13174
rect 258030 13140 258040 13174
rect 257988 13132 258040 13140
rect 262956 13132 263008 13184
rect 263324 13132 263376 13184
rect 266912 13200 266964 13252
rect 267648 13132 267700 13184
rect 268752 13200 268804 13252
rect 270684 13200 270736 13252
rect 270776 13132 270828 13184
rect 270960 13200 271012 13252
rect 281080 13310 281132 13320
rect 281080 13276 281088 13310
rect 281088 13276 281122 13310
rect 281122 13276 281132 13310
rect 281080 13268 281132 13276
rect 284760 13310 284812 13320
rect 284760 13276 284768 13310
rect 284768 13276 284802 13310
rect 284802 13276 284812 13310
rect 284760 13268 284812 13276
rect 290280 13310 290332 13320
rect 290280 13276 290288 13310
rect 290288 13276 290322 13310
rect 290322 13276 290332 13310
rect 290280 13268 290332 13276
rect 305000 13336 305052 13388
rect 271788 13132 271840 13184
rect 272892 13132 272944 13184
rect 299480 13310 299532 13320
rect 299480 13276 299488 13310
rect 299488 13276 299522 13310
rect 299522 13276 299532 13310
rect 299480 13268 299532 13276
rect 303528 13268 303580 13320
rect 295892 13174 295944 13184
rect 295892 13140 295900 13174
rect 295900 13140 295934 13174
rect 295934 13140 295944 13174
rect 295892 13132 295944 13140
rect 77148 13030 77200 13082
rect 77212 13030 77264 13082
rect 77276 13030 77328 13082
rect 77340 13030 77392 13082
rect 77404 13030 77456 13082
rect 153346 13030 153398 13082
rect 153410 13030 153462 13082
rect 153474 13030 153526 13082
rect 153538 13030 153590 13082
rect 153602 13030 153654 13082
rect 229544 13030 229596 13082
rect 229608 13030 229660 13082
rect 229672 13030 229724 13082
rect 229736 13030 229788 13082
rect 229800 13030 229852 13082
rect 26056 12970 26108 12980
rect 26056 12936 26064 12970
rect 26064 12936 26098 12970
rect 26098 12936 26108 12970
rect 26056 12928 26108 12936
rect 20168 12860 20220 12912
rect 27344 12860 27396 12912
rect 32220 12928 32272 12980
rect 34152 12928 34204 12980
rect 35532 12970 35584 12980
rect 35532 12936 35540 12970
rect 35540 12936 35574 12970
rect 35574 12936 35584 12970
rect 35532 12928 35584 12936
rect 29000 12902 29052 12912
rect 23204 12724 23256 12776
rect 29000 12868 29008 12902
rect 29008 12868 29042 12902
rect 29042 12868 29052 12902
rect 29000 12860 29052 12868
rect 27988 12792 28040 12844
rect 28080 12766 28132 12776
rect 27160 12656 27212 12708
rect 28080 12732 28088 12766
rect 28088 12732 28122 12766
rect 28122 12732 28132 12766
rect 28080 12724 28132 12732
rect 30380 12860 30432 12912
rect 31576 12860 31628 12912
rect 34428 12860 34480 12912
rect 33692 12792 33744 12844
rect 37464 12860 37516 12912
rect 39672 12860 39724 12912
rect 41052 12860 41104 12912
rect 43260 12928 43312 12980
rect 44272 12928 44324 12980
rect 44548 12970 44600 12980
rect 44548 12936 44556 12970
rect 44556 12936 44590 12970
rect 44590 12936 44600 12970
rect 44548 12928 44600 12936
rect 53288 12928 53340 12980
rect 42984 12860 43036 12912
rect 54668 12928 54720 12980
rect 55864 12928 55916 12980
rect 57980 12928 58032 12980
rect 59636 12928 59688 12980
rect 72148 12970 72200 12980
rect 72148 12936 72156 12970
rect 72156 12936 72190 12970
rect 72190 12936 72200 12970
rect 72148 12928 72200 12936
rect 72332 12928 72384 12980
rect 74724 12928 74776 12980
rect 29644 12724 29696 12776
rect 29828 12766 29880 12776
rect 29828 12732 29836 12766
rect 29836 12732 29870 12766
rect 29870 12732 29880 12766
rect 29828 12724 29880 12732
rect 30104 12766 30156 12776
rect 30104 12732 30112 12766
rect 30112 12732 30146 12766
rect 30146 12732 30156 12766
rect 30104 12724 30156 12732
rect 28908 12588 28960 12640
rect 33048 12724 33100 12776
rect 33416 12724 33468 12776
rect 34336 12724 34388 12776
rect 39304 12792 39356 12844
rect 41512 12792 41564 12844
rect 34888 12766 34940 12776
rect 34888 12732 34896 12766
rect 34896 12732 34930 12766
rect 34930 12732 34940 12766
rect 34888 12724 34940 12732
rect 35348 12724 35400 12776
rect 39396 12724 39448 12776
rect 40960 12724 41012 12776
rect 43076 12724 43128 12776
rect 43168 12724 43220 12776
rect 45376 12792 45428 12844
rect 55496 12860 55548 12912
rect 57336 12860 57388 12912
rect 60648 12860 60700 12912
rect 65892 12860 65944 12912
rect 53748 12792 53800 12844
rect 54024 12834 54076 12844
rect 43812 12724 43864 12776
rect 45468 12724 45520 12776
rect 51356 12724 51408 12776
rect 54024 12800 54032 12834
rect 54032 12800 54066 12834
rect 54066 12800 54076 12834
rect 54024 12792 54076 12800
rect 54760 12834 54812 12844
rect 54116 12766 54168 12776
rect 54116 12732 54124 12766
rect 54124 12732 54158 12766
rect 54158 12732 54168 12766
rect 54116 12724 54168 12732
rect 54760 12800 54768 12834
rect 54768 12800 54802 12834
rect 54802 12800 54812 12834
rect 54760 12792 54812 12800
rect 57428 12792 57480 12844
rect 74816 12792 74868 12844
rect 75460 12792 75512 12844
rect 78404 12860 78456 12912
rect 79692 12792 79744 12844
rect 83924 12928 83976 12980
rect 80520 12860 80572 12912
rect 82912 12860 82964 12912
rect 86500 12928 86552 12980
rect 87144 12928 87196 12980
rect 90456 12928 90508 12980
rect 91652 12928 91704 12980
rect 98000 12928 98052 12980
rect 55036 12766 55088 12776
rect 55036 12732 55044 12766
rect 55044 12732 55078 12766
rect 55078 12732 55088 12766
rect 55036 12724 55088 12732
rect 78588 12724 78640 12776
rect 31392 12588 31444 12640
rect 32404 12588 32456 12640
rect 34152 12588 34204 12640
rect 38016 12630 38068 12640
rect 38016 12596 38024 12630
rect 38024 12596 38058 12630
rect 38058 12596 38068 12630
rect 38016 12588 38068 12596
rect 41236 12630 41288 12640
rect 41236 12596 41244 12630
rect 41244 12596 41278 12630
rect 41278 12596 41288 12630
rect 41236 12588 41288 12596
rect 41788 12630 41840 12640
rect 41788 12596 41796 12630
rect 41796 12596 41830 12630
rect 41830 12596 41840 12630
rect 41788 12588 41840 12596
rect 42800 12588 42852 12640
rect 43260 12588 43312 12640
rect 43812 12588 43864 12640
rect 53104 12588 53156 12640
rect 54116 12588 54168 12640
rect 55588 12588 55640 12640
rect 56324 12588 56376 12640
rect 56508 12630 56560 12640
rect 56508 12596 56516 12630
rect 56516 12596 56550 12630
rect 56550 12596 56560 12630
rect 56508 12588 56560 12596
rect 57244 12588 57296 12640
rect 72700 12588 72752 12640
rect 75000 12588 75052 12640
rect 75184 12588 75236 12640
rect 77852 12656 77904 12708
rect 78128 12656 78180 12708
rect 80796 12724 80848 12776
rect 77208 12588 77260 12640
rect 81440 12656 81492 12708
rect 81624 12588 81676 12640
rect 84844 12724 84896 12776
rect 85764 12630 85816 12640
rect 85764 12596 85772 12630
rect 85772 12596 85806 12630
rect 85806 12596 85816 12630
rect 85764 12588 85816 12596
rect 90548 12860 90600 12912
rect 90732 12860 90784 12912
rect 99472 12902 99524 12912
rect 99472 12868 99480 12902
rect 99480 12868 99514 12902
rect 99514 12868 99524 12902
rect 99472 12860 99524 12868
rect 99932 12860 99984 12912
rect 104624 12902 104676 12912
rect 104624 12868 104632 12902
rect 104632 12868 104666 12902
rect 104666 12868 104676 12902
rect 104624 12860 104676 12868
rect 104716 12902 104768 12912
rect 104716 12868 104724 12902
rect 104724 12868 104758 12902
rect 104758 12868 104768 12902
rect 104716 12860 104768 12868
rect 90180 12792 90232 12844
rect 90456 12834 90508 12844
rect 90456 12800 90464 12834
rect 90464 12800 90498 12834
rect 90498 12800 90508 12834
rect 90456 12792 90508 12800
rect 90640 12792 90692 12844
rect 86500 12766 86552 12776
rect 86500 12732 86508 12766
rect 86508 12732 86542 12766
rect 86542 12732 86552 12766
rect 86500 12724 86552 12732
rect 88248 12724 88300 12776
rect 89720 12724 89772 12776
rect 90088 12724 90140 12776
rect 105176 12792 105228 12844
rect 99196 12766 99248 12776
rect 99196 12732 99204 12766
rect 99204 12732 99238 12766
rect 99238 12732 99248 12766
rect 101404 12766 101456 12776
rect 99196 12724 99248 12732
rect 101404 12732 101412 12766
rect 101412 12732 101446 12766
rect 101446 12732 101456 12766
rect 101404 12724 101456 12732
rect 101680 12766 101732 12776
rect 101680 12732 101688 12766
rect 101688 12732 101722 12766
rect 101722 12732 101732 12766
rect 101680 12724 101732 12732
rect 87788 12588 87840 12640
rect 87972 12630 88024 12640
rect 87972 12596 87980 12630
rect 87980 12596 88014 12630
rect 88014 12596 88024 12630
rect 87972 12588 88024 12596
rect 88432 12588 88484 12640
rect 89904 12588 89956 12640
rect 99196 12588 99248 12640
rect 101036 12656 101088 12708
rect 103244 12656 103296 12708
rect 105912 12698 105964 12708
rect 105912 12664 105920 12698
rect 105920 12664 105954 12698
rect 105954 12664 105964 12698
rect 105912 12656 105964 12664
rect 111432 12928 111484 12980
rect 114560 12928 114612 12980
rect 114744 12928 114796 12980
rect 117412 12928 117464 12980
rect 118240 12970 118292 12980
rect 118240 12936 118248 12970
rect 118248 12936 118282 12970
rect 118282 12936 118292 12970
rect 118240 12928 118292 12936
rect 118700 12970 118752 12980
rect 118700 12936 118708 12970
rect 118708 12936 118742 12970
rect 118742 12936 118752 12970
rect 118700 12928 118752 12936
rect 126888 12928 126940 12980
rect 128084 12970 128136 12980
rect 128084 12936 128092 12970
rect 128092 12936 128126 12970
rect 128126 12936 128136 12970
rect 128084 12928 128136 12936
rect 128636 12928 128688 12980
rect 129188 12970 129240 12980
rect 129188 12936 129196 12970
rect 129196 12936 129230 12970
rect 129230 12936 129240 12970
rect 129188 12928 129240 12936
rect 133328 12928 133380 12980
rect 109592 12860 109644 12912
rect 113088 12834 113140 12844
rect 113088 12800 113096 12834
rect 113096 12800 113130 12834
rect 113130 12800 113140 12834
rect 113088 12792 113140 12800
rect 113824 12834 113876 12844
rect 113824 12800 113832 12834
rect 113832 12800 113866 12834
rect 113866 12800 113876 12834
rect 113824 12792 113876 12800
rect 114652 12834 114704 12844
rect 114652 12800 114660 12834
rect 114660 12800 114694 12834
rect 114694 12800 114704 12834
rect 115756 12860 115808 12912
rect 117320 12860 117372 12912
rect 126520 12860 126572 12912
rect 114652 12792 114704 12800
rect 118056 12792 118108 12844
rect 132408 12860 132460 12912
rect 133604 12902 133656 12912
rect 133604 12868 133612 12902
rect 133612 12868 133646 12902
rect 133646 12868 133656 12902
rect 133604 12860 133656 12868
rect 133880 12928 133932 12980
rect 147680 12928 147732 12980
rect 134156 12860 134208 12912
rect 143080 12860 143132 12912
rect 145932 12902 145984 12912
rect 127440 12834 127492 12844
rect 127440 12800 127448 12834
rect 127448 12800 127482 12834
rect 127482 12800 127492 12834
rect 127440 12792 127492 12800
rect 113916 12724 113968 12776
rect 114744 12724 114796 12776
rect 115664 12724 115716 12776
rect 115848 12766 115900 12776
rect 115848 12732 115856 12766
rect 115856 12732 115890 12766
rect 115890 12732 115900 12766
rect 115848 12724 115900 12732
rect 116768 12766 116820 12776
rect 114836 12656 114888 12708
rect 116768 12732 116776 12766
rect 116776 12732 116810 12766
rect 116810 12732 116820 12766
rect 116768 12724 116820 12732
rect 100760 12588 100812 12640
rect 103060 12588 103112 12640
rect 103612 12588 103664 12640
rect 111892 12630 111944 12640
rect 111892 12596 111900 12630
rect 111900 12596 111934 12630
rect 111934 12596 111944 12630
rect 111892 12588 111944 12596
rect 113088 12588 113140 12640
rect 114744 12630 114796 12640
rect 114744 12596 114752 12630
rect 114752 12596 114786 12630
rect 114786 12596 114796 12630
rect 114744 12588 114796 12596
rect 115848 12588 115900 12640
rect 127532 12724 127584 12776
rect 128084 12588 128136 12640
rect 129096 12834 129148 12844
rect 129096 12800 129104 12834
rect 129104 12800 129138 12834
rect 129138 12800 129148 12834
rect 129096 12792 129148 12800
rect 128360 12724 128412 12776
rect 130292 12792 130344 12844
rect 129740 12724 129792 12776
rect 131120 12766 131172 12776
rect 131120 12732 131128 12766
rect 131128 12732 131162 12766
rect 131162 12732 131172 12766
rect 131120 12724 131172 12732
rect 132592 12766 132644 12776
rect 132592 12732 132600 12766
rect 132600 12732 132634 12766
rect 132634 12732 132644 12766
rect 133696 12792 133748 12844
rect 145932 12868 145940 12902
rect 145940 12868 145974 12902
rect 145974 12868 145984 12902
rect 145932 12860 145984 12868
rect 152648 12928 152700 12980
rect 152832 12928 152884 12980
rect 157156 12970 157208 12980
rect 157156 12936 157164 12970
rect 157164 12936 157198 12970
rect 157198 12936 157208 12970
rect 157156 12928 157208 12936
rect 158628 12928 158680 12980
rect 145840 12834 145892 12844
rect 132592 12724 132644 12732
rect 143264 12766 143316 12776
rect 130292 12656 130344 12708
rect 133696 12656 133748 12708
rect 133144 12630 133196 12640
rect 133144 12596 133152 12630
rect 133152 12596 133186 12630
rect 133186 12596 133196 12630
rect 133144 12588 133196 12596
rect 133236 12588 133288 12640
rect 143264 12732 143272 12766
rect 143272 12732 143306 12766
rect 143306 12732 143316 12766
rect 143264 12724 143316 12732
rect 145840 12800 145848 12834
rect 145848 12800 145882 12834
rect 145882 12800 145892 12834
rect 145840 12792 145892 12800
rect 156604 12860 156656 12912
rect 147312 12792 147364 12844
rect 149336 12792 149388 12844
rect 147404 12724 147456 12776
rect 147772 12766 147824 12776
rect 133880 12656 133932 12708
rect 145748 12656 145800 12708
rect 147772 12732 147780 12766
rect 147780 12732 147814 12766
rect 147814 12732 147824 12766
rect 147772 12724 147824 12732
rect 148968 12724 149020 12776
rect 149244 12766 149296 12776
rect 149244 12732 149252 12766
rect 149252 12732 149286 12766
rect 149286 12732 149296 12766
rect 149244 12724 149296 12732
rect 150440 12792 150492 12844
rect 155868 12792 155920 12844
rect 157800 12792 157852 12844
rect 160376 12860 160428 12912
rect 161664 12792 161716 12844
rect 151544 12766 151596 12776
rect 151544 12732 151552 12766
rect 151552 12732 151586 12766
rect 151586 12732 151596 12766
rect 151544 12724 151596 12732
rect 150348 12656 150400 12708
rect 151636 12656 151688 12708
rect 148508 12588 148560 12640
rect 149980 12630 150032 12640
rect 149980 12596 149988 12630
rect 149988 12596 150022 12630
rect 150022 12596 150032 12630
rect 149980 12588 150032 12596
rect 151268 12588 151320 12640
rect 151360 12588 151412 12640
rect 152740 12724 152792 12776
rect 152832 12656 152884 12708
rect 153108 12656 153160 12708
rect 155040 12766 155092 12776
rect 155040 12732 155048 12766
rect 155048 12732 155082 12766
rect 155082 12732 155092 12766
rect 159456 12766 159508 12776
rect 155040 12724 155092 12732
rect 158812 12698 158864 12708
rect 158812 12664 158820 12698
rect 158820 12664 158854 12698
rect 158854 12664 158864 12698
rect 158812 12656 158864 12664
rect 159456 12732 159464 12766
rect 159464 12732 159498 12766
rect 159498 12732 159508 12766
rect 159456 12724 159508 12732
rect 159548 12724 159600 12776
rect 161572 12724 161624 12776
rect 154120 12588 154172 12640
rect 157892 12588 157944 12640
rect 160284 12588 160336 12640
rect 163504 12928 163556 12980
rect 163412 12860 163464 12912
rect 165252 12928 165304 12980
rect 162124 12766 162176 12776
rect 162124 12732 162132 12766
rect 162132 12732 162166 12766
rect 162166 12732 162176 12766
rect 162124 12724 162176 12732
rect 162860 12724 162912 12776
rect 167184 12928 167236 12980
rect 175004 12970 175056 12980
rect 175004 12936 175012 12970
rect 175012 12936 175046 12970
rect 175046 12936 175056 12970
rect 175004 12928 175056 12936
rect 175740 12928 175792 12980
rect 176384 12928 176436 12980
rect 165436 12792 165488 12844
rect 166172 12792 166224 12844
rect 166540 12834 166592 12844
rect 166540 12800 166548 12834
rect 166548 12800 166582 12834
rect 166582 12800 166592 12834
rect 166540 12792 166592 12800
rect 173808 12860 173860 12912
rect 175924 12860 175976 12912
rect 176936 12860 176988 12912
rect 177948 12860 178000 12912
rect 176384 12834 176436 12844
rect 164608 12766 164660 12776
rect 164608 12732 164616 12766
rect 164616 12732 164650 12766
rect 164650 12732 164660 12766
rect 164608 12724 164660 12732
rect 163688 12588 163740 12640
rect 164240 12656 164292 12708
rect 176384 12800 176392 12834
rect 176392 12800 176426 12834
rect 176426 12800 176436 12834
rect 176384 12792 176436 12800
rect 180156 12928 180208 12980
rect 180248 12928 180300 12980
rect 180340 12792 180392 12844
rect 181536 12834 181588 12844
rect 181536 12800 181544 12834
rect 181544 12800 181578 12834
rect 181578 12800 181588 12834
rect 188344 12928 188396 12980
rect 191380 12928 191432 12980
rect 192484 12928 192536 12980
rect 188528 12860 188580 12912
rect 190920 12902 190972 12912
rect 181536 12792 181588 12800
rect 188344 12792 188396 12844
rect 188804 12792 188856 12844
rect 189356 12834 189408 12844
rect 189356 12800 189364 12834
rect 189364 12800 189398 12834
rect 189398 12800 189408 12834
rect 189356 12792 189408 12800
rect 176752 12724 176804 12776
rect 180156 12724 180208 12776
rect 189540 12724 189592 12776
rect 190920 12868 190928 12902
rect 190928 12868 190962 12902
rect 190962 12868 190972 12902
rect 190920 12860 190972 12868
rect 191748 12860 191800 12912
rect 193956 12928 194008 12980
rect 194876 12928 194928 12980
rect 195980 12970 196032 12980
rect 195980 12936 195988 12970
rect 195988 12936 196022 12970
rect 196022 12936 196032 12970
rect 195980 12928 196032 12936
rect 197728 12928 197780 12980
rect 192576 12792 192628 12844
rect 195060 12834 195112 12844
rect 195060 12800 195068 12834
rect 195068 12800 195102 12834
rect 195102 12800 195112 12834
rect 195060 12792 195112 12800
rect 197360 12834 197412 12844
rect 197360 12800 197368 12834
rect 197368 12800 197402 12834
rect 197402 12800 197412 12834
rect 197360 12792 197412 12800
rect 197452 12834 197504 12844
rect 197452 12800 197460 12834
rect 197460 12800 197494 12834
rect 197494 12800 197504 12834
rect 198372 12834 198424 12844
rect 197452 12792 197504 12800
rect 192668 12724 192720 12776
rect 193036 12766 193088 12776
rect 193036 12732 193044 12766
rect 193044 12732 193078 12766
rect 193078 12732 193088 12766
rect 193036 12724 193088 12732
rect 166172 12588 166224 12640
rect 166632 12630 166684 12640
rect 166632 12596 166640 12630
rect 166640 12596 166674 12630
rect 166674 12596 166684 12630
rect 166632 12588 166684 12596
rect 180248 12656 180300 12708
rect 180524 12656 180576 12708
rect 182088 12656 182140 12708
rect 188620 12656 188672 12708
rect 189172 12656 189224 12708
rect 191748 12656 191800 12708
rect 191932 12656 191984 12708
rect 192484 12656 192536 12708
rect 194784 12724 194836 12776
rect 195796 12724 195848 12776
rect 197636 12766 197688 12776
rect 197636 12732 197644 12766
rect 197644 12732 197678 12766
rect 197678 12732 197688 12766
rect 197636 12724 197688 12732
rect 198372 12800 198380 12834
rect 198380 12800 198414 12834
rect 198414 12800 198424 12834
rect 198372 12792 198424 12800
rect 200672 12792 200724 12844
rect 201316 12834 201368 12844
rect 201316 12800 201324 12834
rect 201324 12800 201358 12834
rect 201358 12800 201368 12834
rect 201316 12792 201368 12800
rect 198556 12724 198608 12776
rect 200396 12724 200448 12776
rect 202972 12860 203024 12912
rect 203340 12860 203392 12912
rect 205640 12860 205692 12912
rect 206560 12970 206612 12980
rect 206560 12936 206568 12970
rect 206568 12936 206602 12970
rect 206602 12936 206612 12970
rect 206560 12928 206612 12936
rect 207388 12928 207440 12980
rect 207848 12928 207900 12980
rect 202880 12766 202932 12776
rect 177396 12588 177448 12640
rect 177856 12588 177908 12640
rect 179880 12588 179932 12640
rect 180616 12588 180668 12640
rect 181444 12588 181496 12640
rect 187792 12588 187844 12640
rect 188988 12588 189040 12640
rect 190552 12630 190604 12640
rect 190552 12596 190560 12630
rect 190560 12596 190594 12630
rect 190594 12596 190604 12630
rect 190552 12588 190604 12596
rect 192024 12588 192076 12640
rect 192116 12588 192168 12640
rect 193036 12588 193088 12640
rect 202144 12656 202196 12708
rect 202880 12732 202888 12766
rect 202888 12732 202922 12766
rect 202922 12732 202932 12766
rect 202880 12724 202932 12732
rect 202972 12724 203024 12776
rect 204168 12724 204220 12776
rect 205088 12766 205140 12776
rect 205088 12732 205096 12766
rect 205096 12732 205130 12766
rect 205130 12732 205140 12766
rect 205088 12724 205140 12732
rect 205180 12724 205232 12776
rect 210608 12860 210660 12912
rect 219808 12928 219860 12980
rect 207664 12792 207716 12844
rect 216588 12792 216640 12844
rect 228272 12860 228324 12912
rect 230388 12860 230440 12912
rect 219808 12792 219860 12844
rect 223672 12792 223724 12844
rect 226800 12792 226852 12844
rect 227904 12834 227956 12844
rect 227904 12800 227912 12834
rect 227912 12800 227946 12834
rect 227946 12800 227956 12834
rect 227904 12792 227956 12800
rect 230296 12834 230348 12844
rect 230296 12800 230304 12834
rect 230304 12800 230338 12834
rect 230338 12800 230348 12834
rect 230296 12792 230348 12800
rect 238208 12928 238260 12980
rect 231032 12902 231084 12912
rect 231032 12868 231040 12902
rect 231040 12868 231074 12902
rect 231074 12868 231084 12902
rect 231032 12860 231084 12868
rect 232320 12860 232372 12912
rect 238300 12860 238352 12912
rect 233056 12834 233108 12844
rect 207296 12698 207348 12708
rect 194416 12588 194468 12640
rect 195980 12588 196032 12640
rect 198188 12630 198240 12640
rect 198188 12596 198196 12630
rect 198196 12596 198230 12630
rect 198230 12596 198240 12630
rect 198188 12588 198240 12596
rect 201132 12630 201184 12640
rect 201132 12596 201140 12630
rect 201140 12596 201174 12630
rect 201174 12596 201184 12630
rect 201132 12588 201184 12596
rect 201960 12588 202012 12640
rect 204260 12588 204312 12640
rect 204536 12588 204588 12640
rect 205180 12588 205232 12640
rect 205272 12588 205324 12640
rect 207296 12664 207304 12698
rect 207304 12664 207338 12698
rect 207338 12664 207348 12698
rect 207296 12656 207348 12664
rect 210608 12588 210660 12640
rect 219808 12656 219860 12708
rect 226892 12588 226944 12640
rect 228272 12724 228324 12776
rect 230204 12724 230256 12776
rect 233056 12800 233064 12834
rect 233064 12800 233098 12834
rect 233098 12800 233108 12834
rect 233056 12792 233108 12800
rect 237012 12834 237064 12844
rect 237012 12800 237020 12834
rect 237020 12800 237054 12834
rect 237054 12800 237064 12834
rect 237012 12792 237064 12800
rect 238392 12792 238444 12844
rect 239036 12860 239088 12912
rect 240048 12860 240100 12912
rect 251088 12928 251140 12980
rect 254676 12928 254728 12980
rect 256240 12928 256292 12980
rect 264612 12970 264664 12980
rect 240968 12902 241020 12912
rect 240968 12868 240976 12902
rect 240976 12868 241010 12902
rect 241010 12868 241020 12902
rect 240968 12860 241020 12868
rect 242072 12792 242124 12844
rect 242256 12792 242308 12844
rect 244648 12860 244700 12912
rect 244924 12860 244976 12912
rect 245384 12860 245436 12912
rect 251640 12860 251692 12912
rect 252468 12902 252520 12912
rect 252468 12868 252476 12902
rect 252476 12868 252510 12902
rect 252510 12868 252520 12902
rect 252468 12860 252520 12868
rect 244556 12834 244608 12844
rect 244556 12800 244564 12834
rect 244564 12800 244598 12834
rect 244598 12800 244608 12834
rect 244556 12792 244608 12800
rect 244832 12792 244884 12844
rect 251180 12792 251232 12844
rect 251548 12834 251600 12844
rect 251548 12800 251556 12834
rect 251556 12800 251590 12834
rect 251590 12800 251600 12834
rect 251548 12792 251600 12800
rect 256608 12792 256660 12844
rect 237840 12656 237892 12708
rect 237932 12656 237984 12708
rect 229560 12588 229612 12640
rect 230112 12630 230164 12640
rect 230112 12596 230120 12630
rect 230120 12596 230154 12630
rect 230154 12596 230164 12630
rect 230112 12588 230164 12596
rect 230204 12588 230256 12640
rect 232320 12588 232372 12640
rect 232504 12630 232556 12640
rect 232504 12596 232512 12630
rect 232512 12596 232546 12630
rect 232546 12596 232556 12630
rect 232504 12588 232556 12596
rect 233148 12588 233200 12640
rect 238484 12588 238536 12640
rect 238852 12588 238904 12640
rect 239128 12588 239180 12640
rect 240324 12588 240376 12640
rect 242164 12656 242216 12708
rect 242440 12630 242492 12640
rect 242440 12596 242448 12630
rect 242448 12596 242482 12630
rect 242482 12596 242492 12630
rect 242440 12588 242492 12596
rect 242900 12588 242952 12640
rect 244648 12656 244700 12708
rect 248328 12656 248380 12708
rect 250168 12698 250220 12708
rect 250168 12664 250176 12698
rect 250176 12664 250210 12698
rect 250210 12664 250220 12698
rect 250168 12656 250220 12664
rect 252100 12724 252152 12776
rect 253664 12766 253716 12776
rect 253664 12732 253672 12766
rect 253672 12732 253706 12766
rect 253706 12732 253716 12766
rect 253664 12724 253716 12732
rect 253940 12766 253992 12776
rect 253940 12732 253948 12766
rect 253948 12732 253982 12766
rect 253982 12732 253992 12766
rect 253940 12724 253992 12732
rect 255136 12724 255188 12776
rect 256332 12766 256384 12776
rect 256332 12732 256340 12766
rect 256340 12732 256374 12766
rect 256374 12732 256384 12766
rect 256332 12724 256384 12732
rect 256424 12766 256476 12776
rect 256424 12732 256432 12766
rect 256432 12732 256466 12766
rect 256466 12732 256476 12766
rect 256424 12724 256476 12732
rect 251824 12656 251876 12708
rect 255044 12656 255096 12708
rect 251916 12588 251968 12640
rect 252008 12630 252060 12640
rect 252008 12596 252016 12630
rect 252016 12596 252050 12630
rect 252050 12596 252060 12630
rect 257252 12860 257304 12912
rect 261760 12902 261812 12912
rect 261760 12868 261768 12902
rect 261768 12868 261802 12902
rect 261802 12868 261812 12902
rect 261760 12860 261812 12868
rect 263324 12860 263376 12912
rect 264612 12936 264620 12970
rect 264620 12936 264654 12970
rect 264654 12936 264664 12970
rect 264612 12928 264664 12936
rect 268384 12928 268436 12980
rect 302608 12970 302660 12980
rect 265532 12902 265584 12912
rect 261852 12792 261904 12844
rect 264336 12792 264388 12844
rect 264428 12792 264480 12844
rect 265532 12868 265540 12902
rect 265540 12868 265574 12902
rect 265574 12868 265584 12902
rect 265532 12860 265584 12868
rect 266544 12860 266596 12912
rect 257160 12724 257212 12776
rect 262312 12724 262364 12776
rect 271052 12860 271104 12912
rect 271788 12902 271840 12912
rect 271788 12868 271796 12902
rect 271796 12868 271830 12902
rect 271830 12868 271840 12902
rect 271788 12860 271840 12868
rect 272800 12860 272852 12912
rect 273168 12860 273220 12912
rect 268292 12792 268344 12844
rect 269028 12792 269080 12844
rect 257068 12656 257120 12708
rect 262680 12698 262732 12708
rect 252008 12588 252060 12596
rect 262220 12588 262272 12640
rect 262680 12664 262688 12698
rect 262688 12664 262722 12698
rect 262722 12664 262732 12698
rect 262680 12656 262732 12664
rect 267004 12724 267056 12776
rect 267556 12724 267608 12776
rect 268016 12766 268068 12776
rect 268016 12732 268024 12766
rect 268024 12732 268058 12766
rect 268058 12732 268068 12766
rect 268016 12724 268068 12732
rect 268384 12724 268436 12776
rect 270868 12792 270920 12844
rect 272616 12792 272668 12844
rect 295892 12860 295944 12912
rect 302608 12936 302616 12970
rect 302616 12936 302650 12970
rect 302650 12936 302660 12970
rect 302608 12928 302660 12936
rect 305368 12928 305420 12980
rect 305000 12902 305052 12912
rect 269396 12766 269448 12776
rect 269396 12732 269404 12766
rect 269404 12732 269438 12766
rect 269438 12732 269448 12766
rect 269396 12724 269448 12732
rect 263508 12656 263560 12708
rect 263968 12630 264020 12640
rect 263968 12596 263976 12630
rect 263976 12596 264010 12630
rect 264010 12596 264020 12630
rect 263968 12588 264020 12596
rect 267004 12630 267056 12640
rect 267004 12596 267012 12630
rect 267012 12596 267046 12630
rect 267046 12596 267056 12630
rect 267004 12588 267056 12596
rect 267096 12588 267148 12640
rect 267556 12588 267608 12640
rect 269120 12588 269172 12640
rect 272248 12724 272300 12776
rect 272892 12724 272944 12776
rect 272800 12656 272852 12708
rect 273168 12724 273220 12776
rect 290280 12792 290332 12844
rect 302792 12834 302844 12844
rect 302792 12800 302800 12834
rect 302800 12800 302834 12834
rect 302834 12800 302844 12834
rect 302792 12792 302844 12800
rect 305000 12868 305008 12902
rect 305008 12868 305042 12902
rect 305042 12868 305052 12902
rect 305460 12902 305512 12912
rect 305000 12860 305052 12868
rect 305460 12868 305468 12902
rect 305468 12868 305502 12902
rect 305502 12868 305512 12902
rect 305460 12860 305512 12868
rect 270868 12630 270920 12640
rect 270868 12596 270876 12630
rect 270876 12596 270910 12630
rect 270910 12596 270920 12630
rect 270868 12588 270920 12596
rect 271144 12588 271196 12640
rect 272524 12630 272576 12640
rect 272524 12596 272532 12630
rect 272532 12596 272566 12630
rect 272566 12596 272576 12630
rect 272524 12588 272576 12596
rect 272616 12588 272668 12640
rect 281080 12588 281132 12640
rect 39048 12486 39100 12538
rect 39112 12486 39164 12538
rect 39176 12486 39228 12538
rect 39240 12486 39292 12538
rect 39304 12486 39356 12538
rect 115246 12486 115298 12538
rect 115310 12486 115362 12538
rect 115374 12486 115426 12538
rect 115438 12486 115490 12538
rect 115502 12486 115554 12538
rect 191444 12486 191496 12538
rect 191508 12486 191560 12538
rect 191572 12486 191624 12538
rect 191636 12486 191688 12538
rect 191700 12486 191752 12538
rect 267642 12486 267694 12538
rect 267706 12486 267758 12538
rect 267770 12486 267822 12538
rect 267834 12486 267886 12538
rect 267898 12486 267950 12538
rect 26976 12384 27028 12436
rect 28080 12384 28132 12436
rect 14280 12316 14332 12368
rect 28816 12384 28868 12436
rect 32588 12384 32640 12436
rect 34520 12384 34572 12436
rect 35992 12384 36044 12436
rect 4804 12044 4856 12096
rect 26884 12248 26936 12300
rect 28080 12248 28132 12300
rect 28724 12290 28776 12300
rect 28724 12256 28732 12290
rect 28732 12256 28766 12290
rect 28766 12256 28776 12290
rect 28724 12248 28776 12256
rect 34888 12316 34940 12368
rect 37832 12384 37884 12436
rect 38936 12384 38988 12436
rect 39396 12384 39448 12436
rect 40960 12384 41012 12436
rect 43168 12426 43220 12436
rect 43168 12392 43176 12426
rect 43176 12392 43210 12426
rect 43210 12392 43220 12426
rect 43168 12384 43220 12392
rect 43812 12426 43864 12436
rect 43812 12392 43820 12426
rect 43820 12392 43854 12426
rect 43854 12392 43864 12426
rect 43812 12384 43864 12392
rect 54024 12384 54076 12436
rect 55496 12384 55548 12436
rect 56692 12384 56744 12436
rect 57980 12426 58032 12436
rect 57980 12392 57988 12426
rect 57988 12392 58022 12426
rect 58022 12392 58032 12426
rect 57980 12384 58032 12392
rect 75092 12384 75144 12436
rect 79324 12426 79376 12436
rect 29000 12248 29052 12300
rect 29552 12290 29604 12300
rect 29552 12256 29560 12290
rect 29560 12256 29594 12290
rect 29594 12256 29604 12290
rect 29552 12248 29604 12256
rect 17040 12180 17092 12232
rect 27436 12222 27488 12232
rect 27436 12188 27444 12222
rect 27444 12188 27478 12222
rect 27478 12188 27488 12222
rect 27436 12180 27488 12188
rect 29368 12180 29420 12232
rect 34152 12222 34204 12232
rect 34152 12188 34160 12222
rect 34160 12188 34194 12222
rect 34194 12188 34204 12222
rect 34152 12180 34204 12188
rect 34704 12222 34756 12232
rect 34704 12188 34712 12222
rect 34712 12188 34746 12222
rect 34746 12188 34756 12222
rect 35348 12222 35400 12232
rect 34704 12180 34756 12188
rect 35348 12188 35356 12222
rect 35356 12188 35390 12222
rect 35390 12188 35400 12222
rect 35348 12180 35400 12188
rect 27068 12086 27120 12096
rect 27068 12052 27076 12086
rect 27076 12052 27110 12086
rect 27110 12052 27120 12086
rect 27068 12044 27120 12052
rect 27160 12044 27212 12096
rect 27988 12044 28040 12096
rect 29460 12112 29512 12164
rect 29828 12154 29880 12164
rect 29828 12120 29836 12154
rect 29836 12120 29870 12154
rect 29870 12120 29880 12154
rect 29828 12112 29880 12120
rect 31208 12112 31260 12164
rect 32036 12154 32088 12164
rect 32036 12120 32044 12154
rect 32044 12120 32078 12154
rect 32078 12120 32088 12154
rect 32036 12112 32088 12120
rect 43720 12316 43772 12368
rect 40960 12248 41012 12300
rect 38016 12180 38068 12232
rect 40316 12180 40368 12232
rect 40592 12222 40644 12232
rect 40592 12188 40600 12222
rect 40600 12188 40634 12222
rect 40634 12188 40644 12222
rect 40592 12180 40644 12188
rect 76012 12316 76064 12368
rect 53840 12248 53892 12300
rect 43720 12222 43772 12232
rect 43720 12188 43728 12222
rect 43728 12188 43762 12222
rect 43762 12188 43772 12222
rect 43720 12180 43772 12188
rect 41604 12112 41656 12164
rect 41788 12112 41840 12164
rect 28908 12044 28960 12096
rect 31116 12044 31168 12096
rect 32312 12044 32364 12096
rect 32956 12044 33008 12096
rect 36452 12086 36504 12096
rect 36452 12052 36460 12086
rect 36460 12052 36494 12086
rect 36494 12052 36504 12086
rect 36452 12044 36504 12052
rect 40500 12044 40552 12096
rect 40684 12086 40736 12096
rect 40684 12052 40692 12086
rect 40692 12052 40726 12086
rect 40726 12052 40736 12086
rect 40684 12044 40736 12052
rect 56416 12248 56468 12300
rect 74816 12248 74868 12300
rect 77208 12316 77260 12368
rect 78404 12316 78456 12368
rect 55312 12180 55364 12232
rect 56508 12180 56560 12232
rect 76932 12290 76984 12300
rect 76932 12256 76940 12290
rect 76940 12256 76974 12290
rect 76974 12256 76984 12290
rect 78128 12290 78180 12300
rect 76932 12248 76984 12256
rect 78128 12256 78136 12290
rect 78136 12256 78170 12290
rect 78170 12256 78180 12290
rect 78128 12248 78180 12256
rect 52644 12154 52696 12164
rect 52644 12120 52652 12154
rect 52652 12120 52686 12154
rect 52686 12120 52696 12154
rect 52644 12112 52696 12120
rect 53104 12112 53156 12164
rect 77944 12222 77996 12232
rect 77944 12188 77952 12222
rect 77952 12188 77986 12222
rect 77986 12188 77996 12222
rect 77944 12180 77996 12188
rect 79324 12392 79332 12426
rect 79332 12392 79366 12426
rect 79366 12392 79376 12426
rect 79324 12384 79376 12392
rect 80520 12384 80572 12436
rect 85488 12384 85540 12436
rect 86408 12426 86460 12436
rect 86408 12392 86416 12426
rect 86416 12392 86450 12426
rect 86450 12392 86460 12426
rect 86408 12384 86460 12392
rect 87880 12384 87932 12436
rect 90180 12426 90232 12436
rect 90180 12392 90188 12426
rect 90188 12392 90222 12426
rect 90222 12392 90232 12426
rect 90180 12384 90232 12392
rect 99472 12384 99524 12436
rect 99932 12384 99984 12436
rect 104992 12384 105044 12436
rect 105176 12426 105228 12436
rect 105176 12392 105184 12426
rect 105184 12392 105218 12426
rect 105218 12392 105228 12426
rect 105176 12384 105228 12392
rect 112536 12384 112588 12436
rect 115020 12384 115072 12436
rect 116952 12384 117004 12436
rect 127808 12384 127860 12436
rect 129096 12384 129148 12436
rect 130936 12384 130988 12436
rect 132408 12384 132460 12436
rect 147772 12384 147824 12436
rect 152464 12384 152516 12436
rect 78588 12180 78640 12232
rect 86132 12316 86184 12368
rect 87420 12316 87472 12368
rect 81440 12248 81492 12300
rect 84660 12290 84712 12300
rect 84660 12256 84668 12290
rect 84668 12256 84702 12290
rect 84702 12256 84712 12290
rect 84660 12248 84712 12256
rect 83832 12180 83884 12232
rect 85764 12248 85816 12300
rect 86316 12248 86368 12300
rect 88156 12290 88208 12300
rect 88156 12256 88164 12290
rect 88164 12256 88198 12290
rect 88198 12256 88208 12290
rect 88156 12248 88208 12256
rect 85488 12222 85540 12232
rect 85488 12188 85496 12222
rect 85496 12188 85530 12222
rect 85530 12188 85540 12222
rect 85488 12180 85540 12188
rect 86040 12180 86092 12232
rect 88248 12180 88300 12232
rect 89168 12248 89220 12300
rect 88984 12180 89036 12232
rect 92020 12180 92072 12232
rect 99104 12248 99156 12300
rect 102048 12248 102100 12300
rect 103244 12248 103296 12300
rect 103336 12248 103388 12300
rect 115756 12316 115808 12368
rect 97540 12180 97592 12232
rect 103704 12180 103756 12232
rect 100760 12154 100812 12164
rect 55864 12044 55916 12096
rect 56048 12086 56100 12096
rect 56048 12052 56056 12086
rect 56056 12052 56090 12086
rect 56090 12052 56100 12086
rect 56048 12044 56100 12052
rect 57336 12044 57388 12096
rect 76288 12086 76340 12096
rect 76288 12052 76296 12086
rect 76296 12052 76330 12086
rect 76330 12052 76340 12086
rect 76288 12044 76340 12052
rect 80244 12044 80296 12096
rect 84016 12086 84068 12096
rect 84016 12052 84024 12086
rect 84024 12052 84058 12086
rect 84058 12052 84068 12086
rect 84016 12044 84068 12052
rect 84660 12044 84712 12096
rect 86316 12044 86368 12096
rect 87512 12044 87564 12096
rect 87788 12044 87840 12096
rect 87972 12044 88024 12096
rect 88708 12044 88760 12096
rect 100760 12120 100768 12154
rect 100768 12120 100802 12154
rect 100802 12120 100812 12154
rect 100760 12112 100812 12120
rect 101036 12112 101088 12164
rect 101956 12154 102008 12164
rect 101956 12120 101964 12154
rect 101964 12120 101998 12154
rect 101998 12120 102008 12154
rect 101956 12112 102008 12120
rect 102140 12154 102192 12164
rect 102140 12120 102148 12154
rect 102148 12120 102182 12154
rect 102182 12120 102192 12154
rect 111892 12180 111944 12232
rect 114284 12180 114336 12232
rect 118884 12248 118936 12300
rect 141976 12316 142028 12368
rect 147588 12316 147640 12368
rect 151636 12316 151688 12368
rect 102140 12112 102192 12120
rect 113824 12112 113876 12164
rect 100392 12086 100444 12096
rect 100392 12052 100400 12086
rect 100400 12052 100434 12086
rect 100434 12052 100444 12086
rect 100392 12044 100444 12052
rect 102324 12044 102376 12096
rect 102600 12086 102652 12096
rect 102600 12052 102608 12086
rect 102608 12052 102642 12086
rect 102642 12052 102652 12086
rect 102600 12044 102652 12052
rect 103060 12086 103112 12096
rect 103060 12052 103068 12086
rect 103068 12052 103102 12086
rect 103102 12052 103112 12086
rect 103060 12044 103112 12052
rect 113916 12044 113968 12096
rect 115664 12044 115716 12096
rect 116400 12044 116452 12096
rect 118056 12180 118108 12232
rect 118332 12222 118384 12232
rect 118332 12188 118340 12222
rect 118340 12188 118374 12222
rect 118374 12188 118384 12222
rect 118332 12180 118384 12188
rect 126152 12180 126204 12232
rect 128636 12222 128688 12232
rect 128636 12188 128644 12222
rect 128644 12188 128678 12222
rect 128678 12188 128688 12222
rect 128636 12180 128688 12188
rect 131028 12248 131080 12300
rect 133236 12248 133288 12300
rect 149060 12248 149112 12300
rect 118240 12112 118292 12164
rect 130476 12180 130528 12232
rect 132408 12180 132460 12232
rect 132592 12222 132644 12232
rect 132592 12188 132600 12222
rect 132600 12188 132634 12222
rect 132634 12188 132644 12222
rect 132592 12180 132644 12188
rect 137744 12222 137796 12232
rect 137744 12188 137752 12222
rect 137752 12188 137786 12222
rect 137786 12188 137796 12222
rect 137744 12180 137796 12188
rect 148048 12180 148100 12232
rect 149336 12180 149388 12232
rect 149428 12222 149480 12232
rect 149428 12188 149436 12222
rect 149436 12188 149470 12222
rect 149470 12188 149480 12222
rect 149428 12180 149480 12188
rect 151360 12180 151412 12232
rect 152740 12316 152792 12368
rect 132500 12112 132552 12164
rect 138020 12154 138072 12164
rect 138020 12120 138028 12154
rect 138028 12120 138062 12154
rect 138062 12120 138072 12154
rect 138020 12112 138072 12120
rect 153752 12384 153804 12436
rect 157248 12384 157300 12436
rect 160928 12384 160980 12436
rect 161572 12384 161624 12436
rect 155040 12316 155092 12368
rect 158904 12316 158956 12368
rect 166448 12384 166500 12436
rect 176476 12384 176528 12436
rect 179512 12384 179564 12436
rect 189172 12384 189224 12436
rect 189632 12384 189684 12436
rect 190828 12384 190880 12436
rect 194048 12384 194100 12436
rect 165436 12316 165488 12368
rect 166080 12358 166132 12368
rect 166080 12324 166088 12358
rect 166088 12324 166122 12358
rect 166122 12324 166132 12358
rect 166080 12316 166132 12324
rect 154120 12248 154172 12300
rect 160376 12248 160428 12300
rect 161480 12290 161532 12300
rect 161480 12256 161488 12290
rect 161488 12256 161522 12290
rect 161522 12256 161532 12290
rect 162492 12290 162544 12300
rect 161480 12248 161532 12256
rect 162492 12256 162500 12290
rect 162500 12256 162534 12290
rect 162534 12256 162544 12290
rect 162492 12248 162544 12256
rect 162676 12290 162728 12300
rect 162676 12256 162684 12290
rect 162684 12256 162718 12290
rect 162718 12256 162728 12290
rect 162676 12248 162728 12256
rect 163596 12290 163648 12300
rect 163596 12256 163604 12290
rect 163604 12256 163638 12290
rect 163638 12256 163648 12290
rect 163596 12248 163648 12256
rect 177764 12316 177816 12368
rect 180892 12358 180944 12368
rect 180892 12324 180900 12358
rect 180900 12324 180934 12358
rect 180934 12324 180944 12358
rect 180892 12316 180944 12324
rect 192576 12358 192628 12368
rect 177120 12290 177172 12300
rect 177120 12256 177128 12290
rect 177128 12256 177162 12290
rect 177162 12256 177172 12290
rect 177120 12248 177172 12256
rect 158812 12180 158864 12232
rect 161756 12180 161808 12232
rect 187976 12248 188028 12300
rect 177856 12180 177908 12232
rect 179144 12222 179196 12232
rect 179144 12188 179152 12222
rect 179152 12188 179186 12222
rect 179186 12188 179196 12222
rect 179144 12180 179196 12188
rect 180708 12180 180760 12232
rect 189540 12222 189592 12232
rect 131580 12044 131632 12096
rect 155868 12112 155920 12164
rect 156420 12112 156472 12164
rect 162584 12112 162636 12164
rect 162676 12112 162728 12164
rect 164332 12112 164384 12164
rect 165896 12154 165948 12164
rect 165896 12120 165904 12154
rect 165904 12120 165938 12154
rect 165938 12120 165948 12154
rect 165896 12112 165948 12120
rect 166540 12112 166592 12164
rect 179420 12154 179472 12164
rect 149520 12044 149572 12096
rect 151636 12086 151688 12096
rect 151636 12052 151644 12086
rect 151644 12052 151678 12086
rect 151678 12052 151688 12086
rect 151636 12044 151688 12052
rect 151728 12044 151780 12096
rect 152188 12044 152240 12096
rect 152556 12044 152608 12096
rect 161112 12044 161164 12096
rect 162216 12044 162268 12096
rect 162860 12044 162912 12096
rect 176660 12044 176712 12096
rect 178040 12086 178092 12096
rect 178040 12052 178048 12086
rect 178048 12052 178082 12086
rect 178082 12052 178092 12086
rect 178040 12044 178092 12052
rect 179420 12120 179428 12154
rect 179428 12120 179462 12154
rect 179462 12120 179472 12154
rect 179420 12112 179472 12120
rect 181444 12112 181496 12164
rect 189540 12188 189548 12222
rect 189548 12188 189582 12222
rect 189582 12188 189592 12222
rect 189540 12180 189592 12188
rect 192576 12324 192584 12358
rect 192584 12324 192618 12358
rect 192618 12324 192628 12358
rect 192576 12316 192628 12324
rect 191840 12248 191892 12300
rect 192668 12248 192720 12300
rect 194416 12222 194468 12232
rect 190828 12112 190880 12164
rect 191104 12154 191156 12164
rect 191104 12120 191112 12154
rect 191112 12120 191146 12154
rect 191146 12120 191156 12154
rect 191104 12112 191156 12120
rect 191196 12112 191248 12164
rect 180156 12044 180208 12096
rect 193404 12154 193456 12164
rect 193404 12120 193412 12154
rect 193412 12120 193446 12154
rect 193446 12120 193456 12154
rect 193404 12112 193456 12120
rect 193036 12086 193088 12096
rect 193036 12052 193044 12086
rect 193044 12052 193078 12086
rect 193078 12052 193088 12086
rect 193036 12044 193088 12052
rect 193680 12044 193732 12096
rect 194416 12188 194424 12222
rect 194424 12188 194458 12222
rect 194458 12188 194468 12222
rect 194416 12180 194468 12188
rect 194692 12154 194744 12164
rect 194692 12120 194700 12154
rect 194700 12120 194734 12154
rect 194734 12120 194744 12154
rect 194692 12112 194744 12120
rect 197452 12316 197504 12368
rect 202420 12384 202472 12436
rect 205640 12384 205692 12436
rect 207664 12384 207716 12436
rect 230112 12384 230164 12436
rect 231860 12384 231912 12436
rect 239036 12384 239088 12436
rect 240140 12384 240192 12436
rect 228824 12316 228876 12368
rect 231124 12316 231176 12368
rect 232504 12316 232556 12368
rect 194968 12044 195020 12096
rect 200488 12248 200540 12300
rect 197452 12222 197504 12232
rect 197452 12188 197460 12222
rect 197460 12188 197494 12222
rect 197494 12188 197504 12222
rect 197452 12180 197504 12188
rect 198372 12180 198424 12232
rect 200580 12180 200632 12232
rect 201040 12222 201092 12232
rect 201040 12188 201048 12222
rect 201048 12188 201082 12222
rect 201082 12188 201092 12222
rect 201040 12180 201092 12188
rect 202052 12248 202104 12300
rect 203524 12290 203576 12300
rect 203524 12256 203532 12290
rect 203532 12256 203566 12290
rect 203566 12256 203576 12290
rect 203524 12248 203576 12256
rect 204536 12180 204588 12232
rect 229928 12222 229980 12232
rect 229928 12188 229936 12222
rect 229936 12188 229970 12222
rect 229970 12188 229980 12222
rect 229928 12180 229980 12188
rect 231308 12180 231360 12232
rect 204996 12154 205048 12164
rect 204996 12120 205004 12154
rect 205004 12120 205038 12154
rect 205038 12120 205048 12154
rect 204996 12112 205048 12120
rect 196808 12086 196860 12096
rect 196808 12052 196816 12086
rect 196816 12052 196850 12086
rect 196850 12052 196860 12086
rect 196808 12044 196860 12052
rect 196992 12086 197044 12096
rect 196992 12052 197000 12086
rect 197000 12052 197034 12086
rect 197034 12052 197044 12086
rect 196992 12044 197044 12052
rect 197360 12086 197412 12096
rect 197360 12052 197368 12086
rect 197368 12052 197402 12086
rect 197402 12052 197412 12086
rect 197360 12044 197412 12052
rect 203064 12044 203116 12096
rect 203432 12044 203484 12096
rect 204260 12044 204312 12096
rect 230848 12112 230900 12164
rect 231124 12112 231176 12164
rect 231676 12248 231728 12300
rect 238852 12248 238904 12300
rect 239312 12290 239364 12300
rect 239312 12256 239320 12290
rect 239320 12256 239354 12290
rect 239354 12256 239364 12290
rect 239312 12248 239364 12256
rect 232136 12222 232188 12232
rect 232136 12188 232144 12222
rect 232144 12188 232178 12222
rect 232178 12188 232188 12222
rect 232136 12180 232188 12188
rect 233056 12180 233108 12232
rect 238024 12222 238076 12232
rect 238024 12188 238032 12222
rect 238032 12188 238066 12222
rect 238066 12188 238076 12222
rect 238024 12180 238076 12188
rect 238392 12180 238444 12232
rect 239128 12222 239180 12232
rect 239128 12188 239136 12222
rect 239136 12188 239170 12222
rect 239170 12188 239180 12222
rect 239128 12180 239180 12188
rect 239496 12180 239548 12232
rect 239956 12248 240008 12300
rect 242256 12316 242308 12368
rect 242440 12248 242492 12300
rect 242992 12316 243044 12368
rect 242900 12290 242952 12300
rect 242900 12256 242908 12290
rect 242908 12256 242942 12290
rect 242942 12256 242952 12290
rect 242900 12248 242952 12256
rect 242164 12180 242216 12232
rect 243636 12384 243688 12436
rect 244188 12426 244240 12436
rect 244188 12392 244196 12426
rect 244196 12392 244230 12426
rect 244230 12392 244240 12426
rect 244188 12384 244240 12392
rect 251364 12384 251416 12436
rect 251916 12384 251968 12436
rect 251456 12316 251508 12368
rect 252100 12358 252152 12368
rect 252100 12324 252108 12358
rect 252108 12324 252142 12358
rect 252142 12324 252152 12358
rect 252100 12316 252152 12324
rect 254308 12358 254360 12368
rect 254308 12324 254316 12358
rect 254316 12324 254350 12358
rect 254350 12324 254360 12358
rect 254308 12316 254360 12324
rect 255228 12316 255280 12368
rect 243176 12248 243228 12300
rect 248328 12248 248380 12300
rect 249248 12248 249300 12300
rect 251272 12222 251324 12232
rect 251272 12188 251280 12222
rect 251280 12188 251314 12222
rect 251314 12188 251324 12222
rect 251916 12222 251968 12232
rect 251272 12180 251324 12188
rect 251916 12188 251924 12222
rect 251924 12188 251958 12222
rect 251958 12188 251968 12222
rect 251916 12180 251968 12188
rect 255136 12222 255188 12232
rect 255136 12188 255144 12222
rect 255144 12188 255178 12222
rect 255178 12188 255188 12222
rect 255136 12180 255188 12188
rect 249064 12154 249116 12164
rect 228824 12044 228876 12096
rect 231216 12044 231268 12096
rect 249064 12120 249072 12154
rect 249072 12120 249106 12154
rect 249106 12120 249116 12154
rect 249064 12112 249116 12120
rect 249248 12154 249300 12164
rect 249248 12120 249256 12154
rect 249256 12120 249290 12154
rect 249290 12120 249300 12154
rect 249248 12112 249300 12120
rect 253112 12112 253164 12164
rect 255596 12248 255648 12300
rect 256516 12384 256568 12436
rect 262496 12426 262548 12436
rect 262496 12392 262504 12426
rect 262504 12392 262538 12426
rect 262538 12392 262548 12426
rect 262496 12384 262548 12392
rect 265532 12384 265584 12436
rect 256976 12316 257028 12368
rect 264980 12316 265032 12368
rect 268016 12384 268068 12436
rect 268384 12384 268436 12436
rect 271052 12426 271104 12436
rect 271052 12392 271060 12426
rect 271060 12392 271094 12426
rect 271094 12392 271104 12426
rect 271052 12384 271104 12392
rect 305460 12426 305512 12436
rect 305460 12392 305468 12426
rect 305468 12392 305502 12426
rect 305502 12392 305512 12426
rect 305460 12384 305512 12392
rect 261852 12248 261904 12300
rect 262404 12248 262456 12300
rect 256240 12222 256292 12232
rect 256240 12188 256248 12222
rect 256248 12188 256282 12222
rect 256282 12188 256292 12222
rect 256240 12180 256292 12188
rect 256332 12180 256384 12232
rect 263048 12180 263100 12232
rect 264152 12248 264204 12300
rect 265164 12248 265216 12300
rect 264336 12180 264388 12232
rect 265624 12248 265676 12300
rect 269120 12248 269172 12300
rect 269672 12248 269724 12300
rect 271144 12248 271196 12300
rect 272248 12290 272300 12300
rect 272248 12256 272256 12290
rect 272256 12256 272290 12290
rect 272290 12256 272300 12290
rect 272248 12248 272300 12256
rect 272800 12248 272852 12300
rect 231400 12086 231452 12096
rect 231400 12052 231408 12086
rect 231408 12052 231442 12086
rect 231442 12052 231452 12086
rect 231400 12044 231452 12052
rect 231768 12044 231820 12096
rect 233056 12044 233108 12096
rect 240876 12086 240928 12096
rect 240876 12052 240884 12086
rect 240884 12052 240918 12086
rect 240918 12052 240928 12086
rect 240876 12044 240928 12052
rect 241520 12044 241572 12096
rect 242532 12044 242584 12096
rect 244096 12044 244148 12096
rect 254400 12044 254452 12096
rect 255044 12044 255096 12096
rect 255228 12086 255280 12096
rect 255228 12052 255236 12086
rect 255236 12052 255270 12086
rect 255270 12052 255280 12086
rect 255228 12044 255280 12052
rect 256332 12044 256384 12096
rect 265164 12112 265216 12164
rect 268108 12180 268160 12232
rect 268660 12180 268712 12232
rect 266820 12154 266872 12164
rect 266820 12120 266828 12154
rect 266828 12120 266862 12154
rect 266862 12120 266872 12154
rect 266820 12112 266872 12120
rect 267280 12112 267332 12164
rect 268200 12112 268252 12164
rect 269488 12112 269540 12164
rect 267004 12044 267056 12096
rect 268476 12044 268528 12096
rect 268660 12044 268712 12096
rect 271328 12180 271380 12232
rect 272892 12180 272944 12232
rect 270408 12044 270460 12096
rect 284760 12044 284812 12096
rect 77148 11942 77200 11994
rect 77212 11942 77264 11994
rect 77276 11942 77328 11994
rect 77340 11942 77392 11994
rect 77404 11942 77456 11994
rect 153346 11942 153398 11994
rect 153410 11942 153462 11994
rect 153474 11942 153526 11994
rect 153538 11942 153590 11994
rect 153602 11942 153654 11994
rect 229544 11942 229596 11994
rect 229608 11942 229660 11994
rect 229672 11942 229724 11994
rect 229736 11942 229788 11994
rect 229800 11942 229852 11994
rect 29092 11840 29144 11892
rect 29460 11840 29512 11892
rect 30932 11840 30984 11892
rect 32220 11840 32272 11892
rect 33784 11882 33836 11892
rect 33784 11848 33792 11882
rect 33792 11848 33826 11882
rect 33826 11848 33836 11882
rect 33784 11840 33836 11848
rect 34428 11882 34480 11892
rect 34428 11848 34436 11882
rect 34436 11848 34470 11882
rect 34470 11848 34480 11882
rect 34428 11840 34480 11848
rect 38384 11882 38436 11892
rect 27712 11772 27764 11824
rect 28724 11772 28776 11824
rect 29000 11772 29052 11824
rect 28908 11678 28960 11688
rect 28908 11644 28916 11678
rect 28916 11644 28950 11678
rect 28950 11644 28960 11678
rect 28908 11636 28960 11644
rect 30012 11772 30064 11824
rect 32036 11772 32088 11824
rect 38384 11848 38392 11882
rect 38392 11848 38426 11882
rect 38426 11848 38436 11882
rect 38384 11840 38436 11848
rect 39580 11840 39632 11892
rect 29552 11704 29604 11756
rect 32404 11704 32456 11756
rect 29920 11678 29972 11688
rect 29920 11644 29928 11678
rect 29928 11644 29962 11678
rect 29962 11644 29972 11678
rect 29920 11636 29972 11644
rect 28448 11542 28500 11552
rect 28448 11508 28456 11542
rect 28456 11508 28490 11542
rect 28490 11508 28500 11542
rect 28448 11500 28500 11508
rect 32588 11636 32640 11688
rect 34704 11704 34756 11756
rect 39948 11840 40000 11892
rect 41420 11840 41472 11892
rect 42892 11840 42944 11892
rect 52644 11840 52696 11892
rect 53656 11882 53708 11892
rect 53656 11848 53664 11882
rect 53664 11848 53698 11882
rect 53698 11848 53708 11882
rect 53656 11840 53708 11848
rect 54392 11882 54444 11892
rect 54392 11848 54400 11882
rect 54400 11848 54434 11882
rect 54434 11848 54444 11882
rect 54392 11840 54444 11848
rect 55312 11882 55364 11892
rect 55312 11848 55320 11882
rect 55320 11848 55354 11882
rect 55354 11848 55364 11882
rect 55312 11840 55364 11848
rect 56600 11840 56652 11892
rect 58624 11840 58676 11892
rect 75460 11840 75512 11892
rect 75644 11840 75696 11892
rect 76472 11840 76524 11892
rect 77852 11882 77904 11892
rect 77852 11848 77860 11882
rect 77860 11848 77894 11882
rect 77894 11848 77904 11882
rect 77852 11840 77904 11848
rect 78496 11882 78548 11892
rect 78496 11848 78504 11882
rect 78504 11848 78538 11882
rect 78538 11848 78548 11882
rect 78496 11840 78548 11848
rect 84292 11840 84344 11892
rect 86040 11882 86092 11892
rect 34060 11636 34112 11688
rect 31116 11568 31168 11620
rect 40684 11772 40736 11824
rect 41236 11772 41288 11824
rect 53748 11772 53800 11824
rect 40316 11704 40368 11756
rect 42800 11704 42852 11756
rect 42984 11704 43036 11756
rect 53012 11746 53064 11756
rect 40960 11636 41012 11688
rect 41420 11636 41472 11688
rect 53012 11712 53020 11746
rect 53020 11712 53054 11746
rect 53054 11712 53064 11746
rect 53012 11704 53064 11712
rect 57428 11772 57480 11824
rect 84936 11772 84988 11824
rect 54668 11636 54720 11688
rect 55588 11678 55640 11688
rect 55588 11644 55596 11678
rect 55596 11644 55630 11678
rect 55630 11644 55640 11678
rect 55588 11636 55640 11644
rect 55864 11636 55916 11688
rect 76012 11704 76064 11756
rect 76288 11704 76340 11756
rect 78588 11704 78640 11756
rect 81440 11704 81492 11756
rect 86040 11848 86048 11882
rect 86048 11848 86082 11882
rect 86082 11848 86092 11882
rect 86040 11840 86092 11848
rect 86132 11840 86184 11892
rect 87880 11882 87932 11892
rect 87880 11848 87888 11882
rect 87888 11848 87922 11882
rect 87922 11848 87932 11882
rect 87880 11840 87932 11848
rect 89536 11840 89588 11892
rect 99656 11840 99708 11892
rect 100944 11882 100996 11892
rect 100944 11848 100952 11882
rect 100952 11848 100986 11882
rect 100986 11848 100996 11882
rect 100944 11840 100996 11848
rect 103060 11840 103112 11892
rect 103520 11840 103572 11892
rect 113824 11882 113876 11892
rect 85304 11772 85356 11824
rect 113824 11848 113832 11882
rect 113832 11848 113866 11882
rect 113866 11848 113876 11882
rect 113824 11840 113876 11848
rect 114284 11840 114336 11892
rect 115664 11840 115716 11892
rect 116768 11840 116820 11892
rect 117320 11840 117372 11892
rect 118792 11840 118844 11892
rect 129372 11882 129424 11892
rect 129372 11848 129380 11882
rect 129380 11848 129414 11882
rect 129414 11848 129424 11882
rect 129372 11840 129424 11848
rect 130292 11840 130344 11892
rect 130936 11882 130988 11892
rect 130936 11848 130944 11882
rect 130944 11848 130978 11882
rect 130978 11848 130988 11882
rect 130936 11840 130988 11848
rect 131120 11840 131172 11892
rect 137744 11840 137796 11892
rect 151084 11882 151136 11892
rect 75000 11636 75052 11688
rect 76932 11636 76984 11688
rect 84016 11636 84068 11688
rect 85764 11704 85816 11756
rect 86960 11746 87012 11756
rect 86960 11712 86968 11746
rect 86968 11712 87002 11746
rect 87002 11712 87012 11746
rect 86960 11704 87012 11712
rect 86316 11678 86368 11688
rect 86316 11644 86324 11678
rect 86324 11644 86358 11678
rect 86358 11644 86368 11678
rect 86316 11636 86368 11644
rect 89168 11704 89220 11756
rect 100392 11746 100444 11756
rect 100392 11712 100400 11746
rect 100400 11712 100434 11746
rect 100434 11712 100444 11746
rect 100392 11704 100444 11712
rect 102140 11704 102192 11756
rect 103612 11704 103664 11756
rect 56048 11568 56100 11620
rect 90456 11636 90508 11688
rect 100760 11636 100812 11688
rect 102048 11678 102100 11688
rect 102048 11644 102056 11678
rect 102056 11644 102090 11678
rect 102090 11644 102100 11678
rect 102048 11636 102100 11644
rect 102324 11636 102376 11688
rect 103520 11636 103572 11688
rect 114560 11772 114612 11824
rect 114008 11746 114060 11756
rect 114008 11712 114016 11746
rect 114016 11712 114050 11746
rect 114050 11712 114060 11746
rect 114008 11704 114060 11712
rect 138020 11772 138072 11824
rect 149980 11772 150032 11824
rect 151084 11848 151092 11882
rect 151092 11848 151126 11882
rect 151126 11848 151136 11882
rect 151084 11840 151136 11848
rect 152004 11882 152056 11892
rect 152004 11848 152012 11882
rect 152012 11848 152046 11882
rect 152046 11848 152056 11882
rect 152004 11840 152056 11848
rect 154212 11840 154264 11892
rect 115020 11704 115072 11756
rect 116400 11746 116452 11756
rect 116400 11712 116408 11746
rect 116408 11712 116442 11746
rect 116442 11712 116452 11746
rect 116400 11704 116452 11712
rect 115664 11636 115716 11688
rect 115756 11636 115808 11688
rect 118332 11704 118384 11756
rect 128360 11704 128412 11756
rect 130292 11704 130344 11756
rect 131580 11704 131632 11756
rect 129740 11636 129792 11688
rect 131028 11678 131080 11688
rect 131028 11644 131036 11678
rect 131036 11644 131070 11678
rect 131070 11644 131080 11678
rect 131028 11636 131080 11644
rect 132500 11704 132552 11756
rect 147680 11704 147732 11756
rect 151268 11746 151320 11756
rect 151268 11712 151276 11746
rect 151276 11712 151310 11746
rect 151310 11712 151320 11746
rect 151268 11704 151320 11712
rect 152188 11746 152240 11756
rect 152188 11712 152196 11746
rect 152196 11712 152230 11746
rect 152230 11712 152240 11746
rect 152188 11704 152240 11712
rect 152740 11704 152792 11756
rect 161112 11746 161164 11756
rect 161112 11712 161120 11746
rect 161120 11712 161154 11746
rect 161154 11712 161164 11746
rect 161112 11704 161164 11712
rect 161756 11746 161808 11756
rect 161756 11712 161764 11746
rect 161764 11712 161798 11746
rect 161798 11712 161808 11746
rect 161756 11704 161808 11712
rect 137744 11636 137796 11688
rect 148324 11678 148376 11688
rect 148324 11644 148332 11678
rect 148332 11644 148366 11678
rect 148366 11644 148376 11678
rect 148324 11636 148376 11644
rect 148600 11678 148652 11688
rect 148600 11644 148608 11678
rect 148608 11644 148642 11678
rect 148642 11644 148652 11678
rect 148600 11636 148652 11644
rect 143264 11568 143316 11620
rect 146024 11568 146076 11620
rect 161204 11568 161256 11620
rect 161296 11568 161348 11620
rect 162032 11840 162084 11892
rect 162768 11840 162820 11892
rect 163780 11840 163832 11892
rect 164332 11840 164384 11892
rect 164884 11882 164936 11892
rect 164884 11848 164892 11882
rect 164892 11848 164926 11882
rect 164926 11848 164936 11882
rect 164884 11840 164936 11848
rect 176752 11840 176804 11892
rect 177396 11840 177448 11892
rect 177856 11840 177908 11892
rect 179880 11840 179932 11892
rect 179972 11840 180024 11892
rect 180156 11840 180208 11892
rect 188344 11840 188396 11892
rect 191748 11840 191800 11892
rect 191840 11840 191892 11892
rect 162584 11772 162636 11824
rect 189540 11772 189592 11824
rect 193864 11772 193916 11824
rect 163688 11746 163740 11756
rect 163688 11712 163696 11746
rect 163696 11712 163730 11746
rect 163730 11712 163740 11746
rect 163688 11704 163740 11712
rect 163504 11636 163556 11688
rect 166632 11704 166684 11756
rect 176660 11746 176712 11756
rect 176660 11712 176668 11746
rect 176668 11712 176702 11746
rect 176702 11712 176712 11746
rect 176660 11704 176712 11712
rect 179880 11704 179932 11756
rect 177120 11636 177172 11688
rect 165896 11568 165948 11620
rect 31392 11542 31444 11552
rect 31392 11508 31400 11542
rect 31400 11508 31434 11542
rect 31434 11508 31444 11542
rect 31392 11500 31444 11508
rect 32956 11500 33008 11552
rect 55496 11500 55548 11552
rect 84844 11500 84896 11552
rect 86408 11500 86460 11552
rect 101864 11500 101916 11552
rect 104072 11500 104124 11552
rect 114008 11500 114060 11552
rect 131856 11542 131908 11552
rect 131856 11508 131864 11542
rect 131864 11508 131898 11542
rect 131898 11508 131908 11542
rect 131856 11500 131908 11508
rect 147312 11500 147364 11552
rect 151728 11500 151780 11552
rect 180064 11704 180116 11756
rect 180616 11704 180668 11756
rect 180800 11636 180852 11688
rect 181536 11636 181588 11688
rect 189632 11746 189684 11756
rect 189632 11712 189640 11746
rect 189640 11712 189674 11746
rect 189674 11712 189684 11746
rect 189632 11704 189684 11712
rect 190828 11704 190880 11756
rect 191840 11746 191892 11756
rect 191840 11712 191848 11746
rect 191848 11712 191882 11746
rect 191882 11712 191892 11746
rect 191840 11704 191892 11712
rect 194416 11840 194468 11892
rect 194692 11840 194744 11892
rect 202880 11882 202932 11892
rect 202880 11848 202888 11882
rect 202888 11848 202922 11882
rect 202922 11848 202932 11882
rect 202880 11840 202932 11848
rect 204536 11840 204588 11892
rect 206560 11840 206612 11892
rect 227812 11840 227864 11892
rect 228824 11840 228876 11892
rect 196808 11772 196860 11824
rect 203156 11772 203208 11824
rect 205548 11772 205600 11824
rect 227720 11772 227772 11824
rect 229928 11840 229980 11892
rect 230388 11882 230440 11892
rect 230388 11848 230396 11882
rect 230396 11848 230430 11882
rect 230430 11848 230440 11882
rect 230388 11840 230440 11848
rect 231032 11840 231084 11892
rect 231676 11840 231728 11892
rect 240324 11882 240376 11892
rect 240324 11848 240332 11882
rect 240332 11848 240366 11882
rect 240366 11848 240376 11882
rect 240324 11840 240376 11848
rect 241060 11882 241112 11892
rect 241060 11848 241068 11882
rect 241068 11848 241102 11882
rect 241102 11848 241112 11882
rect 241060 11840 241112 11848
rect 241796 11882 241848 11892
rect 241796 11848 241804 11882
rect 241804 11848 241838 11882
rect 241838 11848 241848 11882
rect 241796 11840 241848 11848
rect 252928 11840 252980 11892
rect 254676 11840 254728 11892
rect 254768 11840 254820 11892
rect 255044 11840 255096 11892
rect 266820 11840 266872 11892
rect 197912 11704 197964 11756
rect 201040 11704 201092 11756
rect 203064 11746 203116 11756
rect 203064 11712 203072 11746
rect 203072 11712 203106 11746
rect 203106 11712 203116 11746
rect 203064 11704 203116 11712
rect 192116 11678 192168 11688
rect 192116 11644 192124 11678
rect 192124 11644 192158 11678
rect 192158 11644 192168 11678
rect 192116 11636 192168 11644
rect 194324 11678 194376 11688
rect 194324 11644 194332 11678
rect 194332 11644 194366 11678
rect 194366 11644 194376 11678
rect 194324 11636 194376 11644
rect 194416 11636 194468 11688
rect 180340 11568 180392 11620
rect 197360 11636 197412 11688
rect 201316 11636 201368 11688
rect 202880 11636 202932 11688
rect 206376 11704 206428 11756
rect 230848 11772 230900 11824
rect 229376 11704 229428 11756
rect 240140 11772 240192 11824
rect 203524 11636 203576 11688
rect 207848 11636 207900 11688
rect 227260 11636 227312 11688
rect 180524 11500 180576 11552
rect 189448 11542 189500 11552
rect 189448 11508 189456 11542
rect 189456 11508 189490 11542
rect 189490 11508 189500 11542
rect 189448 11500 189500 11508
rect 197452 11568 197504 11620
rect 203432 11568 203484 11620
rect 204904 11568 204956 11620
rect 230296 11568 230348 11620
rect 193312 11500 193364 11552
rect 193496 11500 193548 11552
rect 195796 11500 195848 11552
rect 195888 11500 195940 11552
rect 196992 11500 197044 11552
rect 201500 11500 201552 11552
rect 204812 11542 204864 11552
rect 204812 11508 204820 11542
rect 204820 11508 204854 11542
rect 204854 11508 204864 11542
rect 204812 11500 204864 11508
rect 229376 11500 229428 11552
rect 231216 11704 231268 11756
rect 241520 11772 241572 11824
rect 239312 11636 239364 11688
rect 239956 11636 240008 11688
rect 232136 11568 232188 11620
rect 242532 11746 242584 11756
rect 242532 11712 242540 11746
rect 242540 11712 242574 11746
rect 242574 11712 242584 11746
rect 242532 11704 242584 11712
rect 241980 11636 242032 11688
rect 244832 11772 244884 11824
rect 254308 11772 254360 11824
rect 270684 11840 270736 11892
rect 270776 11840 270828 11892
rect 268292 11772 268344 11824
rect 269856 11772 269908 11824
rect 252008 11746 252060 11756
rect 252008 11712 252016 11746
rect 252016 11712 252050 11746
rect 252050 11712 252060 11746
rect 252008 11704 252060 11712
rect 252744 11746 252796 11756
rect 252744 11712 252752 11746
rect 252752 11712 252786 11746
rect 252786 11712 252796 11746
rect 252744 11704 252796 11712
rect 253020 11704 253072 11756
rect 256240 11704 256292 11756
rect 257252 11704 257304 11756
rect 264336 11746 264388 11756
rect 264336 11712 264344 11746
rect 264344 11712 264378 11746
rect 264378 11712 264388 11746
rect 264336 11704 264388 11712
rect 265164 11746 265216 11756
rect 265164 11712 265172 11746
rect 265172 11712 265206 11746
rect 265206 11712 265216 11746
rect 265164 11704 265216 11712
rect 265256 11704 265308 11756
rect 242716 11636 242768 11688
rect 244556 11636 244608 11688
rect 252100 11636 252152 11688
rect 255596 11636 255648 11688
rect 256424 11636 256476 11688
rect 263968 11636 264020 11688
rect 268476 11704 268528 11756
rect 269120 11746 269172 11756
rect 269120 11712 269128 11746
rect 269128 11712 269162 11746
rect 269162 11712 269172 11746
rect 269120 11704 269172 11712
rect 271328 11746 271380 11756
rect 271328 11712 271336 11746
rect 271336 11712 271370 11746
rect 271370 11712 271380 11746
rect 271328 11704 271380 11712
rect 231676 11500 231728 11552
rect 239404 11500 239456 11552
rect 241244 11500 241296 11552
rect 251640 11568 251692 11620
rect 249064 11500 249116 11552
rect 253296 11500 253348 11552
rect 268016 11568 268068 11620
rect 261760 11500 261812 11552
rect 262680 11500 262732 11552
rect 266268 11500 266320 11552
rect 266360 11500 266412 11552
rect 269396 11678 269448 11688
rect 269396 11644 269404 11678
rect 269404 11644 269438 11678
rect 269438 11644 269448 11678
rect 269396 11636 269448 11644
rect 269948 11636 270000 11688
rect 273168 11636 273220 11688
rect 275100 11500 275152 11552
rect 39048 11398 39100 11450
rect 39112 11398 39164 11450
rect 39176 11398 39228 11450
rect 39240 11398 39292 11450
rect 39304 11398 39356 11450
rect 115246 11398 115298 11450
rect 115310 11398 115362 11450
rect 115374 11398 115426 11450
rect 115438 11398 115490 11450
rect 115502 11398 115554 11450
rect 191444 11398 191496 11450
rect 191508 11398 191560 11450
rect 191572 11398 191624 11450
rect 191636 11398 191688 11450
rect 191700 11398 191752 11450
rect 267642 11398 267694 11450
rect 267706 11398 267758 11450
rect 267770 11398 267822 11450
rect 267834 11398 267886 11450
rect 267898 11398 267950 11450
rect 29920 11296 29972 11348
rect 30012 11296 30064 11348
rect 28908 11228 28960 11280
rect 32404 11296 32456 11348
rect 33324 11296 33376 11348
rect 33600 11338 33652 11348
rect 33600 11304 33608 11338
rect 33608 11304 33642 11338
rect 33642 11304 33652 11338
rect 33600 11296 33652 11304
rect 40408 11296 40460 11348
rect 41052 11338 41104 11348
rect 41052 11304 41060 11338
rect 41060 11304 41094 11338
rect 41094 11304 41104 11338
rect 41052 11296 41104 11304
rect 41604 11338 41656 11348
rect 41604 11304 41612 11338
rect 41612 11304 41646 11338
rect 41646 11304 41656 11338
rect 41604 11296 41656 11304
rect 55036 11296 55088 11348
rect 57704 11296 57756 11348
rect 76380 11296 76432 11348
rect 78772 11296 78824 11348
rect 84476 11296 84528 11348
rect 87144 11296 87196 11348
rect 89076 11296 89128 11348
rect 102876 11338 102928 11348
rect 102876 11304 102884 11338
rect 102884 11304 102918 11338
rect 102918 11304 102928 11338
rect 102876 11296 102928 11304
rect 115112 11296 115164 11348
rect 117688 11296 117740 11348
rect 130384 11296 130436 11348
rect 131212 11338 131264 11348
rect 131212 11304 131220 11338
rect 131220 11304 131254 11338
rect 131254 11304 131264 11338
rect 131212 11296 131264 11304
rect 132868 11296 132920 11348
rect 148048 11338 148100 11348
rect 148048 11304 148056 11338
rect 148056 11304 148090 11338
rect 148090 11304 148100 11338
rect 148048 11296 148100 11304
rect 150808 11338 150860 11348
rect 150808 11304 150816 11338
rect 150816 11304 150850 11338
rect 150850 11304 150860 11338
rect 150808 11296 150860 11304
rect 157248 11296 157300 11348
rect 162124 11296 162176 11348
rect 162676 11338 162728 11348
rect 162676 11304 162684 11338
rect 162684 11304 162718 11338
rect 162718 11304 162728 11338
rect 162676 11296 162728 11304
rect 163412 11296 163464 11348
rect 165896 11296 165948 11348
rect 239404 11296 239456 11348
rect 239772 11296 239824 11348
rect 240048 11296 240100 11348
rect 240968 11296 241020 11348
rect 242072 11296 242124 11348
rect 252468 11296 252520 11348
rect 253112 11338 253164 11348
rect 253112 11304 253120 11338
rect 253120 11304 253154 11338
rect 253154 11304 253164 11338
rect 253112 11296 253164 11304
rect 254032 11296 254084 11348
rect 265440 11296 265492 11348
rect 266268 11296 266320 11348
rect 27068 11160 27120 11212
rect 29460 11160 29512 11212
rect 29552 11160 29604 11212
rect 36452 11228 36504 11280
rect 41328 11228 41380 11280
rect 86776 11228 86828 11280
rect 102232 11228 102284 11280
rect 114192 11228 114244 11280
rect 147404 11228 147456 11280
rect 31392 11160 31444 11212
rect 32312 11202 32364 11212
rect 32312 11168 32320 11202
rect 32320 11168 32354 11202
rect 32354 11168 32364 11202
rect 32312 11160 32364 11168
rect 27620 11092 27672 11144
rect 32220 11134 32272 11144
rect 32220 11100 32228 11134
rect 32228 11100 32262 11134
rect 32262 11100 32272 11134
rect 32220 11092 32272 11100
rect 27988 11024 28040 11076
rect 29920 11066 29972 11076
rect 29920 11032 29928 11066
rect 29928 11032 29962 11066
rect 29962 11032 29972 11066
rect 29920 11024 29972 11032
rect 31668 11024 31720 11076
rect 31760 11024 31812 11076
rect 32588 11160 32640 11212
rect 34704 11092 34756 11144
rect 40500 11134 40552 11144
rect 40500 11100 40508 11134
rect 40508 11100 40542 11134
rect 40542 11100 40552 11134
rect 40500 11092 40552 11100
rect 41420 11092 41472 11144
rect 45008 11160 45060 11212
rect 85488 11160 85540 11212
rect 42432 11134 42484 11144
rect 42432 11100 42440 11134
rect 42440 11100 42474 11134
rect 42474 11100 42484 11134
rect 42432 11092 42484 11100
rect 55496 11134 55548 11144
rect 55496 11100 55504 11134
rect 55504 11100 55538 11134
rect 55538 11100 55548 11134
rect 55496 11092 55548 11100
rect 57244 11092 57296 11144
rect 74724 11092 74776 11144
rect 78404 11134 78456 11144
rect 78404 11100 78412 11134
rect 78412 11100 78446 11134
rect 78446 11100 78456 11134
rect 78404 11092 78456 11100
rect 86408 11134 86460 11144
rect 86408 11100 86416 11134
rect 86416 11100 86450 11134
rect 86450 11100 86460 11134
rect 86408 11092 86460 11100
rect 89168 11160 89220 11212
rect 102048 11160 102100 11212
rect 102600 11160 102652 11212
rect 87788 11134 87840 11144
rect 87788 11100 87796 11134
rect 87796 11100 87830 11134
rect 87830 11100 87840 11134
rect 87788 11092 87840 11100
rect 88432 11134 88484 11144
rect 88432 11100 88440 11134
rect 88440 11100 88474 11134
rect 88474 11100 88484 11134
rect 88432 11092 88484 11100
rect 102416 11092 102468 11144
rect 103060 11134 103112 11144
rect 103060 11100 103068 11134
rect 103068 11100 103102 11134
rect 103102 11100 103112 11134
rect 103060 11092 103112 11100
rect 130292 11160 130344 11212
rect 114744 11092 114796 11144
rect 115756 11092 115808 11144
rect 115848 11092 115900 11144
rect 119712 11092 119764 11144
rect 130936 11092 130988 11144
rect 132592 11160 132644 11212
rect 143264 11160 143316 11212
rect 133144 11092 133196 11144
rect 142068 11134 142120 11144
rect 142068 11100 142076 11134
rect 142076 11100 142110 11134
rect 142110 11100 142120 11134
rect 142068 11092 142120 11100
rect 145748 11092 145800 11144
rect 147496 11160 147548 11212
rect 156420 11228 156472 11280
rect 165436 11228 165488 11280
rect 151360 11160 151412 11212
rect 81624 11024 81676 11076
rect 87880 11024 87932 11076
rect 113732 11024 113784 11076
rect 140688 11024 140740 11076
rect 153108 11092 153160 11144
rect 162216 11134 162268 11144
rect 162216 11100 162224 11134
rect 162224 11100 162258 11134
rect 162258 11100 162268 11134
rect 162216 11092 162268 11100
rect 165344 11160 165396 11212
rect 177672 11160 177724 11212
rect 177948 11160 178000 11212
rect 163504 11134 163556 11144
rect 163504 11100 163512 11134
rect 163512 11100 163546 11134
rect 163546 11100 163556 11134
rect 163504 11092 163556 11100
rect 178040 11092 178092 11144
rect 180800 11160 180852 11212
rect 191196 11160 191248 11212
rect 191840 11160 191892 11212
rect 252744 11228 252796 11280
rect 253204 11228 253256 11280
rect 265164 11228 265216 11280
rect 269304 11296 269356 11348
rect 193496 11160 193548 11212
rect 194416 11160 194468 11212
rect 194600 11160 194652 11212
rect 180432 11092 180484 11144
rect 188988 11092 189040 11144
rect 190644 11092 190696 11144
rect 190828 11134 190880 11144
rect 190828 11100 190836 11134
rect 190836 11100 190870 11134
rect 190870 11100 190880 11134
rect 190828 11092 190880 11100
rect 191932 11092 191984 11144
rect 194876 11092 194928 11144
rect 196440 11160 196492 11212
rect 201040 11160 201092 11212
rect 195796 11134 195848 11144
rect 31852 10998 31904 11008
rect 31852 10964 31860 10998
rect 31860 10964 31894 10998
rect 31894 10964 31904 10998
rect 31852 10956 31904 10964
rect 149060 10956 149112 11008
rect 149520 10956 149572 11008
rect 156144 11024 156196 11076
rect 179420 11024 179472 11076
rect 189448 11024 189500 11076
rect 193312 11024 193364 11076
rect 195796 11100 195804 11134
rect 195804 11100 195838 11134
rect 195838 11100 195848 11134
rect 195796 11092 195848 11100
rect 202696 11092 202748 11144
rect 203340 11160 203392 11212
rect 194416 10998 194468 11008
rect 194416 10964 194424 10998
rect 194424 10964 194458 10998
rect 194458 10964 194468 10998
rect 194416 10956 194468 10964
rect 195244 11024 195296 11076
rect 204996 11160 205048 11212
rect 238024 11160 238076 11212
rect 242716 11160 242768 11212
rect 267280 11160 267332 11212
rect 268016 11160 268068 11212
rect 204076 11024 204128 11076
rect 204904 11134 204956 11144
rect 204904 11100 204912 11134
rect 204912 11100 204946 11134
rect 204946 11100 204956 11134
rect 229376 11134 229428 11144
rect 204904 11092 204956 11100
rect 229376 11100 229384 11134
rect 229384 11100 229418 11134
rect 229418 11100 229428 11134
rect 229376 11092 229428 11100
rect 205456 11024 205508 11076
rect 230756 11024 230808 11076
rect 240876 11092 240928 11144
rect 241980 11092 242032 11144
rect 251548 11092 251600 11144
rect 253020 11092 253072 11144
rect 253296 11134 253348 11144
rect 253296 11100 253304 11134
rect 253304 11100 253338 11134
rect 253338 11100 253348 11134
rect 253296 11092 253348 11100
rect 254400 11092 254452 11144
rect 254676 11092 254728 11144
rect 264336 11092 264388 11144
rect 264888 11134 264940 11144
rect 264888 11100 264896 11134
rect 264896 11100 264930 11134
rect 264930 11100 264940 11134
rect 264888 11092 264940 11100
rect 265624 11092 265676 11144
rect 268476 11160 268528 11212
rect 268936 11160 268988 11212
rect 272248 11160 272300 11212
rect 269672 11092 269724 11144
rect 270408 11134 270460 11144
rect 270408 11100 270416 11134
rect 270416 11100 270450 11134
rect 270450 11100 270460 11134
rect 270408 11092 270460 11100
rect 270868 11092 270920 11144
rect 268292 11024 268344 11076
rect 268936 11024 268988 11076
rect 269948 11024 270000 11076
rect 268844 10998 268896 11008
rect 268844 10964 268852 10998
rect 268852 10964 268886 10998
rect 268886 10964 268896 10998
rect 268844 10956 268896 10964
rect 270040 10998 270092 11008
rect 270040 10964 270048 10998
rect 270048 10964 270082 10998
rect 270082 10964 270092 10998
rect 270040 10956 270092 10964
rect 77148 10854 77200 10906
rect 77212 10854 77264 10906
rect 77276 10854 77328 10906
rect 77340 10854 77392 10906
rect 77404 10854 77456 10906
rect 153346 10854 153398 10906
rect 153410 10854 153462 10906
rect 153474 10854 153526 10906
rect 153538 10854 153590 10906
rect 153602 10854 153654 10906
rect 229544 10854 229596 10906
rect 229608 10854 229660 10906
rect 229672 10854 229724 10906
rect 229736 10854 229788 10906
rect 229800 10854 229852 10906
rect 29828 10752 29880 10804
rect 30472 10752 30524 10804
rect 30748 10794 30800 10804
rect 30748 10760 30756 10794
rect 30756 10760 30790 10794
rect 30790 10760 30800 10794
rect 30748 10752 30800 10760
rect 29736 10684 29788 10736
rect 28448 10616 28500 10668
rect 30196 10684 30248 10736
rect 32680 10752 32732 10804
rect 33048 10752 33100 10804
rect 101680 10794 101732 10804
rect 101680 10760 101688 10794
rect 101688 10760 101722 10794
rect 101722 10760 101732 10794
rect 101680 10752 101732 10760
rect 130476 10794 130528 10804
rect 130476 10760 130484 10794
rect 130484 10760 130518 10794
rect 130518 10760 130528 10794
rect 130476 10752 130528 10760
rect 141976 10794 142028 10804
rect 141976 10760 141984 10794
rect 141984 10760 142018 10794
rect 142018 10760 142028 10794
rect 141976 10752 142028 10760
rect 148600 10752 148652 10804
rect 148968 10752 149020 10804
rect 191104 10752 191156 10804
rect 31760 10684 31812 10736
rect 31852 10684 31904 10736
rect 140688 10726 140740 10736
rect 32956 10658 33008 10668
rect 32956 10624 32964 10658
rect 32964 10624 32998 10658
rect 32998 10624 33008 10658
rect 32956 10616 33008 10624
rect 140688 10692 140696 10726
rect 140696 10692 140730 10726
rect 140730 10692 140740 10726
rect 140688 10684 140740 10692
rect 101864 10658 101916 10668
rect 101864 10624 101872 10658
rect 101872 10624 101906 10658
rect 101906 10624 101916 10658
rect 101864 10616 101916 10624
rect 130292 10616 130344 10668
rect 151636 10684 151688 10736
rect 156144 10726 156196 10736
rect 156144 10692 156152 10726
rect 156152 10692 156186 10726
rect 156186 10692 156196 10726
rect 156144 10684 156196 10692
rect 150348 10616 150400 10668
rect 192208 10684 192260 10736
rect 190552 10616 190604 10668
rect 192300 10616 192352 10668
rect 193220 10684 193272 10736
rect 193864 10752 193916 10804
rect 205088 10752 205140 10804
rect 255228 10752 255280 10804
rect 266544 10794 266596 10804
rect 266544 10760 266552 10794
rect 266552 10760 266586 10794
rect 266586 10760 266596 10794
rect 266544 10752 266596 10760
rect 268200 10752 268252 10804
rect 269396 10752 269448 10804
rect 195060 10684 195112 10736
rect 264888 10684 264940 10736
rect 194140 10658 194192 10668
rect 194140 10624 194148 10658
rect 194148 10624 194182 10658
rect 194182 10624 194192 10658
rect 194140 10616 194192 10624
rect 194968 10616 195020 10668
rect 204812 10616 204864 10668
rect 254952 10616 255004 10668
rect 266360 10616 266412 10668
rect 270040 10684 270092 10736
rect 187516 10590 187568 10600
rect 187516 10556 187524 10590
rect 187524 10556 187558 10590
rect 187558 10556 187568 10590
rect 187516 10548 187568 10556
rect 192116 10480 192168 10532
rect 201040 10548 201092 10600
rect 269028 10616 269080 10668
rect 270316 10616 270368 10668
rect 272524 10548 272576 10600
rect 179144 10412 179196 10464
rect 268752 10480 268804 10532
rect 203524 10412 203576 10464
rect 269580 10412 269632 10464
rect 39048 10310 39100 10362
rect 39112 10310 39164 10362
rect 39176 10310 39228 10362
rect 39240 10310 39292 10362
rect 39304 10310 39356 10362
rect 115246 10310 115298 10362
rect 115310 10310 115362 10362
rect 115374 10310 115426 10362
rect 115438 10310 115490 10362
rect 115502 10310 115554 10362
rect 191444 10310 191496 10362
rect 191508 10310 191560 10362
rect 191572 10310 191624 10362
rect 191636 10310 191688 10362
rect 191700 10310 191752 10362
rect 267642 10310 267694 10362
rect 267706 10310 267758 10362
rect 267770 10310 267822 10362
rect 267834 10310 267886 10362
rect 267898 10310 267950 10362
rect 30104 10208 30156 10260
rect 31668 10250 31720 10260
rect 31668 10216 31676 10250
rect 31676 10216 31710 10250
rect 31710 10216 31720 10250
rect 31668 10208 31720 10216
rect 32128 10208 32180 10260
rect 33324 10208 33376 10260
rect 191288 10208 191340 10260
rect 192484 10208 192536 10260
rect 266912 10208 266964 10260
rect 268568 10208 268620 10260
rect 27528 10140 27580 10192
rect 31576 10140 31628 10192
rect 163596 10072 163648 10124
rect 29460 10004 29512 10056
rect 30932 10004 30984 10056
rect 33416 10004 33468 10056
rect 33692 10004 33744 10056
rect 140688 10004 140740 10056
rect 156144 10004 156196 10056
rect 192576 10004 192628 10056
rect 195888 10072 195940 10124
rect 267740 10072 267792 10124
rect 194416 10004 194468 10056
rect 268384 10140 268436 10192
rect 269488 10140 269540 10192
rect 268844 10072 268896 10124
rect 268108 10004 268160 10056
rect 269028 10004 269080 10056
rect 269212 10046 269264 10056
rect 269212 10012 269220 10046
rect 269220 10012 269254 10046
rect 269254 10012 269264 10046
rect 269212 10004 269264 10012
rect 304448 10046 304500 10056
rect 304448 10012 304456 10046
rect 304456 10012 304490 10046
rect 304490 10012 304500 10046
rect 304448 10004 304500 10012
rect 252744 9936 252796 9988
rect 117412 9868 117464 9920
rect 194324 9868 194376 9920
rect 267740 9868 267792 9920
rect 270960 9868 271012 9920
rect 77148 9766 77200 9818
rect 77212 9766 77264 9818
rect 77276 9766 77328 9818
rect 77340 9766 77392 9818
rect 77404 9766 77456 9818
rect 153346 9766 153398 9818
rect 153410 9766 153462 9818
rect 153474 9766 153526 9818
rect 153538 9766 153590 9818
rect 153602 9766 153654 9818
rect 229544 9766 229596 9818
rect 229608 9766 229660 9818
rect 229672 9766 229724 9818
rect 229736 9766 229788 9818
rect 229800 9766 229852 9818
rect 31208 9596 31260 9648
rect 140688 9638 140740 9648
rect 140688 9604 140696 9638
rect 140696 9604 140730 9638
rect 140730 9604 140740 9638
rect 140688 9596 140740 9604
rect 156144 9638 156196 9648
rect 156144 9604 156152 9638
rect 156152 9604 156186 9638
rect 156186 9604 156196 9638
rect 156144 9596 156196 9604
rect 158628 9596 158680 9648
rect 190644 9596 190696 9648
rect 27344 9528 27396 9580
rect 33692 9528 33744 9580
rect 193312 9596 193364 9648
rect 269856 9596 269908 9648
rect 30564 9460 30616 9512
rect 194140 9528 194192 9580
rect 268108 9528 268160 9580
rect 195980 9460 196032 9512
rect 29920 9392 29972 9444
rect 194508 9392 194560 9444
rect 104256 9324 104308 9376
rect 148324 9324 148376 9376
rect 39048 9222 39100 9274
rect 39112 9222 39164 9274
rect 39176 9222 39228 9274
rect 39240 9222 39292 9274
rect 39304 9222 39356 9274
rect 115246 9222 115298 9274
rect 115310 9222 115362 9274
rect 115374 9222 115426 9274
rect 115438 9222 115490 9274
rect 115502 9222 115554 9274
rect 191444 9222 191496 9274
rect 191508 9222 191560 9274
rect 191572 9222 191624 9274
rect 191636 9222 191688 9274
rect 191700 9222 191752 9274
rect 267642 9222 267694 9274
rect 267706 9222 267758 9274
rect 267770 9222 267822 9274
rect 267834 9222 267886 9274
rect 267898 9222 267950 9274
rect 77148 8678 77200 8730
rect 77212 8678 77264 8730
rect 77276 8678 77328 8730
rect 77340 8678 77392 8730
rect 77404 8678 77456 8730
rect 153346 8678 153398 8730
rect 153410 8678 153462 8730
rect 153474 8678 153526 8730
rect 153538 8678 153590 8730
rect 153602 8678 153654 8730
rect 229544 8678 229596 8730
rect 229608 8678 229660 8730
rect 229672 8678 229724 8730
rect 229736 8678 229788 8730
rect 229800 8678 229852 8730
rect 1400 8346 1452 8356
rect 1400 8312 1408 8346
rect 1408 8312 1442 8346
rect 1442 8312 1452 8346
rect 1400 8304 1452 8312
rect 187516 8304 187568 8356
rect 39048 8134 39100 8186
rect 39112 8134 39164 8186
rect 39176 8134 39228 8186
rect 39240 8134 39292 8186
rect 39304 8134 39356 8186
rect 115246 8134 115298 8186
rect 115310 8134 115362 8186
rect 115374 8134 115426 8186
rect 115438 8134 115490 8186
rect 115502 8134 115554 8186
rect 191444 8134 191496 8186
rect 191508 8134 191560 8186
rect 191572 8134 191624 8186
rect 191636 8134 191688 8186
rect 191700 8134 191752 8186
rect 267642 8134 267694 8186
rect 267706 8134 267758 8186
rect 267770 8134 267822 8186
rect 267834 8134 267886 8186
rect 267898 8134 267950 8186
rect 77148 7590 77200 7642
rect 77212 7590 77264 7642
rect 77276 7590 77328 7642
rect 77340 7590 77392 7642
rect 77404 7590 77456 7642
rect 153346 7590 153398 7642
rect 153410 7590 153462 7642
rect 153474 7590 153526 7642
rect 153538 7590 153590 7642
rect 153602 7590 153654 7642
rect 229544 7590 229596 7642
rect 229608 7590 229660 7642
rect 229672 7590 229724 7642
rect 229736 7590 229788 7642
rect 229800 7590 229852 7642
rect 39048 7046 39100 7098
rect 39112 7046 39164 7098
rect 39176 7046 39228 7098
rect 39240 7046 39292 7098
rect 39304 7046 39356 7098
rect 115246 7046 115298 7098
rect 115310 7046 115362 7098
rect 115374 7046 115426 7098
rect 115438 7046 115490 7098
rect 115502 7046 115554 7098
rect 191444 7046 191496 7098
rect 191508 7046 191560 7098
rect 191572 7046 191624 7098
rect 191636 7046 191688 7098
rect 191700 7046 191752 7098
rect 267642 7046 267694 7098
rect 267706 7046 267758 7098
rect 267770 7046 267822 7098
rect 267834 7046 267886 7098
rect 267898 7046 267950 7098
rect 77148 6502 77200 6554
rect 77212 6502 77264 6554
rect 77276 6502 77328 6554
rect 77340 6502 77392 6554
rect 77404 6502 77456 6554
rect 153346 6502 153398 6554
rect 153410 6502 153462 6554
rect 153474 6502 153526 6554
rect 153538 6502 153590 6554
rect 153602 6502 153654 6554
rect 229544 6502 229596 6554
rect 229608 6502 229660 6554
rect 229672 6502 229724 6554
rect 229736 6502 229788 6554
rect 229800 6502 229852 6554
rect 303988 6306 304040 6316
rect 303988 6272 303996 6306
rect 303996 6272 304030 6306
rect 304030 6272 304040 6306
rect 303988 6264 304040 6272
rect 249064 6196 249116 6248
rect 39048 5958 39100 6010
rect 39112 5958 39164 6010
rect 39176 5958 39228 6010
rect 39240 5958 39292 6010
rect 39304 5958 39356 6010
rect 115246 5958 115298 6010
rect 115310 5958 115362 6010
rect 115374 5958 115426 6010
rect 115438 5958 115490 6010
rect 115502 5958 115554 6010
rect 191444 5958 191496 6010
rect 191508 5958 191560 6010
rect 191572 5958 191624 6010
rect 191636 5958 191688 6010
rect 191700 5958 191752 6010
rect 267642 5958 267694 6010
rect 267706 5958 267758 6010
rect 267770 5958 267822 6010
rect 267834 5958 267886 6010
rect 267898 5958 267950 6010
rect 77148 5414 77200 5466
rect 77212 5414 77264 5466
rect 77276 5414 77328 5466
rect 77340 5414 77392 5466
rect 77404 5414 77456 5466
rect 153346 5414 153398 5466
rect 153410 5414 153462 5466
rect 153474 5414 153526 5466
rect 153538 5414 153590 5466
rect 153602 5414 153654 5466
rect 229544 5414 229596 5466
rect 229608 5414 229660 5466
rect 229672 5414 229724 5466
rect 229736 5414 229788 5466
rect 229800 5414 229852 5466
rect 39048 4870 39100 4922
rect 39112 4870 39164 4922
rect 39176 4870 39228 4922
rect 39240 4870 39292 4922
rect 39304 4870 39356 4922
rect 115246 4870 115298 4922
rect 115310 4870 115362 4922
rect 115374 4870 115426 4922
rect 115438 4870 115490 4922
rect 115502 4870 115554 4922
rect 191444 4870 191496 4922
rect 191508 4870 191560 4922
rect 191572 4870 191624 4922
rect 191636 4870 191688 4922
rect 191700 4870 191752 4922
rect 267642 4870 267694 4922
rect 267706 4870 267758 4922
rect 267770 4870 267822 4922
rect 267834 4870 267886 4922
rect 267898 4870 267950 4922
rect 77148 4326 77200 4378
rect 77212 4326 77264 4378
rect 77276 4326 77328 4378
rect 77340 4326 77392 4378
rect 77404 4326 77456 4378
rect 153346 4326 153398 4378
rect 153410 4326 153462 4378
rect 153474 4326 153526 4378
rect 153538 4326 153590 4378
rect 153602 4326 153654 4378
rect 229544 4326 229596 4378
rect 229608 4326 229660 4378
rect 229672 4326 229724 4378
rect 229736 4326 229788 4378
rect 229800 4326 229852 4378
rect 39048 3782 39100 3834
rect 39112 3782 39164 3834
rect 39176 3782 39228 3834
rect 39240 3782 39292 3834
rect 39304 3782 39356 3834
rect 115246 3782 115298 3834
rect 115310 3782 115362 3834
rect 115374 3782 115426 3834
rect 115438 3782 115490 3834
rect 115502 3782 115554 3834
rect 191444 3782 191496 3834
rect 191508 3782 191560 3834
rect 191572 3782 191624 3834
rect 191636 3782 191688 3834
rect 191700 3782 191752 3834
rect 267642 3782 267694 3834
rect 267706 3782 267758 3834
rect 267770 3782 267822 3834
rect 267834 3782 267886 3834
rect 267898 3782 267950 3834
rect 77148 3238 77200 3290
rect 77212 3238 77264 3290
rect 77276 3238 77328 3290
rect 77340 3238 77392 3290
rect 77404 3238 77456 3290
rect 153346 3238 153398 3290
rect 153410 3238 153462 3290
rect 153474 3238 153526 3290
rect 153538 3238 153590 3290
rect 153602 3238 153654 3290
rect 229544 3238 229596 3290
rect 229608 3238 229660 3290
rect 229672 3238 229724 3290
rect 229736 3238 229788 3290
rect 229800 3238 229852 3290
rect 39048 2694 39100 2746
rect 39112 2694 39164 2746
rect 39176 2694 39228 2746
rect 39240 2694 39292 2746
rect 39304 2694 39356 2746
rect 115246 2694 115298 2746
rect 115310 2694 115362 2746
rect 115374 2694 115426 2746
rect 115438 2694 115490 2746
rect 115502 2694 115554 2746
rect 191444 2694 191496 2746
rect 191508 2694 191560 2746
rect 191572 2694 191624 2746
rect 191636 2694 191688 2746
rect 191700 2694 191752 2746
rect 267642 2694 267694 2746
rect 267706 2694 267758 2746
rect 267770 2694 267822 2746
rect 267834 2694 267886 2746
rect 267898 2694 267950 2746
rect 149428 2592 149480 2644
rect 302240 2592 302292 2644
rect 77148 2150 77200 2202
rect 77212 2150 77264 2202
rect 77276 2150 77328 2202
rect 77340 2150 77392 2202
rect 77404 2150 77456 2202
rect 153346 2150 153398 2202
rect 153410 2150 153462 2202
rect 153474 2150 153526 2202
rect 153538 2150 153590 2202
rect 153602 2150 153654 2202
rect 229544 2150 229596 2202
rect 229608 2150 229660 2202
rect 229672 2150 229724 2202
rect 229736 2150 229788 2202
rect 229800 2150 229852 2202
<< metal2 >>
rect 1490 15314 1546 16000
rect 4526 15314 4582 16000
rect 7562 15314 7618 16000
rect 10690 15314 10746 16000
rect 1490 15286 1624 15314
rect 1490 15200 1546 15286
rect 1596 13530 1624 15286
rect 4526 15286 4660 15314
rect 4526 15200 4582 15286
rect 4632 13530 4660 15286
rect 7562 15286 7696 15314
rect 7562 15200 7618 15286
rect 7668 13530 7696 15286
rect 10690 15286 10824 15314
rect 10690 15200 10746 15286
rect 10796 13530 10824 15286
rect 13726 15200 13782 16000
rect 16762 15314 16818 16000
rect 19890 15314 19946 16000
rect 22926 15314 22982 16000
rect 25962 15314 26018 16000
rect 16762 15286 16896 15314
rect 16762 15200 16818 15286
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 10784 13524 10836 13530
rect 13740 13512 13768 15200
rect 16868 13530 16896 15286
rect 19890 15286 20024 15314
rect 19890 15200 19946 15286
rect 19996 13530 20024 15286
rect 22926 15286 23060 15314
rect 22926 15200 22982 15286
rect 23032 13530 23060 15286
rect 25962 15286 26096 15314
rect 25962 15200 26018 15286
rect 13820 13524 13872 13530
rect 13740 13484 13820 13512
rect 10784 13466 10836 13472
rect 13820 13466 13872 13472
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 4816 12102 4844 13262
rect 14292 12374 14320 13262
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 17052 12238 17080 13262
rect 20180 12918 20208 13262
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 23216 12782 23244 13262
rect 26068 12986 26096 15286
rect 29090 15200 29146 16000
rect 32126 15200 32182 16000
rect 35254 15314 35310 16000
rect 38290 15314 38346 16000
rect 35254 15286 35572 15314
rect 35254 15200 35310 15286
rect 29000 13796 29052 13802
rect 29000 13738 29052 13744
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27172 13462 27200 13670
rect 27448 13654 27752 13682
rect 27160 13456 27212 13462
rect 27160 13398 27212 13404
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 26988 12442 27016 13330
rect 27172 12714 27200 13398
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27264 13002 27292 13126
rect 27448 13002 27476 13654
rect 27724 13530 27752 13654
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27528 13252 27580 13258
rect 27528 13194 27580 13200
rect 27264 12974 27476 13002
rect 27344 12912 27396 12918
rect 27344 12854 27396 12860
rect 27160 12708 27212 12714
rect 27160 12650 27212 12656
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 26896 12186 26924 12242
rect 26896 12158 27200 12186
rect 27172 12102 27200 12158
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 27068 12096 27120 12102
rect 27068 12038 27120 12044
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27080 11218 27108 12038
rect 27068 11212 27120 11218
rect 27068 11154 27120 11160
rect 27356 9586 27384 12854
rect 27448 12238 27476 12974
rect 27436 12232 27488 12238
rect 27436 12174 27488 12180
rect 27540 10198 27568 13194
rect 27632 11150 27660 13466
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27724 11830 27752 13126
rect 29012 12918 29040 13738
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 28000 12102 28028 12786
rect 28080 12776 28132 12782
rect 28080 12718 28132 12724
rect 28092 12442 28120 12718
rect 28908 12640 28960 12646
rect 28908 12582 28960 12588
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 28816 12436 28868 12442
rect 28816 12378 28868 12384
rect 28092 12306 28120 12378
rect 28828 12322 28856 12378
rect 28736 12306 28856 12322
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 28724 12300 28856 12306
rect 28776 12294 28856 12300
rect 28724 12242 28776 12248
rect 27988 12096 28040 12102
rect 27988 12038 28040 12044
rect 27712 11824 27764 11830
rect 27712 11766 27764 11772
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 28000 11082 28028 12038
rect 28736 11830 28764 12242
rect 28920 12102 28948 12582
rect 29000 12300 29052 12306
rect 29000 12242 29052 12248
rect 28908 12096 28960 12102
rect 28908 12038 28960 12044
rect 29012 11830 29040 12242
rect 29104 11898 29132 15200
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30484 13410 30512 13466
rect 30392 13382 30512 13410
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29840 12782 29868 13262
rect 30196 13252 30248 13258
rect 30196 13194 30248 13200
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29828 12776 29880 12782
rect 29828 12718 29880 12724
rect 30104 12776 30156 12782
rect 30104 12718 30156 12724
rect 29656 12434 29684 12718
rect 29656 12406 29776 12434
rect 29552 12300 29604 12306
rect 29552 12242 29604 12248
rect 29368 12232 29420 12238
rect 29366 12200 29368 12208
rect 29420 12200 29422 12208
rect 29366 12134 29422 12144
rect 29460 12164 29512 12170
rect 29460 12106 29512 12112
rect 29472 11898 29500 12106
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 29460 11892 29512 11898
rect 29460 11834 29512 11840
rect 28724 11824 28776 11830
rect 28724 11766 28776 11772
rect 29000 11824 29052 11830
rect 29000 11766 29052 11772
rect 29564 11762 29592 12242
rect 29552 11756 29604 11762
rect 29552 11698 29604 11704
rect 28908 11688 28960 11694
rect 28908 11630 28960 11636
rect 28448 11552 28500 11558
rect 28448 11494 28500 11500
rect 27988 11076 28040 11082
rect 27988 11018 28040 11024
rect 28460 10674 28488 11494
rect 28920 11286 28948 11630
rect 28908 11280 28960 11286
rect 28908 11222 28960 11228
rect 29564 11218 29592 11698
rect 29460 11212 29512 11218
rect 29460 11154 29512 11160
rect 29552 11212 29604 11218
rect 29552 11154 29604 11160
rect 28448 10668 28500 10674
rect 28448 10610 28500 10616
rect 27528 10192 27580 10198
rect 27528 10134 27580 10140
rect 29472 10062 29500 11154
rect 29748 10742 29776 12406
rect 29828 12164 29880 12170
rect 29828 12106 29880 12112
rect 29840 10810 29868 12106
rect 30012 11824 30064 11830
rect 30012 11766 30064 11772
rect 29920 11688 29972 11694
rect 29920 11630 29972 11636
rect 29932 11354 29960 11630
rect 30024 11354 30052 11766
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 30012 11348 30064 11354
rect 30012 11290 30064 11296
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 29828 10804 29880 10810
rect 29828 10746 29880 10752
rect 29736 10736 29788 10742
rect 29736 10678 29788 10684
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 29932 9450 29960 11018
rect 30116 10266 30144 12718
rect 30208 10742 30236 13194
rect 30392 12918 30420 13382
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 30392 11370 30420 12854
rect 30484 12434 30512 13126
rect 31576 12912 31628 12918
rect 31576 12854 31628 12860
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 30484 12406 30604 12434
rect 30392 11342 30512 11370
rect 30484 10810 30512 11342
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30196 10736 30248 10742
rect 30196 10678 30248 10684
rect 30104 10260 30156 10266
rect 30104 10202 30156 10208
rect 30576 9518 30604 12406
rect 31404 12208 31432 12582
rect 30746 12200 30802 12208
rect 31390 12200 31446 12208
rect 30746 12134 30802 12144
rect 31208 12164 31260 12170
rect 30760 10810 30788 12134
rect 31390 12134 31446 12144
rect 31208 12106 31260 12112
rect 31116 12096 31168 12102
rect 31116 12038 31168 12044
rect 30932 11892 30984 11898
rect 30932 11834 30984 11840
rect 30748 10804 30800 10810
rect 30748 10746 30800 10752
rect 30944 10062 30972 11834
rect 31128 11626 31156 12038
rect 31116 11620 31168 11626
rect 31116 11562 31168 11568
rect 30932 10056 30984 10062
rect 30932 9998 30984 10004
rect 31220 9654 31248 12106
rect 31392 11552 31444 11558
rect 31392 11494 31444 11500
rect 31404 11218 31432 11494
rect 31392 11212 31444 11218
rect 31392 11154 31444 11160
rect 31588 10198 31616 12854
rect 32036 12164 32088 12170
rect 32036 12106 32088 12112
rect 32048 11830 32076 12106
rect 32036 11824 32088 11830
rect 32036 11766 32088 11772
rect 31668 11076 31720 11082
rect 31668 11018 31720 11024
rect 31760 11076 31812 11082
rect 31760 11018 31812 11024
rect 31680 10266 31708 11018
rect 31772 10742 31800 11018
rect 31852 11008 31904 11014
rect 31852 10950 31904 10956
rect 31864 10742 31892 10950
rect 31760 10736 31812 10742
rect 31760 10678 31812 10684
rect 31852 10736 31904 10742
rect 31852 10678 31904 10684
rect 32140 10266 32168 15200
rect 32956 13796 33008 13802
rect 32956 13738 33008 13744
rect 32404 13320 32456 13326
rect 32404 13262 32456 13268
rect 32220 12980 32272 12986
rect 32220 12922 32272 12928
rect 32232 11898 32260 12922
rect 32416 12646 32444 13262
rect 32680 13252 32732 13258
rect 32680 13194 32732 13200
rect 32404 12640 32456 12646
rect 32404 12582 32456 12588
rect 32588 12436 32640 12442
rect 32588 12378 32640 12384
rect 32312 12096 32364 12102
rect 32312 12038 32364 12044
rect 32220 11892 32272 11898
rect 32220 11834 32272 11840
rect 32232 11150 32260 11834
rect 32324 11218 32352 12038
rect 32404 11756 32456 11762
rect 32404 11698 32456 11704
rect 32416 11354 32444 11698
rect 32600 11694 32628 12378
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32404 11348 32456 11354
rect 32404 11290 32456 11296
rect 32600 11218 32628 11630
rect 32312 11212 32364 11218
rect 32312 11154 32364 11160
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32692 10810 32720 13194
rect 32968 12102 32996 13738
rect 33784 13320 33836 13326
rect 33784 13262 33836 13268
rect 33600 13184 33652 13190
rect 33600 13126 33652 13132
rect 33048 12776 33100 12782
rect 33048 12718 33100 12724
rect 33416 12776 33468 12782
rect 33416 12718 33468 12724
rect 32956 12096 33008 12102
rect 32956 12038 33008 12044
rect 32956 11552 33008 11558
rect 32956 11494 33008 11500
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32968 10674 32996 11494
rect 33060 10810 33088 12718
rect 33324 11348 33376 11354
rect 33324 11290 33376 11296
rect 33048 10804 33100 10810
rect 33048 10746 33100 10752
rect 32956 10668 33008 10674
rect 32956 10610 33008 10616
rect 33336 10266 33364 11290
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 32128 10260 32180 10266
rect 32128 10202 32180 10208
rect 33324 10260 33376 10266
rect 33324 10202 33376 10208
rect 31576 10192 31628 10198
rect 31576 10134 31628 10140
rect 33428 10062 33456 12718
rect 33612 11354 33640 13126
rect 33692 12844 33744 12850
rect 33692 12786 33744 12792
rect 33600 11348 33652 11354
rect 33600 11290 33652 11296
rect 33704 10062 33732 12786
rect 33796 11898 33824 13262
rect 34520 13252 34572 13258
rect 34520 13194 34572 13200
rect 34152 13184 34204 13190
rect 34152 13126 34204 13132
rect 34336 13184 34388 13190
rect 34336 13126 34388 13132
rect 34164 12986 34192 13126
rect 34152 12980 34204 12986
rect 34152 12922 34204 12928
rect 34164 12832 34192 12922
rect 34072 12804 34192 12832
rect 33784 11892 33836 11898
rect 33784 11834 33836 11840
rect 34072 11694 34100 12804
rect 34348 12782 34376 13126
rect 34428 12912 34480 12918
rect 34428 12854 34480 12860
rect 34336 12776 34388 12782
rect 34336 12718 34388 12724
rect 34152 12640 34204 12646
rect 34152 12582 34204 12588
rect 34164 12238 34192 12582
rect 34152 12232 34204 12238
rect 34152 12174 34204 12180
rect 34440 11898 34468 12854
rect 34532 12442 34560 13194
rect 35544 12986 35572 15286
rect 38290 15286 38424 15314
rect 38290 15200 38346 15286
rect 36544 13728 36596 13734
rect 36544 13670 36596 13676
rect 36556 13530 36584 13670
rect 36544 13524 36596 13530
rect 36544 13466 36596 13472
rect 35992 13252 36044 13258
rect 35992 13194 36044 13200
rect 37832 13252 37884 13258
rect 37832 13194 37884 13200
rect 35532 12980 35584 12986
rect 35532 12922 35584 12928
rect 34888 12776 34940 12782
rect 34888 12718 34940 12724
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 34520 12436 34572 12442
rect 34520 12378 34572 12384
rect 34900 12374 34928 12718
rect 34888 12368 34940 12374
rect 34888 12310 34940 12316
rect 35360 12238 35388 12718
rect 36004 12442 36032 13194
rect 37464 13184 37516 13190
rect 37464 13126 37516 13132
rect 37476 12918 37504 13126
rect 37464 12912 37516 12918
rect 37464 12854 37516 12860
rect 37844 12442 37872 13194
rect 38016 12640 38068 12646
rect 38016 12582 38068 12588
rect 35992 12436 36044 12442
rect 35992 12378 36044 12384
rect 37832 12436 37884 12442
rect 37832 12378 37884 12384
rect 38028 12238 38056 12582
rect 34704 12232 34756 12238
rect 34704 12174 34756 12180
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 38016 12232 38068 12238
rect 38016 12174 38068 12180
rect 34428 11892 34480 11898
rect 34428 11834 34480 11840
rect 34716 11762 34744 12174
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 34704 11756 34756 11762
rect 34704 11698 34756 11704
rect 34060 11688 34112 11694
rect 34060 11630 34112 11636
rect 34716 11150 34744 11698
rect 36464 11286 36492 12038
rect 38396 11898 38424 15286
rect 41326 15200 41382 16000
rect 44454 15314 44510 16000
rect 47490 15314 47546 16000
rect 44454 15286 44588 15314
rect 44454 15200 44510 15286
rect 39048 13628 39356 13636
rect 39048 13626 39054 13628
rect 39110 13626 39134 13628
rect 39190 13626 39214 13628
rect 39270 13626 39294 13628
rect 39350 13626 39356 13628
rect 39110 13574 39112 13626
rect 39292 13574 39294 13626
rect 39048 13572 39054 13574
rect 39110 13572 39134 13574
rect 39190 13572 39214 13574
rect 39270 13572 39294 13574
rect 39350 13572 39356 13574
rect 39048 13562 39356 13572
rect 38936 13320 38988 13326
rect 38936 13262 38988 13268
rect 38948 12442 38976 13262
rect 40408 13252 40460 13258
rect 40408 13194 40460 13200
rect 39304 13184 39356 13190
rect 39304 13126 39356 13132
rect 39948 13184 40000 13190
rect 39948 13126 40000 13132
rect 39316 12850 39344 13126
rect 39672 12912 39724 12918
rect 39672 12854 39724 12860
rect 39304 12844 39356 12850
rect 39304 12786 39356 12792
rect 39396 12776 39448 12782
rect 39396 12718 39448 12724
rect 39048 12540 39356 12548
rect 39048 12538 39054 12540
rect 39110 12538 39134 12540
rect 39190 12538 39214 12540
rect 39270 12538 39294 12540
rect 39350 12538 39356 12540
rect 39110 12486 39112 12538
rect 39292 12486 39294 12538
rect 39048 12484 39054 12486
rect 39110 12484 39134 12486
rect 39190 12484 39214 12486
rect 39270 12484 39294 12486
rect 39350 12484 39356 12486
rect 39048 12474 39356 12484
rect 39408 12442 39436 12718
rect 38936 12436 38988 12442
rect 38936 12378 38988 12384
rect 39396 12436 39448 12442
rect 39396 12378 39448 12384
rect 38384 11892 38436 11898
rect 38384 11834 38436 11840
rect 39580 11892 39632 11898
rect 39684 11880 39712 12854
rect 39960 11898 39988 13126
rect 40316 12232 40368 12238
rect 40316 12174 40368 12180
rect 39632 11852 39712 11880
rect 39948 11892 40000 11898
rect 39580 11834 39632 11840
rect 39948 11834 40000 11840
rect 40328 11762 40356 12174
rect 40316 11756 40368 11762
rect 40316 11698 40368 11704
rect 39048 11452 39356 11460
rect 39048 11450 39054 11452
rect 39110 11450 39134 11452
rect 39190 11450 39214 11452
rect 39270 11450 39294 11452
rect 39350 11450 39356 11452
rect 39110 11398 39112 11450
rect 39292 11398 39294 11450
rect 39048 11396 39054 11398
rect 39110 11396 39134 11398
rect 39190 11396 39214 11398
rect 39270 11396 39294 11398
rect 39350 11396 39356 11398
rect 39048 11386 39356 11396
rect 40420 11354 40448 13194
rect 41052 12912 41104 12918
rect 41052 12854 41104 12860
rect 40960 12776 41012 12782
rect 40960 12718 41012 12724
rect 40972 12442 41000 12718
rect 40960 12436 41012 12442
rect 40960 12378 41012 12384
rect 40972 12306 41000 12378
rect 40960 12300 41012 12306
rect 40960 12242 41012 12248
rect 40592 12232 40644 12238
rect 40590 12200 40592 12208
rect 40644 12200 40646 12208
rect 40590 12134 40646 12144
rect 40500 12096 40552 12102
rect 40500 12038 40552 12044
rect 40684 12096 40736 12102
rect 40684 12038 40736 12044
rect 40408 11348 40460 11354
rect 40408 11290 40460 11296
rect 36452 11280 36504 11286
rect 36452 11222 36504 11228
rect 40512 11150 40540 12038
rect 40696 11830 40724 12038
rect 40684 11824 40736 11830
rect 40684 11766 40736 11772
rect 40972 11694 41000 12242
rect 40960 11688 41012 11694
rect 40960 11630 41012 11636
rect 41064 11354 41092 12854
rect 41236 12640 41288 12646
rect 41236 12582 41288 12588
rect 41248 11830 41276 12582
rect 41236 11824 41288 11830
rect 41236 11766 41288 11772
rect 41052 11348 41104 11354
rect 41052 11290 41104 11296
rect 41340 11286 41368 15200
rect 42524 13728 42576 13734
rect 42524 13670 42576 13676
rect 42536 13326 42564 13670
rect 44180 13456 44232 13462
rect 44364 13456 44416 13462
rect 44232 13416 44364 13444
rect 44180 13398 44232 13404
rect 44364 13398 44416 13404
rect 42524 13320 42576 13326
rect 42524 13262 42576 13268
rect 44272 13320 44324 13326
rect 44272 13262 44324 13268
rect 41420 13252 41472 13258
rect 41420 13194 41472 13200
rect 42892 13252 42944 13258
rect 42892 13194 42944 13200
rect 43260 13252 43312 13258
rect 43260 13194 43312 13200
rect 41432 11898 41460 13194
rect 42432 13184 42484 13190
rect 42432 13126 42484 13132
rect 41512 12844 41564 12850
rect 41512 12786 41564 12792
rect 41420 11892 41472 11898
rect 41420 11834 41472 11840
rect 41420 11688 41472 11694
rect 41524 11676 41552 12786
rect 41788 12640 41840 12646
rect 41788 12582 41840 12588
rect 41800 12170 41828 12582
rect 42444 12208 42472 13126
rect 42800 12640 42852 12646
rect 42800 12582 42852 12588
rect 42430 12200 42486 12208
rect 41604 12164 41656 12170
rect 41604 12106 41656 12112
rect 41788 12164 41840 12170
rect 42430 12134 42486 12144
rect 41788 12106 41840 12112
rect 41472 11648 41552 11676
rect 41420 11630 41472 11636
rect 41328 11280 41380 11286
rect 41328 11222 41380 11228
rect 41432 11150 41460 11630
rect 41616 11354 41644 12106
rect 41604 11348 41656 11354
rect 41604 11290 41656 11296
rect 42444 11150 42472 12134
rect 42812 11762 42840 12582
rect 42904 11898 42932 13194
rect 43272 12986 43300 13194
rect 44284 12986 44312 13262
rect 44560 12986 44588 15286
rect 47490 15286 47624 15314
rect 47490 15200 47546 15286
rect 46204 13796 46256 13802
rect 46204 13738 46256 13744
rect 46216 13530 46244 13738
rect 47596 13530 47624 15286
rect 50526 15200 50582 16000
rect 53654 15200 53710 16000
rect 56690 15200 56746 16000
rect 59818 15200 59874 16000
rect 62854 15314 62910 16000
rect 65890 15314 65946 16000
rect 69018 15314 69074 16000
rect 72054 15314 72110 16000
rect 62854 15286 63080 15314
rect 62854 15200 62910 15286
rect 47860 13728 47912 13734
rect 47860 13670 47912 13676
rect 46204 13524 46256 13530
rect 46204 13466 46256 13472
rect 47584 13524 47636 13530
rect 47584 13466 47636 13472
rect 45560 13388 45612 13394
rect 45560 13330 45612 13336
rect 45008 13184 45060 13190
rect 45008 13126 45060 13132
rect 45376 13184 45428 13190
rect 45376 13126 45428 13132
rect 43260 12980 43312 12986
rect 43260 12922 43312 12928
rect 44272 12980 44324 12986
rect 44272 12922 44324 12928
rect 44548 12980 44600 12986
rect 44548 12922 44600 12928
rect 42984 12912 43036 12918
rect 42984 12854 43036 12860
rect 42892 11892 42944 11898
rect 42892 11834 42944 11840
rect 42996 11762 43024 12854
rect 43088 12838 43300 12866
rect 43088 12782 43116 12838
rect 43076 12776 43128 12782
rect 43076 12718 43128 12724
rect 43168 12776 43220 12782
rect 43168 12718 43220 12724
rect 43180 12442 43208 12718
rect 43272 12646 43300 12838
rect 43812 12776 43864 12782
rect 43812 12718 43864 12724
rect 43824 12646 43852 12718
rect 43260 12640 43312 12646
rect 43260 12582 43312 12588
rect 43812 12640 43864 12646
rect 43812 12582 43864 12588
rect 43824 12442 43852 12582
rect 43168 12436 43220 12442
rect 43168 12378 43220 12384
rect 43812 12436 43864 12442
rect 43812 12378 43864 12384
rect 43720 12368 43772 12374
rect 43720 12310 43772 12316
rect 43732 12238 43760 12310
rect 43720 12232 43772 12238
rect 43720 12174 43772 12180
rect 42800 11756 42852 11762
rect 42800 11698 42852 11704
rect 42984 11756 43036 11762
rect 42984 11698 43036 11704
rect 45020 11218 45048 13126
rect 45388 12850 45416 13126
rect 45376 12844 45428 12850
rect 45376 12786 45428 12792
rect 45468 12776 45520 12782
rect 45572 12764 45600 13330
rect 47872 13258 47900 13670
rect 50540 13530 50568 15200
rect 51632 13728 51684 13734
rect 51632 13670 51684 13676
rect 50528 13524 50580 13530
rect 50528 13466 50580 13472
rect 51644 13394 51672 13670
rect 53012 13524 53064 13530
rect 53012 13466 53064 13472
rect 51632 13388 51684 13394
rect 51632 13330 51684 13336
rect 51356 13320 51408 13326
rect 51356 13262 51408 13268
rect 47860 13252 47912 13258
rect 47860 13194 47912 13200
rect 51368 12782 51396 13262
rect 45520 12736 45600 12764
rect 51356 12776 51408 12782
rect 45468 12718 45520 12724
rect 51356 12718 51408 12724
rect 52644 12164 52696 12170
rect 52644 12106 52696 12112
rect 52656 11898 52684 12106
rect 52644 11892 52696 11898
rect 52644 11834 52696 11840
rect 53024 11762 53052 13466
rect 53288 13252 53340 13258
rect 53288 13194 53340 13200
rect 53300 12986 53328 13194
rect 53288 12980 53340 12986
rect 53288 12922 53340 12928
rect 53104 12640 53156 12646
rect 53104 12582 53156 12588
rect 53116 12170 53144 12582
rect 53104 12164 53156 12170
rect 53104 12106 53156 12112
rect 53668 11898 53696 15200
rect 54116 13728 54168 13734
rect 54116 13670 54168 13676
rect 53748 12844 53800 12850
rect 53748 12786 53800 12792
rect 54024 12844 54076 12850
rect 54024 12786 54076 12792
rect 53760 12322 53788 12786
rect 54036 12442 54064 12786
rect 54128 12782 54156 13670
rect 55588 13524 55640 13530
rect 55588 13466 55640 13472
rect 55600 13326 55628 13466
rect 54392 13320 54444 13326
rect 54392 13262 54444 13268
rect 54760 13320 54812 13326
rect 54760 13262 54812 13268
rect 55588 13320 55640 13326
rect 55588 13262 55640 13268
rect 54116 12776 54168 12782
rect 54116 12718 54168 12724
rect 54128 12646 54156 12718
rect 54116 12640 54168 12646
rect 54116 12582 54168 12588
rect 54024 12436 54076 12442
rect 54024 12378 54076 12384
rect 53760 12306 53880 12322
rect 53760 12300 53892 12306
rect 53760 12294 53840 12300
rect 53656 11892 53708 11898
rect 53656 11834 53708 11840
rect 53760 11830 53788 12294
rect 53840 12242 53892 12248
rect 54404 11898 54432 13262
rect 54668 13184 54720 13190
rect 54668 13126 54720 13132
rect 54680 12986 54708 13126
rect 54668 12980 54720 12986
rect 54668 12922 54720 12928
rect 54392 11892 54444 11898
rect 54392 11834 54444 11840
rect 53748 11824 53800 11830
rect 53748 11766 53800 11772
rect 53012 11756 53064 11762
rect 53012 11698 53064 11704
rect 54680 11694 54708 12922
rect 54772 12850 54800 13262
rect 55864 13252 55916 13258
rect 55864 13194 55916 13200
rect 56600 13252 56652 13258
rect 56600 13194 56652 13200
rect 55876 12986 55904 13194
rect 55864 12980 55916 12986
rect 55864 12922 55916 12928
rect 55496 12912 55548 12918
rect 55496 12854 55548 12860
rect 54760 12844 54812 12850
rect 54760 12786 54812 12792
rect 55036 12776 55088 12782
rect 55036 12718 55088 12724
rect 54668 11688 54720 11694
rect 54668 11630 54720 11636
rect 55048 11354 55076 12718
rect 55508 12442 55536 12854
rect 55588 12640 55640 12646
rect 55588 12582 55640 12588
rect 56324 12640 56376 12646
rect 56324 12582 56376 12588
rect 56508 12640 56560 12646
rect 56508 12582 56560 12588
rect 55496 12436 55548 12442
rect 55496 12378 55548 12384
rect 55312 12232 55364 12238
rect 55312 12174 55364 12180
rect 55324 11898 55352 12174
rect 55312 11892 55364 11898
rect 55312 11834 55364 11840
rect 55600 11694 55628 12582
rect 56336 12434 56364 12582
rect 56336 12406 56456 12434
rect 56428 12306 56456 12406
rect 56416 12300 56468 12306
rect 56416 12242 56468 12248
rect 56520 12238 56548 12582
rect 56508 12232 56560 12238
rect 56508 12174 56560 12180
rect 55864 12096 55916 12102
rect 55864 12038 55916 12044
rect 56048 12096 56100 12102
rect 56048 12038 56100 12044
rect 55876 11694 55904 12038
rect 55588 11688 55640 11694
rect 55588 11630 55640 11636
rect 55864 11688 55916 11694
rect 55864 11630 55916 11636
rect 56060 11626 56088 12038
rect 56612 11898 56640 13194
rect 56704 12442 56732 15200
rect 57888 13524 57940 13530
rect 57888 13466 57940 13472
rect 57900 13326 57928 13466
rect 59832 13462 59860 15200
rect 61752 13524 61804 13530
rect 61752 13466 61804 13472
rect 59820 13456 59872 13462
rect 59820 13398 59872 13404
rect 57888 13320 57940 13326
rect 57888 13262 57940 13268
rect 60648 13320 60700 13326
rect 60648 13262 60700 13268
rect 57704 13252 57756 13258
rect 57704 13194 57756 13200
rect 58624 13252 58676 13258
rect 58624 13194 58676 13200
rect 57336 13184 57388 13190
rect 57336 13126 57388 13132
rect 57348 12918 57376 13126
rect 57336 12912 57388 12918
rect 57336 12854 57388 12860
rect 57244 12640 57296 12646
rect 57244 12582 57296 12588
rect 56692 12436 56744 12442
rect 56692 12378 56744 12384
rect 56600 11892 56652 11898
rect 56600 11834 56652 11840
rect 56048 11620 56100 11626
rect 56048 11562 56100 11568
rect 55496 11552 55548 11558
rect 55496 11494 55548 11500
rect 55036 11348 55088 11354
rect 55036 11290 55088 11296
rect 45008 11212 45060 11218
rect 45008 11154 45060 11160
rect 55508 11150 55536 11494
rect 57256 11150 57284 12582
rect 57348 12102 57376 12854
rect 57428 12844 57480 12850
rect 57428 12786 57480 12792
rect 57336 12096 57388 12102
rect 57336 12038 57388 12044
rect 57440 11830 57468 12786
rect 57428 11824 57480 11830
rect 57428 11766 57480 11772
rect 57716 11354 57744 13194
rect 57980 12980 58032 12986
rect 57980 12922 58032 12928
rect 57992 12442 58020 12922
rect 57980 12436 58032 12442
rect 57980 12378 58032 12384
rect 58636 11898 58664 13194
rect 59636 13184 59688 13190
rect 59636 13126 59688 13132
rect 59648 12986 59676 13126
rect 59636 12980 59688 12986
rect 59636 12922 59688 12928
rect 60660 12918 60688 13262
rect 61488 13258 61700 13274
rect 61764 13258 61792 13466
rect 63052 13462 63080 15286
rect 65890 15286 66024 15314
rect 65890 15200 65946 15286
rect 63408 13796 63460 13802
rect 63408 13738 63460 13744
rect 63420 13530 63448 13738
rect 63408 13524 63460 13530
rect 63408 13466 63460 13472
rect 63040 13456 63092 13462
rect 63040 13398 63092 13404
rect 61476 13252 61700 13258
rect 61528 13246 61700 13252
rect 61476 13194 61528 13200
rect 61672 13190 61700 13246
rect 61752 13252 61804 13258
rect 61752 13194 61804 13200
rect 65996 13190 66024 15286
rect 69018 15286 69152 15314
rect 69018 15200 69074 15286
rect 66168 13728 66220 13734
rect 66168 13670 66220 13676
rect 66180 13326 66208 13670
rect 66168 13320 66220 13326
rect 66168 13262 66220 13268
rect 69124 13190 69152 15286
rect 72054 15286 72188 15314
rect 72054 15200 72110 15286
rect 69296 13796 69348 13802
rect 69296 13738 69348 13744
rect 69308 13326 69336 13738
rect 69296 13320 69348 13326
rect 69296 13262 69348 13268
rect 61660 13184 61712 13190
rect 61660 13126 61712 13132
rect 65892 13184 65944 13190
rect 65892 13126 65944 13132
rect 65984 13184 66036 13190
rect 65984 13126 66036 13132
rect 69112 13184 69164 13190
rect 69112 13126 69164 13132
rect 65904 12918 65932 13126
rect 72160 12986 72188 15286
rect 75090 15200 75146 16000
rect 78218 15314 78274 16000
rect 81254 15314 81310 16000
rect 78218 15286 78536 15314
rect 78218 15200 78274 15286
rect 72424 13728 72476 13734
rect 72424 13670 72476 13676
rect 73896 13728 73948 13734
rect 73896 13670 73948 13676
rect 72436 13190 72464 13670
rect 72700 13388 72752 13394
rect 72700 13330 72752 13336
rect 72332 13184 72384 13190
rect 72332 13126 72384 13132
rect 72424 13184 72476 13190
rect 72424 13126 72476 13132
rect 72344 12986 72372 13126
rect 72148 12980 72200 12986
rect 72148 12922 72200 12928
rect 72332 12980 72384 12986
rect 72332 12922 72384 12928
rect 60648 12912 60700 12918
rect 60648 12854 60700 12860
rect 65892 12912 65944 12918
rect 65892 12854 65944 12860
rect 72712 12646 72740 13330
rect 73908 13258 73936 13670
rect 73896 13252 73948 13258
rect 73896 13194 73948 13200
rect 74724 12980 74776 12986
rect 74724 12922 74776 12928
rect 72700 12640 72752 12646
rect 72700 12582 72752 12588
rect 58624 11892 58676 11898
rect 58624 11834 58676 11840
rect 57704 11348 57756 11354
rect 57704 11290 57756 11296
rect 74736 11150 74764 12922
rect 74816 12844 74868 12850
rect 74816 12786 74868 12792
rect 74828 12306 74856 12786
rect 75000 12640 75052 12646
rect 75000 12582 75052 12588
rect 74816 12300 74868 12306
rect 74816 12242 74868 12248
rect 75012 11694 75040 12582
rect 75104 12442 75132 15200
rect 75368 13796 75420 13802
rect 75368 13738 75420 13744
rect 76012 13796 76064 13802
rect 76012 13738 76064 13744
rect 75380 13462 75408 13738
rect 75368 13456 75420 13462
rect 75368 13398 75420 13404
rect 75644 13456 75696 13462
rect 75644 13398 75696 13404
rect 75184 13252 75236 13258
rect 75184 13194 75236 13200
rect 75196 12646 75224 13194
rect 75460 12844 75512 12850
rect 75460 12786 75512 12792
rect 75184 12640 75236 12646
rect 75184 12582 75236 12588
rect 75092 12436 75144 12442
rect 75092 12378 75144 12384
rect 75472 11898 75500 12786
rect 75656 11898 75684 13398
rect 76024 12374 76052 13738
rect 76380 13728 76432 13734
rect 76380 13670 76432 13676
rect 76012 12368 76064 12374
rect 76012 12310 76064 12316
rect 75460 11892 75512 11898
rect 75460 11834 75512 11840
rect 75644 11892 75696 11898
rect 75644 11834 75696 11840
rect 76024 11762 76052 12310
rect 76288 12096 76340 12102
rect 76288 12038 76340 12044
rect 76300 11762 76328 12038
rect 76012 11756 76064 11762
rect 76012 11698 76064 11704
rect 76288 11756 76340 11762
rect 76288 11698 76340 11704
rect 75000 11688 75052 11694
rect 75000 11630 75052 11636
rect 76392 11354 76420 13670
rect 78404 13320 78456 13326
rect 78404 13262 78456 13268
rect 76472 13252 76524 13258
rect 76472 13194 76524 13200
rect 76484 11898 76512 13194
rect 77944 13184 77996 13190
rect 77944 13126 77996 13132
rect 77148 13084 77456 13092
rect 77148 13082 77154 13084
rect 77210 13082 77234 13084
rect 77290 13082 77314 13084
rect 77370 13082 77394 13084
rect 77450 13082 77456 13084
rect 77210 13030 77212 13082
rect 77392 13030 77394 13082
rect 77148 13028 77154 13030
rect 77210 13028 77234 13030
rect 77290 13028 77314 13030
rect 77370 13028 77394 13030
rect 77450 13028 77456 13030
rect 77148 13018 77456 13028
rect 77852 12708 77904 12714
rect 77852 12650 77904 12656
rect 77208 12640 77260 12646
rect 77208 12582 77260 12588
rect 77220 12374 77248 12582
rect 77208 12368 77260 12374
rect 77208 12310 77260 12316
rect 76932 12300 76984 12306
rect 76932 12242 76984 12248
rect 76472 11892 76524 11898
rect 76472 11834 76524 11840
rect 76944 11694 76972 12242
rect 77148 11996 77456 12004
rect 77148 11994 77154 11996
rect 77210 11994 77234 11996
rect 77290 11994 77314 11996
rect 77370 11994 77394 11996
rect 77450 11994 77456 11996
rect 77210 11942 77212 11994
rect 77392 11942 77394 11994
rect 77148 11940 77154 11942
rect 77210 11940 77234 11942
rect 77290 11940 77314 11942
rect 77370 11940 77394 11942
rect 77450 11940 77456 11942
rect 77148 11930 77456 11940
rect 77864 11898 77892 12650
rect 77956 12238 77984 13126
rect 78416 12918 78444 13262
rect 78404 12912 78456 12918
rect 78404 12854 78456 12860
rect 78128 12708 78180 12714
rect 78128 12650 78180 12656
rect 78140 12306 78168 12650
rect 78404 12368 78456 12374
rect 78404 12310 78456 12316
rect 78128 12300 78180 12306
rect 78128 12242 78180 12248
rect 77944 12232 77996 12238
rect 77944 12174 77996 12180
rect 77852 11892 77904 11898
rect 77852 11834 77904 11840
rect 76932 11688 76984 11694
rect 76932 11630 76984 11636
rect 76380 11348 76432 11354
rect 76380 11290 76432 11296
rect 78416 11150 78444 12310
rect 78508 11898 78536 15286
rect 81254 15286 81388 15314
rect 81254 15200 81310 15286
rect 81360 13410 81388 15286
rect 84290 15200 84346 16000
rect 87418 15200 87474 16000
rect 90454 15200 90510 16000
rect 93582 15314 93638 16000
rect 96618 15314 96674 16000
rect 93582 15286 93808 15314
rect 93582 15200 93638 15286
rect 83096 13728 83148 13734
rect 83096 13670 83148 13676
rect 80244 13388 80296 13394
rect 81360 13382 81480 13410
rect 80244 13330 80296 13336
rect 79980 13258 80100 13274
rect 78772 13252 78824 13258
rect 78772 13194 78824 13200
rect 79324 13252 79376 13258
rect 79324 13194 79376 13200
rect 79980 13252 80112 13258
rect 79980 13246 80060 13252
rect 78588 12776 78640 12782
rect 78588 12718 78640 12724
rect 78600 12238 78628 12718
rect 78588 12232 78640 12238
rect 78588 12174 78640 12180
rect 78496 11892 78548 11898
rect 78496 11834 78548 11840
rect 78600 11762 78628 12174
rect 78588 11756 78640 11762
rect 78588 11698 78640 11704
rect 78784 11354 78812 13194
rect 79336 12442 79364 13194
rect 79980 12866 80008 13246
rect 80060 13194 80112 13200
rect 79704 12850 80008 12866
rect 79692 12844 80008 12850
rect 79744 12838 80008 12844
rect 79692 12786 79744 12792
rect 79324 12436 79376 12442
rect 79324 12378 79376 12384
rect 80256 12102 80284 13330
rect 81452 13326 81480 13382
rect 81624 13388 81676 13394
rect 81624 13330 81676 13336
rect 81440 13320 81492 13326
rect 81440 13262 81492 13268
rect 80796 13184 80848 13190
rect 80796 13126 80848 13132
rect 81440 13184 81492 13190
rect 81440 13126 81492 13132
rect 80520 12912 80572 12918
rect 80520 12854 80572 12860
rect 80532 12442 80560 12854
rect 80808 12782 80836 13126
rect 80796 12776 80848 12782
rect 80796 12718 80848 12724
rect 81452 12714 81480 13126
rect 81440 12708 81492 12714
rect 81440 12650 81492 12656
rect 80520 12436 80572 12442
rect 80520 12378 80572 12384
rect 81452 12306 81480 12650
rect 81636 12646 81664 13330
rect 83108 13326 83136 13670
rect 83096 13320 83148 13326
rect 83096 13262 83148 13268
rect 83924 13320 83976 13326
rect 83924 13262 83976 13268
rect 83832 13252 83884 13258
rect 83832 13194 83884 13200
rect 82912 13184 82964 13190
rect 82912 13126 82964 13132
rect 82924 12918 82952 13126
rect 82912 12912 82964 12918
rect 82912 12854 82964 12860
rect 81624 12640 81676 12646
rect 81624 12582 81676 12588
rect 81440 12300 81492 12306
rect 81440 12242 81492 12248
rect 80244 12096 80296 12102
rect 80244 12038 80296 12044
rect 81452 11762 81480 12242
rect 81440 11756 81492 11762
rect 81440 11698 81492 11704
rect 78772 11348 78824 11354
rect 78772 11290 78824 11296
rect 34704 11144 34756 11150
rect 34704 11086 34756 11092
rect 40500 11144 40552 11150
rect 40500 11086 40552 11092
rect 41420 11144 41472 11150
rect 41420 11086 41472 11092
rect 42432 11144 42484 11150
rect 42432 11086 42484 11092
rect 55496 11144 55548 11150
rect 55496 11086 55548 11092
rect 57244 11144 57296 11150
rect 57244 11086 57296 11092
rect 74724 11144 74776 11150
rect 74724 11086 74776 11092
rect 78404 11144 78456 11150
rect 78404 11086 78456 11092
rect 81636 11082 81664 12582
rect 83844 12238 83872 13194
rect 83936 13190 83964 13262
rect 83924 13184 83976 13190
rect 83924 13126 83976 13132
rect 83936 12986 83964 13126
rect 83924 12980 83976 12986
rect 83924 12922 83976 12928
rect 83832 12232 83884 12238
rect 83832 12174 83884 12180
rect 84016 12096 84068 12102
rect 84016 12038 84068 12044
rect 84028 11694 84056 12038
rect 84304 11898 84332 15200
rect 86408 13728 86460 13734
rect 86408 13670 86460 13676
rect 84476 13252 84528 13258
rect 84476 13194 84528 13200
rect 85488 13252 85540 13258
rect 85488 13194 85540 13200
rect 84292 11892 84344 11898
rect 84292 11834 84344 11840
rect 84016 11688 84068 11694
rect 84016 11630 84068 11636
rect 84488 11354 84516 13194
rect 84844 12776 84896 12782
rect 84844 12718 84896 12724
rect 84660 12300 84712 12306
rect 84660 12242 84712 12248
rect 84672 12102 84700 12242
rect 84660 12096 84712 12102
rect 84660 12038 84712 12044
rect 84856 11558 84884 12718
rect 85500 12442 85528 13194
rect 86040 13184 86092 13190
rect 86040 13126 86092 13132
rect 85764 12640 85816 12646
rect 85764 12582 85816 12588
rect 85488 12436 85540 12442
rect 85488 12378 85540 12384
rect 85776 12306 85804 12582
rect 85764 12300 85816 12306
rect 85764 12242 85816 12248
rect 85488 12232 85540 12238
rect 85488 12174 85540 12180
rect 84936 11824 84988 11830
rect 85304 11824 85356 11830
rect 84988 11772 85304 11778
rect 84936 11766 85356 11772
rect 84948 11750 85344 11766
rect 84844 11552 84896 11558
rect 84844 11494 84896 11500
rect 84476 11348 84528 11354
rect 84476 11290 84528 11296
rect 85500 11218 85528 12174
rect 85776 11762 85804 12242
rect 86052 12238 86080 13126
rect 86420 12442 86448 13670
rect 86776 13252 86828 13258
rect 86776 13194 86828 13200
rect 86500 12980 86552 12986
rect 86500 12922 86552 12928
rect 86512 12782 86540 12922
rect 86500 12776 86552 12782
rect 86500 12718 86552 12724
rect 86408 12436 86460 12442
rect 86408 12378 86460 12384
rect 86132 12368 86184 12374
rect 86132 12310 86184 12316
rect 86040 12232 86092 12238
rect 86040 12174 86092 12180
rect 86052 11898 86080 12174
rect 86144 11898 86172 12310
rect 86316 12300 86368 12306
rect 86316 12242 86368 12248
rect 86328 12102 86356 12242
rect 86316 12096 86368 12102
rect 86316 12038 86368 12044
rect 86040 11892 86092 11898
rect 86040 11834 86092 11840
rect 86132 11892 86184 11898
rect 86132 11834 86184 11840
rect 85764 11756 85816 11762
rect 85764 11698 85816 11704
rect 86328 11694 86356 12038
rect 86316 11688 86368 11694
rect 86316 11630 86368 11636
rect 86408 11552 86460 11558
rect 86408 11494 86460 11500
rect 85488 11212 85540 11218
rect 85488 11154 85540 11160
rect 86420 11150 86448 11494
rect 86788 11286 86816 13194
rect 86958 13152 87014 13160
rect 86958 13086 87014 13096
rect 86972 11762 87000 13086
rect 87144 12980 87196 12986
rect 87144 12922 87196 12928
rect 86960 11756 87012 11762
rect 86960 11698 87012 11704
rect 87156 11354 87184 12922
rect 87432 12374 87460 15200
rect 87880 13320 87932 13326
rect 87880 13262 87932 13268
rect 87786 12744 87842 12752
rect 87786 12678 87842 12688
rect 87800 12646 87828 12678
rect 87788 12640 87840 12646
rect 87788 12582 87840 12588
rect 87892 12442 87920 13262
rect 89076 13252 89128 13258
rect 89076 13194 89128 13200
rect 89536 13252 89588 13258
rect 89536 13194 89588 13200
rect 88248 13184 88300 13190
rect 88248 13126 88300 13132
rect 88260 12782 88288 13126
rect 88248 12776 88300 12782
rect 88248 12718 88300 12724
rect 87972 12640 88024 12646
rect 87972 12582 88024 12588
rect 87880 12436 87932 12442
rect 87880 12378 87932 12384
rect 87420 12368 87472 12374
rect 87420 12310 87472 12316
rect 87984 12186 88012 12582
rect 88154 12336 88210 12344
rect 88154 12270 88156 12280
rect 88208 12270 88210 12280
rect 88156 12242 88208 12248
rect 88260 12238 88288 12718
rect 88432 12640 88484 12646
rect 88432 12582 88484 12588
rect 87524 12158 88012 12186
rect 88248 12232 88300 12238
rect 88248 12174 88300 12180
rect 87524 12102 87552 12158
rect 87984 12102 88012 12158
rect 87512 12096 87564 12102
rect 87512 12038 87564 12044
rect 87788 12096 87840 12102
rect 87788 12038 87840 12044
rect 87972 12096 88024 12102
rect 87972 12038 88024 12044
rect 87144 11348 87196 11354
rect 87144 11290 87196 11296
rect 86776 11280 86828 11286
rect 86776 11222 86828 11228
rect 87800 11150 87828 12038
rect 87880 11892 87932 11898
rect 87880 11834 87932 11840
rect 86408 11144 86460 11150
rect 86408 11086 86460 11092
rect 87788 11144 87840 11150
rect 87788 11086 87840 11092
rect 87892 11082 87920 11834
rect 88444 11150 88472 12582
rect 88984 12232 89036 12238
rect 88720 12180 88984 12186
rect 88720 12174 89036 12180
rect 88720 12158 89024 12174
rect 88720 12102 88748 12158
rect 88708 12096 88760 12102
rect 88708 12038 88760 12044
rect 89088 11354 89116 13194
rect 89168 12300 89220 12306
rect 89168 12242 89220 12248
rect 89180 11762 89208 12242
rect 89548 11898 89576 13194
rect 90468 12986 90496 15200
rect 90640 13796 90692 13802
rect 90640 13738 90692 13744
rect 90548 13184 90600 13190
rect 90548 13126 90600 13132
rect 90456 12980 90508 12986
rect 90456 12922 90508 12928
rect 90560 12918 90588 13126
rect 90548 12912 90600 12918
rect 90548 12854 90600 12860
rect 90652 12850 90680 13738
rect 91836 13728 91888 13734
rect 91836 13670 91888 13676
rect 91848 13258 91876 13670
rect 93780 13546 93808 15286
rect 96618 15286 96752 15314
rect 96618 15200 96674 15286
rect 93780 13518 93900 13546
rect 93872 13462 93900 13518
rect 93860 13456 93912 13462
rect 93860 13398 93912 13404
rect 91652 13252 91704 13258
rect 91652 13194 91704 13200
rect 91836 13252 91888 13258
rect 91836 13194 91888 13200
rect 92020 13252 92072 13258
rect 92020 13194 92072 13200
rect 91664 12986 91692 13194
rect 91848 13160 91876 13194
rect 91834 13152 91890 13160
rect 91834 13086 91890 13096
rect 91652 12980 91704 12986
rect 91652 12922 91704 12928
rect 90732 12912 90784 12918
rect 90732 12854 90784 12860
rect 90180 12844 90232 12850
rect 90180 12786 90232 12792
rect 90456 12844 90508 12850
rect 90456 12786 90508 12792
rect 90640 12844 90692 12850
rect 90640 12786 90692 12792
rect 89720 12776 89772 12782
rect 90088 12776 90140 12782
rect 89772 12736 90088 12764
rect 89720 12718 89772 12724
rect 90088 12718 90140 12724
rect 89904 12640 89956 12646
rect 89904 12582 89956 12588
rect 89916 12344 89944 12582
rect 90192 12442 90220 12786
rect 90180 12436 90232 12442
rect 90180 12378 90232 12384
rect 89902 12336 89958 12344
rect 89902 12270 89958 12280
rect 89536 11892 89588 11898
rect 89536 11834 89588 11840
rect 89168 11756 89220 11762
rect 89168 11698 89220 11704
rect 89076 11348 89128 11354
rect 89076 11290 89128 11296
rect 89180 11218 89208 11698
rect 90468 11694 90496 12786
rect 90744 12752 90772 12854
rect 90730 12744 90786 12752
rect 90730 12678 90786 12688
rect 92032 12238 92060 13194
rect 96724 13190 96752 15286
rect 99654 15200 99710 16000
rect 102782 15314 102838 16000
rect 105818 15314 105874 16000
rect 108854 15314 108910 16000
rect 111982 15314 112038 16000
rect 102782 15286 102916 15314
rect 102782 15200 102838 15286
rect 99668 13410 99696 15200
rect 102416 13796 102468 13802
rect 102416 13738 102468 13744
rect 101956 13728 102008 13734
rect 101956 13670 102008 13676
rect 99104 13388 99156 13394
rect 99104 13330 99156 13336
rect 99392 13382 99696 13410
rect 100760 13456 100812 13462
rect 100760 13398 100812 13404
rect 98000 13252 98052 13258
rect 98000 13194 98052 13200
rect 96712 13184 96764 13190
rect 96712 13126 96764 13132
rect 97540 13184 97592 13190
rect 97540 13126 97592 13132
rect 97552 12238 97580 13126
rect 98012 12986 98040 13194
rect 98000 12980 98052 12986
rect 98000 12922 98052 12928
rect 99116 12306 99144 13330
rect 99196 13252 99248 13258
rect 99196 13194 99248 13200
rect 99208 12782 99236 13194
rect 99196 12776 99248 12782
rect 99196 12718 99248 12724
rect 99196 12640 99248 12646
rect 99392 12628 99420 13382
rect 99656 13252 99708 13258
rect 99656 13194 99708 13200
rect 99472 12912 99524 12918
rect 99472 12854 99524 12860
rect 99248 12600 99420 12628
rect 99196 12582 99248 12588
rect 99484 12442 99512 12854
rect 99472 12436 99524 12442
rect 99472 12378 99524 12384
rect 99104 12300 99156 12306
rect 99104 12242 99156 12248
rect 92020 12232 92072 12238
rect 92020 12174 92072 12180
rect 97540 12232 97592 12238
rect 97540 12174 97592 12180
rect 99668 11898 99696 13194
rect 99932 12912 99984 12918
rect 99932 12854 99984 12860
rect 99944 12442 99972 12854
rect 100772 12646 100800 13398
rect 101404 13320 101456 13326
rect 101404 13262 101456 13268
rect 100944 13252 100996 13258
rect 100944 13194 100996 13200
rect 100760 12640 100812 12646
rect 100760 12582 100812 12588
rect 99932 12436 99984 12442
rect 99932 12378 99984 12384
rect 100772 12170 100800 12582
rect 100760 12164 100812 12170
rect 100760 12106 100812 12112
rect 100392 12096 100444 12102
rect 100392 12038 100444 12044
rect 99656 11892 99708 11898
rect 99656 11834 99708 11840
rect 100404 11762 100432 12038
rect 100392 11756 100444 11762
rect 100392 11698 100444 11704
rect 100772 11694 100800 12106
rect 100956 11898 100984 13194
rect 101036 13184 101088 13190
rect 101036 13126 101088 13132
rect 101048 12714 101076 13126
rect 101416 12782 101444 13262
rect 101404 12776 101456 12782
rect 101404 12718 101456 12724
rect 101680 12776 101732 12782
rect 101680 12718 101732 12724
rect 101036 12708 101088 12714
rect 101036 12650 101088 12656
rect 101048 12170 101076 12650
rect 101036 12164 101088 12170
rect 101036 12106 101088 12112
rect 100944 11892 100996 11898
rect 100944 11834 100996 11840
rect 90456 11688 90508 11694
rect 90456 11630 90508 11636
rect 100760 11688 100812 11694
rect 100760 11630 100812 11636
rect 89168 11212 89220 11218
rect 89168 11154 89220 11160
rect 88432 11144 88484 11150
rect 88432 11086 88484 11092
rect 81624 11076 81676 11082
rect 81624 11018 81676 11024
rect 87880 11076 87932 11082
rect 87880 11018 87932 11024
rect 77148 10908 77456 10916
rect 77148 10906 77154 10908
rect 77210 10906 77234 10908
rect 77290 10906 77314 10908
rect 77370 10906 77394 10908
rect 77450 10906 77456 10908
rect 77210 10854 77212 10906
rect 77392 10854 77394 10906
rect 77148 10852 77154 10854
rect 77210 10852 77234 10854
rect 77290 10852 77314 10854
rect 77370 10852 77394 10854
rect 77450 10852 77456 10854
rect 77148 10842 77456 10852
rect 101692 10810 101720 12718
rect 101968 12170 101996 13670
rect 102232 13252 102284 13258
rect 102232 13194 102284 13200
rect 102048 12300 102100 12306
rect 102048 12242 102100 12248
rect 101956 12164 102008 12170
rect 101956 12106 102008 12112
rect 102060 11694 102088 12242
rect 102140 12164 102192 12170
rect 102140 12106 102192 12112
rect 102152 11762 102180 12106
rect 102140 11756 102192 11762
rect 102140 11698 102192 11704
rect 102048 11688 102100 11694
rect 102048 11630 102100 11636
rect 101864 11552 101916 11558
rect 101864 11494 101916 11500
rect 101680 10804 101732 10810
rect 101680 10746 101732 10752
rect 101876 10674 101904 11494
rect 102060 11218 102088 11630
rect 102244 11286 102272 13194
rect 102324 12096 102376 12102
rect 102324 12038 102376 12044
rect 102336 11694 102364 12038
rect 102324 11688 102376 11694
rect 102324 11630 102376 11636
rect 102232 11280 102284 11286
rect 102232 11222 102284 11228
rect 102048 11212 102100 11218
rect 102048 11154 102100 11160
rect 102428 11150 102456 13738
rect 102600 12096 102652 12102
rect 102600 12038 102652 12044
rect 102612 11218 102640 12038
rect 102888 11354 102916 15286
rect 105818 15286 105952 15314
rect 105818 15200 105874 15286
rect 103336 13320 103388 13326
rect 103336 13262 103388 13268
rect 104256 13320 104308 13326
rect 104256 13262 104308 13268
rect 103244 12708 103296 12714
rect 103244 12650 103296 12656
rect 103060 12640 103112 12646
rect 103060 12582 103112 12588
rect 103072 12102 103100 12582
rect 103256 12306 103284 12650
rect 103348 12306 103376 13262
rect 104072 13252 104124 13258
rect 104072 13194 104124 13200
rect 103704 13184 103756 13190
rect 103704 13126 103756 13132
rect 103612 12640 103664 12646
rect 103612 12582 103664 12588
rect 103244 12300 103296 12306
rect 103244 12242 103296 12248
rect 103336 12300 103388 12306
rect 103336 12242 103388 12248
rect 103060 12096 103112 12102
rect 103060 12038 103112 12044
rect 103072 11898 103100 12038
rect 103060 11892 103112 11898
rect 103060 11834 103112 11840
rect 103520 11892 103572 11898
rect 103520 11834 103572 11840
rect 102876 11348 102928 11354
rect 102876 11290 102928 11296
rect 102600 11212 102652 11218
rect 102600 11154 102652 11160
rect 103072 11150 103100 11834
rect 103532 11694 103560 11834
rect 103624 11762 103652 12582
rect 103716 12238 103744 13126
rect 103704 12232 103756 12238
rect 103704 12174 103756 12180
rect 103612 11756 103664 11762
rect 103612 11698 103664 11704
rect 103520 11688 103572 11694
rect 103520 11630 103572 11636
rect 104084 11558 104112 13194
rect 104072 11552 104124 11558
rect 104072 11494 104124 11500
rect 102416 11144 102468 11150
rect 102416 11086 102468 11092
rect 103060 11144 103112 11150
rect 103060 11086 103112 11092
rect 101864 10668 101916 10674
rect 101864 10610 101916 10616
rect 39048 10364 39356 10372
rect 39048 10362 39054 10364
rect 39110 10362 39134 10364
rect 39190 10362 39214 10364
rect 39270 10362 39294 10364
rect 39350 10362 39356 10364
rect 39110 10310 39112 10362
rect 39292 10310 39294 10362
rect 39048 10308 39054 10310
rect 39110 10308 39134 10310
rect 39190 10308 39214 10310
rect 39270 10308 39294 10310
rect 39350 10308 39356 10310
rect 39048 10298 39356 10308
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33692 10056 33744 10062
rect 33692 9998 33744 10004
rect 31208 9648 31260 9654
rect 31208 9590 31260 9596
rect 33704 9586 33732 9998
rect 77148 9820 77456 9828
rect 77148 9818 77154 9820
rect 77210 9818 77234 9820
rect 77290 9818 77314 9820
rect 77370 9818 77394 9820
rect 77450 9818 77456 9820
rect 77210 9766 77212 9818
rect 77392 9766 77394 9818
rect 77148 9764 77154 9766
rect 77210 9764 77234 9766
rect 77290 9764 77314 9766
rect 77370 9764 77394 9766
rect 77450 9764 77456 9766
rect 77148 9754 77456 9764
rect 33692 9580 33744 9586
rect 33692 9522 33744 9528
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 29920 9444 29972 9450
rect 29920 9386 29972 9392
rect 104268 9382 104296 13262
rect 104452 13246 104756 13274
rect 104452 13190 104480 13246
rect 104440 13184 104492 13190
rect 104440 13126 104492 13132
rect 104624 13184 104676 13190
rect 104624 13126 104676 13132
rect 104636 12918 104664 13126
rect 104728 12918 104756 13246
rect 104992 13252 105044 13258
rect 104992 13194 105044 13200
rect 104624 12912 104676 12918
rect 104624 12854 104676 12860
rect 104716 12912 104768 12918
rect 104716 12854 104768 12860
rect 105004 12442 105032 13194
rect 105176 12844 105228 12850
rect 105176 12786 105228 12792
rect 105188 12442 105216 12786
rect 105924 12714 105952 15286
rect 108854 15286 108988 15314
rect 108854 15200 108910 15286
rect 108960 13546 108988 15286
rect 111812 15286 112038 15314
rect 111812 13546 111840 15286
rect 111982 15200 112038 15286
rect 115018 15200 115074 16000
rect 118146 15314 118202 16000
rect 121182 15314 121238 16000
rect 118146 15286 118648 15314
rect 118146 15200 118202 15286
rect 113824 13796 113876 13802
rect 113824 13738 113876 13744
rect 108960 13518 109080 13546
rect 109052 13462 109080 13518
rect 111720 13518 111840 13546
rect 111720 13462 111748 13518
rect 109040 13456 109092 13462
rect 109040 13398 109092 13404
rect 111708 13456 111760 13462
rect 111708 13398 111760 13404
rect 109592 13320 109644 13326
rect 109592 13262 109644 13268
rect 111432 13320 111484 13326
rect 111432 13262 111484 13268
rect 109604 13190 109632 13262
rect 109592 13184 109644 13190
rect 109592 13126 109644 13132
rect 109604 12918 109632 13126
rect 111444 12986 111472 13262
rect 112536 13252 112588 13258
rect 112536 13194 112588 13200
rect 111432 12980 111484 12986
rect 111432 12922 111484 12928
rect 109592 12912 109644 12918
rect 109592 12854 109644 12860
rect 105912 12708 105964 12714
rect 105912 12650 105964 12656
rect 111892 12640 111944 12646
rect 111892 12582 111944 12588
rect 104992 12436 105044 12442
rect 104992 12378 105044 12384
rect 105176 12436 105228 12442
rect 105176 12378 105228 12384
rect 111904 12238 111932 12582
rect 112548 12442 112576 13194
rect 113836 12850 113864 13738
rect 114652 13728 114704 13734
rect 114652 13670 114704 13676
rect 114192 13252 114244 13258
rect 114192 13194 114244 13200
rect 113088 12844 113140 12850
rect 113088 12786 113140 12792
rect 113824 12844 113876 12850
rect 113824 12786 113876 12792
rect 113100 12646 113128 12786
rect 113088 12640 113140 12646
rect 113088 12582 113140 12588
rect 112536 12436 112588 12442
rect 112536 12378 112588 12384
rect 113836 12322 113864 12786
rect 113916 12776 113968 12782
rect 113916 12718 113968 12724
rect 113744 12294 113864 12322
rect 111892 12232 111944 12238
rect 111892 12174 111944 12180
rect 113744 11082 113772 12294
rect 113824 12164 113876 12170
rect 113824 12106 113876 12112
rect 113836 11898 113864 12106
rect 113928 12102 113956 12718
rect 113916 12096 113968 12102
rect 113916 12038 113968 12044
rect 113824 11892 113876 11898
rect 113824 11834 113876 11840
rect 114008 11756 114060 11762
rect 114008 11698 114060 11704
rect 114020 11558 114048 11698
rect 114008 11552 114060 11558
rect 114008 11494 114060 11500
rect 114204 11286 114232 13194
rect 114560 13184 114612 13190
rect 114560 13126 114612 13132
rect 114572 12986 114600 13126
rect 114560 12980 114612 12986
rect 114560 12922 114612 12928
rect 114664 12850 114692 13670
rect 114836 13320 114888 13326
rect 114836 13262 114888 13268
rect 114744 12980 114796 12986
rect 114744 12922 114796 12928
rect 114652 12844 114704 12850
rect 114652 12786 114704 12792
rect 114664 12322 114692 12786
rect 114756 12782 114784 12922
rect 114744 12776 114796 12782
rect 114744 12718 114796 12724
rect 114848 12714 114876 13262
rect 114928 13184 114980 13190
rect 114928 13126 114980 13132
rect 114836 12708 114888 12714
rect 114836 12650 114888 12656
rect 114744 12640 114796 12646
rect 114744 12582 114796 12588
rect 114572 12294 114692 12322
rect 114284 12232 114336 12238
rect 114284 12174 114336 12180
rect 114296 11898 114324 12174
rect 114284 11892 114336 11898
rect 114284 11834 114336 11840
rect 114572 11830 114600 12294
rect 114560 11824 114612 11830
rect 114560 11766 114612 11772
rect 114192 11280 114244 11286
rect 114192 11222 114244 11228
rect 114756 11150 114784 12582
rect 114940 12322 114968 13126
rect 115032 12442 115060 15200
rect 118620 13682 118648 15286
rect 121182 15286 121316 15314
rect 121182 15200 121238 15286
rect 118620 13654 118740 13682
rect 115246 13628 115554 13636
rect 115246 13626 115252 13628
rect 115308 13626 115332 13628
rect 115388 13626 115412 13628
rect 115468 13626 115492 13628
rect 115548 13626 115554 13628
rect 115308 13574 115310 13626
rect 115490 13574 115492 13626
rect 115246 13572 115252 13574
rect 115308 13572 115332 13574
rect 115388 13572 115412 13574
rect 115468 13572 115492 13574
rect 115548 13572 115554 13574
rect 115246 13562 115554 13572
rect 118240 13388 118292 13394
rect 118240 13330 118292 13336
rect 117412 13320 117464 13326
rect 117412 13262 117464 13268
rect 115112 13252 115164 13258
rect 115112 13194 115164 13200
rect 116952 13252 117004 13258
rect 116952 13194 117004 13200
rect 115020 12436 115072 12442
rect 115020 12378 115072 12384
rect 114940 12294 115060 12322
rect 115032 11762 115060 12294
rect 115020 11756 115072 11762
rect 115020 11698 115072 11704
rect 115124 11354 115152 13194
rect 115756 13184 115808 13190
rect 115756 13126 115808 13132
rect 115768 12918 115796 13126
rect 115756 12912 115808 12918
rect 115756 12854 115808 12860
rect 115664 12776 115716 12782
rect 115848 12776 115900 12782
rect 115664 12718 115716 12724
rect 115768 12724 115848 12730
rect 115768 12718 115900 12724
rect 116768 12776 116820 12782
rect 116768 12718 116820 12724
rect 115246 12540 115554 12548
rect 115246 12538 115252 12540
rect 115308 12538 115332 12540
rect 115388 12538 115412 12540
rect 115468 12538 115492 12540
rect 115548 12538 115554 12540
rect 115308 12486 115310 12538
rect 115490 12486 115492 12538
rect 115246 12484 115252 12486
rect 115308 12484 115332 12486
rect 115388 12484 115412 12486
rect 115468 12484 115492 12486
rect 115548 12484 115554 12486
rect 115246 12474 115554 12484
rect 115676 12102 115704 12718
rect 115768 12702 115888 12718
rect 115768 12374 115796 12702
rect 115848 12640 115900 12646
rect 115848 12582 115900 12588
rect 115756 12368 115808 12374
rect 115756 12310 115808 12316
rect 115664 12096 115716 12102
rect 115664 12038 115716 12044
rect 115676 11898 115704 12038
rect 115664 11892 115716 11898
rect 115664 11834 115716 11840
rect 115768 11778 115796 12310
rect 115676 11750 115796 11778
rect 115676 11694 115704 11750
rect 115664 11688 115716 11694
rect 115664 11630 115716 11636
rect 115756 11688 115808 11694
rect 115756 11630 115808 11636
rect 115246 11452 115554 11460
rect 115246 11450 115252 11452
rect 115308 11450 115332 11452
rect 115388 11450 115412 11452
rect 115468 11450 115492 11452
rect 115548 11450 115554 11452
rect 115308 11398 115310 11450
rect 115490 11398 115492 11450
rect 115246 11396 115252 11398
rect 115308 11396 115332 11398
rect 115388 11396 115412 11398
rect 115468 11396 115492 11398
rect 115548 11396 115554 11398
rect 115246 11386 115554 11396
rect 115112 11348 115164 11354
rect 115112 11290 115164 11296
rect 115768 11150 115796 11630
rect 115860 11150 115888 12582
rect 116400 12096 116452 12102
rect 116400 12038 116452 12044
rect 116412 11762 116440 12038
rect 116780 11898 116808 12718
rect 116964 12442 116992 13194
rect 117424 12986 117452 13262
rect 117688 13252 117740 13258
rect 117688 13194 117740 13200
rect 117412 12980 117464 12986
rect 117412 12922 117464 12928
rect 117320 12912 117372 12918
rect 117320 12854 117372 12860
rect 116952 12436 117004 12442
rect 116952 12378 117004 12384
rect 117332 11898 117360 12854
rect 116768 11892 116820 11898
rect 116768 11834 116820 11840
rect 117320 11892 117372 11898
rect 117320 11834 117372 11840
rect 116400 11756 116452 11762
rect 116400 11698 116452 11704
rect 114744 11144 114796 11150
rect 114744 11086 114796 11092
rect 115756 11144 115808 11150
rect 115756 11086 115808 11092
rect 115848 11144 115900 11150
rect 115848 11086 115900 11092
rect 113732 11076 113784 11082
rect 113732 11018 113784 11024
rect 115246 10364 115554 10372
rect 115246 10362 115252 10364
rect 115308 10362 115332 10364
rect 115388 10362 115412 10364
rect 115468 10362 115492 10364
rect 115548 10362 115554 10364
rect 115308 10310 115310 10362
rect 115490 10310 115492 10362
rect 115246 10308 115252 10310
rect 115308 10308 115332 10310
rect 115388 10308 115412 10310
rect 115468 10308 115492 10310
rect 115548 10308 115554 10310
rect 115246 10298 115554 10308
rect 117424 9926 117452 12922
rect 117700 11354 117728 13194
rect 118056 13184 118108 13190
rect 118056 13126 118108 13132
rect 118068 12850 118096 13126
rect 118252 12986 118280 13330
rect 118712 12986 118740 13654
rect 121288 13462 121316 15286
rect 124218 15200 124274 16000
rect 127346 15314 127402 16000
rect 126992 15286 127402 15314
rect 124232 13682 124260 15200
rect 125508 13796 125560 13802
rect 125508 13738 125560 13744
rect 124140 13654 124260 13682
rect 124140 13462 124168 13654
rect 118884 13456 118936 13462
rect 118884 13398 118936 13404
rect 121276 13456 121328 13462
rect 121276 13398 121328 13404
rect 124128 13456 124180 13462
rect 124128 13398 124180 13404
rect 118792 13320 118844 13326
rect 118792 13262 118844 13268
rect 118240 12980 118292 12986
rect 118240 12922 118292 12928
rect 118700 12980 118752 12986
rect 118700 12922 118752 12928
rect 118056 12844 118108 12850
rect 118056 12786 118108 12792
rect 118068 12238 118096 12786
rect 118056 12232 118108 12238
rect 118056 12174 118108 12180
rect 118252 12170 118280 12922
rect 118332 12232 118384 12238
rect 118332 12174 118384 12180
rect 118240 12164 118292 12170
rect 118240 12106 118292 12112
rect 118344 11762 118372 12174
rect 118804 11898 118832 13262
rect 118896 12306 118924 13398
rect 125520 13258 125548 13738
rect 125508 13252 125560 13258
rect 125508 13194 125560 13200
rect 119712 13184 119764 13190
rect 119712 13126 119764 13132
rect 126152 13184 126204 13190
rect 126152 13126 126204 13132
rect 126520 13184 126572 13190
rect 126520 13126 126572 13132
rect 118884 12300 118936 12306
rect 118884 12242 118936 12248
rect 118792 11892 118844 11898
rect 118792 11834 118844 11840
rect 118332 11756 118384 11762
rect 118332 11698 118384 11704
rect 117688 11348 117740 11354
rect 117688 11290 117740 11296
rect 119724 11150 119752 13126
rect 126164 12238 126192 13126
rect 126532 12918 126560 13126
rect 126992 13002 127020 15286
rect 127346 15200 127402 15286
rect 130382 15200 130438 16000
rect 133418 15314 133474 16000
rect 133418 15286 133828 15314
rect 133418 15200 133474 15286
rect 127440 13728 127492 13734
rect 127440 13670 127492 13676
rect 127532 13728 127584 13734
rect 127532 13670 127584 13676
rect 129740 13728 129792 13734
rect 129740 13670 129792 13676
rect 126900 12986 127020 13002
rect 126888 12980 127020 12986
rect 126940 12974 127020 12980
rect 126888 12922 126940 12928
rect 126520 12912 126572 12918
rect 126520 12854 126572 12860
rect 127452 12850 127480 13670
rect 127544 13462 127572 13670
rect 127532 13456 127584 13462
rect 127532 13398 127584 13404
rect 127532 13320 127584 13326
rect 127532 13262 127584 13268
rect 129372 13320 129424 13326
rect 129372 13262 129424 13268
rect 127440 12844 127492 12850
rect 127440 12786 127492 12792
rect 127544 12782 127572 13262
rect 127808 13252 127860 13258
rect 127808 13194 127860 13200
rect 127532 12776 127584 12782
rect 127532 12718 127584 12724
rect 127820 12442 127848 13194
rect 128084 13184 128136 13190
rect 128084 13126 128136 13132
rect 129188 13184 129240 13190
rect 129188 13126 129240 13132
rect 128096 12986 128124 13126
rect 129200 12986 129228 13126
rect 128084 12980 128136 12986
rect 128084 12922 128136 12928
rect 128636 12980 128688 12986
rect 128636 12922 128688 12928
rect 129188 12980 129240 12986
rect 129188 12922 129240 12928
rect 128360 12776 128412 12782
rect 128360 12718 128412 12724
rect 128084 12640 128136 12646
rect 128372 12594 128400 12718
rect 128136 12588 128400 12594
rect 128084 12582 128400 12588
rect 128096 12566 128400 12582
rect 127808 12436 127860 12442
rect 127808 12378 127860 12384
rect 126152 12232 126204 12238
rect 126152 12174 126204 12180
rect 128372 11762 128400 12566
rect 128648 12238 128676 12922
rect 129096 12844 129148 12850
rect 129096 12786 129148 12792
rect 129108 12442 129136 12786
rect 129096 12436 129148 12442
rect 129096 12378 129148 12384
rect 128636 12232 128688 12238
rect 128636 12174 128688 12180
rect 129384 11898 129412 13262
rect 129752 12782 129780 13670
rect 130292 13388 130344 13394
rect 130292 13330 130344 13336
rect 130304 12850 130332 13330
rect 130292 12844 130344 12850
rect 130292 12786 130344 12792
rect 129740 12776 129792 12782
rect 129740 12718 129792 12724
rect 129372 11892 129424 11898
rect 129372 11834 129424 11840
rect 128360 11756 128412 11762
rect 128360 11698 128412 11704
rect 129752 11694 129780 12718
rect 130292 12708 130344 12714
rect 130292 12650 130344 12656
rect 130304 11898 130332 12650
rect 130292 11892 130344 11898
rect 130292 11834 130344 11840
rect 130292 11756 130344 11762
rect 130292 11698 130344 11704
rect 129740 11688 129792 11694
rect 129740 11630 129792 11636
rect 130304 11218 130332 11698
rect 130396 11354 130424 15200
rect 131856 13796 131908 13802
rect 131856 13738 131908 13744
rect 131212 13252 131264 13258
rect 131212 13194 131264 13200
rect 131120 12776 131172 12782
rect 131120 12718 131172 12724
rect 130936 12436 130988 12442
rect 130936 12378 130988 12384
rect 130476 12232 130528 12238
rect 130476 12174 130528 12180
rect 130384 11348 130436 11354
rect 130384 11290 130436 11296
rect 130292 11212 130344 11218
rect 130292 11154 130344 11160
rect 119712 11144 119764 11150
rect 119712 11086 119764 11092
rect 130304 10674 130332 11154
rect 130488 10810 130516 12174
rect 130948 11898 130976 12378
rect 131028 12300 131080 12306
rect 131028 12242 131080 12248
rect 130936 11892 130988 11898
rect 130936 11834 130988 11840
rect 130948 11150 130976 11834
rect 131040 11694 131068 12242
rect 131132 11898 131160 12718
rect 131120 11892 131172 11898
rect 131120 11834 131172 11840
rect 131028 11688 131080 11694
rect 131028 11630 131080 11636
rect 131224 11354 131252 13194
rect 131580 13184 131632 13190
rect 131580 13126 131632 13132
rect 131592 12102 131620 13126
rect 131580 12096 131632 12102
rect 131580 12038 131632 12044
rect 131592 11762 131620 12038
rect 131580 11756 131632 11762
rect 131580 11698 131632 11704
rect 131868 11558 131896 13738
rect 133604 13728 133656 13734
rect 133604 13670 133656 13676
rect 132868 13252 132920 13258
rect 132868 13194 132920 13200
rect 133328 13252 133380 13258
rect 133328 13194 133380 13200
rect 132408 12912 132460 12918
rect 132408 12854 132460 12860
rect 132420 12442 132448 12854
rect 132592 12776 132644 12782
rect 132592 12718 132644 12724
rect 132408 12436 132460 12442
rect 132408 12378 132460 12384
rect 132604 12322 132632 12718
rect 132420 12294 132632 12322
rect 132420 12238 132448 12294
rect 132408 12232 132460 12238
rect 132408 12174 132460 12180
rect 132592 12232 132644 12238
rect 132592 12174 132644 12180
rect 132500 12164 132552 12170
rect 132500 12106 132552 12112
rect 132512 11762 132540 12106
rect 132500 11756 132552 11762
rect 132500 11698 132552 11704
rect 131856 11552 131908 11558
rect 131856 11494 131908 11500
rect 131212 11348 131264 11354
rect 131212 11290 131264 11296
rect 132604 11218 132632 12174
rect 132880 11354 132908 13194
rect 133340 12986 133368 13194
rect 133328 12980 133380 12986
rect 133328 12922 133380 12928
rect 133616 12918 133644 13670
rect 133800 13274 133828 15286
rect 136546 15200 136602 16000
rect 139582 15200 139638 16000
rect 142710 15314 142766 16000
rect 142710 15286 142936 15314
rect 142710 15200 142766 15286
rect 136560 13682 136588 15200
rect 136824 13728 136876 13734
rect 136560 13654 136680 13682
rect 136824 13670 136876 13676
rect 136652 13462 136680 13654
rect 136640 13456 136692 13462
rect 136640 13398 136692 13404
rect 136836 13326 136864 13670
rect 139596 13462 139624 15200
rect 142908 13530 142936 15286
rect 145746 15200 145802 16000
rect 148782 15314 148838 16000
rect 148520 15286 148838 15314
rect 145760 13530 145788 15200
rect 148140 13728 148192 13734
rect 148140 13670 148192 13676
rect 148152 13530 148180 13670
rect 142896 13524 142948 13530
rect 142896 13466 142948 13472
rect 145748 13524 145800 13530
rect 145748 13466 145800 13472
rect 148140 13524 148192 13530
rect 148140 13466 148192 13472
rect 139584 13456 139636 13462
rect 139584 13398 139636 13404
rect 142068 13388 142120 13394
rect 142068 13330 142120 13336
rect 136824 13320 136876 13326
rect 133800 13246 133920 13274
rect 136824 13262 136876 13268
rect 133696 13184 133748 13190
rect 133696 13126 133748 13132
rect 133604 12912 133656 12918
rect 133604 12854 133656 12860
rect 133708 12850 133736 13126
rect 133892 12986 133920 13246
rect 134156 13184 134208 13190
rect 134156 13126 134208 13132
rect 133880 12980 133932 12986
rect 133880 12922 133932 12928
rect 134168 12918 134196 13126
rect 134156 12912 134208 12918
rect 134156 12854 134208 12860
rect 133696 12844 133748 12850
rect 133696 12786 133748 12792
rect 133708 12714 133920 12730
rect 133696 12708 133932 12714
rect 133748 12702 133880 12708
rect 133696 12650 133748 12656
rect 133880 12650 133932 12656
rect 133144 12640 133196 12646
rect 133144 12582 133196 12588
rect 133236 12640 133288 12646
rect 133236 12582 133288 12588
rect 132868 11348 132920 11354
rect 132868 11290 132920 11296
rect 132592 11212 132644 11218
rect 132592 11154 132644 11160
rect 133156 11150 133184 12582
rect 133248 12306 133276 12582
rect 141976 12368 142028 12374
rect 141976 12310 142028 12316
rect 133236 12300 133288 12306
rect 133236 12242 133288 12248
rect 137744 12232 137796 12238
rect 137744 12174 137796 12180
rect 137756 11898 137784 12174
rect 138020 12164 138072 12170
rect 138020 12106 138072 12112
rect 137744 11892 137796 11898
rect 137744 11834 137796 11840
rect 137756 11694 137784 11834
rect 138032 11830 138060 12106
rect 138020 11824 138072 11830
rect 138020 11766 138072 11772
rect 137744 11688 137796 11694
rect 137744 11630 137796 11636
rect 130936 11144 130988 11150
rect 130936 11086 130988 11092
rect 133144 11144 133196 11150
rect 133144 11086 133196 11092
rect 140688 11076 140740 11082
rect 140688 11018 140740 11024
rect 130476 10804 130528 10810
rect 130476 10746 130528 10752
rect 140700 10742 140728 11018
rect 141988 10810 142016 12310
rect 142080 11150 142108 13330
rect 143080 13320 143132 13326
rect 143080 13262 143132 13268
rect 145748 13320 145800 13326
rect 145748 13262 145800 13268
rect 143092 12918 143120 13262
rect 143080 12912 143132 12918
rect 143080 12854 143132 12860
rect 143264 12776 143316 12782
rect 143264 12718 143316 12724
rect 143276 11626 143304 12718
rect 145760 12714 145788 13262
rect 145932 13252 145984 13258
rect 145932 13194 145984 13200
rect 146024 13252 146076 13258
rect 146024 13194 146076 13200
rect 147588 13252 147640 13258
rect 147588 13194 147640 13200
rect 145840 13184 145892 13190
rect 145840 13126 145892 13132
rect 145852 12850 145880 13126
rect 145944 12918 145972 13194
rect 145932 12912 145984 12918
rect 145932 12854 145984 12860
rect 145840 12844 145892 12850
rect 145840 12786 145892 12792
rect 145748 12708 145800 12714
rect 145748 12650 145800 12656
rect 143264 11620 143316 11626
rect 143264 11562 143316 11568
rect 143276 11218 143304 11562
rect 143264 11212 143316 11218
rect 143264 11154 143316 11160
rect 145760 11150 145788 12650
rect 146036 11626 146064 13194
rect 147496 13184 147548 13190
rect 147496 13126 147548 13132
rect 147312 12844 147364 12850
rect 147312 12786 147364 12792
rect 146024 11620 146076 11626
rect 146024 11562 146076 11568
rect 147324 11558 147352 12786
rect 147404 12776 147456 12782
rect 147404 12718 147456 12724
rect 147312 11552 147364 11558
rect 147312 11494 147364 11500
rect 147416 11286 147444 12718
rect 147404 11280 147456 11286
rect 147404 11222 147456 11228
rect 147508 11218 147536 13126
rect 147600 12374 147628 13194
rect 147680 12980 147732 12986
rect 147680 12922 147732 12928
rect 147588 12368 147640 12374
rect 147588 12310 147640 12316
rect 147692 11762 147720 12922
rect 147772 12776 147824 12782
rect 147772 12718 147824 12724
rect 147784 12442 147812 12718
rect 148520 12646 148548 15286
rect 148782 15200 148838 15286
rect 151910 15314 151966 16000
rect 151910 15286 152044 15314
rect 151910 15200 151966 15286
rect 150440 13728 150492 13734
rect 150440 13670 150492 13676
rect 150452 13258 150480 13670
rect 150808 13524 150860 13530
rect 150808 13466 150860 13472
rect 150440 13252 150492 13258
rect 150440 13194 150492 13200
rect 149244 13184 149296 13190
rect 149244 13126 149296 13132
rect 149256 12782 149284 13126
rect 150452 12850 150480 13194
rect 149336 12844 149388 12850
rect 149336 12786 149388 12792
rect 150440 12844 150492 12850
rect 150440 12786 150492 12792
rect 148968 12776 149020 12782
rect 149244 12776 149296 12782
rect 148968 12718 149020 12724
rect 149072 12736 149244 12764
rect 148508 12640 148560 12646
rect 148508 12582 148560 12588
rect 147772 12436 147824 12442
rect 147772 12378 147824 12384
rect 148048 12232 148100 12238
rect 148048 12174 148100 12180
rect 147680 11756 147732 11762
rect 147680 11698 147732 11704
rect 148060 11354 148088 12174
rect 148324 11688 148376 11694
rect 148324 11630 148376 11636
rect 148600 11688 148652 11694
rect 148600 11630 148652 11636
rect 148048 11348 148100 11354
rect 148048 11290 148100 11296
rect 147496 11212 147548 11218
rect 147496 11154 147548 11160
rect 142068 11144 142120 11150
rect 142068 11086 142120 11092
rect 145748 11144 145800 11150
rect 145748 11086 145800 11092
rect 141976 10804 142028 10810
rect 141976 10746 142028 10752
rect 140688 10736 140740 10742
rect 140688 10678 140740 10684
rect 130292 10668 130344 10674
rect 130292 10610 130344 10616
rect 140700 10062 140728 10678
rect 140688 10056 140740 10062
rect 140688 9998 140740 10004
rect 117412 9920 117464 9926
rect 117412 9862 117464 9868
rect 140700 9654 140728 9998
rect 140688 9648 140740 9654
rect 140688 9590 140740 9596
rect 148336 9382 148364 11630
rect 148612 10810 148640 11630
rect 148980 10810 149008 12718
rect 149072 12306 149100 12736
rect 149244 12718 149296 12724
rect 149060 12300 149112 12306
rect 149060 12242 149112 12248
rect 149072 11014 149100 12242
rect 149348 12238 149376 12786
rect 150348 12708 150400 12714
rect 150348 12650 150400 12656
rect 149980 12640 150032 12646
rect 149980 12582 150032 12588
rect 149336 12232 149388 12238
rect 149336 12174 149388 12180
rect 149428 12232 149480 12238
rect 149428 12174 149480 12180
rect 149060 11008 149112 11014
rect 149060 10950 149112 10956
rect 148600 10804 148652 10810
rect 148600 10746 148652 10752
rect 148968 10804 149020 10810
rect 148968 10746 149020 10752
rect 104256 9376 104308 9382
rect 104256 9318 104308 9324
rect 148324 9376 148376 9382
rect 148324 9318 148376 9324
rect 39048 9276 39356 9284
rect 39048 9274 39054 9276
rect 39110 9274 39134 9276
rect 39190 9274 39214 9276
rect 39270 9274 39294 9276
rect 39350 9274 39356 9276
rect 39110 9222 39112 9274
rect 39292 9222 39294 9274
rect 39048 9220 39054 9222
rect 39110 9220 39134 9222
rect 39190 9220 39214 9222
rect 39270 9220 39294 9222
rect 39350 9220 39356 9222
rect 39048 9210 39356 9220
rect 115246 9276 115554 9284
rect 115246 9274 115252 9276
rect 115308 9274 115332 9276
rect 115388 9274 115412 9276
rect 115468 9274 115492 9276
rect 115548 9274 115554 9276
rect 115308 9222 115310 9274
rect 115490 9222 115492 9274
rect 115246 9220 115252 9222
rect 115308 9220 115332 9222
rect 115388 9220 115412 9222
rect 115468 9220 115492 9222
rect 115548 9220 115554 9222
rect 115246 9210 115554 9220
rect 77148 8732 77456 8740
rect 77148 8730 77154 8732
rect 77210 8730 77234 8732
rect 77290 8730 77314 8732
rect 77370 8730 77394 8732
rect 77450 8730 77456 8732
rect 77210 8678 77212 8730
rect 77392 8678 77394 8730
rect 77148 8676 77154 8678
rect 77210 8676 77234 8678
rect 77290 8676 77314 8678
rect 77370 8676 77394 8678
rect 77450 8676 77456 8678
rect 77148 8666 77456 8676
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 8130 1440 8298
rect 39048 8188 39356 8196
rect 39048 8186 39054 8188
rect 39110 8186 39134 8188
rect 39190 8186 39214 8188
rect 39270 8186 39294 8188
rect 39350 8186 39356 8188
rect 39110 8134 39112 8186
rect 39292 8134 39294 8186
rect 39048 8132 39054 8134
rect 39110 8132 39134 8134
rect 39190 8132 39214 8134
rect 39270 8132 39294 8134
rect 39350 8132 39356 8134
rect 1398 8120 1454 8130
rect 39048 8122 39356 8132
rect 115246 8188 115554 8196
rect 115246 8186 115252 8188
rect 115308 8186 115332 8188
rect 115388 8186 115412 8188
rect 115468 8186 115492 8188
rect 115548 8186 115554 8188
rect 115308 8134 115310 8186
rect 115490 8134 115492 8186
rect 115246 8132 115252 8134
rect 115308 8132 115332 8134
rect 115388 8132 115412 8134
rect 115468 8132 115492 8134
rect 115548 8132 115554 8134
rect 115246 8122 115554 8132
rect 1398 8054 1454 8064
rect 77148 7644 77456 7652
rect 77148 7642 77154 7644
rect 77210 7642 77234 7644
rect 77290 7642 77314 7644
rect 77370 7642 77394 7644
rect 77450 7642 77456 7644
rect 77210 7590 77212 7642
rect 77392 7590 77394 7642
rect 77148 7588 77154 7590
rect 77210 7588 77234 7590
rect 77290 7588 77314 7590
rect 77370 7588 77394 7590
rect 77450 7588 77456 7590
rect 77148 7578 77456 7588
rect 39048 7100 39356 7108
rect 39048 7098 39054 7100
rect 39110 7098 39134 7100
rect 39190 7098 39214 7100
rect 39270 7098 39294 7100
rect 39350 7098 39356 7100
rect 39110 7046 39112 7098
rect 39292 7046 39294 7098
rect 39048 7044 39054 7046
rect 39110 7044 39134 7046
rect 39190 7044 39214 7046
rect 39270 7044 39294 7046
rect 39350 7044 39356 7046
rect 39048 7034 39356 7044
rect 115246 7100 115554 7108
rect 115246 7098 115252 7100
rect 115308 7098 115332 7100
rect 115388 7098 115412 7100
rect 115468 7098 115492 7100
rect 115548 7098 115554 7100
rect 115308 7046 115310 7098
rect 115490 7046 115492 7098
rect 115246 7044 115252 7046
rect 115308 7044 115332 7046
rect 115388 7044 115412 7046
rect 115468 7044 115492 7046
rect 115548 7044 115554 7046
rect 115246 7034 115554 7044
rect 77148 6556 77456 6564
rect 77148 6554 77154 6556
rect 77210 6554 77234 6556
rect 77290 6554 77314 6556
rect 77370 6554 77394 6556
rect 77450 6554 77456 6556
rect 77210 6502 77212 6554
rect 77392 6502 77394 6554
rect 77148 6500 77154 6502
rect 77210 6500 77234 6502
rect 77290 6500 77314 6502
rect 77370 6500 77394 6502
rect 77450 6500 77456 6502
rect 77148 6490 77456 6500
rect 39048 6012 39356 6020
rect 39048 6010 39054 6012
rect 39110 6010 39134 6012
rect 39190 6010 39214 6012
rect 39270 6010 39294 6012
rect 39350 6010 39356 6012
rect 39110 5958 39112 6010
rect 39292 5958 39294 6010
rect 39048 5956 39054 5958
rect 39110 5956 39134 5958
rect 39190 5956 39214 5958
rect 39270 5956 39294 5958
rect 39350 5956 39356 5958
rect 39048 5946 39356 5956
rect 115246 6012 115554 6020
rect 115246 6010 115252 6012
rect 115308 6010 115332 6012
rect 115388 6010 115412 6012
rect 115468 6010 115492 6012
rect 115548 6010 115554 6012
rect 115308 5958 115310 6010
rect 115490 5958 115492 6010
rect 115246 5956 115252 5958
rect 115308 5956 115332 5958
rect 115388 5956 115412 5958
rect 115468 5956 115492 5958
rect 115548 5956 115554 5958
rect 115246 5946 115554 5956
rect 77148 5468 77456 5476
rect 77148 5466 77154 5468
rect 77210 5466 77234 5468
rect 77290 5466 77314 5468
rect 77370 5466 77394 5468
rect 77450 5466 77456 5468
rect 77210 5414 77212 5466
rect 77392 5414 77394 5466
rect 77148 5412 77154 5414
rect 77210 5412 77234 5414
rect 77290 5412 77314 5414
rect 77370 5412 77394 5414
rect 77450 5412 77456 5414
rect 77148 5402 77456 5412
rect 39048 4924 39356 4932
rect 39048 4922 39054 4924
rect 39110 4922 39134 4924
rect 39190 4922 39214 4924
rect 39270 4922 39294 4924
rect 39350 4922 39356 4924
rect 39110 4870 39112 4922
rect 39292 4870 39294 4922
rect 39048 4868 39054 4870
rect 39110 4868 39134 4870
rect 39190 4868 39214 4870
rect 39270 4868 39294 4870
rect 39350 4868 39356 4870
rect 39048 4858 39356 4868
rect 115246 4924 115554 4932
rect 115246 4922 115252 4924
rect 115308 4922 115332 4924
rect 115388 4922 115412 4924
rect 115468 4922 115492 4924
rect 115548 4922 115554 4924
rect 115308 4870 115310 4922
rect 115490 4870 115492 4922
rect 115246 4868 115252 4870
rect 115308 4868 115332 4870
rect 115388 4868 115412 4870
rect 115468 4868 115492 4870
rect 115548 4868 115554 4870
rect 115246 4858 115554 4868
rect 77148 4380 77456 4388
rect 77148 4378 77154 4380
rect 77210 4378 77234 4380
rect 77290 4378 77314 4380
rect 77370 4378 77394 4380
rect 77450 4378 77456 4380
rect 77210 4326 77212 4378
rect 77392 4326 77394 4378
rect 77148 4324 77154 4326
rect 77210 4324 77234 4326
rect 77290 4324 77314 4326
rect 77370 4324 77394 4326
rect 77450 4324 77456 4326
rect 77148 4314 77456 4324
rect 39048 3836 39356 3844
rect 39048 3834 39054 3836
rect 39110 3834 39134 3836
rect 39190 3834 39214 3836
rect 39270 3834 39294 3836
rect 39350 3834 39356 3836
rect 39110 3782 39112 3834
rect 39292 3782 39294 3834
rect 39048 3780 39054 3782
rect 39110 3780 39134 3782
rect 39190 3780 39214 3782
rect 39270 3780 39294 3782
rect 39350 3780 39356 3782
rect 39048 3770 39356 3780
rect 115246 3836 115554 3844
rect 115246 3834 115252 3836
rect 115308 3834 115332 3836
rect 115388 3834 115412 3836
rect 115468 3834 115492 3836
rect 115548 3834 115554 3836
rect 115308 3782 115310 3834
rect 115490 3782 115492 3834
rect 115246 3780 115252 3782
rect 115308 3780 115332 3782
rect 115388 3780 115412 3782
rect 115468 3780 115492 3782
rect 115548 3780 115554 3782
rect 115246 3770 115554 3780
rect 77148 3292 77456 3300
rect 77148 3290 77154 3292
rect 77210 3290 77234 3292
rect 77290 3290 77314 3292
rect 77370 3290 77394 3292
rect 77450 3290 77456 3292
rect 77210 3238 77212 3290
rect 77392 3238 77394 3290
rect 77148 3236 77154 3238
rect 77210 3236 77234 3238
rect 77290 3236 77314 3238
rect 77370 3236 77394 3238
rect 77450 3236 77456 3238
rect 77148 3226 77456 3236
rect 39048 2748 39356 2756
rect 39048 2746 39054 2748
rect 39110 2746 39134 2748
rect 39190 2746 39214 2748
rect 39270 2746 39294 2748
rect 39350 2746 39356 2748
rect 39110 2694 39112 2746
rect 39292 2694 39294 2746
rect 39048 2692 39054 2694
rect 39110 2692 39134 2694
rect 39190 2692 39214 2694
rect 39270 2692 39294 2694
rect 39350 2692 39356 2694
rect 39048 2682 39356 2692
rect 115246 2748 115554 2756
rect 115246 2746 115252 2748
rect 115308 2746 115332 2748
rect 115388 2746 115412 2748
rect 115468 2746 115492 2748
rect 115548 2746 115554 2748
rect 115308 2694 115310 2746
rect 115490 2694 115492 2746
rect 115246 2692 115252 2694
rect 115308 2692 115332 2694
rect 115388 2692 115412 2694
rect 115468 2692 115492 2694
rect 115548 2692 115554 2694
rect 115246 2682 115554 2692
rect 149440 2650 149468 12174
rect 149520 12096 149572 12102
rect 149520 12038 149572 12044
rect 149532 11014 149560 12038
rect 149992 11830 150020 12582
rect 149980 11824 150032 11830
rect 149980 11766 150032 11772
rect 149520 11008 149572 11014
rect 149520 10950 149572 10956
rect 150360 10674 150388 12650
rect 150820 11354 150848 13466
rect 151084 13252 151136 13258
rect 151084 13194 151136 13200
rect 151096 11898 151124 13194
rect 151544 12776 151596 12782
rect 151544 12718 151596 12724
rect 151268 12640 151320 12646
rect 151268 12582 151320 12588
rect 151360 12640 151412 12646
rect 151360 12582 151412 12588
rect 151084 11892 151136 11898
rect 151084 11834 151136 11840
rect 151280 11762 151308 12582
rect 151372 12238 151400 12582
rect 151360 12232 151412 12238
rect 151360 12174 151412 12180
rect 151556 12186 151584 12718
rect 151636 12708 151688 12714
rect 151636 12650 151688 12656
rect 151648 12374 151676 12650
rect 151636 12368 151688 12374
rect 151636 12310 151688 12316
rect 151268 11756 151320 11762
rect 151268 11698 151320 11704
rect 150808 11348 150860 11354
rect 150808 11290 150860 11296
rect 151372 11218 151400 12174
rect 151556 12158 151768 12186
rect 151740 12102 151768 12158
rect 151636 12096 151688 12102
rect 151636 12038 151688 12044
rect 151728 12096 151780 12102
rect 151728 12038 151780 12044
rect 151360 11212 151412 11218
rect 151360 11154 151412 11160
rect 151648 10742 151676 12038
rect 151740 11558 151768 12038
rect 152016 11898 152044 15286
rect 154946 15200 155002 16000
rect 157982 15200 158038 16000
rect 161110 15314 161166 16000
rect 161110 15286 161336 15314
rect 161110 15200 161166 15286
rect 154960 13462 154988 15200
rect 157156 13728 157208 13734
rect 157156 13670 157208 13676
rect 154948 13456 155000 13462
rect 154948 13398 155000 13404
rect 155224 13320 155276 13326
rect 155224 13262 155276 13268
rect 155868 13320 155920 13326
rect 155868 13262 155920 13268
rect 156420 13320 156472 13326
rect 156420 13262 156472 13268
rect 152464 13252 152516 13258
rect 152464 13194 152516 13200
rect 153752 13252 153804 13258
rect 153752 13194 153804 13200
rect 154212 13252 154264 13258
rect 154212 13194 154264 13200
rect 152476 12442 152504 13194
rect 152648 13184 152700 13190
rect 152648 13126 152700 13132
rect 152660 12986 152688 13126
rect 153346 13084 153654 13092
rect 153346 13082 153352 13084
rect 153408 13082 153432 13084
rect 153488 13082 153512 13084
rect 153568 13082 153592 13084
rect 153648 13082 153654 13084
rect 153408 13030 153410 13082
rect 153590 13030 153592 13082
rect 153346 13028 153352 13030
rect 153408 13028 153432 13030
rect 153488 13028 153512 13030
rect 153568 13028 153592 13030
rect 153648 13028 153654 13030
rect 153346 13018 153654 13028
rect 152648 12980 152700 12986
rect 152648 12922 152700 12928
rect 152832 12980 152884 12986
rect 152832 12922 152884 12928
rect 152660 12832 152688 12922
rect 152568 12804 152688 12832
rect 152464 12436 152516 12442
rect 152464 12378 152516 12384
rect 152568 12102 152596 12804
rect 152740 12776 152792 12782
rect 152740 12718 152792 12724
rect 152752 12374 152780 12718
rect 152844 12714 152872 12922
rect 152832 12708 152884 12714
rect 152832 12650 152884 12656
rect 153108 12708 153160 12714
rect 153108 12650 153160 12656
rect 152740 12368 152792 12374
rect 152740 12310 152792 12316
rect 152188 12096 152240 12102
rect 152188 12038 152240 12044
rect 152556 12096 152608 12102
rect 152556 12038 152608 12044
rect 152004 11892 152056 11898
rect 152004 11834 152056 11840
rect 152200 11762 152228 12038
rect 152752 11762 152780 12310
rect 152188 11756 152240 11762
rect 152188 11698 152240 11704
rect 152740 11756 152792 11762
rect 152740 11698 152792 11704
rect 151728 11552 151780 11558
rect 151728 11494 151780 11500
rect 153120 11150 153148 12650
rect 153764 12442 153792 13194
rect 154120 12640 154172 12646
rect 154120 12582 154172 12588
rect 153752 12436 153804 12442
rect 153752 12378 153804 12384
rect 154132 12306 154160 12582
rect 154120 12300 154172 12306
rect 154120 12242 154172 12248
rect 153346 11996 153654 12004
rect 153346 11994 153352 11996
rect 153408 11994 153432 11996
rect 153488 11994 153512 11996
rect 153568 11994 153592 11996
rect 153648 11994 153654 11996
rect 153408 11942 153410 11994
rect 153590 11942 153592 11994
rect 153346 11940 153352 11942
rect 153408 11940 153432 11942
rect 153488 11940 153512 11942
rect 153568 11940 153592 11942
rect 153648 11940 153654 11942
rect 153346 11930 153654 11940
rect 154224 11898 154252 13194
rect 155236 13190 155264 13262
rect 155224 13184 155276 13190
rect 155224 13126 155276 13132
rect 155038 12880 155094 12888
rect 155880 12850 155908 13262
rect 155038 12814 155094 12824
rect 155868 12844 155920 12850
rect 155052 12782 155080 12814
rect 155868 12786 155920 12792
rect 155040 12776 155092 12782
rect 155040 12718 155092 12724
rect 155052 12374 155080 12718
rect 155040 12368 155092 12374
rect 155040 12310 155092 12316
rect 155880 12170 155908 12786
rect 156432 12170 156460 13262
rect 156604 13252 156656 13258
rect 156604 13194 156656 13200
rect 156616 12918 156644 13194
rect 157168 12986 157196 13670
rect 157996 13530 158024 15200
rect 157248 13524 157300 13530
rect 157248 13466 157300 13472
rect 157984 13524 158036 13530
rect 157984 13466 158036 13472
rect 159456 13524 159508 13530
rect 159456 13466 159508 13472
rect 157156 12980 157208 12986
rect 157156 12922 157208 12928
rect 156604 12912 156656 12918
rect 156604 12854 156656 12860
rect 157260 12442 157288 13466
rect 157800 13320 157852 13326
rect 157800 13262 157852 13268
rect 158628 13320 158680 13326
rect 158628 13262 158680 13268
rect 157812 12850 157840 13262
rect 158640 12986 158668 13262
rect 158904 13252 158956 13258
rect 158904 13194 158956 13200
rect 158628 12980 158680 12986
rect 158628 12922 158680 12928
rect 157800 12844 157852 12850
rect 157800 12786 157852 12792
rect 157892 12640 157944 12646
rect 157890 12608 157892 12616
rect 157944 12608 157946 12616
rect 157890 12542 157946 12552
rect 157248 12436 157300 12442
rect 157248 12378 157300 12384
rect 155868 12164 155920 12170
rect 155868 12106 155920 12112
rect 156420 12164 156472 12170
rect 156420 12106 156472 12112
rect 154212 11892 154264 11898
rect 154212 11834 154264 11840
rect 156432 11286 156460 12106
rect 157260 11354 157288 12378
rect 157248 11348 157300 11354
rect 157248 11290 157300 11296
rect 156420 11280 156472 11286
rect 156420 11222 156472 11228
rect 153108 11144 153160 11150
rect 153108 11086 153160 11092
rect 156144 11076 156196 11082
rect 156144 11018 156196 11024
rect 153346 10908 153654 10916
rect 153346 10906 153352 10908
rect 153408 10906 153432 10908
rect 153488 10906 153512 10908
rect 153568 10906 153592 10908
rect 153648 10906 153654 10908
rect 153408 10854 153410 10906
rect 153590 10854 153592 10906
rect 153346 10852 153352 10854
rect 153408 10852 153432 10854
rect 153488 10852 153512 10854
rect 153568 10852 153592 10854
rect 153648 10852 153654 10854
rect 153346 10842 153654 10852
rect 156156 10742 156184 11018
rect 151636 10736 151688 10742
rect 151636 10678 151688 10684
rect 156144 10736 156196 10742
rect 156144 10678 156196 10684
rect 150348 10668 150400 10674
rect 150348 10610 150400 10616
rect 156156 10062 156184 10678
rect 156144 10056 156196 10062
rect 156144 9998 156196 10004
rect 153346 9820 153654 9828
rect 153346 9818 153352 9820
rect 153408 9818 153432 9820
rect 153488 9818 153512 9820
rect 153568 9818 153592 9820
rect 153648 9818 153654 9820
rect 153408 9766 153410 9818
rect 153590 9766 153592 9818
rect 153346 9764 153352 9766
rect 153408 9764 153432 9766
rect 153488 9764 153512 9766
rect 153568 9764 153592 9766
rect 153648 9764 153654 9766
rect 153346 9754 153654 9764
rect 156156 9654 156184 9998
rect 158640 9654 158668 12922
rect 158812 12708 158864 12714
rect 158812 12650 158864 12656
rect 158824 12238 158852 12650
rect 158916 12374 158944 13194
rect 159468 12782 159496 13466
rect 160928 13388 160980 13394
rect 160928 13330 160980 13336
rect 159548 13184 159600 13190
rect 159548 13126 159600 13132
rect 160376 13184 160428 13190
rect 160376 13126 160428 13132
rect 159560 12782 159588 13126
rect 160388 12918 160416 13126
rect 160376 12912 160428 12918
rect 160376 12854 160428 12860
rect 159456 12776 159508 12782
rect 159456 12718 159508 12724
rect 159548 12776 159600 12782
rect 159548 12718 159600 12724
rect 160284 12640 160336 12646
rect 160282 12608 160284 12616
rect 160336 12608 160338 12616
rect 160282 12542 160338 12552
rect 158904 12368 158956 12374
rect 158904 12310 158956 12316
rect 160388 12306 160416 12854
rect 160940 12442 160968 13330
rect 161204 13252 161256 13258
rect 161204 13194 161256 13200
rect 160928 12436 160980 12442
rect 160928 12378 160980 12384
rect 160376 12300 160428 12306
rect 160376 12242 160428 12248
rect 158812 12232 158864 12238
rect 158812 12174 158864 12180
rect 161112 12096 161164 12102
rect 161112 12038 161164 12044
rect 161124 11762 161152 12038
rect 161112 11756 161164 11762
rect 161112 11698 161164 11704
rect 161216 11626 161244 13194
rect 161308 11626 161336 15286
rect 164146 15200 164202 16000
rect 167182 15200 167238 16000
rect 170310 15314 170366 16000
rect 173346 15314 173402 16000
rect 170310 15286 170444 15314
rect 170310 15200 170366 15286
rect 161664 13796 161716 13802
rect 161664 13738 161716 13744
rect 161572 13524 161624 13530
rect 161492 13484 161572 13512
rect 161492 12306 161520 13484
rect 161572 13466 161624 13472
rect 161676 12850 161704 13738
rect 162676 13524 162728 13530
rect 162676 13466 162728 13472
rect 163504 13524 163556 13530
rect 163504 13466 163556 13472
rect 162688 13326 162716 13466
rect 163516 13326 163544 13466
rect 162676 13320 162728 13326
rect 162676 13262 162728 13268
rect 163504 13320 163556 13326
rect 163504 13262 163556 13268
rect 162032 13184 162084 13190
rect 162032 13126 162084 13132
rect 162492 13184 162544 13190
rect 162492 13126 162544 13132
rect 161664 12844 161716 12850
rect 161664 12786 161716 12792
rect 161572 12776 161624 12782
rect 161572 12718 161624 12724
rect 161584 12442 161612 12718
rect 161572 12436 161624 12442
rect 161572 12378 161624 12384
rect 161480 12300 161532 12306
rect 161480 12242 161532 12248
rect 161756 12232 161808 12238
rect 161756 12174 161808 12180
rect 161768 11762 161796 12174
rect 162044 11898 162072 13126
rect 162124 12776 162176 12782
rect 162124 12718 162176 12724
rect 162032 11892 162084 11898
rect 162032 11834 162084 11840
rect 161756 11756 161808 11762
rect 161756 11698 161808 11704
rect 161204 11620 161256 11626
rect 161204 11562 161256 11568
rect 161296 11620 161348 11626
rect 161296 11562 161348 11568
rect 162136 11354 162164 12718
rect 162504 12306 162532 13126
rect 162688 12306 162716 13262
rect 162768 13252 162820 13258
rect 162768 13194 162820 13200
rect 162492 12300 162544 12306
rect 162492 12242 162544 12248
rect 162676 12300 162728 12306
rect 162676 12242 162728 12248
rect 162584 12164 162636 12170
rect 162584 12106 162636 12112
rect 162676 12164 162728 12170
rect 162676 12106 162728 12112
rect 162216 12096 162268 12102
rect 162216 12038 162268 12044
rect 162124 11348 162176 11354
rect 162124 11290 162176 11296
rect 162228 11150 162256 12038
rect 162596 11830 162624 12106
rect 162584 11824 162636 11830
rect 162584 11766 162636 11772
rect 162688 11354 162716 12106
rect 162780 11898 162808 13194
rect 163516 12986 163544 13262
rect 163780 13252 163832 13258
rect 163780 13194 163832 13200
rect 163504 12980 163556 12986
rect 163504 12922 163556 12928
rect 163412 12912 163464 12918
rect 163412 12854 163464 12860
rect 162860 12776 162912 12782
rect 162860 12718 162912 12724
rect 162872 12102 162900 12718
rect 162860 12096 162912 12102
rect 162860 12038 162912 12044
rect 162768 11892 162820 11898
rect 162768 11834 162820 11840
rect 163424 11354 163452 12854
rect 163688 12640 163740 12646
rect 163688 12582 163740 12588
rect 163594 12336 163650 12344
rect 163594 12270 163596 12280
rect 163648 12270 163650 12280
rect 163596 12242 163648 12248
rect 163504 11688 163556 11694
rect 163504 11630 163556 11636
rect 162676 11348 162728 11354
rect 162676 11290 162728 11296
rect 163412 11348 163464 11354
rect 163412 11290 163464 11296
rect 163516 11150 163544 11630
rect 162216 11144 162268 11150
rect 162216 11086 162268 11092
rect 163504 11144 163556 11150
rect 163504 11086 163556 11092
rect 163608 10130 163636 12242
rect 163700 11762 163728 12582
rect 163792 11898 163820 13194
rect 164160 12730 164188 15200
rect 166080 13796 166132 13802
rect 166080 13738 166132 13744
rect 165252 13388 165304 13394
rect 165252 13330 165304 13336
rect 164884 13320 164936 13326
rect 165264 13274 165292 13330
rect 164884 13262 164936 13268
rect 164608 13184 164660 13190
rect 164608 13126 164660 13132
rect 164620 12782 164648 13126
rect 164608 12776 164660 12782
rect 164160 12714 164280 12730
rect 164608 12718 164660 12724
rect 164160 12708 164292 12714
rect 164160 12702 164240 12708
rect 164240 12650 164292 12656
rect 164332 12164 164384 12170
rect 164332 12106 164384 12112
rect 164344 11898 164372 12106
rect 164896 11898 164924 13262
rect 165172 13258 165292 13274
rect 165160 13252 165292 13258
rect 165212 13246 165292 13252
rect 165160 13194 165212 13200
rect 165252 13184 165304 13190
rect 165252 13126 165304 13132
rect 165344 13184 165396 13190
rect 165344 13126 165396 13132
rect 165264 12986 165292 13126
rect 165252 12980 165304 12986
rect 165252 12922 165304 12928
rect 163780 11892 163832 11898
rect 163780 11834 163832 11840
rect 164332 11892 164384 11898
rect 164332 11834 164384 11840
rect 164884 11892 164936 11898
rect 164884 11834 164936 11840
rect 163688 11756 163740 11762
rect 163688 11698 163740 11704
rect 165356 11218 165384 13126
rect 165436 12844 165488 12850
rect 165436 12786 165488 12792
rect 165448 12374 165476 12786
rect 166092 12374 166120 13738
rect 166448 13456 166500 13462
rect 166448 13398 166500 13404
rect 166460 13190 166488 13398
rect 166448 13184 166500 13190
rect 166448 13126 166500 13132
rect 166172 12844 166224 12850
rect 166172 12786 166224 12792
rect 166184 12646 166212 12786
rect 166172 12640 166224 12646
rect 166172 12582 166224 12588
rect 166460 12442 166488 13126
rect 167196 12986 167224 15200
rect 167368 13796 167420 13802
rect 167368 13738 167420 13744
rect 167380 13258 167408 13738
rect 170416 13462 170444 15286
rect 173084 15286 173402 15314
rect 173084 13462 173112 15286
rect 173346 15200 173402 15286
rect 176474 15200 176530 16000
rect 179510 15200 179566 16000
rect 182546 15314 182602 16000
rect 185674 15314 185730 16000
rect 182546 15286 182772 15314
rect 182546 15200 182602 15286
rect 174176 13796 174228 13802
rect 174176 13738 174228 13744
rect 170404 13456 170456 13462
rect 170404 13398 170456 13404
rect 173072 13456 173124 13462
rect 173072 13398 173124 13404
rect 173808 13456 173860 13462
rect 173808 13398 173860 13404
rect 167368 13252 167420 13258
rect 167368 13194 167420 13200
rect 167184 12980 167236 12986
rect 167184 12922 167236 12928
rect 173820 12918 173848 13398
rect 174188 13326 174216 13738
rect 175844 13518 176056 13546
rect 175844 13326 175872 13518
rect 176028 13462 176056 13518
rect 176384 13524 176436 13530
rect 176384 13466 176436 13472
rect 175924 13456 175976 13462
rect 175924 13398 175976 13404
rect 176016 13456 176068 13462
rect 176016 13398 176068 13404
rect 174176 13320 174228 13326
rect 174176 13262 174228 13268
rect 175832 13320 175884 13326
rect 175832 13262 175884 13268
rect 175740 13252 175792 13258
rect 175740 13194 175792 13200
rect 175004 13184 175056 13190
rect 175004 13126 175056 13132
rect 175016 12986 175044 13126
rect 175752 12986 175780 13194
rect 175004 12980 175056 12986
rect 175004 12922 175056 12928
rect 175740 12980 175792 12986
rect 175740 12922 175792 12928
rect 175936 12918 175964 13398
rect 176396 13326 176424 13466
rect 176384 13320 176436 13326
rect 176384 13262 176436 13268
rect 176396 12986 176424 13262
rect 176384 12980 176436 12986
rect 176384 12922 176436 12928
rect 173808 12912 173860 12918
rect 173808 12854 173860 12860
rect 175924 12912 175976 12918
rect 175924 12854 175976 12860
rect 176396 12850 176424 12922
rect 166540 12844 166592 12850
rect 166540 12786 166592 12792
rect 176384 12844 176436 12850
rect 176384 12786 176436 12792
rect 166448 12436 166500 12442
rect 166448 12378 166500 12384
rect 165436 12368 165488 12374
rect 165436 12310 165488 12316
rect 166080 12368 166132 12374
rect 166080 12310 166132 12316
rect 165448 11286 165476 12310
rect 166552 12170 166580 12786
rect 166632 12640 166684 12646
rect 166632 12582 166684 12588
rect 165896 12164 165948 12170
rect 165896 12106 165948 12112
rect 166540 12164 166592 12170
rect 166540 12106 166592 12112
rect 165908 11626 165936 12106
rect 166644 11762 166672 12582
rect 176488 12442 176516 15200
rect 177764 13796 177816 13802
rect 177764 13738 177816 13744
rect 177776 13462 177804 13738
rect 177764 13456 177816 13462
rect 177764 13398 177816 13404
rect 177672 13252 177724 13258
rect 177672 13194 177724 13200
rect 176936 12912 176988 12918
rect 176936 12854 176988 12860
rect 176752 12776 176804 12782
rect 176752 12718 176804 12724
rect 176476 12436 176528 12442
rect 176476 12378 176528 12384
rect 176660 12096 176712 12102
rect 176660 12038 176712 12044
rect 176672 11762 176700 12038
rect 176764 11898 176792 12718
rect 176948 12458 176976 12854
rect 177396 12640 177448 12646
rect 177396 12582 177448 12588
rect 176948 12430 177160 12458
rect 177132 12306 177160 12430
rect 177120 12300 177172 12306
rect 177120 12242 177172 12248
rect 176752 11892 176804 11898
rect 176752 11834 176804 11840
rect 166632 11756 166684 11762
rect 166632 11698 166684 11704
rect 176660 11756 176712 11762
rect 176660 11698 176712 11704
rect 177132 11694 177160 12242
rect 177408 11898 177436 12582
rect 177396 11892 177448 11898
rect 177396 11834 177448 11840
rect 177120 11688 177172 11694
rect 177120 11630 177172 11636
rect 165896 11620 165948 11626
rect 165896 11562 165948 11568
rect 165908 11354 165936 11562
rect 165896 11348 165948 11354
rect 165896 11290 165948 11296
rect 165436 11280 165488 11286
rect 165436 11222 165488 11228
rect 177684 11218 177712 13194
rect 177776 12374 177804 13398
rect 177948 12912 178000 12918
rect 177948 12854 178000 12860
rect 177856 12640 177908 12646
rect 177856 12582 177908 12588
rect 177764 12368 177816 12374
rect 177764 12310 177816 12316
rect 177868 12238 177896 12582
rect 177856 12232 177908 12238
rect 177856 12174 177908 12180
rect 177868 11898 177896 12174
rect 177856 11892 177908 11898
rect 177856 11834 177908 11840
rect 177960 11218 177988 12854
rect 179524 12442 179552 15200
rect 181904 13796 181956 13802
rect 181904 13738 181956 13744
rect 180432 13456 180484 13462
rect 180432 13398 180484 13404
rect 179972 13252 180024 13258
rect 179972 13194 180024 13200
rect 179880 12640 179932 12646
rect 179880 12582 179932 12588
rect 179512 12436 179564 12442
rect 179512 12378 179564 12384
rect 179144 12232 179196 12238
rect 179144 12174 179196 12180
rect 178040 12096 178092 12102
rect 178040 12038 178092 12044
rect 165344 11212 165396 11218
rect 165344 11154 165396 11160
rect 177672 11212 177724 11218
rect 177672 11154 177724 11160
rect 177948 11212 178000 11218
rect 177948 11154 178000 11160
rect 178052 11150 178080 12038
rect 178040 11144 178092 11150
rect 178040 11086 178092 11092
rect 179156 10470 179184 12174
rect 179420 12164 179472 12170
rect 179420 12106 179472 12112
rect 179432 11082 179460 12106
rect 179892 11898 179920 12582
rect 179984 11898 180012 13194
rect 180156 12980 180208 12986
rect 180156 12922 180208 12928
rect 180248 12980 180300 12986
rect 180248 12922 180300 12928
rect 180168 12782 180196 12922
rect 180156 12776 180208 12782
rect 180156 12718 180208 12724
rect 180260 12714 180288 12922
rect 180340 12844 180392 12850
rect 180340 12786 180392 12792
rect 180248 12708 180300 12714
rect 180248 12650 180300 12656
rect 180156 12096 180208 12102
rect 180156 12038 180208 12044
rect 180168 11898 180196 12038
rect 179880 11892 179932 11898
rect 179880 11834 179932 11840
rect 179972 11892 180024 11898
rect 179972 11834 180024 11840
rect 180156 11892 180208 11898
rect 180156 11834 180208 11840
rect 179880 11756 179932 11762
rect 180064 11756 180116 11762
rect 179932 11716 180064 11744
rect 179880 11698 179932 11704
rect 180064 11698 180116 11704
rect 180352 11626 180380 12786
rect 180340 11620 180392 11626
rect 180340 11562 180392 11568
rect 180444 11150 180472 13398
rect 181916 13394 181944 13738
rect 182744 13530 182772 15286
rect 185674 15286 185808 15314
rect 185674 15200 185730 15286
rect 185780 13530 185808 15286
rect 188710 15200 188766 16000
rect 191746 15314 191802 16000
rect 191300 15286 191802 15314
rect 182732 13524 182784 13530
rect 182732 13466 182784 13472
rect 185768 13524 185820 13530
rect 185768 13466 185820 13472
rect 181904 13388 181956 13394
rect 181904 13330 181956 13336
rect 182088 13388 182140 13394
rect 182088 13330 182140 13336
rect 188528 13388 188580 13394
rect 188528 13330 188580 13336
rect 180616 13320 180668 13326
rect 180616 13262 180668 13268
rect 180524 12708 180576 12714
rect 180524 12650 180576 12656
rect 180536 11558 180564 12650
rect 180628 12646 180656 13262
rect 180892 13252 180944 13258
rect 180892 13194 180944 13200
rect 180708 13184 180760 13190
rect 180708 13126 180760 13132
rect 180616 12640 180668 12646
rect 180616 12582 180668 12588
rect 180720 12238 180748 13126
rect 180904 12374 180932 13194
rect 181536 12844 181588 12850
rect 181536 12786 181588 12792
rect 181444 12640 181496 12646
rect 181444 12582 181496 12588
rect 180892 12368 180944 12374
rect 180892 12310 180944 12316
rect 180708 12232 180760 12238
rect 180708 12174 180760 12180
rect 180616 11756 180668 11762
rect 180720 11744 180748 12174
rect 181456 12170 181484 12582
rect 181444 12164 181496 12170
rect 181444 12106 181496 12112
rect 180668 11716 180748 11744
rect 180616 11698 180668 11704
rect 181548 11694 181576 12786
rect 182100 12714 182128 13330
rect 187792 13184 187844 13190
rect 187792 13126 187844 13132
rect 187976 13184 188028 13190
rect 187976 13126 188028 13132
rect 188344 13184 188396 13190
rect 188344 13126 188396 13132
rect 182088 12708 182140 12714
rect 182088 12650 182140 12656
rect 187804 12646 187832 13126
rect 187792 12640 187844 12646
rect 187792 12582 187844 12588
rect 187988 12306 188016 13126
rect 188356 12986 188384 13126
rect 188344 12980 188396 12986
rect 188344 12922 188396 12928
rect 188540 12918 188568 13330
rect 188528 12912 188580 12918
rect 188528 12854 188580 12860
rect 188344 12844 188396 12850
rect 188344 12786 188396 12792
rect 187976 12300 188028 12306
rect 187976 12242 188028 12248
rect 188356 11898 188384 12786
rect 188620 12708 188672 12714
rect 188724 12696 188752 15200
rect 189908 13864 189960 13870
rect 189908 13806 189960 13812
rect 189356 13796 189408 13802
rect 189356 13738 189408 13744
rect 189368 13530 189396 13738
rect 189356 13524 189408 13530
rect 189356 13466 189408 13472
rect 188804 13456 188856 13462
rect 188804 13398 188856 13404
rect 188816 12850 188844 13398
rect 189368 12850 189396 13466
rect 189540 13456 189592 13462
rect 189592 13416 189672 13444
rect 189540 13398 189592 13404
rect 189540 13320 189592 13326
rect 189540 13262 189592 13268
rect 189552 13190 189580 13262
rect 189540 13184 189592 13190
rect 189540 13126 189592 13132
rect 188804 12844 188856 12850
rect 188804 12786 188856 12792
rect 189356 12844 189408 12850
rect 189356 12786 189408 12792
rect 189552 12782 189580 13126
rect 189540 12776 189592 12782
rect 189540 12718 189592 12724
rect 188672 12668 188752 12696
rect 189172 12708 189224 12714
rect 188620 12650 188672 12656
rect 189172 12650 189224 12656
rect 188988 12640 189040 12646
rect 188988 12582 189040 12588
rect 188344 11892 188396 11898
rect 188344 11834 188396 11840
rect 180800 11688 180852 11694
rect 180800 11630 180852 11636
rect 181536 11688 181588 11694
rect 181536 11630 181588 11636
rect 180524 11552 180576 11558
rect 180524 11494 180576 11500
rect 180812 11218 180840 11630
rect 180800 11212 180852 11218
rect 180800 11154 180852 11160
rect 189000 11150 189028 12582
rect 189184 12442 189212 12650
rect 189644 12442 189672 13416
rect 189920 13394 189948 13806
rect 190920 13524 190972 13530
rect 190920 13466 190972 13472
rect 189908 13388 189960 13394
rect 189908 13330 189960 13336
rect 190932 12918 190960 13466
rect 190920 12912 190972 12918
rect 190920 12854 190972 12860
rect 190552 12640 190604 12646
rect 190552 12582 190604 12588
rect 189172 12436 189224 12442
rect 189172 12378 189224 12384
rect 189632 12436 189684 12442
rect 189632 12378 189684 12384
rect 189540 12232 189592 12238
rect 189540 12174 189592 12180
rect 189552 11830 189580 12174
rect 189540 11824 189592 11830
rect 189540 11766 189592 11772
rect 189630 11792 189686 11800
rect 189630 11726 189632 11736
rect 189684 11726 189686 11736
rect 189632 11698 189684 11704
rect 189448 11552 189500 11558
rect 189448 11494 189500 11500
rect 180432 11144 180484 11150
rect 180432 11086 180484 11092
rect 188988 11144 189040 11150
rect 188988 11086 189040 11092
rect 189460 11082 189488 11494
rect 179420 11076 179472 11082
rect 179420 11018 179472 11024
rect 189448 11076 189500 11082
rect 189448 11018 189500 11024
rect 190564 10674 190592 12582
rect 190828 12436 190880 12442
rect 190828 12378 190880 12384
rect 190840 12170 190868 12378
rect 190828 12164 190880 12170
rect 190828 12106 190880 12112
rect 191104 12164 191156 12170
rect 191104 12106 191156 12112
rect 191196 12164 191248 12170
rect 191196 12106 191248 12112
rect 190828 11756 190880 11762
rect 190828 11698 190880 11704
rect 190840 11150 190868 11698
rect 190644 11144 190696 11150
rect 190644 11086 190696 11092
rect 190828 11144 190880 11150
rect 190828 11086 190880 11092
rect 190552 10668 190604 10674
rect 190552 10610 190604 10616
rect 187516 10600 187568 10606
rect 187516 10542 187568 10548
rect 179144 10464 179196 10470
rect 179144 10406 179196 10412
rect 163596 10124 163648 10130
rect 163596 10066 163648 10072
rect 156144 9648 156196 9654
rect 156144 9590 156196 9596
rect 158628 9648 158680 9654
rect 158628 9590 158680 9596
rect 153346 8732 153654 8740
rect 153346 8730 153352 8732
rect 153408 8730 153432 8732
rect 153488 8730 153512 8732
rect 153568 8730 153592 8732
rect 153648 8730 153654 8732
rect 153408 8678 153410 8730
rect 153590 8678 153592 8730
rect 153346 8676 153352 8678
rect 153408 8676 153432 8678
rect 153488 8676 153512 8678
rect 153568 8676 153592 8678
rect 153648 8676 153654 8678
rect 153346 8666 153654 8676
rect 187528 8362 187556 10542
rect 190656 9654 190684 11086
rect 191116 10810 191144 12106
rect 191208 11218 191236 12106
rect 191196 11212 191248 11218
rect 191196 11154 191248 11160
rect 191104 10804 191156 10810
rect 191104 10746 191156 10752
rect 191300 10266 191328 15286
rect 191746 15200 191802 15286
rect 194874 15314 194930 16000
rect 197910 15314 197966 16000
rect 201038 15314 201094 16000
rect 194874 15286 195284 15314
rect 194874 15200 194930 15286
rect 193220 13796 193272 13802
rect 193220 13738 193272 13744
rect 191444 13628 191752 13636
rect 191444 13626 191450 13628
rect 191506 13626 191530 13628
rect 191586 13626 191610 13628
rect 191666 13626 191690 13628
rect 191746 13626 191752 13628
rect 191506 13574 191508 13626
rect 191688 13574 191690 13626
rect 191444 13572 191450 13574
rect 191506 13572 191530 13574
rect 191586 13572 191610 13574
rect 191666 13572 191690 13574
rect 191746 13572 191752 13574
rect 191444 13562 191752 13572
rect 191840 13456 191892 13462
rect 191840 13398 191892 13404
rect 191380 13184 191432 13190
rect 191380 13126 191432 13132
rect 191392 12986 191420 13126
rect 191380 12980 191432 12986
rect 191380 12922 191432 12928
rect 191748 12912 191800 12918
rect 191748 12854 191800 12860
rect 191760 12714 191788 12854
rect 191748 12708 191800 12714
rect 191748 12650 191800 12656
rect 191852 12616 191880 13398
rect 192392 13252 192444 13258
rect 192392 13194 192444 13200
rect 191932 12708 191984 12714
rect 191932 12650 191984 12656
rect 192036 12702 192340 12730
rect 191838 12608 191894 12616
rect 191444 12540 191752 12548
rect 191838 12542 191894 12552
rect 191444 12538 191450 12540
rect 191506 12538 191530 12540
rect 191586 12538 191610 12540
rect 191666 12538 191690 12540
rect 191746 12538 191752 12540
rect 191506 12486 191508 12538
rect 191688 12486 191690 12538
rect 191444 12484 191450 12486
rect 191506 12484 191530 12486
rect 191586 12484 191610 12486
rect 191666 12484 191690 12486
rect 191746 12484 191752 12486
rect 191444 12474 191752 12484
rect 191944 12434 191972 12650
rect 192036 12646 192064 12702
rect 192024 12640 192076 12646
rect 192024 12582 192076 12588
rect 192116 12640 192168 12646
rect 192116 12582 192168 12588
rect 192206 12608 192262 12616
rect 192128 12434 192156 12582
rect 192206 12542 192262 12552
rect 191760 12406 191972 12434
rect 192036 12406 192156 12434
rect 191760 11898 191788 12406
rect 191840 12300 191892 12306
rect 191840 12242 191892 12248
rect 191852 11898 191880 12242
rect 191748 11892 191800 11898
rect 191748 11834 191800 11840
rect 191840 11892 191892 11898
rect 191840 11834 191892 11840
rect 191852 11762 191880 11834
rect 191840 11756 191892 11762
rect 191840 11698 191892 11704
rect 191444 11452 191752 11460
rect 191444 11450 191450 11452
rect 191506 11450 191530 11452
rect 191586 11450 191610 11452
rect 191666 11450 191690 11452
rect 191746 11450 191752 11452
rect 191506 11398 191508 11450
rect 191688 11398 191690 11450
rect 191444 11396 191450 11398
rect 191506 11396 191530 11398
rect 191586 11396 191610 11398
rect 191666 11396 191690 11398
rect 191746 11396 191752 11398
rect 191444 11386 191752 11396
rect 191852 11218 191880 11698
rect 192036 11234 192064 12406
rect 192116 11688 192168 11694
rect 192116 11630 192168 11636
rect 191840 11212 191892 11218
rect 191840 11154 191892 11160
rect 191944 11206 192064 11234
rect 191944 11150 191972 11206
rect 191932 11144 191984 11150
rect 191932 11086 191984 11092
rect 192128 10538 192156 11630
rect 192220 10742 192248 12542
rect 192208 10736 192260 10742
rect 192208 10678 192260 10684
rect 192312 10674 192340 12702
rect 192404 12434 192432 13194
rect 192484 12980 192536 12986
rect 192484 12922 192536 12928
rect 192496 12714 192524 12922
rect 192576 12844 192628 12850
rect 192576 12786 192628 12792
rect 192484 12708 192536 12714
rect 192484 12650 192536 12656
rect 192404 12406 192524 12434
rect 192300 10668 192352 10674
rect 192300 10610 192352 10616
rect 192116 10532 192168 10538
rect 192116 10474 192168 10480
rect 191444 10364 191752 10372
rect 191444 10362 191450 10364
rect 191506 10362 191530 10364
rect 191586 10362 191610 10364
rect 191666 10362 191690 10364
rect 191746 10362 191752 10364
rect 191506 10310 191508 10362
rect 191688 10310 191690 10362
rect 191444 10308 191450 10310
rect 191506 10308 191530 10310
rect 191586 10308 191610 10310
rect 191666 10308 191690 10310
rect 191746 10308 191752 10310
rect 191444 10298 191752 10308
rect 192496 10266 192524 12406
rect 192588 12374 192616 12786
rect 192668 12776 192720 12782
rect 192668 12718 192720 12724
rect 193036 12776 193088 12782
rect 193036 12718 193088 12724
rect 192576 12368 192628 12374
rect 192576 12310 192628 12316
rect 191288 10260 191340 10266
rect 191288 10202 191340 10208
rect 192484 10260 192536 10266
rect 192484 10202 192536 10208
rect 192588 10062 192616 12310
rect 192680 12306 192708 12718
rect 193048 12646 193076 12718
rect 193036 12640 193088 12646
rect 193036 12582 193088 12588
rect 193048 12344 193076 12582
rect 193034 12336 193090 12344
rect 192668 12300 192720 12306
rect 193034 12270 193090 12280
rect 192668 12242 192720 12248
rect 193036 12096 193088 12102
rect 193036 12038 193088 12044
rect 193048 11800 193076 12038
rect 193034 11792 193090 11800
rect 193034 11726 193090 11736
rect 193232 10742 193260 13738
rect 193496 13524 193548 13530
rect 193496 13466 193548 13472
rect 193404 13252 193456 13258
rect 193404 13194 193456 13200
rect 193416 12434 193444 13194
rect 193324 12406 193444 12434
rect 193324 11558 193352 12406
rect 193404 12164 193456 12170
rect 193404 12106 193456 12112
rect 193312 11552 193364 11558
rect 193312 11494 193364 11500
rect 193416 11370 193444 12106
rect 193508 12050 193536 13466
rect 193956 13252 194008 13258
rect 193956 13194 194008 13200
rect 194600 13252 194652 13258
rect 194600 13194 194652 13200
rect 194784 13252 194836 13258
rect 194784 13194 194836 13200
rect 193968 12986 193996 13194
rect 194612 13138 194640 13194
rect 194520 13110 194640 13138
rect 193956 12980 194008 12986
rect 193956 12922 194008 12928
rect 194416 12640 194468 12646
rect 194416 12582 194468 12588
rect 194048 12436 194100 12442
rect 194428 12434 194456 12582
rect 194100 12406 194456 12434
rect 194048 12378 194100 12384
rect 194416 12232 194468 12238
rect 194416 12174 194468 12180
rect 193680 12096 193732 12102
rect 193508 12044 193680 12050
rect 193508 12038 193732 12044
rect 193508 12022 193720 12038
rect 193508 11558 193536 12022
rect 194428 11898 194456 12174
rect 194416 11892 194468 11898
rect 194416 11834 194468 11840
rect 193864 11824 193916 11830
rect 193864 11766 193916 11772
rect 193496 11552 193548 11558
rect 193496 11494 193548 11500
rect 193416 11342 193536 11370
rect 193508 11218 193536 11342
rect 193496 11212 193548 11218
rect 193496 11154 193548 11160
rect 193312 11076 193364 11082
rect 193312 11018 193364 11024
rect 193220 10736 193272 10742
rect 193220 10678 193272 10684
rect 192576 10056 192628 10062
rect 192576 9998 192628 10004
rect 193324 9654 193352 11018
rect 193876 10810 193904 11766
rect 194324 11688 194376 11694
rect 194324 11630 194376 11636
rect 194416 11688 194468 11694
rect 194416 11630 194468 11636
rect 193864 10804 193916 10810
rect 193864 10746 193916 10752
rect 194140 10668 194192 10674
rect 194140 10610 194192 10616
rect 190644 9648 190696 9654
rect 190644 9590 190696 9596
rect 193312 9648 193364 9654
rect 193312 9590 193364 9596
rect 194152 9586 194180 10610
rect 194336 9926 194364 11630
rect 194428 11218 194456 11630
rect 194416 11212 194468 11218
rect 194416 11154 194468 11160
rect 194416 11008 194468 11014
rect 194416 10950 194468 10956
rect 194428 10062 194456 10950
rect 194416 10056 194468 10062
rect 194416 9998 194468 10004
rect 194324 9920 194376 9926
rect 194324 9862 194376 9868
rect 194140 9580 194192 9586
rect 194140 9522 194192 9528
rect 194520 9450 194548 13110
rect 194598 12880 194654 12888
rect 194598 12814 194654 12824
rect 194612 11218 194640 12814
rect 194796 12782 194824 13194
rect 194876 12980 194928 12986
rect 194876 12922 194928 12928
rect 194784 12776 194836 12782
rect 194784 12718 194836 12724
rect 194692 12164 194744 12170
rect 194692 12106 194744 12112
rect 194704 11898 194732 12106
rect 194692 11892 194744 11898
rect 194692 11834 194744 11840
rect 194600 11212 194652 11218
rect 194600 11154 194652 11160
rect 194888 11150 194916 12922
rect 195060 12844 195112 12850
rect 195060 12786 195112 12792
rect 195072 12752 195100 12786
rect 195058 12744 195114 12752
rect 195058 12678 195114 12688
rect 194968 12096 195020 12102
rect 194968 12038 195020 12044
rect 194876 11144 194928 11150
rect 194876 11086 194928 11092
rect 194980 10674 195008 12038
rect 195072 10742 195100 12678
rect 195256 11082 195284 15286
rect 197910 15286 198228 15314
rect 197910 15200 197966 15286
rect 195980 13796 196032 13802
rect 195980 13738 196032 13744
rect 195992 12986 196020 13738
rect 197636 13388 197688 13394
rect 197636 13330 197688 13336
rect 196440 13252 196492 13258
rect 196440 13194 196492 13200
rect 197360 13252 197412 13258
rect 197360 13194 197412 13200
rect 195980 12980 196032 12986
rect 195980 12922 196032 12928
rect 195794 12880 195850 12888
rect 195794 12814 195850 12824
rect 195808 12782 195836 12814
rect 195796 12776 195848 12782
rect 195796 12718 195848 12724
rect 195980 12640 196032 12646
rect 195980 12582 196032 12588
rect 195796 11552 195848 11558
rect 195796 11494 195848 11500
rect 195888 11552 195940 11558
rect 195888 11494 195940 11500
rect 195808 11150 195836 11494
rect 195796 11144 195848 11150
rect 195796 11086 195848 11092
rect 195244 11076 195296 11082
rect 195244 11018 195296 11024
rect 195060 10736 195112 10742
rect 195060 10678 195112 10684
rect 194968 10668 195020 10674
rect 194968 10610 195020 10616
rect 195900 10130 195928 11494
rect 195888 10124 195940 10130
rect 195888 10066 195940 10072
rect 195992 9518 196020 12582
rect 196452 11218 196480 13194
rect 197372 12888 197400 13194
rect 197358 12880 197414 12888
rect 197358 12814 197360 12824
rect 197412 12814 197414 12824
rect 197452 12844 197504 12850
rect 197360 12786 197412 12792
rect 197452 12786 197504 12792
rect 197464 12374 197492 12786
rect 197648 12782 197676 13330
rect 197728 13184 197780 13190
rect 197728 13126 197780 13132
rect 197912 13184 197964 13190
rect 197912 13126 197964 13132
rect 197740 12986 197768 13126
rect 197728 12980 197780 12986
rect 197728 12922 197780 12928
rect 197636 12776 197688 12782
rect 197636 12718 197688 12724
rect 197452 12368 197504 12374
rect 197452 12310 197504 12316
rect 197452 12232 197504 12238
rect 197452 12174 197504 12180
rect 196808 12096 196860 12102
rect 196808 12038 196860 12044
rect 196992 12096 197044 12102
rect 196992 12038 197044 12044
rect 197360 12096 197412 12102
rect 197360 12038 197412 12044
rect 196820 11830 196848 12038
rect 196808 11824 196860 11830
rect 196808 11766 196860 11772
rect 197004 11558 197032 12038
rect 197372 11694 197400 12038
rect 197360 11688 197412 11694
rect 197360 11630 197412 11636
rect 197464 11626 197492 12174
rect 197924 11762 197952 13126
rect 198200 12646 198228 15286
rect 201038 15286 201172 15314
rect 201038 15200 201094 15286
rect 200854 13288 200910 13296
rect 200854 13222 200910 13232
rect 200868 13190 200896 13222
rect 198556 13184 198608 13190
rect 198556 13126 198608 13132
rect 200488 13184 200540 13190
rect 200488 13126 200540 13132
rect 200856 13184 200908 13190
rect 200856 13126 200908 13132
rect 198372 12844 198424 12850
rect 198372 12786 198424 12792
rect 198188 12640 198240 12646
rect 198188 12582 198240 12588
rect 198384 12238 198412 12786
rect 198568 12782 198596 13126
rect 198556 12776 198608 12782
rect 198556 12718 198608 12724
rect 200396 12776 200448 12782
rect 200396 12718 200448 12724
rect 200408 12616 200436 12718
rect 200394 12608 200450 12616
rect 200394 12542 200450 12552
rect 200500 12306 200528 13126
rect 200672 12844 200724 12850
rect 200672 12786 200724 12792
rect 200684 12434 200712 12786
rect 201144 12646 201172 15286
rect 204074 15200 204130 16000
rect 207110 15314 207166 16000
rect 210238 15314 210294 16000
rect 213274 15314 213330 16000
rect 216310 15314 216366 16000
rect 207110 15286 207336 15314
rect 207110 15200 207166 15286
rect 201960 13456 202012 13462
rect 201960 13398 202012 13404
rect 203432 13456 203484 13462
rect 203432 13398 203484 13404
rect 201500 13320 201552 13326
rect 201500 13262 201552 13268
rect 201316 13184 201368 13190
rect 201316 13126 201368 13132
rect 201328 12850 201356 13126
rect 201316 12844 201368 12850
rect 201316 12786 201368 12792
rect 201132 12640 201184 12646
rect 201132 12582 201184 12588
rect 200592 12406 200712 12434
rect 200488 12300 200540 12306
rect 200488 12242 200540 12248
rect 200592 12238 200620 12406
rect 198372 12232 198424 12238
rect 198372 12174 198424 12180
rect 200580 12232 200632 12238
rect 200580 12174 200632 12180
rect 201040 12232 201092 12238
rect 201040 12174 201092 12180
rect 201052 11762 201080 12174
rect 197912 11756 197964 11762
rect 197912 11698 197964 11704
rect 201040 11756 201092 11762
rect 201040 11698 201092 11704
rect 197452 11620 197504 11626
rect 197452 11562 197504 11568
rect 196992 11552 197044 11558
rect 196992 11494 197044 11500
rect 201052 11218 201080 11698
rect 201328 11694 201356 12786
rect 201316 11688 201368 11694
rect 201316 11630 201368 11636
rect 201512 11558 201540 13262
rect 201972 12646 202000 13398
rect 202052 13388 202104 13394
rect 202052 13330 202104 13336
rect 201960 12640 202012 12646
rect 201960 12582 202012 12588
rect 202064 12306 202092 13330
rect 202144 13320 202196 13326
rect 203444 13296 203472 13398
rect 202144 13262 202196 13268
rect 203430 13288 203486 13296
rect 202156 12714 202184 13262
rect 202420 13252 202472 13258
rect 202420 13194 202472 13200
rect 203156 13252 203208 13258
rect 203430 13222 203486 13232
rect 203156 13194 203208 13200
rect 202144 12708 202196 12714
rect 202144 12650 202196 12656
rect 202432 12442 202460 13194
rect 202972 12912 203024 12918
rect 202972 12854 203024 12860
rect 202984 12782 203012 12854
rect 202880 12776 202932 12782
rect 202880 12718 202932 12724
rect 202972 12776 203024 12782
rect 202972 12718 203024 12724
rect 202420 12436 202472 12442
rect 202420 12378 202472 12384
rect 202052 12300 202104 12306
rect 202052 12242 202104 12248
rect 202892 11898 202920 12718
rect 203064 12096 203116 12102
rect 203064 12038 203116 12044
rect 202880 11892 202932 11898
rect 202880 11834 202932 11840
rect 203076 11762 203104 12038
rect 203168 11830 203196 13194
rect 203340 12912 203392 12918
rect 203340 12854 203392 12860
rect 203156 11824 203208 11830
rect 203156 11766 203208 11772
rect 203064 11756 203116 11762
rect 203064 11698 203116 11704
rect 202880 11688 202932 11694
rect 202880 11630 202932 11636
rect 201500 11552 201552 11558
rect 201500 11494 201552 11500
rect 196440 11212 196492 11218
rect 196440 11154 196492 11160
rect 201040 11212 201092 11218
rect 201040 11154 201092 11160
rect 201052 10606 201080 11154
rect 202696 11144 202748 11150
rect 202892 11098 202920 11630
rect 203352 11218 203380 12854
rect 203444 12102 203472 13222
rect 203524 12300 203576 12306
rect 203524 12242 203576 12248
rect 203432 12096 203484 12102
rect 203432 12038 203484 12044
rect 203444 11626 203472 12038
rect 203536 11694 203564 12242
rect 203524 11688 203576 11694
rect 203524 11630 203576 11636
rect 203432 11620 203484 11626
rect 203432 11562 203484 11568
rect 203340 11212 203392 11218
rect 203340 11154 203392 11160
rect 202748 11092 202920 11098
rect 202696 11086 202920 11092
rect 202708 11070 202920 11086
rect 201040 10600 201092 10606
rect 201040 10542 201092 10548
rect 203536 10470 203564 11630
rect 204088 11082 204116 15200
rect 207110 13560 207166 13568
rect 207110 13494 207112 13504
rect 207164 13494 207166 13504
rect 207112 13466 207164 13472
rect 206008 13456 206060 13462
rect 205652 13404 206008 13410
rect 205652 13398 206060 13404
rect 205652 13382 206048 13398
rect 205546 13288 205602 13296
rect 204260 13252 204312 13258
rect 204260 13194 204312 13200
rect 205456 13252 205508 13258
rect 205546 13222 205602 13232
rect 205456 13194 205508 13200
rect 204168 12776 204220 12782
rect 204168 12718 204220 12724
rect 204180 12434 204208 12718
rect 204272 12646 204300 13194
rect 205088 12776 205140 12782
rect 205088 12718 205140 12724
rect 205180 12776 205232 12782
rect 205180 12718 205232 12724
rect 204260 12640 204312 12646
rect 204260 12582 204312 12588
rect 204536 12640 204588 12646
rect 204536 12582 204588 12588
rect 204180 12406 204300 12434
rect 204272 12102 204300 12406
rect 204548 12238 204576 12582
rect 204536 12232 204588 12238
rect 204536 12174 204588 12180
rect 204260 12096 204312 12102
rect 204260 12038 204312 12044
rect 204548 11898 204576 12174
rect 204996 12164 205048 12170
rect 204996 12106 205048 12112
rect 204536 11892 204588 11898
rect 204536 11834 204588 11840
rect 204904 11620 204956 11626
rect 204904 11562 204956 11568
rect 204812 11552 204864 11558
rect 204812 11494 204864 11500
rect 204076 11076 204128 11082
rect 204076 11018 204128 11024
rect 204824 10674 204852 11494
rect 204916 11150 204944 11562
rect 205008 11218 205036 12106
rect 204996 11212 205048 11218
rect 204996 11154 205048 11160
rect 204904 11144 204956 11150
rect 204904 11086 204956 11092
rect 205100 10810 205128 12718
rect 205192 12646 205220 12718
rect 205180 12640 205232 12646
rect 205272 12640 205324 12646
rect 205180 12582 205232 12588
rect 205270 12608 205272 12616
rect 205324 12608 205326 12616
rect 205270 12542 205326 12552
rect 205468 11082 205496 13194
rect 205560 11830 205588 13222
rect 205652 13190 205680 13382
rect 207204 13320 207256 13326
rect 205730 13288 205786 13296
rect 207202 13288 207204 13296
rect 207256 13288 207258 13296
rect 205730 13222 205786 13232
rect 206376 13252 206428 13258
rect 205744 13190 205772 13222
rect 207202 13222 207258 13232
rect 206376 13194 206428 13200
rect 205640 13184 205692 13190
rect 205640 13126 205692 13132
rect 205732 13184 205784 13190
rect 205732 13126 205784 13132
rect 205640 12912 205692 12918
rect 205640 12854 205692 12860
rect 205652 12442 205680 12854
rect 205640 12436 205692 12442
rect 205640 12378 205692 12384
rect 205548 11824 205600 11830
rect 205548 11766 205600 11772
rect 206388 11762 206416 13194
rect 206560 12980 206612 12986
rect 206560 12922 206612 12928
rect 206572 11898 206600 12922
rect 207308 12714 207336 15286
rect 210238 15286 210372 15314
rect 210238 15200 210294 15286
rect 208030 13560 208086 13568
rect 210344 13530 210372 15286
rect 213274 15286 213408 15314
rect 213274 15200 213330 15286
rect 213380 13530 213408 15286
rect 216310 15286 216444 15314
rect 216310 15200 216366 15286
rect 208030 13494 208086 13504
rect 210332 13524 210384 13530
rect 208044 13462 208072 13494
rect 210332 13466 210384 13472
rect 213368 13524 213420 13530
rect 213368 13466 213420 13472
rect 216416 13462 216444 15286
rect 219438 15200 219494 16000
rect 222474 15314 222530 16000
rect 225602 15314 225658 16000
rect 228638 15314 228694 16000
rect 231674 15314 231730 16000
rect 234802 15314 234858 16000
rect 222474 15286 222792 15314
rect 222474 15200 222530 15286
rect 219452 13462 219480 15200
rect 207756 13456 207808 13462
rect 207756 13398 207808 13404
rect 208032 13456 208084 13462
rect 213276 13456 213328 13462
rect 208032 13398 208084 13404
rect 213274 13424 213276 13432
rect 216404 13456 216456 13462
rect 213328 13424 213330 13432
rect 207572 13252 207624 13258
rect 207624 13212 207704 13240
rect 207572 13194 207624 13200
rect 207388 13184 207440 13190
rect 207388 13126 207440 13132
rect 207400 12986 207428 13126
rect 207388 12980 207440 12986
rect 207388 12922 207440 12928
rect 207676 12850 207704 13212
rect 207664 12844 207716 12850
rect 207664 12786 207716 12792
rect 207296 12708 207348 12714
rect 207296 12650 207348 12656
rect 207676 12442 207704 12786
rect 207664 12436 207716 12442
rect 207768 12434 207796 13398
rect 216404 13398 216456 13404
rect 219440 13456 219492 13462
rect 219440 13398 219492 13404
rect 219806 13424 219862 13432
rect 213274 13358 213330 13368
rect 219806 13358 219862 13368
rect 207940 13320 207992 13326
rect 207938 13288 207940 13296
rect 213552 13320 213604 13326
rect 207992 13288 207994 13296
rect 213552 13262 213604 13268
rect 216588 13320 216640 13326
rect 216588 13262 216640 13268
rect 207938 13222 207994 13232
rect 213564 13190 213592 13262
rect 213552 13184 213604 13190
rect 213552 13126 213604 13132
rect 207848 12980 207900 12986
rect 207848 12922 207900 12928
rect 207860 12752 207888 12922
rect 210608 12912 210660 12918
rect 210608 12854 210660 12860
rect 207846 12744 207902 12752
rect 207846 12678 207902 12688
rect 210620 12646 210648 12854
rect 216600 12850 216628 13262
rect 219820 12986 219848 13358
rect 222764 13190 222792 15286
rect 225602 15286 225736 15314
rect 225602 15200 225658 15286
rect 224052 13518 224448 13546
rect 224052 13394 224080 13518
rect 224132 13456 224184 13462
rect 224132 13398 224184 13404
rect 224040 13388 224092 13394
rect 224040 13330 224092 13336
rect 224052 13190 224080 13330
rect 224144 13190 224172 13398
rect 224420 13394 224448 13518
rect 224408 13388 224460 13394
rect 224408 13330 224460 13336
rect 224236 13258 224448 13274
rect 224224 13252 224460 13258
rect 224276 13246 224408 13252
rect 224224 13194 224276 13200
rect 224408 13194 224460 13200
rect 225708 13190 225736 15286
rect 228638 15286 228864 15314
rect 228638 15200 228694 15286
rect 226444 13518 227208 13546
rect 226444 13462 226472 13518
rect 226432 13456 226484 13462
rect 226432 13398 226484 13404
rect 226616 13456 226668 13462
rect 226616 13398 226668 13404
rect 226892 13456 226944 13462
rect 226892 13398 226944 13404
rect 227074 13424 227130 13432
rect 222752 13184 222804 13190
rect 222752 13126 222804 13132
rect 223672 13184 223724 13190
rect 223672 13126 223724 13132
rect 224040 13184 224092 13190
rect 224040 13126 224092 13132
rect 224132 13184 224184 13190
rect 225420 13184 225472 13190
rect 224132 13126 224184 13132
rect 225418 13152 225420 13160
rect 225696 13184 225748 13190
rect 225472 13152 225474 13160
rect 219808 12980 219860 12986
rect 219808 12922 219860 12928
rect 223684 12850 223712 13126
rect 225696 13126 225748 13132
rect 225418 13086 225474 13096
rect 226628 12866 226656 13398
rect 226628 12850 226840 12866
rect 216588 12844 216640 12850
rect 216588 12786 216640 12792
rect 219808 12844 219860 12850
rect 219808 12786 219860 12792
rect 223672 12844 223724 12850
rect 226628 12844 226852 12850
rect 226628 12838 226800 12844
rect 223672 12786 223724 12792
rect 226800 12786 226852 12792
rect 219820 12714 219848 12786
rect 219808 12708 219860 12714
rect 219808 12650 219860 12656
rect 226904 12646 226932 13398
rect 227180 13394 227208 13518
rect 227904 13456 227956 13462
rect 227956 13404 228036 13410
rect 227904 13398 228036 13404
rect 227074 13358 227076 13368
rect 227128 13358 227130 13368
rect 227168 13388 227220 13394
rect 227076 13330 227128 13336
rect 227916 13382 228036 13398
rect 227168 13330 227220 13336
rect 227076 13184 227128 13190
rect 227074 13152 227076 13160
rect 227128 13152 227130 13160
rect 227180 13138 227208 13330
rect 227720 13320 227772 13326
rect 227720 13262 227772 13268
rect 228008 13274 228036 13382
rect 227628 13184 227680 13190
rect 227180 13110 227300 13138
rect 227628 13126 227680 13132
rect 227074 13086 227130 13096
rect 210608 12640 210660 12646
rect 210608 12582 210660 12588
rect 226892 12640 226944 12646
rect 226892 12582 226944 12588
rect 207768 12406 207888 12434
rect 207664 12378 207716 12384
rect 206560 11892 206612 11898
rect 206560 11834 206612 11840
rect 206376 11756 206428 11762
rect 206376 11698 206428 11704
rect 207860 11694 207888 12406
rect 227272 11694 227300 13110
rect 227640 12730 227668 13126
rect 227732 12866 227760 13262
rect 228008 13258 228128 13274
rect 228008 13252 228140 13258
rect 228008 13246 228088 13252
rect 228088 13194 228140 13200
rect 227904 13184 227956 13190
rect 227904 13126 227956 13132
rect 227732 12838 227852 12866
rect 227916 12850 227944 13126
rect 228272 12912 228324 12918
rect 228272 12854 228324 12860
rect 227640 12702 227760 12730
rect 227732 11830 227760 12702
rect 227824 11898 227852 12838
rect 227904 12844 227956 12850
rect 227904 12786 227956 12792
rect 228284 12782 228312 12854
rect 228272 12776 228324 12782
rect 228272 12718 228324 12724
rect 228836 12374 228864 15286
rect 231674 15286 231808 15314
rect 231674 15200 231730 15286
rect 231780 13682 231808 15286
rect 234802 15286 234936 15314
rect 234802 15200 234858 15286
rect 231780 13654 232084 13682
rect 229192 13456 229244 13462
rect 229190 13424 229192 13432
rect 229244 13424 229246 13432
rect 229190 13358 229246 13368
rect 231780 13394 231992 13410
rect 231780 13388 232004 13394
rect 231780 13382 231952 13388
rect 230388 13320 230440 13326
rect 230386 13288 230388 13296
rect 230440 13288 230442 13296
rect 230386 13222 230442 13232
rect 230756 13252 230808 13258
rect 230756 13194 230808 13200
rect 229544 13084 229852 13092
rect 229544 13082 229550 13084
rect 229606 13082 229630 13084
rect 229686 13082 229710 13084
rect 229766 13082 229790 13084
rect 229846 13082 229852 13084
rect 229606 13030 229608 13082
rect 229788 13030 229790 13082
rect 229544 13028 229550 13030
rect 229606 13028 229630 13030
rect 229686 13028 229710 13030
rect 229766 13028 229790 13030
rect 229846 13028 229852 13030
rect 229544 13018 229852 13028
rect 230388 12912 230440 12918
rect 230388 12854 230440 12860
rect 230296 12844 230348 12850
rect 230296 12786 230348 12792
rect 230204 12776 230256 12782
rect 230204 12718 230256 12724
rect 230216 12646 230244 12718
rect 229560 12640 229612 12646
rect 229560 12582 229612 12588
rect 230112 12640 230164 12646
rect 230112 12582 230164 12588
rect 230204 12640 230256 12646
rect 230204 12582 230256 12588
rect 228824 12368 228876 12374
rect 228824 12310 228876 12316
rect 228824 12096 228876 12102
rect 229572 12084 229600 12582
rect 230124 12442 230152 12582
rect 230112 12436 230164 12442
rect 230112 12378 230164 12384
rect 229928 12232 229980 12238
rect 229928 12174 229980 12180
rect 228824 12038 228876 12044
rect 229480 12056 229600 12084
rect 228836 11898 228864 12038
rect 227812 11892 227864 11898
rect 227812 11834 227864 11840
rect 228824 11892 228876 11898
rect 228824 11834 228876 11840
rect 227720 11824 227772 11830
rect 229480 11778 229508 12056
rect 229544 11996 229852 12004
rect 229544 11994 229550 11996
rect 229606 11994 229630 11996
rect 229686 11994 229710 11996
rect 229766 11994 229790 11996
rect 229846 11994 229852 11996
rect 229606 11942 229608 11994
rect 229788 11942 229790 11994
rect 229544 11940 229550 11942
rect 229606 11940 229630 11942
rect 229686 11940 229710 11942
rect 229766 11940 229790 11942
rect 229846 11940 229852 11942
rect 229544 11930 229852 11940
rect 229940 11898 229968 12174
rect 229928 11892 229980 11898
rect 229928 11834 229980 11840
rect 227720 11766 227772 11772
rect 229388 11762 229508 11778
rect 229376 11756 229508 11762
rect 229428 11750 229508 11756
rect 229376 11698 229428 11704
rect 207848 11688 207900 11694
rect 207848 11630 207900 11636
rect 227260 11688 227312 11694
rect 227260 11630 227312 11636
rect 230308 11626 230336 12786
rect 230400 11898 230428 12854
rect 230388 11892 230440 11898
rect 230388 11834 230440 11840
rect 230296 11620 230348 11626
rect 230296 11562 230348 11568
rect 229376 11552 229428 11558
rect 229376 11494 229428 11500
rect 229388 11150 229416 11494
rect 229376 11144 229428 11150
rect 229376 11086 229428 11092
rect 230768 11082 230796 13194
rect 231032 12912 231084 12918
rect 231032 12854 231084 12860
rect 230848 12164 230900 12170
rect 230848 12106 230900 12112
rect 230860 11830 230888 12106
rect 231044 11898 231072 12854
rect 231124 12368 231176 12374
rect 231124 12310 231176 12316
rect 231136 12170 231164 12310
rect 231676 12300 231728 12306
rect 231676 12242 231728 12248
rect 231308 12232 231360 12238
rect 231308 12174 231360 12180
rect 231124 12164 231176 12170
rect 231124 12106 231176 12112
rect 231216 12096 231268 12102
rect 231320 12084 231348 12174
rect 231400 12096 231452 12102
rect 231320 12056 231400 12084
rect 231216 12038 231268 12044
rect 231400 12038 231452 12044
rect 231032 11892 231084 11898
rect 231032 11834 231084 11840
rect 230848 11824 230900 11830
rect 230848 11766 230900 11772
rect 231228 11762 231256 12038
rect 231688 11898 231716 12242
rect 231780 12102 231808 13382
rect 231952 13330 232004 13336
rect 232056 13326 232084 13654
rect 233148 13388 233200 13394
rect 233148 13330 233200 13336
rect 233332 13388 233384 13394
rect 233332 13330 233384 13336
rect 231860 13320 231912 13326
rect 231860 13262 231912 13268
rect 232044 13320 232096 13326
rect 233056 13320 233108 13326
rect 232044 13262 232096 13268
rect 232134 13288 232190 13296
rect 231872 12442 231900 13262
rect 233056 13262 233108 13268
rect 232134 13222 232190 13232
rect 232148 13190 232176 13222
rect 232136 13184 232188 13190
rect 232136 13126 232188 13132
rect 232320 12912 232372 12918
rect 232320 12854 232372 12860
rect 232332 12646 232360 12854
rect 233068 12850 233096 13262
rect 233160 13172 233188 13330
rect 233240 13184 233292 13190
rect 233160 13144 233240 13172
rect 233240 13126 233292 13132
rect 233344 13002 233372 13330
rect 234908 13190 234936 15286
rect 237838 15200 237894 16000
rect 240874 15314 240930 16000
rect 244002 15314 244058 16000
rect 247038 15314 247094 16000
rect 250074 15314 250130 16000
rect 240874 15286 241284 15314
rect 240874 15200 240930 15286
rect 234896 13184 234948 13190
rect 234896 13126 234948 13132
rect 237012 13184 237064 13190
rect 237012 13126 237064 13132
rect 233160 12974 233372 13002
rect 233056 12844 233108 12850
rect 233056 12786 233108 12792
rect 232320 12640 232372 12646
rect 232320 12582 232372 12588
rect 232504 12640 232556 12646
rect 232504 12582 232556 12588
rect 231860 12436 231912 12442
rect 231860 12378 231912 12384
rect 232516 12374 232544 12582
rect 232504 12368 232556 12374
rect 232504 12310 232556 12316
rect 233068 12238 233096 12786
rect 233160 12646 233188 12974
rect 237024 12850 237052 13126
rect 237012 12844 237064 12850
rect 237012 12786 237064 12792
rect 237852 12714 237880 15200
rect 239496 13456 239548 13462
rect 238114 13424 238170 13432
rect 237932 13388 237984 13394
rect 238114 13358 238116 13368
rect 237932 13330 237984 13336
rect 238168 13358 238170 13368
rect 239494 13424 239496 13432
rect 239548 13424 239550 13432
rect 239494 13358 239550 13368
rect 238116 13330 238168 13336
rect 237944 12714 237972 13330
rect 238208 13320 238260 13326
rect 238208 13262 238260 13268
rect 238220 12986 238248 13262
rect 238484 13252 238536 13258
rect 238484 13194 238536 13200
rect 238208 12980 238260 12986
rect 238208 12922 238260 12928
rect 238300 12912 238352 12918
rect 238300 12854 238352 12860
rect 238312 12752 238340 12854
rect 238392 12844 238444 12850
rect 238392 12786 238444 12792
rect 238298 12744 238354 12752
rect 237840 12708 237892 12714
rect 237840 12650 237892 12656
rect 237932 12708 237984 12714
rect 238298 12678 238354 12688
rect 237932 12650 237984 12656
rect 233148 12640 233200 12646
rect 233148 12582 233200 12588
rect 238404 12238 238432 12786
rect 238496 12646 238524 13194
rect 239036 12912 239088 12918
rect 239036 12854 239088 12860
rect 238484 12640 238536 12646
rect 238484 12582 238536 12588
rect 238852 12640 238904 12646
rect 238852 12582 238904 12588
rect 238864 12306 238892 12582
rect 239048 12442 239076 12854
rect 239128 12640 239180 12646
rect 239128 12582 239180 12588
rect 239036 12436 239088 12442
rect 239036 12378 239088 12384
rect 238852 12300 238904 12306
rect 238852 12242 238904 12248
rect 239140 12238 239168 12582
rect 239312 12300 239364 12306
rect 239312 12242 239364 12248
rect 232136 12232 232188 12238
rect 232136 12174 232188 12180
rect 233056 12232 233108 12238
rect 233056 12174 233108 12180
rect 238024 12232 238076 12238
rect 238024 12174 238076 12180
rect 238392 12232 238444 12238
rect 238392 12174 238444 12180
rect 239128 12232 239180 12238
rect 239128 12174 239180 12180
rect 231768 12096 231820 12102
rect 231768 12038 231820 12044
rect 231676 11892 231728 11898
rect 231676 11834 231728 11840
rect 231216 11756 231268 11762
rect 231216 11698 231268 11704
rect 231688 11558 231716 11834
rect 232148 11626 232176 12174
rect 233068 12102 233096 12174
rect 233056 12096 233108 12102
rect 233056 12038 233108 12044
rect 232136 11620 232188 11626
rect 232136 11562 232188 11568
rect 231676 11552 231728 11558
rect 231676 11494 231728 11500
rect 238036 11218 238064 12174
rect 239324 11694 239352 12242
rect 239508 12238 239536 13358
rect 239772 13320 239824 13326
rect 239772 13262 239824 13268
rect 239496 12232 239548 12238
rect 239496 12174 239548 12180
rect 239312 11688 239364 11694
rect 239312 11630 239364 11636
rect 239404 11552 239456 11558
rect 239404 11494 239456 11500
rect 239416 11354 239444 11494
rect 239784 11354 239812 13262
rect 241060 13252 241112 13258
rect 241060 13194 241112 13200
rect 240048 12912 240100 12918
rect 240048 12854 240100 12860
rect 240968 12912 241020 12918
rect 240968 12854 241020 12860
rect 239956 12300 240008 12306
rect 239956 12242 240008 12248
rect 239968 11694 239996 12242
rect 239956 11688 240008 11694
rect 239956 11630 240008 11636
rect 240060 11354 240088 12854
rect 240324 12640 240376 12646
rect 240324 12582 240376 12588
rect 240140 12436 240192 12442
rect 240140 12378 240192 12384
rect 240152 11830 240180 12378
rect 240336 11898 240364 12582
rect 240876 12096 240928 12102
rect 240876 12038 240928 12044
rect 240324 11892 240376 11898
rect 240324 11834 240376 11840
rect 240140 11824 240192 11830
rect 240140 11766 240192 11772
rect 239404 11348 239456 11354
rect 239404 11290 239456 11296
rect 239772 11348 239824 11354
rect 239772 11290 239824 11296
rect 240048 11348 240100 11354
rect 240048 11290 240100 11296
rect 238024 11212 238076 11218
rect 238024 11154 238076 11160
rect 240888 11150 240916 12038
rect 240980 11354 241008 12854
rect 241072 11898 241100 13194
rect 241060 11892 241112 11898
rect 241060 11834 241112 11840
rect 241256 11558 241284 15286
rect 244002 15286 244228 15314
rect 244002 15200 244058 15286
rect 244096 13388 244148 13394
rect 244096 13330 244148 13336
rect 241796 13252 241848 13258
rect 241796 13194 241848 13200
rect 243636 13252 243688 13258
rect 243636 13194 243688 13200
rect 241520 12096 241572 12102
rect 241520 12038 241572 12044
rect 241532 11830 241560 12038
rect 241808 11898 241836 13194
rect 242532 13184 242584 13190
rect 242532 13126 242584 13132
rect 242072 12844 242124 12850
rect 242072 12786 242124 12792
rect 242256 12844 242308 12850
rect 242256 12786 242308 12792
rect 241796 11892 241848 11898
rect 241796 11834 241848 11840
rect 241520 11824 241572 11830
rect 241520 11766 241572 11772
rect 241980 11688 242032 11694
rect 241980 11630 242032 11636
rect 241244 11552 241296 11558
rect 241244 11494 241296 11500
rect 240968 11348 241020 11354
rect 240968 11290 241020 11296
rect 241992 11150 242020 11630
rect 242084 11354 242112 12786
rect 242162 12744 242218 12752
rect 242162 12678 242164 12688
rect 242216 12678 242218 12688
rect 242164 12650 242216 12656
rect 242268 12374 242296 12786
rect 242440 12640 242492 12646
rect 242440 12582 242492 12588
rect 242256 12368 242308 12374
rect 242256 12310 242308 12316
rect 242452 12306 242480 12582
rect 242440 12300 242492 12306
rect 242440 12242 242492 12248
rect 242164 12232 242216 12238
rect 242452 12186 242480 12242
rect 242216 12180 242480 12186
rect 242164 12174 242480 12180
rect 242176 12158 242480 12174
rect 242544 12102 242572 13126
rect 242900 12640 242952 12646
rect 242900 12582 242952 12588
rect 242912 12306 242940 12582
rect 243648 12442 243676 13194
rect 243636 12436 243688 12442
rect 243636 12378 243688 12384
rect 242992 12368 243044 12374
rect 243044 12316 243216 12322
rect 242992 12310 243216 12316
rect 243004 12306 243216 12310
rect 242900 12300 242952 12306
rect 243004 12300 243228 12306
rect 243004 12294 243176 12300
rect 242900 12242 242952 12248
rect 243176 12242 243228 12248
rect 244108 12102 244136 13330
rect 244200 12442 244228 15286
rect 247038 15286 247172 15314
rect 247038 15200 247094 15286
rect 247144 13462 247172 15286
rect 250074 15286 250208 15314
rect 250074 15200 250130 15286
rect 244648 13456 244700 13462
rect 244648 13398 244700 13404
rect 245384 13456 245436 13462
rect 245384 13398 245436 13404
rect 247132 13456 247184 13462
rect 247132 13398 247184 13404
rect 244660 13002 244688 13398
rect 244924 13252 244976 13258
rect 244924 13194 244976 13200
rect 244568 12974 244688 13002
rect 244568 12850 244596 12974
rect 244936 12918 244964 13194
rect 245396 12918 245424 13398
rect 244648 12912 244700 12918
rect 244648 12854 244700 12860
rect 244924 12912 244976 12918
rect 244924 12854 244976 12860
rect 245384 12912 245436 12918
rect 245384 12854 245436 12860
rect 244556 12844 244608 12850
rect 244556 12786 244608 12792
rect 244188 12436 244240 12442
rect 244188 12378 244240 12384
rect 242532 12096 242584 12102
rect 242532 12038 242584 12044
rect 244096 12096 244148 12102
rect 244096 12038 244148 12044
rect 242544 11762 242572 12038
rect 242532 11756 242584 11762
rect 242532 11698 242584 11704
rect 244568 11694 244596 12786
rect 244660 12714 244688 12854
rect 244832 12844 244884 12850
rect 244832 12786 244884 12792
rect 244648 12708 244700 12714
rect 244648 12650 244700 12656
rect 244844 11830 244872 12786
rect 250180 12714 250208 15286
rect 253202 15200 253258 16000
rect 256238 15200 256294 16000
rect 259366 15200 259422 16000
rect 262402 15314 262458 16000
rect 262402 15286 262536 15314
rect 262402 15200 262458 15286
rect 251008 13518 251496 13546
rect 251008 13394 251036 13518
rect 251088 13456 251140 13462
rect 251140 13404 251312 13410
rect 251088 13398 251312 13404
rect 250996 13388 251048 13394
rect 251100 13382 251312 13398
rect 250996 13330 251048 13336
rect 251088 13320 251140 13326
rect 251088 13262 251140 13268
rect 251100 12986 251128 13262
rect 251180 13184 251232 13190
rect 251180 13126 251232 13132
rect 251088 12980 251140 12986
rect 251088 12922 251140 12928
rect 251192 12850 251220 13126
rect 251180 12844 251232 12850
rect 251180 12786 251232 12792
rect 248328 12708 248380 12714
rect 248328 12650 248380 12656
rect 250168 12708 250220 12714
rect 250168 12650 250220 12656
rect 248340 12306 248368 12650
rect 248328 12300 248380 12306
rect 248328 12242 248380 12248
rect 249248 12300 249300 12306
rect 249248 12242 249300 12248
rect 249260 12170 249288 12242
rect 251284 12238 251312 13382
rect 251364 13252 251416 13258
rect 251364 13194 251416 13200
rect 251376 12442 251404 13194
rect 251364 12436 251416 12442
rect 251364 12378 251416 12384
rect 251468 12374 251496 13518
rect 252468 13456 252520 13462
rect 252468 13398 252520 13404
rect 252376 13252 252428 13258
rect 252376 13194 252428 13200
rect 251640 12912 251692 12918
rect 251640 12854 251692 12860
rect 251548 12844 251600 12850
rect 251548 12786 251600 12792
rect 251456 12368 251508 12374
rect 251456 12310 251508 12316
rect 251272 12232 251324 12238
rect 251272 12174 251324 12180
rect 249064 12164 249116 12170
rect 249064 12106 249116 12112
rect 249248 12164 249300 12170
rect 249248 12106 249300 12112
rect 244832 11824 244884 11830
rect 244832 11766 244884 11772
rect 242716 11688 242768 11694
rect 242716 11630 242768 11636
rect 244556 11688 244608 11694
rect 244556 11630 244608 11636
rect 242072 11348 242124 11354
rect 242072 11290 242124 11296
rect 242728 11218 242756 11630
rect 249076 11558 249104 12106
rect 249064 11552 249116 11558
rect 249064 11494 249116 11500
rect 242716 11212 242768 11218
rect 242716 11154 242768 11160
rect 240876 11144 240928 11150
rect 240876 11086 240928 11092
rect 241980 11144 242032 11150
rect 241980 11086 242032 11092
rect 205456 11076 205508 11082
rect 205456 11018 205508 11024
rect 230756 11076 230808 11082
rect 230756 11018 230808 11024
rect 229544 10908 229852 10916
rect 229544 10906 229550 10908
rect 229606 10906 229630 10908
rect 229686 10906 229710 10908
rect 229766 10906 229790 10908
rect 229846 10906 229852 10908
rect 229606 10854 229608 10906
rect 229788 10854 229790 10906
rect 229544 10852 229550 10854
rect 229606 10852 229630 10854
rect 229686 10852 229710 10854
rect 229766 10852 229790 10854
rect 229846 10852 229852 10854
rect 229544 10842 229852 10852
rect 205088 10804 205140 10810
rect 205088 10746 205140 10752
rect 204812 10668 204864 10674
rect 204812 10610 204864 10616
rect 203524 10464 203576 10470
rect 203524 10406 203576 10412
rect 229544 9820 229852 9828
rect 229544 9818 229550 9820
rect 229606 9818 229630 9820
rect 229686 9818 229710 9820
rect 229766 9818 229790 9820
rect 229846 9818 229852 9820
rect 229606 9766 229608 9818
rect 229788 9766 229790 9818
rect 229544 9764 229550 9766
rect 229606 9764 229630 9766
rect 229686 9764 229710 9766
rect 229766 9764 229790 9766
rect 229846 9764 229852 9766
rect 229544 9754 229852 9764
rect 195980 9512 196032 9518
rect 195980 9454 196032 9460
rect 194508 9444 194560 9450
rect 194508 9386 194560 9392
rect 191444 9276 191752 9284
rect 191444 9274 191450 9276
rect 191506 9274 191530 9276
rect 191586 9274 191610 9276
rect 191666 9274 191690 9276
rect 191746 9274 191752 9276
rect 191506 9222 191508 9274
rect 191688 9222 191690 9274
rect 191444 9220 191450 9222
rect 191506 9220 191530 9222
rect 191586 9220 191610 9222
rect 191666 9220 191690 9222
rect 191746 9220 191752 9222
rect 191444 9210 191752 9220
rect 229544 8732 229852 8740
rect 229544 8730 229550 8732
rect 229606 8730 229630 8732
rect 229686 8730 229710 8732
rect 229766 8730 229790 8732
rect 229846 8730 229852 8732
rect 229606 8678 229608 8730
rect 229788 8678 229790 8730
rect 229544 8676 229550 8678
rect 229606 8676 229630 8678
rect 229686 8676 229710 8678
rect 229766 8676 229790 8678
rect 229846 8676 229852 8678
rect 229544 8666 229852 8676
rect 187516 8356 187568 8362
rect 187516 8298 187568 8304
rect 191444 8188 191752 8196
rect 191444 8186 191450 8188
rect 191506 8186 191530 8188
rect 191586 8186 191610 8188
rect 191666 8186 191690 8188
rect 191746 8186 191752 8188
rect 191506 8134 191508 8186
rect 191688 8134 191690 8186
rect 191444 8132 191450 8134
rect 191506 8132 191530 8134
rect 191586 8132 191610 8134
rect 191666 8132 191690 8134
rect 191746 8132 191752 8134
rect 191444 8122 191752 8132
rect 153346 7644 153654 7652
rect 153346 7642 153352 7644
rect 153408 7642 153432 7644
rect 153488 7642 153512 7644
rect 153568 7642 153592 7644
rect 153648 7642 153654 7644
rect 153408 7590 153410 7642
rect 153590 7590 153592 7642
rect 153346 7588 153352 7590
rect 153408 7588 153432 7590
rect 153488 7588 153512 7590
rect 153568 7588 153592 7590
rect 153648 7588 153654 7590
rect 153346 7578 153654 7588
rect 229544 7644 229852 7652
rect 229544 7642 229550 7644
rect 229606 7642 229630 7644
rect 229686 7642 229710 7644
rect 229766 7642 229790 7644
rect 229846 7642 229852 7644
rect 229606 7590 229608 7642
rect 229788 7590 229790 7642
rect 229544 7588 229550 7590
rect 229606 7588 229630 7590
rect 229686 7588 229710 7590
rect 229766 7588 229790 7590
rect 229846 7588 229852 7590
rect 229544 7578 229852 7588
rect 191444 7100 191752 7108
rect 191444 7098 191450 7100
rect 191506 7098 191530 7100
rect 191586 7098 191610 7100
rect 191666 7098 191690 7100
rect 191746 7098 191752 7100
rect 191506 7046 191508 7098
rect 191688 7046 191690 7098
rect 191444 7044 191450 7046
rect 191506 7044 191530 7046
rect 191586 7044 191610 7046
rect 191666 7044 191690 7046
rect 191746 7044 191752 7046
rect 191444 7034 191752 7044
rect 153346 6556 153654 6564
rect 153346 6554 153352 6556
rect 153408 6554 153432 6556
rect 153488 6554 153512 6556
rect 153568 6554 153592 6556
rect 153648 6554 153654 6556
rect 153408 6502 153410 6554
rect 153590 6502 153592 6554
rect 153346 6500 153352 6502
rect 153408 6500 153432 6502
rect 153488 6500 153512 6502
rect 153568 6500 153592 6502
rect 153648 6500 153654 6502
rect 153346 6490 153654 6500
rect 229544 6556 229852 6564
rect 229544 6554 229550 6556
rect 229606 6554 229630 6556
rect 229686 6554 229710 6556
rect 229766 6554 229790 6556
rect 229846 6554 229852 6556
rect 229606 6502 229608 6554
rect 229788 6502 229790 6554
rect 229544 6500 229550 6502
rect 229606 6500 229630 6502
rect 229686 6500 229710 6502
rect 229766 6500 229790 6502
rect 229846 6500 229852 6502
rect 229544 6490 229852 6500
rect 249076 6254 249104 11494
rect 251560 11150 251588 12786
rect 251652 11626 251680 12854
rect 252100 12776 252152 12782
rect 252100 12718 252152 12724
rect 251824 12708 251876 12714
rect 251824 12650 251876 12656
rect 251836 12480 251864 12650
rect 251916 12640 251968 12646
rect 251914 12608 251916 12616
rect 252008 12640 252060 12646
rect 251968 12608 251970 12616
rect 252008 12582 252060 12588
rect 251914 12542 251970 12552
rect 251822 12472 251878 12480
rect 251822 12406 251878 12416
rect 251916 12436 251968 12442
rect 251916 12378 251968 12384
rect 251928 12238 251956 12378
rect 251916 12232 251968 12238
rect 251916 12174 251968 12180
rect 252020 11762 252048 12582
rect 252112 12374 252140 12718
rect 252388 12434 252416 13194
rect 252480 12918 252508 13398
rect 253020 13252 253072 13258
rect 253020 13194 253072 13200
rect 252468 12912 252520 12918
rect 252468 12854 252520 12860
rect 253032 12434 253060 13194
rect 252388 12406 252508 12434
rect 252100 12368 252152 12374
rect 252100 12310 252152 12316
rect 252008 11756 252060 11762
rect 252008 11698 252060 11704
rect 252112 11694 252140 12310
rect 252100 11688 252152 11694
rect 252100 11630 252152 11636
rect 251640 11620 251692 11626
rect 251640 11562 251692 11568
rect 252480 11354 252508 12406
rect 252940 12406 253060 12434
rect 252940 11898 252968 12406
rect 253112 12164 253164 12170
rect 253112 12106 253164 12112
rect 252928 11892 252980 11898
rect 252928 11834 252980 11840
rect 252744 11756 252796 11762
rect 252744 11698 252796 11704
rect 253020 11756 253072 11762
rect 253020 11698 253072 11704
rect 252468 11348 252520 11354
rect 252468 11290 252520 11296
rect 252756 11286 252784 11698
rect 252744 11280 252796 11286
rect 252744 11222 252796 11228
rect 251548 11144 251600 11150
rect 251548 11086 251600 11092
rect 252756 9994 252784 11222
rect 253032 11150 253060 11698
rect 253124 11354 253152 12106
rect 253112 11348 253164 11354
rect 253112 11290 253164 11296
rect 253216 11286 253244 15200
rect 254952 13456 255004 13462
rect 254688 13416 254952 13444
rect 253480 13184 253532 13190
rect 253480 13126 253532 13132
rect 253492 12764 253520 13126
rect 254688 12986 254716 13416
rect 254952 13398 255004 13404
rect 256252 13410 256280 15200
rect 259380 13682 259408 15200
rect 259380 13654 259500 13682
rect 259472 13462 259500 13654
rect 259460 13456 259512 13462
rect 256252 13382 256556 13410
rect 259460 13398 259512 13404
rect 256240 13320 256292 13326
rect 256240 13262 256292 13268
rect 254952 13252 255004 13258
rect 254952 13194 255004 13200
rect 255320 13252 255372 13258
rect 255320 13194 255372 13200
rect 254676 12980 254728 12986
rect 254676 12922 254728 12928
rect 253664 12776 253716 12782
rect 253492 12736 253664 12764
rect 253664 12718 253716 12724
rect 253940 12776 253992 12782
rect 253940 12718 253992 12724
rect 253952 12322 253980 12718
rect 254308 12368 254360 12374
rect 253952 12294 254072 12322
rect 254308 12310 254360 12316
rect 253296 11552 253348 11558
rect 253296 11494 253348 11500
rect 253204 11280 253256 11286
rect 253204 11222 253256 11228
rect 253308 11150 253336 11494
rect 254044 11354 254072 12294
rect 254320 11830 254348 12310
rect 254400 12096 254452 12102
rect 254400 12038 254452 12044
rect 254308 11824 254360 11830
rect 254308 11766 254360 11772
rect 254032 11348 254084 11354
rect 254032 11290 254084 11296
rect 254412 11150 254440 12038
rect 254688 11898 254716 12922
rect 254964 12434 254992 13194
rect 255332 13138 255360 13194
rect 255240 13110 255360 13138
rect 255136 12776 255188 12782
rect 255136 12718 255188 12724
rect 255044 12708 255096 12714
rect 255044 12650 255096 12656
rect 254780 12406 254992 12434
rect 254780 11898 254808 12406
rect 255056 12186 255084 12650
rect 255148 12238 255176 12718
rect 255240 12434 255268 13110
rect 256252 12986 256280 13262
rect 256332 13184 256384 13190
rect 256332 13126 256384 13132
rect 256240 12980 256292 12986
rect 256240 12922 256292 12928
rect 256344 12782 256372 13126
rect 256332 12776 256384 12782
rect 256332 12718 256384 12724
rect 256424 12776 256476 12782
rect 256424 12718 256476 12724
rect 255240 12406 255360 12434
rect 255228 12368 255280 12374
rect 255228 12310 255280 12316
rect 254964 12158 255084 12186
rect 255136 12232 255188 12238
rect 255136 12174 255188 12180
rect 254676 11892 254728 11898
rect 254676 11834 254728 11840
rect 254768 11892 254820 11898
rect 254768 11834 254820 11840
rect 254688 11150 254716 11834
rect 253020 11144 253072 11150
rect 253020 11086 253072 11092
rect 253296 11144 253348 11150
rect 253296 11086 253348 11092
rect 254400 11144 254452 11150
rect 254400 11086 254452 11092
rect 254676 11144 254728 11150
rect 254676 11086 254728 11092
rect 254964 10674 254992 12158
rect 255240 12102 255268 12310
rect 255044 12096 255096 12102
rect 255044 12038 255096 12044
rect 255228 12096 255280 12102
rect 255228 12038 255280 12044
rect 255056 11898 255084 12038
rect 255044 11892 255096 11898
rect 255044 11834 255096 11840
rect 255332 11676 255360 12406
rect 255596 12300 255648 12306
rect 255596 12242 255648 12248
rect 255608 11694 255636 12242
rect 256240 12232 256292 12238
rect 256240 12174 256292 12180
rect 256332 12232 256384 12238
rect 256332 12174 256384 12180
rect 256252 11762 256280 12174
rect 256344 12102 256372 12174
rect 256332 12096 256384 12102
rect 256332 12038 256384 12044
rect 256240 11756 256292 11762
rect 256240 11698 256292 11704
rect 256436 11694 256464 12718
rect 256528 12442 256556 13382
rect 256976 13252 257028 13258
rect 256976 13194 257028 13200
rect 261852 13252 261904 13258
rect 261852 13194 261904 13200
rect 256606 13016 256662 13024
rect 256606 12950 256662 12960
rect 256620 12850 256648 12950
rect 256608 12844 256660 12850
rect 256608 12786 256660 12792
rect 256516 12436 256568 12442
rect 256516 12378 256568 12384
rect 256988 12374 257016 13194
rect 257988 13184 258040 13190
rect 257988 13126 258040 13132
rect 258000 13024 258028 13126
rect 257986 13016 258042 13024
rect 257986 12950 258042 12960
rect 257252 12912 257304 12918
rect 257252 12854 257304 12860
rect 261760 12912 261812 12918
rect 261760 12854 261812 12860
rect 257160 12776 257212 12782
rect 257160 12718 257212 12724
rect 257068 12708 257120 12714
rect 257068 12650 257120 12656
rect 257080 12616 257108 12650
rect 257066 12608 257122 12616
rect 257066 12542 257122 12552
rect 257172 12480 257200 12718
rect 257158 12472 257214 12480
rect 257158 12406 257214 12416
rect 256976 12368 257028 12374
rect 256976 12310 257028 12316
rect 257264 11762 257292 12854
rect 257252 11756 257304 11762
rect 257252 11698 257304 11704
rect 255240 11648 255360 11676
rect 255596 11688 255648 11694
rect 255240 10810 255268 11648
rect 255596 11630 255648 11636
rect 256424 11688 256476 11694
rect 256424 11630 256476 11636
rect 261772 11558 261800 12854
rect 261864 12850 261892 13194
rect 261852 12844 261904 12850
rect 261852 12786 261904 12792
rect 261864 12306 261892 12786
rect 262312 12776 262364 12782
rect 262310 12744 262312 12752
rect 262364 12744 262366 12752
rect 262310 12678 262366 12688
rect 262220 12640 262272 12646
rect 262272 12600 262444 12628
rect 262220 12582 262272 12588
rect 262416 12306 262444 12600
rect 262508 12442 262536 15286
rect 265438 15200 265494 16000
rect 268566 15200 268622 16000
rect 271602 15314 271658 16000
rect 274638 15314 274694 16000
rect 277766 15314 277822 16000
rect 280802 15314 280858 16000
rect 283930 15314 283986 16000
rect 271602 15286 271828 15314
rect 271602 15200 271658 15286
rect 263508 13456 263560 13462
rect 263508 13398 263560 13404
rect 263414 13288 263470 13296
rect 263520 13258 263548 13398
rect 264152 13388 264204 13394
rect 264152 13330 264204 13336
rect 263414 13222 263416 13232
rect 263468 13222 263470 13232
rect 263508 13252 263560 13258
rect 263416 13194 263468 13200
rect 263508 13194 263560 13200
rect 262956 13184 263008 13190
rect 263324 13184 263376 13190
rect 263008 13144 263088 13172
rect 262956 13126 263008 13132
rect 262680 12708 262732 12714
rect 262680 12650 262732 12656
rect 262496 12436 262548 12442
rect 262496 12378 262548 12384
rect 261852 12300 261904 12306
rect 261852 12242 261904 12248
rect 262404 12300 262456 12306
rect 262404 12242 262456 12248
rect 262692 11558 262720 12650
rect 263060 12238 263088 13144
rect 263324 13126 263376 13132
rect 263336 12918 263364 13126
rect 263324 12912 263376 12918
rect 263324 12854 263376 12860
rect 263506 12744 263562 12752
rect 263506 12678 263508 12688
rect 263560 12678 263562 12688
rect 263508 12650 263560 12656
rect 263968 12640 264020 12646
rect 263968 12582 264020 12588
rect 263048 12232 263100 12238
rect 263048 12174 263100 12180
rect 263980 11694 264008 12582
rect 264164 12306 264192 13330
rect 264428 13252 264480 13258
rect 264428 13194 264480 13200
rect 264612 13252 264664 13258
rect 264612 13194 264664 13200
rect 264980 13252 265032 13258
rect 264980 13194 265032 13200
rect 264440 12850 264468 13194
rect 264624 12986 264652 13194
rect 264612 12980 264664 12986
rect 264612 12922 264664 12928
rect 264336 12844 264388 12850
rect 264336 12786 264388 12792
rect 264428 12844 264480 12850
rect 264428 12786 264480 12792
rect 264348 12752 264376 12786
rect 264334 12744 264390 12752
rect 264334 12678 264390 12688
rect 264992 12374 265020 13194
rect 264980 12368 265032 12374
rect 264980 12310 265032 12316
rect 264152 12300 264204 12306
rect 264152 12242 264204 12248
rect 265164 12300 265216 12306
rect 265164 12242 265216 12248
rect 264336 12232 264388 12238
rect 264336 12174 264388 12180
rect 264348 11762 264376 12174
rect 265176 12170 265204 12242
rect 265164 12164 265216 12170
rect 265164 12106 265216 12112
rect 265176 11914 265204 12106
rect 265176 11886 265296 11914
rect 265268 11762 265296 11886
rect 264336 11756 264388 11762
rect 264336 11698 264388 11704
rect 265164 11756 265216 11762
rect 265164 11698 265216 11704
rect 265256 11756 265308 11762
rect 265256 11698 265308 11704
rect 263968 11688 264020 11694
rect 263968 11630 264020 11636
rect 261760 11552 261812 11558
rect 261760 11494 261812 11500
rect 262680 11552 262732 11558
rect 262680 11494 262732 11500
rect 264348 11150 264376 11698
rect 265176 11286 265204 11698
rect 265452 11354 265480 15200
rect 267642 13628 267950 13636
rect 267642 13626 267648 13628
rect 267704 13626 267728 13628
rect 267784 13626 267808 13628
rect 267864 13626 267888 13628
rect 267944 13626 267950 13628
rect 267704 13574 267706 13626
rect 267886 13574 267888 13626
rect 267642 13572 267648 13574
rect 267704 13572 267728 13574
rect 267784 13572 267808 13574
rect 267864 13572 267888 13574
rect 267944 13572 267950 13574
rect 267642 13562 267950 13572
rect 265532 13456 265584 13462
rect 265532 13398 265584 13404
rect 265544 13296 265572 13398
rect 265530 13288 265586 13296
rect 265586 13246 265664 13274
rect 265530 13222 265586 13232
rect 265532 12912 265584 12918
rect 265532 12854 265584 12860
rect 265544 12442 265572 12854
rect 265532 12436 265584 12442
rect 265532 12378 265584 12384
rect 265636 12306 265664 13246
rect 266912 13252 266964 13258
rect 266912 13194 266964 13200
rect 266544 12912 266596 12918
rect 266544 12854 266596 12860
rect 265624 12300 265676 12306
rect 265624 12242 265676 12248
rect 265440 11348 265492 11354
rect 265440 11290 265492 11296
rect 265164 11280 265216 11286
rect 265164 11222 265216 11228
rect 265636 11150 265664 12242
rect 266268 11552 266320 11558
rect 266268 11494 266320 11500
rect 266360 11552 266412 11558
rect 266360 11494 266412 11500
rect 266280 11354 266308 11494
rect 266268 11348 266320 11354
rect 266268 11290 266320 11296
rect 264336 11144 264388 11150
rect 264336 11086 264388 11092
rect 264888 11144 264940 11150
rect 264888 11086 264940 11092
rect 265624 11144 265676 11150
rect 265624 11086 265676 11092
rect 255228 10804 255280 10810
rect 255228 10746 255280 10752
rect 264900 10742 264928 11086
rect 264888 10736 264940 10742
rect 264888 10678 264940 10684
rect 266372 10674 266400 11494
rect 266556 10810 266584 12854
rect 266820 12164 266872 12170
rect 266820 12106 266872 12112
rect 266832 11898 266860 12106
rect 266820 11892 266872 11898
rect 266820 11834 266872 11840
rect 266544 10804 266596 10810
rect 266544 10746 266596 10752
rect 254952 10668 255004 10674
rect 254952 10610 255004 10616
rect 266360 10668 266412 10674
rect 266360 10610 266412 10616
rect 266924 10266 266952 13194
rect 267648 13184 267700 13190
rect 267648 13126 267700 13132
rect 267004 12776 267056 12782
rect 267556 12776 267608 12782
rect 267004 12718 267056 12724
rect 267094 12744 267150 12752
rect 267016 12646 267044 12718
rect 267660 12752 267688 13126
rect 268384 12980 268436 12986
rect 268384 12922 268436 12928
rect 268292 12844 268344 12850
rect 268292 12786 268344 12792
rect 268016 12776 268068 12782
rect 267556 12718 267608 12724
rect 267646 12744 267702 12752
rect 267094 12678 267150 12688
rect 267108 12646 267136 12678
rect 267568 12646 267596 12718
rect 268016 12718 268068 12724
rect 268106 12744 268162 12752
rect 267646 12678 267702 12688
rect 267004 12640 267056 12646
rect 267004 12582 267056 12588
rect 267096 12640 267148 12646
rect 267096 12582 267148 12588
rect 267556 12640 267608 12646
rect 267556 12582 267608 12588
rect 267016 12102 267044 12582
rect 267642 12540 267950 12548
rect 267642 12538 267648 12540
rect 267704 12538 267728 12540
rect 267784 12538 267808 12540
rect 267864 12538 267888 12540
rect 267944 12538 267950 12540
rect 267704 12486 267706 12538
rect 267886 12486 267888 12538
rect 267642 12484 267648 12486
rect 267704 12484 267728 12486
rect 267784 12484 267808 12486
rect 267864 12484 267888 12486
rect 267944 12484 267950 12486
rect 267642 12474 267950 12484
rect 268028 12442 268056 12718
rect 268106 12678 268162 12688
rect 268016 12436 268068 12442
rect 268016 12378 268068 12384
rect 267280 12164 267332 12170
rect 267280 12106 267332 12112
rect 267004 12096 267056 12102
rect 267004 12038 267056 12044
rect 267292 11218 267320 12106
rect 268028 11626 268056 12378
rect 268120 12238 268148 12678
rect 268108 12232 268160 12238
rect 268108 12174 268160 12180
rect 268016 11620 268068 11626
rect 268016 11562 268068 11568
rect 267642 11452 267950 11460
rect 267642 11450 267648 11452
rect 267704 11450 267728 11452
rect 267784 11450 267808 11452
rect 267864 11450 267888 11452
rect 267944 11450 267950 11452
rect 267704 11398 267706 11450
rect 267886 11398 267888 11450
rect 267642 11396 267648 11398
rect 267704 11396 267728 11398
rect 267784 11396 267808 11398
rect 267864 11396 267888 11398
rect 267944 11396 267950 11398
rect 267642 11386 267950 11396
rect 268028 11218 268056 11562
rect 267280 11212 267332 11218
rect 267280 11154 267332 11160
rect 268016 11212 268068 11218
rect 268016 11154 268068 11160
rect 267642 10364 267950 10372
rect 267642 10362 267648 10364
rect 267704 10362 267728 10364
rect 267784 10362 267808 10364
rect 267864 10362 267888 10364
rect 267944 10362 267950 10364
rect 267704 10310 267706 10362
rect 267886 10310 267888 10362
rect 267642 10308 267648 10310
rect 267704 10308 267728 10310
rect 267784 10308 267808 10310
rect 267864 10308 267888 10310
rect 267944 10308 267950 10310
rect 267642 10298 267950 10308
rect 266912 10260 266964 10266
rect 266912 10202 266964 10208
rect 267740 10124 267792 10130
rect 267740 10066 267792 10072
rect 252744 9988 252796 9994
rect 252744 9930 252796 9936
rect 267752 9926 267780 10066
rect 268120 10062 268148 12174
rect 268200 12164 268252 12170
rect 268200 12106 268252 12112
rect 268212 10810 268240 12106
rect 268304 11830 268332 12786
rect 268396 12782 268424 12922
rect 268384 12776 268436 12782
rect 268384 12718 268436 12724
rect 268384 12436 268436 12442
rect 268384 12378 268436 12384
rect 268292 11824 268344 11830
rect 268292 11766 268344 11772
rect 268304 11082 268332 11766
rect 268292 11076 268344 11082
rect 268292 11018 268344 11024
rect 268200 10804 268252 10810
rect 268200 10746 268252 10752
rect 268396 10198 268424 12378
rect 268476 12096 268528 12102
rect 268476 12038 268528 12044
rect 268488 11762 268516 12038
rect 268476 11756 268528 11762
rect 268476 11698 268528 11704
rect 268488 11218 268516 11698
rect 268476 11212 268528 11218
rect 268476 11154 268528 11160
rect 268580 10266 268608 15200
rect 271800 13530 271828 15286
rect 274638 15286 274956 15314
rect 274638 15200 274694 15286
rect 274928 13530 274956 15286
rect 277766 15286 277900 15314
rect 277766 15200 277822 15286
rect 277872 13530 277900 15286
rect 280802 15286 280936 15314
rect 280802 15200 280858 15286
rect 280908 13530 280936 15286
rect 283930 15286 284248 15314
rect 283930 15200 283986 15286
rect 268936 13524 268988 13530
rect 268936 13466 268988 13472
rect 269580 13524 269632 13530
rect 269580 13466 269632 13472
rect 271788 13524 271840 13530
rect 271788 13466 271840 13472
rect 274916 13524 274968 13530
rect 274916 13466 274968 13472
rect 277860 13524 277912 13530
rect 277860 13466 277912 13472
rect 280896 13524 280948 13530
rect 284220 13512 284248 15286
rect 286966 15200 287022 16000
rect 290002 15314 290058 16000
rect 293130 15314 293186 16000
rect 296166 15314 296222 16000
rect 299202 15314 299258 16000
rect 302330 15314 302386 16000
rect 290002 15286 290136 15314
rect 290002 15200 290058 15286
rect 284300 13524 284352 13530
rect 284220 13484 284300 13512
rect 280896 13466 280948 13472
rect 286980 13512 287008 15200
rect 290108 13530 290136 15286
rect 293130 15286 293264 15314
rect 293130 15200 293186 15286
rect 293236 13530 293264 15286
rect 296166 15286 296300 15314
rect 296166 15200 296222 15286
rect 296272 13530 296300 15286
rect 299202 15286 299336 15314
rect 299202 15200 299258 15286
rect 299308 13530 299336 15286
rect 302330 15286 302648 15314
rect 302330 15200 302386 15286
rect 301412 13728 301464 13734
rect 301412 13670 301464 13676
rect 301424 13530 301452 13670
rect 287060 13524 287112 13530
rect 286980 13484 287060 13512
rect 284300 13466 284352 13472
rect 287060 13466 287112 13472
rect 290096 13524 290148 13530
rect 290096 13466 290148 13472
rect 293224 13524 293276 13530
rect 293224 13466 293276 13472
rect 296260 13524 296312 13530
rect 296260 13466 296312 13472
rect 299296 13524 299348 13530
rect 299296 13466 299348 13472
rect 301412 13524 301464 13530
rect 301412 13466 301464 13472
rect 268948 13432 268976 13466
rect 268934 13424 268990 13432
rect 268934 13358 268990 13368
rect 268948 13326 268976 13358
rect 268936 13320 268988 13326
rect 268936 13262 268988 13268
rect 269026 13288 269082 13296
rect 268752 13252 268804 13258
rect 268752 13194 268804 13200
rect 268660 12232 268712 12238
rect 268660 12174 268712 12180
rect 268672 12102 268700 12174
rect 268660 12096 268712 12102
rect 268660 12038 268712 12044
rect 268764 10538 268792 13194
rect 268948 11218 268976 13262
rect 269026 13222 269082 13232
rect 269040 12850 269068 13222
rect 269028 12844 269080 12850
rect 269028 12786 269080 12792
rect 269396 12776 269448 12782
rect 269316 12736 269396 12764
rect 269120 12640 269172 12646
rect 269172 12600 269252 12628
rect 269120 12582 269172 12588
rect 269120 12300 269172 12306
rect 269120 12242 269172 12248
rect 269132 11762 269160 12242
rect 269120 11756 269172 11762
rect 269120 11698 269172 11704
rect 268936 11212 268988 11218
rect 268936 11154 268988 11160
rect 268948 11082 268976 11154
rect 268936 11076 268988 11082
rect 268936 11018 268988 11024
rect 268844 11008 268896 11014
rect 268844 10950 268896 10956
rect 268752 10532 268804 10538
rect 268752 10474 268804 10480
rect 268568 10260 268620 10266
rect 268568 10202 268620 10208
rect 268384 10192 268436 10198
rect 268384 10134 268436 10140
rect 268856 10130 268884 10950
rect 269028 10668 269080 10674
rect 269028 10610 269080 10616
rect 268844 10124 268896 10130
rect 268844 10066 268896 10072
rect 269040 10062 269068 10610
rect 269224 10062 269252 12600
rect 269316 11354 269344 12736
rect 269396 12718 269448 12724
rect 269488 12164 269540 12170
rect 269488 12106 269540 12112
rect 269396 11688 269448 11694
rect 269396 11630 269448 11636
rect 269304 11348 269356 11354
rect 269304 11290 269356 11296
rect 269408 10810 269436 11630
rect 269396 10804 269448 10810
rect 269396 10746 269448 10752
rect 269500 10198 269528 12106
rect 269592 10470 269620 13466
rect 270408 13456 270460 13462
rect 272984 13456 273036 13462
rect 270408 13398 270460 13404
rect 272812 13404 272984 13410
rect 272812 13398 273036 13404
rect 273166 13424 273222 13432
rect 269672 12300 269724 12306
rect 269672 12242 269724 12248
rect 269684 11150 269712 12242
rect 270420 12186 270448 13398
rect 272812 13382 273024 13398
rect 270684 13252 270736 13258
rect 270684 13194 270736 13200
rect 270960 13252 271012 13258
rect 270960 13194 271012 13200
rect 270328 12158 270448 12186
rect 269856 11824 269908 11830
rect 269856 11766 269908 11772
rect 269672 11144 269724 11150
rect 269672 11086 269724 11092
rect 269580 10464 269632 10470
rect 269580 10406 269632 10412
rect 269488 10192 269540 10198
rect 269488 10134 269540 10140
rect 268108 10056 268160 10062
rect 268108 9998 268160 10004
rect 269028 10056 269080 10062
rect 269028 9998 269080 10004
rect 269212 10056 269264 10062
rect 269212 9998 269264 10004
rect 267740 9920 267792 9926
rect 267740 9862 267792 9868
rect 268120 9586 268148 9998
rect 269868 9654 269896 11766
rect 269948 11688 270000 11694
rect 269948 11630 270000 11636
rect 269960 11082 269988 11630
rect 269948 11076 270000 11082
rect 269948 11018 270000 11024
rect 270040 11008 270092 11014
rect 270040 10950 270092 10956
rect 270052 10742 270080 10950
rect 270040 10736 270092 10742
rect 270040 10678 270092 10684
rect 270328 10674 270356 12158
rect 270408 12096 270460 12102
rect 270408 12038 270460 12044
rect 270420 11150 270448 12038
rect 270696 11898 270724 13194
rect 270776 13184 270828 13190
rect 270776 13126 270828 13132
rect 270788 11898 270816 13126
rect 270868 12844 270920 12850
rect 270868 12786 270920 12792
rect 270880 12646 270908 12786
rect 270868 12640 270920 12646
rect 270868 12582 270920 12588
rect 270684 11892 270736 11898
rect 270684 11834 270736 11840
rect 270776 11892 270828 11898
rect 270776 11834 270828 11840
rect 270880 11150 270908 12582
rect 270408 11144 270460 11150
rect 270408 11086 270460 11092
rect 270868 11144 270920 11150
rect 270868 11086 270920 11092
rect 270316 10668 270368 10674
rect 270316 10610 270368 10616
rect 270972 9926 271000 13194
rect 271788 13184 271840 13190
rect 271788 13126 271840 13132
rect 271800 12918 271828 13126
rect 272812 12918 272840 13382
rect 273166 13358 273168 13368
rect 273220 13358 273222 13368
rect 273168 13330 273220 13336
rect 273260 13320 273312 13326
rect 273258 13288 273260 13296
rect 275100 13320 275152 13326
rect 273312 13288 273314 13296
rect 275100 13262 275152 13268
rect 281080 13320 281132 13326
rect 281080 13262 281132 13268
rect 284760 13320 284812 13326
rect 284760 13262 284812 13268
rect 290280 13320 290332 13326
rect 290280 13262 290332 13268
rect 299480 13320 299532 13326
rect 299480 13262 299532 13268
rect 273258 13222 273314 13232
rect 272892 13184 272944 13190
rect 272892 13126 272944 13132
rect 271052 12912 271104 12918
rect 271052 12854 271104 12860
rect 271788 12912 271840 12918
rect 271788 12854 271840 12860
rect 272800 12912 272852 12918
rect 272800 12854 272852 12860
rect 271064 12442 271092 12854
rect 272616 12844 272668 12850
rect 272616 12786 272668 12792
rect 272248 12776 272300 12782
rect 272248 12718 272300 12724
rect 271144 12640 271196 12646
rect 271144 12582 271196 12588
rect 271052 12436 271104 12442
rect 271052 12378 271104 12384
rect 271156 12306 271184 12582
rect 272260 12306 272288 12718
rect 272628 12646 272656 12786
rect 272904 12782 272932 13126
rect 273168 12912 273220 12918
rect 273168 12854 273220 12860
rect 273180 12782 273208 12854
rect 272892 12776 272944 12782
rect 272892 12718 272944 12724
rect 273168 12776 273220 12782
rect 273168 12718 273220 12724
rect 272800 12708 272852 12714
rect 272800 12650 272852 12656
rect 272524 12640 272576 12646
rect 272524 12582 272576 12588
rect 272616 12640 272668 12646
rect 272616 12582 272668 12588
rect 271144 12300 271196 12306
rect 271144 12242 271196 12248
rect 272248 12300 272300 12306
rect 272248 12242 272300 12248
rect 271328 12232 271380 12238
rect 271328 12174 271380 12180
rect 271340 11762 271368 12174
rect 271328 11756 271380 11762
rect 271328 11698 271380 11704
rect 272260 11218 272288 12242
rect 272248 11212 272300 11218
rect 272248 11154 272300 11160
rect 272536 10606 272564 12582
rect 272812 12306 272840 12650
rect 272800 12300 272852 12306
rect 272800 12242 272852 12248
rect 272904 12238 272932 12718
rect 272892 12232 272944 12238
rect 272892 12174 272944 12180
rect 273180 11694 273208 12718
rect 273168 11688 273220 11694
rect 273168 11630 273220 11636
rect 275112 11558 275140 13262
rect 281092 12646 281120 13262
rect 281080 12640 281132 12646
rect 281080 12582 281132 12588
rect 284772 12102 284800 13262
rect 290292 12850 290320 13262
rect 295892 13184 295944 13190
rect 295892 13126 295944 13132
rect 295904 12918 295932 13126
rect 295892 12912 295944 12918
rect 299492 12888 299520 13262
rect 302620 12986 302648 15286
rect 305366 15200 305422 16000
rect 303512 13968 303602 13982
rect 303512 13912 303526 13968
rect 303582 13912 303602 13968
rect 303512 13898 303602 13912
rect 302792 13796 302844 13802
rect 302792 13738 302844 13744
rect 302608 12980 302660 12986
rect 302608 12922 302660 12928
rect 295892 12854 295944 12860
rect 299478 12880 299534 12888
rect 290280 12844 290332 12850
rect 302804 12850 302832 13738
rect 303540 13326 303568 13898
rect 305000 13388 305052 13394
rect 305000 13330 305052 13336
rect 303528 13320 303580 13326
rect 303528 13262 303580 13268
rect 305012 12918 305040 13330
rect 305380 12986 305408 15200
rect 305368 12980 305420 12986
rect 305368 12922 305420 12928
rect 305000 12912 305052 12918
rect 305000 12854 305052 12860
rect 305460 12912 305512 12918
rect 305460 12854 305512 12860
rect 299478 12814 299534 12824
rect 302792 12844 302844 12850
rect 290280 12786 290332 12792
rect 302792 12786 302844 12792
rect 305472 12442 305500 12854
rect 305460 12436 305512 12442
rect 305460 12378 305512 12384
rect 284760 12096 284812 12102
rect 284760 12038 284812 12044
rect 275100 11552 275152 11558
rect 275100 11494 275152 11500
rect 272524 10600 272576 10606
rect 272524 10542 272576 10548
rect 304448 10056 304500 10062
rect 304446 10024 304448 10032
rect 304500 10024 304502 10032
rect 304446 9958 304502 9968
rect 270960 9920 271012 9926
rect 270960 9862 271012 9868
rect 269856 9648 269908 9654
rect 269856 9590 269908 9596
rect 268108 9580 268160 9586
rect 268108 9522 268160 9528
rect 267642 9276 267950 9284
rect 267642 9274 267648 9276
rect 267704 9274 267728 9276
rect 267784 9274 267808 9276
rect 267864 9274 267888 9276
rect 267944 9274 267950 9276
rect 267704 9222 267706 9274
rect 267886 9222 267888 9274
rect 267642 9220 267648 9222
rect 267704 9220 267728 9222
rect 267784 9220 267808 9222
rect 267864 9220 267888 9222
rect 267944 9220 267950 9222
rect 267642 9210 267950 9220
rect 267642 8188 267950 8196
rect 267642 8186 267648 8188
rect 267704 8186 267728 8188
rect 267784 8186 267808 8188
rect 267864 8186 267888 8188
rect 267944 8186 267950 8188
rect 267704 8134 267706 8186
rect 267886 8134 267888 8186
rect 267642 8132 267648 8134
rect 267704 8132 267728 8134
rect 267784 8132 267808 8134
rect 267864 8132 267888 8134
rect 267944 8132 267950 8134
rect 267642 8122 267950 8132
rect 267642 7100 267950 7108
rect 267642 7098 267648 7100
rect 267704 7098 267728 7100
rect 267784 7098 267808 7100
rect 267864 7098 267888 7100
rect 267944 7098 267950 7100
rect 267704 7046 267706 7098
rect 267886 7046 267888 7098
rect 267642 7044 267648 7046
rect 267704 7044 267728 7046
rect 267784 7044 267808 7046
rect 267864 7044 267888 7046
rect 267944 7044 267950 7046
rect 267642 7034 267950 7044
rect 303988 6316 304040 6322
rect 303988 6258 304040 6264
rect 249064 6248 249116 6254
rect 249064 6190 249116 6196
rect 191444 6012 191752 6020
rect 191444 6010 191450 6012
rect 191506 6010 191530 6012
rect 191586 6010 191610 6012
rect 191666 6010 191690 6012
rect 191746 6010 191752 6012
rect 191506 5958 191508 6010
rect 191688 5958 191690 6010
rect 191444 5956 191450 5958
rect 191506 5956 191530 5958
rect 191586 5956 191610 5958
rect 191666 5956 191690 5958
rect 191746 5956 191752 5958
rect 191444 5946 191752 5956
rect 267642 6012 267950 6020
rect 267642 6010 267648 6012
rect 267704 6010 267728 6012
rect 267784 6010 267808 6012
rect 267864 6010 267888 6012
rect 267944 6010 267950 6012
rect 267704 5958 267706 6010
rect 267886 5958 267888 6010
rect 267642 5956 267648 5958
rect 267704 5956 267728 5958
rect 267784 5956 267808 5958
rect 267864 5956 267888 5958
rect 267944 5956 267950 5958
rect 267642 5946 267950 5956
rect 304000 5952 304028 6258
rect 303986 5944 304042 5952
rect 303986 5878 304042 5888
rect 153346 5468 153654 5476
rect 153346 5466 153352 5468
rect 153408 5466 153432 5468
rect 153488 5466 153512 5468
rect 153568 5466 153592 5468
rect 153648 5466 153654 5468
rect 153408 5414 153410 5466
rect 153590 5414 153592 5466
rect 153346 5412 153352 5414
rect 153408 5412 153432 5414
rect 153488 5412 153512 5414
rect 153568 5412 153592 5414
rect 153648 5412 153654 5414
rect 153346 5402 153654 5412
rect 229544 5468 229852 5476
rect 229544 5466 229550 5468
rect 229606 5466 229630 5468
rect 229686 5466 229710 5468
rect 229766 5466 229790 5468
rect 229846 5466 229852 5468
rect 229606 5414 229608 5466
rect 229788 5414 229790 5466
rect 229544 5412 229550 5414
rect 229606 5412 229630 5414
rect 229686 5412 229710 5414
rect 229766 5412 229790 5414
rect 229846 5412 229852 5414
rect 229544 5402 229852 5412
rect 191444 4924 191752 4932
rect 191444 4922 191450 4924
rect 191506 4922 191530 4924
rect 191586 4922 191610 4924
rect 191666 4922 191690 4924
rect 191746 4922 191752 4924
rect 191506 4870 191508 4922
rect 191688 4870 191690 4922
rect 191444 4868 191450 4870
rect 191506 4868 191530 4870
rect 191586 4868 191610 4870
rect 191666 4868 191690 4870
rect 191746 4868 191752 4870
rect 191444 4858 191752 4868
rect 267642 4924 267950 4932
rect 267642 4922 267648 4924
rect 267704 4922 267728 4924
rect 267784 4922 267808 4924
rect 267864 4922 267888 4924
rect 267944 4922 267950 4924
rect 267704 4870 267706 4922
rect 267886 4870 267888 4922
rect 267642 4868 267648 4870
rect 267704 4868 267728 4870
rect 267784 4868 267808 4870
rect 267864 4868 267888 4870
rect 267944 4868 267950 4870
rect 267642 4858 267950 4868
rect 153346 4380 153654 4388
rect 153346 4378 153352 4380
rect 153408 4378 153432 4380
rect 153488 4378 153512 4380
rect 153568 4378 153592 4380
rect 153648 4378 153654 4380
rect 153408 4326 153410 4378
rect 153590 4326 153592 4378
rect 153346 4324 153352 4326
rect 153408 4324 153432 4326
rect 153488 4324 153512 4326
rect 153568 4324 153592 4326
rect 153648 4324 153654 4326
rect 153346 4314 153654 4324
rect 229544 4380 229852 4388
rect 229544 4378 229550 4380
rect 229606 4378 229630 4380
rect 229686 4378 229710 4380
rect 229766 4378 229790 4380
rect 229846 4378 229852 4380
rect 229606 4326 229608 4378
rect 229788 4326 229790 4378
rect 229544 4324 229550 4326
rect 229606 4324 229630 4326
rect 229686 4324 229710 4326
rect 229766 4324 229790 4326
rect 229846 4324 229852 4326
rect 229544 4314 229852 4324
rect 191444 3836 191752 3844
rect 191444 3834 191450 3836
rect 191506 3834 191530 3836
rect 191586 3834 191610 3836
rect 191666 3834 191690 3836
rect 191746 3834 191752 3836
rect 191506 3782 191508 3834
rect 191688 3782 191690 3834
rect 191444 3780 191450 3782
rect 191506 3780 191530 3782
rect 191586 3780 191610 3782
rect 191666 3780 191690 3782
rect 191746 3780 191752 3782
rect 191444 3770 191752 3780
rect 267642 3836 267950 3844
rect 267642 3834 267648 3836
rect 267704 3834 267728 3836
rect 267784 3834 267808 3836
rect 267864 3834 267888 3836
rect 267944 3834 267950 3836
rect 267704 3782 267706 3834
rect 267886 3782 267888 3834
rect 267642 3780 267648 3782
rect 267704 3780 267728 3782
rect 267784 3780 267808 3782
rect 267864 3780 267888 3782
rect 267944 3780 267950 3782
rect 267642 3770 267950 3780
rect 153346 3292 153654 3300
rect 153346 3290 153352 3292
rect 153408 3290 153432 3292
rect 153488 3290 153512 3292
rect 153568 3290 153592 3292
rect 153648 3290 153654 3292
rect 153408 3238 153410 3290
rect 153590 3238 153592 3290
rect 153346 3236 153352 3238
rect 153408 3236 153432 3238
rect 153488 3236 153512 3238
rect 153568 3236 153592 3238
rect 153648 3236 153654 3238
rect 153346 3226 153654 3236
rect 229544 3292 229852 3300
rect 229544 3290 229550 3292
rect 229606 3290 229630 3292
rect 229686 3290 229710 3292
rect 229766 3290 229790 3292
rect 229846 3290 229852 3292
rect 229606 3238 229608 3290
rect 229788 3238 229790 3290
rect 229544 3236 229550 3238
rect 229606 3236 229630 3238
rect 229686 3236 229710 3238
rect 229766 3236 229790 3238
rect 229846 3236 229852 3238
rect 229544 3226 229852 3236
rect 191444 2748 191752 2756
rect 191444 2746 191450 2748
rect 191506 2746 191530 2748
rect 191586 2746 191610 2748
rect 191666 2746 191690 2748
rect 191746 2746 191752 2748
rect 191506 2694 191508 2746
rect 191688 2694 191690 2746
rect 191444 2692 191450 2694
rect 191506 2692 191530 2694
rect 191586 2692 191610 2694
rect 191666 2692 191690 2694
rect 191746 2692 191752 2694
rect 191444 2682 191752 2692
rect 267642 2748 267950 2756
rect 267642 2746 267648 2748
rect 267704 2746 267728 2748
rect 267784 2746 267808 2748
rect 267864 2746 267888 2748
rect 267944 2746 267950 2748
rect 267704 2694 267706 2746
rect 267886 2694 267888 2746
rect 267642 2692 267648 2694
rect 267704 2692 267728 2694
rect 267784 2692 267808 2694
rect 267864 2692 267888 2694
rect 267944 2692 267950 2694
rect 267642 2682 267950 2692
rect 149428 2644 149480 2650
rect 149428 2586 149480 2592
rect 302240 2644 302292 2650
rect 302240 2586 302292 2592
rect 77148 2204 77456 2212
rect 77148 2202 77154 2204
rect 77210 2202 77234 2204
rect 77290 2202 77314 2204
rect 77370 2202 77394 2204
rect 77450 2202 77456 2204
rect 77210 2150 77212 2202
rect 77392 2150 77394 2202
rect 77148 2148 77154 2150
rect 77210 2148 77234 2150
rect 77290 2148 77314 2150
rect 77370 2148 77394 2150
rect 77450 2148 77456 2150
rect 77148 2138 77456 2148
rect 153346 2204 153654 2212
rect 153346 2202 153352 2204
rect 153408 2202 153432 2204
rect 153488 2202 153512 2204
rect 153568 2202 153592 2204
rect 153648 2202 153654 2204
rect 153408 2150 153410 2202
rect 153590 2150 153592 2202
rect 153346 2148 153352 2150
rect 153408 2148 153432 2150
rect 153488 2148 153512 2150
rect 153568 2148 153592 2150
rect 153648 2148 153654 2150
rect 153346 2138 153654 2148
rect 229544 2204 229852 2212
rect 229544 2202 229550 2204
rect 229606 2202 229630 2204
rect 229686 2202 229710 2204
rect 229766 2202 229790 2204
rect 229846 2202 229852 2204
rect 229606 2150 229608 2202
rect 229788 2150 229790 2202
rect 229544 2148 229550 2150
rect 229606 2148 229630 2150
rect 229686 2148 229710 2150
rect 229766 2148 229790 2150
rect 229846 2148 229852 2150
rect 229544 2138 229852 2148
rect 302252 2008 302280 2586
rect 302238 2000 302294 2008
rect 302238 1934 302294 1944
<< via2 >>
rect 29366 12180 29368 12200
rect 29368 12180 29420 12200
rect 29420 12180 29422 12200
rect 29366 12144 29422 12180
rect 30746 12144 30802 12200
rect 31390 12144 31446 12200
rect 39054 13626 39110 13628
rect 39134 13626 39190 13628
rect 39214 13626 39270 13628
rect 39294 13626 39350 13628
rect 39054 13574 39100 13626
rect 39100 13574 39110 13626
rect 39134 13574 39164 13626
rect 39164 13574 39176 13626
rect 39176 13574 39190 13626
rect 39214 13574 39228 13626
rect 39228 13574 39240 13626
rect 39240 13574 39270 13626
rect 39294 13574 39304 13626
rect 39304 13574 39350 13626
rect 39054 13572 39110 13574
rect 39134 13572 39190 13574
rect 39214 13572 39270 13574
rect 39294 13572 39350 13574
rect 39054 12538 39110 12540
rect 39134 12538 39190 12540
rect 39214 12538 39270 12540
rect 39294 12538 39350 12540
rect 39054 12486 39100 12538
rect 39100 12486 39110 12538
rect 39134 12486 39164 12538
rect 39164 12486 39176 12538
rect 39176 12486 39190 12538
rect 39214 12486 39228 12538
rect 39228 12486 39240 12538
rect 39240 12486 39270 12538
rect 39294 12486 39304 12538
rect 39304 12486 39350 12538
rect 39054 12484 39110 12486
rect 39134 12484 39190 12486
rect 39214 12484 39270 12486
rect 39294 12484 39350 12486
rect 39054 11450 39110 11452
rect 39134 11450 39190 11452
rect 39214 11450 39270 11452
rect 39294 11450 39350 11452
rect 39054 11398 39100 11450
rect 39100 11398 39110 11450
rect 39134 11398 39164 11450
rect 39164 11398 39176 11450
rect 39176 11398 39190 11450
rect 39214 11398 39228 11450
rect 39228 11398 39240 11450
rect 39240 11398 39270 11450
rect 39294 11398 39304 11450
rect 39304 11398 39350 11450
rect 39054 11396 39110 11398
rect 39134 11396 39190 11398
rect 39214 11396 39270 11398
rect 39294 11396 39350 11398
rect 40590 12180 40592 12200
rect 40592 12180 40644 12200
rect 40644 12180 40646 12200
rect 40590 12144 40646 12180
rect 42430 12144 42486 12200
rect 77154 13082 77210 13084
rect 77234 13082 77290 13084
rect 77314 13082 77370 13084
rect 77394 13082 77450 13084
rect 77154 13030 77200 13082
rect 77200 13030 77210 13082
rect 77234 13030 77264 13082
rect 77264 13030 77276 13082
rect 77276 13030 77290 13082
rect 77314 13030 77328 13082
rect 77328 13030 77340 13082
rect 77340 13030 77370 13082
rect 77394 13030 77404 13082
rect 77404 13030 77450 13082
rect 77154 13028 77210 13030
rect 77234 13028 77290 13030
rect 77314 13028 77370 13030
rect 77394 13028 77450 13030
rect 77154 11994 77210 11996
rect 77234 11994 77290 11996
rect 77314 11994 77370 11996
rect 77394 11994 77450 11996
rect 77154 11942 77200 11994
rect 77200 11942 77210 11994
rect 77234 11942 77264 11994
rect 77264 11942 77276 11994
rect 77276 11942 77290 11994
rect 77314 11942 77328 11994
rect 77328 11942 77340 11994
rect 77340 11942 77370 11994
rect 77394 11942 77404 11994
rect 77404 11942 77450 11994
rect 77154 11940 77210 11942
rect 77234 11940 77290 11942
rect 77314 11940 77370 11942
rect 77394 11940 77450 11942
rect 86958 13096 87014 13152
rect 87786 12688 87842 12744
rect 88154 12300 88210 12336
rect 88154 12280 88156 12300
rect 88156 12280 88208 12300
rect 88208 12280 88210 12300
rect 91834 13096 91890 13152
rect 89902 12280 89958 12336
rect 90730 12688 90786 12744
rect 77154 10906 77210 10908
rect 77234 10906 77290 10908
rect 77314 10906 77370 10908
rect 77394 10906 77450 10908
rect 77154 10854 77200 10906
rect 77200 10854 77210 10906
rect 77234 10854 77264 10906
rect 77264 10854 77276 10906
rect 77276 10854 77290 10906
rect 77314 10854 77328 10906
rect 77328 10854 77340 10906
rect 77340 10854 77370 10906
rect 77394 10854 77404 10906
rect 77404 10854 77450 10906
rect 77154 10852 77210 10854
rect 77234 10852 77290 10854
rect 77314 10852 77370 10854
rect 77394 10852 77450 10854
rect 39054 10362 39110 10364
rect 39134 10362 39190 10364
rect 39214 10362 39270 10364
rect 39294 10362 39350 10364
rect 39054 10310 39100 10362
rect 39100 10310 39110 10362
rect 39134 10310 39164 10362
rect 39164 10310 39176 10362
rect 39176 10310 39190 10362
rect 39214 10310 39228 10362
rect 39228 10310 39240 10362
rect 39240 10310 39270 10362
rect 39294 10310 39304 10362
rect 39304 10310 39350 10362
rect 39054 10308 39110 10310
rect 39134 10308 39190 10310
rect 39214 10308 39270 10310
rect 39294 10308 39350 10310
rect 77154 9818 77210 9820
rect 77234 9818 77290 9820
rect 77314 9818 77370 9820
rect 77394 9818 77450 9820
rect 77154 9766 77200 9818
rect 77200 9766 77210 9818
rect 77234 9766 77264 9818
rect 77264 9766 77276 9818
rect 77276 9766 77290 9818
rect 77314 9766 77328 9818
rect 77328 9766 77340 9818
rect 77340 9766 77370 9818
rect 77394 9766 77404 9818
rect 77404 9766 77450 9818
rect 77154 9764 77210 9766
rect 77234 9764 77290 9766
rect 77314 9764 77370 9766
rect 77394 9764 77450 9766
rect 115252 13626 115308 13628
rect 115332 13626 115388 13628
rect 115412 13626 115468 13628
rect 115492 13626 115548 13628
rect 115252 13574 115298 13626
rect 115298 13574 115308 13626
rect 115332 13574 115362 13626
rect 115362 13574 115374 13626
rect 115374 13574 115388 13626
rect 115412 13574 115426 13626
rect 115426 13574 115438 13626
rect 115438 13574 115468 13626
rect 115492 13574 115502 13626
rect 115502 13574 115548 13626
rect 115252 13572 115308 13574
rect 115332 13572 115388 13574
rect 115412 13572 115468 13574
rect 115492 13572 115548 13574
rect 115252 12538 115308 12540
rect 115332 12538 115388 12540
rect 115412 12538 115468 12540
rect 115492 12538 115548 12540
rect 115252 12486 115298 12538
rect 115298 12486 115308 12538
rect 115332 12486 115362 12538
rect 115362 12486 115374 12538
rect 115374 12486 115388 12538
rect 115412 12486 115426 12538
rect 115426 12486 115438 12538
rect 115438 12486 115468 12538
rect 115492 12486 115502 12538
rect 115502 12486 115548 12538
rect 115252 12484 115308 12486
rect 115332 12484 115388 12486
rect 115412 12484 115468 12486
rect 115492 12484 115548 12486
rect 115252 11450 115308 11452
rect 115332 11450 115388 11452
rect 115412 11450 115468 11452
rect 115492 11450 115548 11452
rect 115252 11398 115298 11450
rect 115298 11398 115308 11450
rect 115332 11398 115362 11450
rect 115362 11398 115374 11450
rect 115374 11398 115388 11450
rect 115412 11398 115426 11450
rect 115426 11398 115438 11450
rect 115438 11398 115468 11450
rect 115492 11398 115502 11450
rect 115502 11398 115548 11450
rect 115252 11396 115308 11398
rect 115332 11396 115388 11398
rect 115412 11396 115468 11398
rect 115492 11396 115548 11398
rect 115252 10362 115308 10364
rect 115332 10362 115388 10364
rect 115412 10362 115468 10364
rect 115492 10362 115548 10364
rect 115252 10310 115298 10362
rect 115298 10310 115308 10362
rect 115332 10310 115362 10362
rect 115362 10310 115374 10362
rect 115374 10310 115388 10362
rect 115412 10310 115426 10362
rect 115426 10310 115438 10362
rect 115438 10310 115468 10362
rect 115492 10310 115502 10362
rect 115502 10310 115548 10362
rect 115252 10308 115308 10310
rect 115332 10308 115388 10310
rect 115412 10308 115468 10310
rect 115492 10308 115548 10310
rect 39054 9274 39110 9276
rect 39134 9274 39190 9276
rect 39214 9274 39270 9276
rect 39294 9274 39350 9276
rect 39054 9222 39100 9274
rect 39100 9222 39110 9274
rect 39134 9222 39164 9274
rect 39164 9222 39176 9274
rect 39176 9222 39190 9274
rect 39214 9222 39228 9274
rect 39228 9222 39240 9274
rect 39240 9222 39270 9274
rect 39294 9222 39304 9274
rect 39304 9222 39350 9274
rect 39054 9220 39110 9222
rect 39134 9220 39190 9222
rect 39214 9220 39270 9222
rect 39294 9220 39350 9222
rect 115252 9274 115308 9276
rect 115332 9274 115388 9276
rect 115412 9274 115468 9276
rect 115492 9274 115548 9276
rect 115252 9222 115298 9274
rect 115298 9222 115308 9274
rect 115332 9222 115362 9274
rect 115362 9222 115374 9274
rect 115374 9222 115388 9274
rect 115412 9222 115426 9274
rect 115426 9222 115438 9274
rect 115438 9222 115468 9274
rect 115492 9222 115502 9274
rect 115502 9222 115548 9274
rect 115252 9220 115308 9222
rect 115332 9220 115388 9222
rect 115412 9220 115468 9222
rect 115492 9220 115548 9222
rect 77154 8730 77210 8732
rect 77234 8730 77290 8732
rect 77314 8730 77370 8732
rect 77394 8730 77450 8732
rect 77154 8678 77200 8730
rect 77200 8678 77210 8730
rect 77234 8678 77264 8730
rect 77264 8678 77276 8730
rect 77276 8678 77290 8730
rect 77314 8678 77328 8730
rect 77328 8678 77340 8730
rect 77340 8678 77370 8730
rect 77394 8678 77404 8730
rect 77404 8678 77450 8730
rect 77154 8676 77210 8678
rect 77234 8676 77290 8678
rect 77314 8676 77370 8678
rect 77394 8676 77450 8678
rect 39054 8186 39110 8188
rect 39134 8186 39190 8188
rect 39214 8186 39270 8188
rect 39294 8186 39350 8188
rect 39054 8134 39100 8186
rect 39100 8134 39110 8186
rect 39134 8134 39164 8186
rect 39164 8134 39176 8186
rect 39176 8134 39190 8186
rect 39214 8134 39228 8186
rect 39228 8134 39240 8186
rect 39240 8134 39270 8186
rect 39294 8134 39304 8186
rect 39304 8134 39350 8186
rect 39054 8132 39110 8134
rect 39134 8132 39190 8134
rect 39214 8132 39270 8134
rect 39294 8132 39350 8134
rect 115252 8186 115308 8188
rect 115332 8186 115388 8188
rect 115412 8186 115468 8188
rect 115492 8186 115548 8188
rect 115252 8134 115298 8186
rect 115298 8134 115308 8186
rect 115332 8134 115362 8186
rect 115362 8134 115374 8186
rect 115374 8134 115388 8186
rect 115412 8134 115426 8186
rect 115426 8134 115438 8186
rect 115438 8134 115468 8186
rect 115492 8134 115502 8186
rect 115502 8134 115548 8186
rect 115252 8132 115308 8134
rect 115332 8132 115388 8134
rect 115412 8132 115468 8134
rect 115492 8132 115548 8134
rect 1398 8064 1454 8120
rect 77154 7642 77210 7644
rect 77234 7642 77290 7644
rect 77314 7642 77370 7644
rect 77394 7642 77450 7644
rect 77154 7590 77200 7642
rect 77200 7590 77210 7642
rect 77234 7590 77264 7642
rect 77264 7590 77276 7642
rect 77276 7590 77290 7642
rect 77314 7590 77328 7642
rect 77328 7590 77340 7642
rect 77340 7590 77370 7642
rect 77394 7590 77404 7642
rect 77404 7590 77450 7642
rect 77154 7588 77210 7590
rect 77234 7588 77290 7590
rect 77314 7588 77370 7590
rect 77394 7588 77450 7590
rect 39054 7098 39110 7100
rect 39134 7098 39190 7100
rect 39214 7098 39270 7100
rect 39294 7098 39350 7100
rect 39054 7046 39100 7098
rect 39100 7046 39110 7098
rect 39134 7046 39164 7098
rect 39164 7046 39176 7098
rect 39176 7046 39190 7098
rect 39214 7046 39228 7098
rect 39228 7046 39240 7098
rect 39240 7046 39270 7098
rect 39294 7046 39304 7098
rect 39304 7046 39350 7098
rect 39054 7044 39110 7046
rect 39134 7044 39190 7046
rect 39214 7044 39270 7046
rect 39294 7044 39350 7046
rect 115252 7098 115308 7100
rect 115332 7098 115388 7100
rect 115412 7098 115468 7100
rect 115492 7098 115548 7100
rect 115252 7046 115298 7098
rect 115298 7046 115308 7098
rect 115332 7046 115362 7098
rect 115362 7046 115374 7098
rect 115374 7046 115388 7098
rect 115412 7046 115426 7098
rect 115426 7046 115438 7098
rect 115438 7046 115468 7098
rect 115492 7046 115502 7098
rect 115502 7046 115548 7098
rect 115252 7044 115308 7046
rect 115332 7044 115388 7046
rect 115412 7044 115468 7046
rect 115492 7044 115548 7046
rect 77154 6554 77210 6556
rect 77234 6554 77290 6556
rect 77314 6554 77370 6556
rect 77394 6554 77450 6556
rect 77154 6502 77200 6554
rect 77200 6502 77210 6554
rect 77234 6502 77264 6554
rect 77264 6502 77276 6554
rect 77276 6502 77290 6554
rect 77314 6502 77328 6554
rect 77328 6502 77340 6554
rect 77340 6502 77370 6554
rect 77394 6502 77404 6554
rect 77404 6502 77450 6554
rect 77154 6500 77210 6502
rect 77234 6500 77290 6502
rect 77314 6500 77370 6502
rect 77394 6500 77450 6502
rect 39054 6010 39110 6012
rect 39134 6010 39190 6012
rect 39214 6010 39270 6012
rect 39294 6010 39350 6012
rect 39054 5958 39100 6010
rect 39100 5958 39110 6010
rect 39134 5958 39164 6010
rect 39164 5958 39176 6010
rect 39176 5958 39190 6010
rect 39214 5958 39228 6010
rect 39228 5958 39240 6010
rect 39240 5958 39270 6010
rect 39294 5958 39304 6010
rect 39304 5958 39350 6010
rect 39054 5956 39110 5958
rect 39134 5956 39190 5958
rect 39214 5956 39270 5958
rect 39294 5956 39350 5958
rect 115252 6010 115308 6012
rect 115332 6010 115388 6012
rect 115412 6010 115468 6012
rect 115492 6010 115548 6012
rect 115252 5958 115298 6010
rect 115298 5958 115308 6010
rect 115332 5958 115362 6010
rect 115362 5958 115374 6010
rect 115374 5958 115388 6010
rect 115412 5958 115426 6010
rect 115426 5958 115438 6010
rect 115438 5958 115468 6010
rect 115492 5958 115502 6010
rect 115502 5958 115548 6010
rect 115252 5956 115308 5958
rect 115332 5956 115388 5958
rect 115412 5956 115468 5958
rect 115492 5956 115548 5958
rect 77154 5466 77210 5468
rect 77234 5466 77290 5468
rect 77314 5466 77370 5468
rect 77394 5466 77450 5468
rect 77154 5414 77200 5466
rect 77200 5414 77210 5466
rect 77234 5414 77264 5466
rect 77264 5414 77276 5466
rect 77276 5414 77290 5466
rect 77314 5414 77328 5466
rect 77328 5414 77340 5466
rect 77340 5414 77370 5466
rect 77394 5414 77404 5466
rect 77404 5414 77450 5466
rect 77154 5412 77210 5414
rect 77234 5412 77290 5414
rect 77314 5412 77370 5414
rect 77394 5412 77450 5414
rect 39054 4922 39110 4924
rect 39134 4922 39190 4924
rect 39214 4922 39270 4924
rect 39294 4922 39350 4924
rect 39054 4870 39100 4922
rect 39100 4870 39110 4922
rect 39134 4870 39164 4922
rect 39164 4870 39176 4922
rect 39176 4870 39190 4922
rect 39214 4870 39228 4922
rect 39228 4870 39240 4922
rect 39240 4870 39270 4922
rect 39294 4870 39304 4922
rect 39304 4870 39350 4922
rect 39054 4868 39110 4870
rect 39134 4868 39190 4870
rect 39214 4868 39270 4870
rect 39294 4868 39350 4870
rect 115252 4922 115308 4924
rect 115332 4922 115388 4924
rect 115412 4922 115468 4924
rect 115492 4922 115548 4924
rect 115252 4870 115298 4922
rect 115298 4870 115308 4922
rect 115332 4870 115362 4922
rect 115362 4870 115374 4922
rect 115374 4870 115388 4922
rect 115412 4870 115426 4922
rect 115426 4870 115438 4922
rect 115438 4870 115468 4922
rect 115492 4870 115502 4922
rect 115502 4870 115548 4922
rect 115252 4868 115308 4870
rect 115332 4868 115388 4870
rect 115412 4868 115468 4870
rect 115492 4868 115548 4870
rect 77154 4378 77210 4380
rect 77234 4378 77290 4380
rect 77314 4378 77370 4380
rect 77394 4378 77450 4380
rect 77154 4326 77200 4378
rect 77200 4326 77210 4378
rect 77234 4326 77264 4378
rect 77264 4326 77276 4378
rect 77276 4326 77290 4378
rect 77314 4326 77328 4378
rect 77328 4326 77340 4378
rect 77340 4326 77370 4378
rect 77394 4326 77404 4378
rect 77404 4326 77450 4378
rect 77154 4324 77210 4326
rect 77234 4324 77290 4326
rect 77314 4324 77370 4326
rect 77394 4324 77450 4326
rect 39054 3834 39110 3836
rect 39134 3834 39190 3836
rect 39214 3834 39270 3836
rect 39294 3834 39350 3836
rect 39054 3782 39100 3834
rect 39100 3782 39110 3834
rect 39134 3782 39164 3834
rect 39164 3782 39176 3834
rect 39176 3782 39190 3834
rect 39214 3782 39228 3834
rect 39228 3782 39240 3834
rect 39240 3782 39270 3834
rect 39294 3782 39304 3834
rect 39304 3782 39350 3834
rect 39054 3780 39110 3782
rect 39134 3780 39190 3782
rect 39214 3780 39270 3782
rect 39294 3780 39350 3782
rect 115252 3834 115308 3836
rect 115332 3834 115388 3836
rect 115412 3834 115468 3836
rect 115492 3834 115548 3836
rect 115252 3782 115298 3834
rect 115298 3782 115308 3834
rect 115332 3782 115362 3834
rect 115362 3782 115374 3834
rect 115374 3782 115388 3834
rect 115412 3782 115426 3834
rect 115426 3782 115438 3834
rect 115438 3782 115468 3834
rect 115492 3782 115502 3834
rect 115502 3782 115548 3834
rect 115252 3780 115308 3782
rect 115332 3780 115388 3782
rect 115412 3780 115468 3782
rect 115492 3780 115548 3782
rect 77154 3290 77210 3292
rect 77234 3290 77290 3292
rect 77314 3290 77370 3292
rect 77394 3290 77450 3292
rect 77154 3238 77200 3290
rect 77200 3238 77210 3290
rect 77234 3238 77264 3290
rect 77264 3238 77276 3290
rect 77276 3238 77290 3290
rect 77314 3238 77328 3290
rect 77328 3238 77340 3290
rect 77340 3238 77370 3290
rect 77394 3238 77404 3290
rect 77404 3238 77450 3290
rect 77154 3236 77210 3238
rect 77234 3236 77290 3238
rect 77314 3236 77370 3238
rect 77394 3236 77450 3238
rect 39054 2746 39110 2748
rect 39134 2746 39190 2748
rect 39214 2746 39270 2748
rect 39294 2746 39350 2748
rect 39054 2694 39100 2746
rect 39100 2694 39110 2746
rect 39134 2694 39164 2746
rect 39164 2694 39176 2746
rect 39176 2694 39190 2746
rect 39214 2694 39228 2746
rect 39228 2694 39240 2746
rect 39240 2694 39270 2746
rect 39294 2694 39304 2746
rect 39304 2694 39350 2746
rect 39054 2692 39110 2694
rect 39134 2692 39190 2694
rect 39214 2692 39270 2694
rect 39294 2692 39350 2694
rect 115252 2746 115308 2748
rect 115332 2746 115388 2748
rect 115412 2746 115468 2748
rect 115492 2746 115548 2748
rect 115252 2694 115298 2746
rect 115298 2694 115308 2746
rect 115332 2694 115362 2746
rect 115362 2694 115374 2746
rect 115374 2694 115388 2746
rect 115412 2694 115426 2746
rect 115426 2694 115438 2746
rect 115438 2694 115468 2746
rect 115492 2694 115502 2746
rect 115502 2694 115548 2746
rect 115252 2692 115308 2694
rect 115332 2692 115388 2694
rect 115412 2692 115468 2694
rect 115492 2692 115548 2694
rect 153352 13082 153408 13084
rect 153432 13082 153488 13084
rect 153512 13082 153568 13084
rect 153592 13082 153648 13084
rect 153352 13030 153398 13082
rect 153398 13030 153408 13082
rect 153432 13030 153462 13082
rect 153462 13030 153474 13082
rect 153474 13030 153488 13082
rect 153512 13030 153526 13082
rect 153526 13030 153538 13082
rect 153538 13030 153568 13082
rect 153592 13030 153602 13082
rect 153602 13030 153648 13082
rect 153352 13028 153408 13030
rect 153432 13028 153488 13030
rect 153512 13028 153568 13030
rect 153592 13028 153648 13030
rect 153352 11994 153408 11996
rect 153432 11994 153488 11996
rect 153512 11994 153568 11996
rect 153592 11994 153648 11996
rect 153352 11942 153398 11994
rect 153398 11942 153408 11994
rect 153432 11942 153462 11994
rect 153462 11942 153474 11994
rect 153474 11942 153488 11994
rect 153512 11942 153526 11994
rect 153526 11942 153538 11994
rect 153538 11942 153568 11994
rect 153592 11942 153602 11994
rect 153602 11942 153648 11994
rect 153352 11940 153408 11942
rect 153432 11940 153488 11942
rect 153512 11940 153568 11942
rect 153592 11940 153648 11942
rect 155038 12824 155094 12880
rect 157890 12588 157892 12608
rect 157892 12588 157944 12608
rect 157944 12588 157946 12608
rect 157890 12552 157946 12588
rect 153352 10906 153408 10908
rect 153432 10906 153488 10908
rect 153512 10906 153568 10908
rect 153592 10906 153648 10908
rect 153352 10854 153398 10906
rect 153398 10854 153408 10906
rect 153432 10854 153462 10906
rect 153462 10854 153474 10906
rect 153474 10854 153488 10906
rect 153512 10854 153526 10906
rect 153526 10854 153538 10906
rect 153538 10854 153568 10906
rect 153592 10854 153602 10906
rect 153602 10854 153648 10906
rect 153352 10852 153408 10854
rect 153432 10852 153488 10854
rect 153512 10852 153568 10854
rect 153592 10852 153648 10854
rect 153352 9818 153408 9820
rect 153432 9818 153488 9820
rect 153512 9818 153568 9820
rect 153592 9818 153648 9820
rect 153352 9766 153398 9818
rect 153398 9766 153408 9818
rect 153432 9766 153462 9818
rect 153462 9766 153474 9818
rect 153474 9766 153488 9818
rect 153512 9766 153526 9818
rect 153526 9766 153538 9818
rect 153538 9766 153568 9818
rect 153592 9766 153602 9818
rect 153602 9766 153648 9818
rect 153352 9764 153408 9766
rect 153432 9764 153488 9766
rect 153512 9764 153568 9766
rect 153592 9764 153648 9766
rect 160282 12588 160284 12608
rect 160284 12588 160336 12608
rect 160336 12588 160338 12608
rect 160282 12552 160338 12588
rect 163594 12300 163650 12336
rect 163594 12280 163596 12300
rect 163596 12280 163648 12300
rect 163648 12280 163650 12300
rect 189630 11756 189686 11792
rect 189630 11736 189632 11756
rect 189632 11736 189684 11756
rect 189684 11736 189686 11756
rect 153352 8730 153408 8732
rect 153432 8730 153488 8732
rect 153512 8730 153568 8732
rect 153592 8730 153648 8732
rect 153352 8678 153398 8730
rect 153398 8678 153408 8730
rect 153432 8678 153462 8730
rect 153462 8678 153474 8730
rect 153474 8678 153488 8730
rect 153512 8678 153526 8730
rect 153526 8678 153538 8730
rect 153538 8678 153568 8730
rect 153592 8678 153602 8730
rect 153602 8678 153648 8730
rect 153352 8676 153408 8678
rect 153432 8676 153488 8678
rect 153512 8676 153568 8678
rect 153592 8676 153648 8678
rect 191450 13626 191506 13628
rect 191530 13626 191586 13628
rect 191610 13626 191666 13628
rect 191690 13626 191746 13628
rect 191450 13574 191496 13626
rect 191496 13574 191506 13626
rect 191530 13574 191560 13626
rect 191560 13574 191572 13626
rect 191572 13574 191586 13626
rect 191610 13574 191624 13626
rect 191624 13574 191636 13626
rect 191636 13574 191666 13626
rect 191690 13574 191700 13626
rect 191700 13574 191746 13626
rect 191450 13572 191506 13574
rect 191530 13572 191586 13574
rect 191610 13572 191666 13574
rect 191690 13572 191746 13574
rect 191838 12552 191894 12608
rect 191450 12538 191506 12540
rect 191530 12538 191586 12540
rect 191610 12538 191666 12540
rect 191690 12538 191746 12540
rect 191450 12486 191496 12538
rect 191496 12486 191506 12538
rect 191530 12486 191560 12538
rect 191560 12486 191572 12538
rect 191572 12486 191586 12538
rect 191610 12486 191624 12538
rect 191624 12486 191636 12538
rect 191636 12486 191666 12538
rect 191690 12486 191700 12538
rect 191700 12486 191746 12538
rect 191450 12484 191506 12486
rect 191530 12484 191586 12486
rect 191610 12484 191666 12486
rect 191690 12484 191746 12486
rect 192206 12552 192262 12608
rect 191450 11450 191506 11452
rect 191530 11450 191586 11452
rect 191610 11450 191666 11452
rect 191690 11450 191746 11452
rect 191450 11398 191496 11450
rect 191496 11398 191506 11450
rect 191530 11398 191560 11450
rect 191560 11398 191572 11450
rect 191572 11398 191586 11450
rect 191610 11398 191624 11450
rect 191624 11398 191636 11450
rect 191636 11398 191666 11450
rect 191690 11398 191700 11450
rect 191700 11398 191746 11450
rect 191450 11396 191506 11398
rect 191530 11396 191586 11398
rect 191610 11396 191666 11398
rect 191690 11396 191746 11398
rect 191450 10362 191506 10364
rect 191530 10362 191586 10364
rect 191610 10362 191666 10364
rect 191690 10362 191746 10364
rect 191450 10310 191496 10362
rect 191496 10310 191506 10362
rect 191530 10310 191560 10362
rect 191560 10310 191572 10362
rect 191572 10310 191586 10362
rect 191610 10310 191624 10362
rect 191624 10310 191636 10362
rect 191636 10310 191666 10362
rect 191690 10310 191700 10362
rect 191700 10310 191746 10362
rect 191450 10308 191506 10310
rect 191530 10308 191586 10310
rect 191610 10308 191666 10310
rect 191690 10308 191746 10310
rect 193034 12280 193090 12336
rect 193034 11736 193090 11792
rect 194598 12824 194654 12880
rect 195058 12688 195114 12744
rect 195794 12824 195850 12880
rect 197358 12844 197414 12880
rect 197358 12824 197360 12844
rect 197360 12824 197412 12844
rect 197412 12824 197414 12844
rect 200854 13232 200910 13288
rect 200394 12552 200450 12608
rect 203430 13232 203486 13288
rect 207110 13524 207166 13560
rect 207110 13504 207112 13524
rect 207112 13504 207164 13524
rect 207164 13504 207166 13524
rect 205546 13232 205602 13288
rect 205270 12588 205272 12608
rect 205272 12588 205324 12608
rect 205324 12588 205326 12608
rect 205270 12552 205326 12588
rect 205730 13232 205786 13288
rect 207202 13268 207204 13288
rect 207204 13268 207256 13288
rect 207256 13268 207258 13288
rect 207202 13232 207258 13268
rect 208030 13504 208086 13560
rect 213274 13404 213276 13424
rect 213276 13404 213328 13424
rect 213328 13404 213330 13424
rect 213274 13368 213330 13404
rect 219806 13368 219862 13424
rect 207938 13268 207940 13288
rect 207940 13268 207992 13288
rect 207992 13268 207994 13288
rect 207938 13232 207994 13268
rect 207846 12688 207902 12744
rect 225418 13132 225420 13152
rect 225420 13132 225472 13152
rect 225472 13132 225474 13152
rect 225418 13096 225474 13132
rect 227074 13388 227130 13424
rect 227074 13368 227076 13388
rect 227076 13368 227128 13388
rect 227128 13368 227130 13388
rect 227074 13132 227076 13152
rect 227076 13132 227128 13152
rect 227128 13132 227130 13152
rect 227074 13096 227130 13132
rect 229190 13404 229192 13424
rect 229192 13404 229244 13424
rect 229244 13404 229246 13424
rect 229190 13368 229246 13404
rect 230386 13268 230388 13288
rect 230388 13268 230440 13288
rect 230440 13268 230442 13288
rect 230386 13232 230442 13268
rect 229550 13082 229606 13084
rect 229630 13082 229686 13084
rect 229710 13082 229766 13084
rect 229790 13082 229846 13084
rect 229550 13030 229596 13082
rect 229596 13030 229606 13082
rect 229630 13030 229660 13082
rect 229660 13030 229672 13082
rect 229672 13030 229686 13082
rect 229710 13030 229724 13082
rect 229724 13030 229736 13082
rect 229736 13030 229766 13082
rect 229790 13030 229800 13082
rect 229800 13030 229846 13082
rect 229550 13028 229606 13030
rect 229630 13028 229686 13030
rect 229710 13028 229766 13030
rect 229790 13028 229846 13030
rect 229550 11994 229606 11996
rect 229630 11994 229686 11996
rect 229710 11994 229766 11996
rect 229790 11994 229846 11996
rect 229550 11942 229596 11994
rect 229596 11942 229606 11994
rect 229630 11942 229660 11994
rect 229660 11942 229672 11994
rect 229672 11942 229686 11994
rect 229710 11942 229724 11994
rect 229724 11942 229736 11994
rect 229736 11942 229766 11994
rect 229790 11942 229800 11994
rect 229800 11942 229846 11994
rect 229550 11940 229606 11942
rect 229630 11940 229686 11942
rect 229710 11940 229766 11942
rect 229790 11940 229846 11942
rect 232134 13232 232190 13288
rect 238114 13388 238170 13424
rect 238114 13368 238116 13388
rect 238116 13368 238168 13388
rect 238168 13368 238170 13388
rect 239494 13404 239496 13424
rect 239496 13404 239548 13424
rect 239548 13404 239550 13424
rect 239494 13368 239550 13404
rect 238298 12688 238354 12744
rect 242162 12708 242218 12744
rect 242162 12688 242164 12708
rect 242164 12688 242216 12708
rect 242216 12688 242218 12708
rect 229550 10906 229606 10908
rect 229630 10906 229686 10908
rect 229710 10906 229766 10908
rect 229790 10906 229846 10908
rect 229550 10854 229596 10906
rect 229596 10854 229606 10906
rect 229630 10854 229660 10906
rect 229660 10854 229672 10906
rect 229672 10854 229686 10906
rect 229710 10854 229724 10906
rect 229724 10854 229736 10906
rect 229736 10854 229766 10906
rect 229790 10854 229800 10906
rect 229800 10854 229846 10906
rect 229550 10852 229606 10854
rect 229630 10852 229686 10854
rect 229710 10852 229766 10854
rect 229790 10852 229846 10854
rect 229550 9818 229606 9820
rect 229630 9818 229686 9820
rect 229710 9818 229766 9820
rect 229790 9818 229846 9820
rect 229550 9766 229596 9818
rect 229596 9766 229606 9818
rect 229630 9766 229660 9818
rect 229660 9766 229672 9818
rect 229672 9766 229686 9818
rect 229710 9766 229724 9818
rect 229724 9766 229736 9818
rect 229736 9766 229766 9818
rect 229790 9766 229800 9818
rect 229800 9766 229846 9818
rect 229550 9764 229606 9766
rect 229630 9764 229686 9766
rect 229710 9764 229766 9766
rect 229790 9764 229846 9766
rect 191450 9274 191506 9276
rect 191530 9274 191586 9276
rect 191610 9274 191666 9276
rect 191690 9274 191746 9276
rect 191450 9222 191496 9274
rect 191496 9222 191506 9274
rect 191530 9222 191560 9274
rect 191560 9222 191572 9274
rect 191572 9222 191586 9274
rect 191610 9222 191624 9274
rect 191624 9222 191636 9274
rect 191636 9222 191666 9274
rect 191690 9222 191700 9274
rect 191700 9222 191746 9274
rect 191450 9220 191506 9222
rect 191530 9220 191586 9222
rect 191610 9220 191666 9222
rect 191690 9220 191746 9222
rect 229550 8730 229606 8732
rect 229630 8730 229686 8732
rect 229710 8730 229766 8732
rect 229790 8730 229846 8732
rect 229550 8678 229596 8730
rect 229596 8678 229606 8730
rect 229630 8678 229660 8730
rect 229660 8678 229672 8730
rect 229672 8678 229686 8730
rect 229710 8678 229724 8730
rect 229724 8678 229736 8730
rect 229736 8678 229766 8730
rect 229790 8678 229800 8730
rect 229800 8678 229846 8730
rect 229550 8676 229606 8678
rect 229630 8676 229686 8678
rect 229710 8676 229766 8678
rect 229790 8676 229846 8678
rect 191450 8186 191506 8188
rect 191530 8186 191586 8188
rect 191610 8186 191666 8188
rect 191690 8186 191746 8188
rect 191450 8134 191496 8186
rect 191496 8134 191506 8186
rect 191530 8134 191560 8186
rect 191560 8134 191572 8186
rect 191572 8134 191586 8186
rect 191610 8134 191624 8186
rect 191624 8134 191636 8186
rect 191636 8134 191666 8186
rect 191690 8134 191700 8186
rect 191700 8134 191746 8186
rect 191450 8132 191506 8134
rect 191530 8132 191586 8134
rect 191610 8132 191666 8134
rect 191690 8132 191746 8134
rect 153352 7642 153408 7644
rect 153432 7642 153488 7644
rect 153512 7642 153568 7644
rect 153592 7642 153648 7644
rect 153352 7590 153398 7642
rect 153398 7590 153408 7642
rect 153432 7590 153462 7642
rect 153462 7590 153474 7642
rect 153474 7590 153488 7642
rect 153512 7590 153526 7642
rect 153526 7590 153538 7642
rect 153538 7590 153568 7642
rect 153592 7590 153602 7642
rect 153602 7590 153648 7642
rect 153352 7588 153408 7590
rect 153432 7588 153488 7590
rect 153512 7588 153568 7590
rect 153592 7588 153648 7590
rect 229550 7642 229606 7644
rect 229630 7642 229686 7644
rect 229710 7642 229766 7644
rect 229790 7642 229846 7644
rect 229550 7590 229596 7642
rect 229596 7590 229606 7642
rect 229630 7590 229660 7642
rect 229660 7590 229672 7642
rect 229672 7590 229686 7642
rect 229710 7590 229724 7642
rect 229724 7590 229736 7642
rect 229736 7590 229766 7642
rect 229790 7590 229800 7642
rect 229800 7590 229846 7642
rect 229550 7588 229606 7590
rect 229630 7588 229686 7590
rect 229710 7588 229766 7590
rect 229790 7588 229846 7590
rect 191450 7098 191506 7100
rect 191530 7098 191586 7100
rect 191610 7098 191666 7100
rect 191690 7098 191746 7100
rect 191450 7046 191496 7098
rect 191496 7046 191506 7098
rect 191530 7046 191560 7098
rect 191560 7046 191572 7098
rect 191572 7046 191586 7098
rect 191610 7046 191624 7098
rect 191624 7046 191636 7098
rect 191636 7046 191666 7098
rect 191690 7046 191700 7098
rect 191700 7046 191746 7098
rect 191450 7044 191506 7046
rect 191530 7044 191586 7046
rect 191610 7044 191666 7046
rect 191690 7044 191746 7046
rect 153352 6554 153408 6556
rect 153432 6554 153488 6556
rect 153512 6554 153568 6556
rect 153592 6554 153648 6556
rect 153352 6502 153398 6554
rect 153398 6502 153408 6554
rect 153432 6502 153462 6554
rect 153462 6502 153474 6554
rect 153474 6502 153488 6554
rect 153512 6502 153526 6554
rect 153526 6502 153538 6554
rect 153538 6502 153568 6554
rect 153592 6502 153602 6554
rect 153602 6502 153648 6554
rect 153352 6500 153408 6502
rect 153432 6500 153488 6502
rect 153512 6500 153568 6502
rect 153592 6500 153648 6502
rect 229550 6554 229606 6556
rect 229630 6554 229686 6556
rect 229710 6554 229766 6556
rect 229790 6554 229846 6556
rect 229550 6502 229596 6554
rect 229596 6502 229606 6554
rect 229630 6502 229660 6554
rect 229660 6502 229672 6554
rect 229672 6502 229686 6554
rect 229710 6502 229724 6554
rect 229724 6502 229736 6554
rect 229736 6502 229766 6554
rect 229790 6502 229800 6554
rect 229800 6502 229846 6554
rect 229550 6500 229606 6502
rect 229630 6500 229686 6502
rect 229710 6500 229766 6502
rect 229790 6500 229846 6502
rect 251914 12588 251916 12608
rect 251916 12588 251968 12608
rect 251968 12588 251970 12608
rect 251914 12552 251970 12588
rect 251822 12416 251878 12472
rect 256606 12960 256662 13016
rect 257986 12960 258042 13016
rect 257066 12552 257122 12608
rect 257158 12416 257214 12472
rect 262310 12724 262312 12744
rect 262312 12724 262364 12744
rect 262364 12724 262366 12744
rect 262310 12688 262366 12724
rect 263414 13252 263470 13288
rect 263414 13232 263416 13252
rect 263416 13232 263468 13252
rect 263468 13232 263470 13252
rect 263506 12708 263562 12744
rect 263506 12688 263508 12708
rect 263508 12688 263560 12708
rect 263560 12688 263562 12708
rect 264334 12688 264390 12744
rect 267648 13626 267704 13628
rect 267728 13626 267784 13628
rect 267808 13626 267864 13628
rect 267888 13626 267944 13628
rect 267648 13574 267694 13626
rect 267694 13574 267704 13626
rect 267728 13574 267758 13626
rect 267758 13574 267770 13626
rect 267770 13574 267784 13626
rect 267808 13574 267822 13626
rect 267822 13574 267834 13626
rect 267834 13574 267864 13626
rect 267888 13574 267898 13626
rect 267898 13574 267944 13626
rect 267648 13572 267704 13574
rect 267728 13572 267784 13574
rect 267808 13572 267864 13574
rect 267888 13572 267944 13574
rect 265530 13232 265586 13288
rect 267094 12688 267150 12744
rect 267646 12688 267702 12744
rect 267648 12538 267704 12540
rect 267728 12538 267784 12540
rect 267808 12538 267864 12540
rect 267888 12538 267944 12540
rect 267648 12486 267694 12538
rect 267694 12486 267704 12538
rect 267728 12486 267758 12538
rect 267758 12486 267770 12538
rect 267770 12486 267784 12538
rect 267808 12486 267822 12538
rect 267822 12486 267834 12538
rect 267834 12486 267864 12538
rect 267888 12486 267898 12538
rect 267898 12486 267944 12538
rect 267648 12484 267704 12486
rect 267728 12484 267784 12486
rect 267808 12484 267864 12486
rect 267888 12484 267944 12486
rect 268106 12688 268162 12744
rect 267648 11450 267704 11452
rect 267728 11450 267784 11452
rect 267808 11450 267864 11452
rect 267888 11450 267944 11452
rect 267648 11398 267694 11450
rect 267694 11398 267704 11450
rect 267728 11398 267758 11450
rect 267758 11398 267770 11450
rect 267770 11398 267784 11450
rect 267808 11398 267822 11450
rect 267822 11398 267834 11450
rect 267834 11398 267864 11450
rect 267888 11398 267898 11450
rect 267898 11398 267944 11450
rect 267648 11396 267704 11398
rect 267728 11396 267784 11398
rect 267808 11396 267864 11398
rect 267888 11396 267944 11398
rect 267648 10362 267704 10364
rect 267728 10362 267784 10364
rect 267808 10362 267864 10364
rect 267888 10362 267944 10364
rect 267648 10310 267694 10362
rect 267694 10310 267704 10362
rect 267728 10310 267758 10362
rect 267758 10310 267770 10362
rect 267770 10310 267784 10362
rect 267808 10310 267822 10362
rect 267822 10310 267834 10362
rect 267834 10310 267864 10362
rect 267888 10310 267898 10362
rect 267898 10310 267944 10362
rect 267648 10308 267704 10310
rect 267728 10308 267784 10310
rect 267808 10308 267864 10310
rect 267888 10308 267944 10310
rect 268934 13368 268990 13424
rect 269026 13232 269082 13288
rect 273166 13388 273222 13424
rect 273166 13368 273168 13388
rect 273168 13368 273220 13388
rect 273220 13368 273222 13388
rect 273258 13268 273260 13288
rect 273260 13268 273312 13288
rect 273312 13268 273314 13288
rect 273258 13232 273314 13268
rect 303526 13912 303582 13968
rect 299478 12824 299534 12880
rect 304446 10004 304448 10024
rect 304448 10004 304500 10024
rect 304500 10004 304502 10024
rect 304446 9968 304502 10004
rect 267648 9274 267704 9276
rect 267728 9274 267784 9276
rect 267808 9274 267864 9276
rect 267888 9274 267944 9276
rect 267648 9222 267694 9274
rect 267694 9222 267704 9274
rect 267728 9222 267758 9274
rect 267758 9222 267770 9274
rect 267770 9222 267784 9274
rect 267808 9222 267822 9274
rect 267822 9222 267834 9274
rect 267834 9222 267864 9274
rect 267888 9222 267898 9274
rect 267898 9222 267944 9274
rect 267648 9220 267704 9222
rect 267728 9220 267784 9222
rect 267808 9220 267864 9222
rect 267888 9220 267944 9222
rect 267648 8186 267704 8188
rect 267728 8186 267784 8188
rect 267808 8186 267864 8188
rect 267888 8186 267944 8188
rect 267648 8134 267694 8186
rect 267694 8134 267704 8186
rect 267728 8134 267758 8186
rect 267758 8134 267770 8186
rect 267770 8134 267784 8186
rect 267808 8134 267822 8186
rect 267822 8134 267834 8186
rect 267834 8134 267864 8186
rect 267888 8134 267898 8186
rect 267898 8134 267944 8186
rect 267648 8132 267704 8134
rect 267728 8132 267784 8134
rect 267808 8132 267864 8134
rect 267888 8132 267944 8134
rect 267648 7098 267704 7100
rect 267728 7098 267784 7100
rect 267808 7098 267864 7100
rect 267888 7098 267944 7100
rect 267648 7046 267694 7098
rect 267694 7046 267704 7098
rect 267728 7046 267758 7098
rect 267758 7046 267770 7098
rect 267770 7046 267784 7098
rect 267808 7046 267822 7098
rect 267822 7046 267834 7098
rect 267834 7046 267864 7098
rect 267888 7046 267898 7098
rect 267898 7046 267944 7098
rect 267648 7044 267704 7046
rect 267728 7044 267784 7046
rect 267808 7044 267864 7046
rect 267888 7044 267944 7046
rect 191450 6010 191506 6012
rect 191530 6010 191586 6012
rect 191610 6010 191666 6012
rect 191690 6010 191746 6012
rect 191450 5958 191496 6010
rect 191496 5958 191506 6010
rect 191530 5958 191560 6010
rect 191560 5958 191572 6010
rect 191572 5958 191586 6010
rect 191610 5958 191624 6010
rect 191624 5958 191636 6010
rect 191636 5958 191666 6010
rect 191690 5958 191700 6010
rect 191700 5958 191746 6010
rect 191450 5956 191506 5958
rect 191530 5956 191586 5958
rect 191610 5956 191666 5958
rect 191690 5956 191746 5958
rect 267648 6010 267704 6012
rect 267728 6010 267784 6012
rect 267808 6010 267864 6012
rect 267888 6010 267944 6012
rect 267648 5958 267694 6010
rect 267694 5958 267704 6010
rect 267728 5958 267758 6010
rect 267758 5958 267770 6010
rect 267770 5958 267784 6010
rect 267808 5958 267822 6010
rect 267822 5958 267834 6010
rect 267834 5958 267864 6010
rect 267888 5958 267898 6010
rect 267898 5958 267944 6010
rect 267648 5956 267704 5958
rect 267728 5956 267784 5958
rect 267808 5956 267864 5958
rect 267888 5956 267944 5958
rect 303986 5888 304042 5944
rect 153352 5466 153408 5468
rect 153432 5466 153488 5468
rect 153512 5466 153568 5468
rect 153592 5466 153648 5468
rect 153352 5414 153398 5466
rect 153398 5414 153408 5466
rect 153432 5414 153462 5466
rect 153462 5414 153474 5466
rect 153474 5414 153488 5466
rect 153512 5414 153526 5466
rect 153526 5414 153538 5466
rect 153538 5414 153568 5466
rect 153592 5414 153602 5466
rect 153602 5414 153648 5466
rect 153352 5412 153408 5414
rect 153432 5412 153488 5414
rect 153512 5412 153568 5414
rect 153592 5412 153648 5414
rect 229550 5466 229606 5468
rect 229630 5466 229686 5468
rect 229710 5466 229766 5468
rect 229790 5466 229846 5468
rect 229550 5414 229596 5466
rect 229596 5414 229606 5466
rect 229630 5414 229660 5466
rect 229660 5414 229672 5466
rect 229672 5414 229686 5466
rect 229710 5414 229724 5466
rect 229724 5414 229736 5466
rect 229736 5414 229766 5466
rect 229790 5414 229800 5466
rect 229800 5414 229846 5466
rect 229550 5412 229606 5414
rect 229630 5412 229686 5414
rect 229710 5412 229766 5414
rect 229790 5412 229846 5414
rect 191450 4922 191506 4924
rect 191530 4922 191586 4924
rect 191610 4922 191666 4924
rect 191690 4922 191746 4924
rect 191450 4870 191496 4922
rect 191496 4870 191506 4922
rect 191530 4870 191560 4922
rect 191560 4870 191572 4922
rect 191572 4870 191586 4922
rect 191610 4870 191624 4922
rect 191624 4870 191636 4922
rect 191636 4870 191666 4922
rect 191690 4870 191700 4922
rect 191700 4870 191746 4922
rect 191450 4868 191506 4870
rect 191530 4868 191586 4870
rect 191610 4868 191666 4870
rect 191690 4868 191746 4870
rect 267648 4922 267704 4924
rect 267728 4922 267784 4924
rect 267808 4922 267864 4924
rect 267888 4922 267944 4924
rect 267648 4870 267694 4922
rect 267694 4870 267704 4922
rect 267728 4870 267758 4922
rect 267758 4870 267770 4922
rect 267770 4870 267784 4922
rect 267808 4870 267822 4922
rect 267822 4870 267834 4922
rect 267834 4870 267864 4922
rect 267888 4870 267898 4922
rect 267898 4870 267944 4922
rect 267648 4868 267704 4870
rect 267728 4868 267784 4870
rect 267808 4868 267864 4870
rect 267888 4868 267944 4870
rect 153352 4378 153408 4380
rect 153432 4378 153488 4380
rect 153512 4378 153568 4380
rect 153592 4378 153648 4380
rect 153352 4326 153398 4378
rect 153398 4326 153408 4378
rect 153432 4326 153462 4378
rect 153462 4326 153474 4378
rect 153474 4326 153488 4378
rect 153512 4326 153526 4378
rect 153526 4326 153538 4378
rect 153538 4326 153568 4378
rect 153592 4326 153602 4378
rect 153602 4326 153648 4378
rect 153352 4324 153408 4326
rect 153432 4324 153488 4326
rect 153512 4324 153568 4326
rect 153592 4324 153648 4326
rect 229550 4378 229606 4380
rect 229630 4378 229686 4380
rect 229710 4378 229766 4380
rect 229790 4378 229846 4380
rect 229550 4326 229596 4378
rect 229596 4326 229606 4378
rect 229630 4326 229660 4378
rect 229660 4326 229672 4378
rect 229672 4326 229686 4378
rect 229710 4326 229724 4378
rect 229724 4326 229736 4378
rect 229736 4326 229766 4378
rect 229790 4326 229800 4378
rect 229800 4326 229846 4378
rect 229550 4324 229606 4326
rect 229630 4324 229686 4326
rect 229710 4324 229766 4326
rect 229790 4324 229846 4326
rect 191450 3834 191506 3836
rect 191530 3834 191586 3836
rect 191610 3834 191666 3836
rect 191690 3834 191746 3836
rect 191450 3782 191496 3834
rect 191496 3782 191506 3834
rect 191530 3782 191560 3834
rect 191560 3782 191572 3834
rect 191572 3782 191586 3834
rect 191610 3782 191624 3834
rect 191624 3782 191636 3834
rect 191636 3782 191666 3834
rect 191690 3782 191700 3834
rect 191700 3782 191746 3834
rect 191450 3780 191506 3782
rect 191530 3780 191586 3782
rect 191610 3780 191666 3782
rect 191690 3780 191746 3782
rect 267648 3834 267704 3836
rect 267728 3834 267784 3836
rect 267808 3834 267864 3836
rect 267888 3834 267944 3836
rect 267648 3782 267694 3834
rect 267694 3782 267704 3834
rect 267728 3782 267758 3834
rect 267758 3782 267770 3834
rect 267770 3782 267784 3834
rect 267808 3782 267822 3834
rect 267822 3782 267834 3834
rect 267834 3782 267864 3834
rect 267888 3782 267898 3834
rect 267898 3782 267944 3834
rect 267648 3780 267704 3782
rect 267728 3780 267784 3782
rect 267808 3780 267864 3782
rect 267888 3780 267944 3782
rect 153352 3290 153408 3292
rect 153432 3290 153488 3292
rect 153512 3290 153568 3292
rect 153592 3290 153648 3292
rect 153352 3238 153398 3290
rect 153398 3238 153408 3290
rect 153432 3238 153462 3290
rect 153462 3238 153474 3290
rect 153474 3238 153488 3290
rect 153512 3238 153526 3290
rect 153526 3238 153538 3290
rect 153538 3238 153568 3290
rect 153592 3238 153602 3290
rect 153602 3238 153648 3290
rect 153352 3236 153408 3238
rect 153432 3236 153488 3238
rect 153512 3236 153568 3238
rect 153592 3236 153648 3238
rect 229550 3290 229606 3292
rect 229630 3290 229686 3292
rect 229710 3290 229766 3292
rect 229790 3290 229846 3292
rect 229550 3238 229596 3290
rect 229596 3238 229606 3290
rect 229630 3238 229660 3290
rect 229660 3238 229672 3290
rect 229672 3238 229686 3290
rect 229710 3238 229724 3290
rect 229724 3238 229736 3290
rect 229736 3238 229766 3290
rect 229790 3238 229800 3290
rect 229800 3238 229846 3290
rect 229550 3236 229606 3238
rect 229630 3236 229686 3238
rect 229710 3236 229766 3238
rect 229790 3236 229846 3238
rect 191450 2746 191506 2748
rect 191530 2746 191586 2748
rect 191610 2746 191666 2748
rect 191690 2746 191746 2748
rect 191450 2694 191496 2746
rect 191496 2694 191506 2746
rect 191530 2694 191560 2746
rect 191560 2694 191572 2746
rect 191572 2694 191586 2746
rect 191610 2694 191624 2746
rect 191624 2694 191636 2746
rect 191636 2694 191666 2746
rect 191690 2694 191700 2746
rect 191700 2694 191746 2746
rect 191450 2692 191506 2694
rect 191530 2692 191586 2694
rect 191610 2692 191666 2694
rect 191690 2692 191746 2694
rect 267648 2746 267704 2748
rect 267728 2746 267784 2748
rect 267808 2746 267864 2748
rect 267888 2746 267944 2748
rect 267648 2694 267694 2746
rect 267694 2694 267704 2746
rect 267728 2694 267758 2746
rect 267758 2694 267770 2746
rect 267770 2694 267784 2746
rect 267808 2694 267822 2746
rect 267822 2694 267834 2746
rect 267834 2694 267864 2746
rect 267888 2694 267898 2746
rect 267898 2694 267944 2746
rect 267648 2692 267704 2694
rect 267728 2692 267784 2694
rect 267808 2692 267864 2694
rect 267888 2692 267944 2694
rect 77154 2202 77210 2204
rect 77234 2202 77290 2204
rect 77314 2202 77370 2204
rect 77394 2202 77450 2204
rect 77154 2150 77200 2202
rect 77200 2150 77210 2202
rect 77234 2150 77264 2202
rect 77264 2150 77276 2202
rect 77276 2150 77290 2202
rect 77314 2150 77328 2202
rect 77328 2150 77340 2202
rect 77340 2150 77370 2202
rect 77394 2150 77404 2202
rect 77404 2150 77450 2202
rect 77154 2148 77210 2150
rect 77234 2148 77290 2150
rect 77314 2148 77370 2150
rect 77394 2148 77450 2150
rect 153352 2202 153408 2204
rect 153432 2202 153488 2204
rect 153512 2202 153568 2204
rect 153592 2202 153648 2204
rect 153352 2150 153398 2202
rect 153398 2150 153408 2202
rect 153432 2150 153462 2202
rect 153462 2150 153474 2202
rect 153474 2150 153488 2202
rect 153512 2150 153526 2202
rect 153526 2150 153538 2202
rect 153538 2150 153568 2202
rect 153592 2150 153602 2202
rect 153602 2150 153648 2202
rect 153352 2148 153408 2150
rect 153432 2148 153488 2150
rect 153512 2148 153568 2150
rect 153592 2148 153648 2150
rect 229550 2202 229606 2204
rect 229630 2202 229686 2204
rect 229710 2202 229766 2204
rect 229790 2202 229846 2204
rect 229550 2150 229596 2202
rect 229596 2150 229606 2202
rect 229630 2150 229660 2202
rect 229660 2150 229672 2202
rect 229672 2150 229686 2202
rect 229710 2150 229724 2202
rect 229724 2150 229736 2202
rect 229736 2150 229766 2202
rect 229790 2150 229800 2202
rect 229800 2150 229846 2202
rect 229550 2148 229606 2150
rect 229630 2148 229686 2150
rect 229710 2148 229766 2150
rect 229790 2148 229846 2150
rect 302238 1944 302294 2000
<< metal3 >>
rect 303512 13970 303602 13982
rect 306200 13970 307000 14000
rect 303512 13968 307000 13970
rect 303512 13912 303526 13968
rect 303582 13912 307000 13968
rect 303512 13910 307000 13912
rect 303512 13898 303602 13910
rect 306200 13880 307000 13910
rect 39044 13568 39050 13632
rect 39114 13568 39130 13632
rect 39194 13568 39210 13632
rect 39274 13568 39290 13632
rect 39354 13568 39360 13632
rect 39044 13566 39360 13568
rect 115242 13568 115248 13632
rect 115312 13568 115328 13632
rect 115392 13568 115408 13632
rect 115472 13568 115488 13632
rect 115552 13568 115558 13632
rect 115242 13566 115558 13568
rect 191440 13568 191446 13632
rect 191510 13568 191526 13632
rect 191590 13568 191606 13632
rect 191670 13568 191686 13632
rect 191750 13568 191756 13632
rect 191440 13566 191756 13568
rect 267638 13568 267644 13632
rect 267708 13568 267724 13632
rect 267788 13568 267804 13632
rect 267868 13568 267884 13632
rect 267948 13568 267954 13632
rect 267638 13566 267954 13568
rect 207104 13562 207170 13564
rect 208024 13562 208090 13564
rect 207104 13560 208090 13562
rect 207104 13504 207110 13560
rect 207166 13504 208030 13560
rect 208086 13504 208090 13560
rect 207104 13502 208090 13504
rect 207104 13498 207170 13502
rect 208024 13498 208090 13502
rect 213268 13426 213334 13428
rect 219800 13426 219866 13428
rect 213268 13424 219866 13426
rect 213268 13368 213274 13424
rect 213330 13368 219806 13424
rect 219862 13368 219866 13424
rect 213268 13366 219866 13368
rect 213268 13362 213334 13366
rect 219800 13362 219866 13366
rect 227068 13426 227134 13428
rect 229184 13426 229250 13428
rect 227068 13424 229250 13426
rect 227068 13368 227074 13424
rect 227130 13368 229190 13424
rect 229246 13368 229250 13424
rect 227068 13366 229250 13368
rect 227068 13362 227134 13366
rect 229184 13362 229250 13366
rect 238108 13426 238174 13428
rect 239488 13426 239554 13428
rect 238108 13424 239554 13426
rect 238108 13368 238114 13424
rect 238170 13368 239494 13424
rect 239550 13368 239554 13424
rect 238108 13366 239554 13368
rect 238108 13362 238174 13366
rect 239488 13362 239554 13366
rect 268928 13426 268994 13428
rect 273160 13426 273226 13428
rect 268928 13424 273226 13426
rect 268928 13368 268934 13424
rect 268990 13368 273166 13424
rect 273222 13368 273226 13424
rect 268928 13366 273226 13368
rect 268928 13362 268994 13366
rect 273160 13362 273226 13366
rect 200848 13290 200914 13292
rect 203424 13290 203490 13292
rect 200848 13288 203490 13290
rect 200848 13232 200854 13288
rect 200910 13232 203430 13288
rect 203486 13232 203490 13288
rect 200848 13230 203490 13232
rect 200848 13226 200914 13230
rect 203424 13226 203490 13230
rect 205540 13290 205606 13292
rect 205724 13290 205790 13292
rect 205540 13288 205790 13290
rect 205540 13232 205546 13288
rect 205602 13232 205730 13288
rect 205786 13232 205790 13288
rect 205540 13230 205790 13232
rect 205540 13226 205606 13230
rect 205724 13226 205790 13230
rect 207196 13290 207262 13292
rect 207932 13290 207998 13292
rect 207196 13288 207998 13290
rect 207196 13232 207202 13288
rect 207258 13232 207938 13288
rect 207994 13232 207998 13288
rect 207196 13230 207998 13232
rect 207196 13226 207262 13230
rect 207932 13226 207998 13230
rect 230380 13290 230446 13292
rect 232128 13290 232194 13292
rect 230380 13288 232194 13290
rect 230380 13232 230386 13288
rect 230442 13232 232134 13288
rect 232190 13232 232194 13288
rect 230380 13230 232194 13232
rect 230380 13226 230446 13230
rect 232128 13226 232194 13230
rect 263408 13290 263474 13292
rect 265524 13290 265590 13292
rect 263408 13288 265590 13290
rect 263408 13232 263414 13288
rect 263470 13232 265530 13288
rect 265586 13232 265590 13288
rect 263408 13230 265590 13232
rect 263408 13226 263474 13230
rect 265524 13226 265590 13230
rect 269020 13290 269086 13292
rect 273252 13290 273318 13292
rect 269020 13288 273318 13290
rect 269020 13232 269026 13288
rect 269082 13232 273258 13288
rect 273314 13232 273318 13288
rect 269020 13230 273318 13232
rect 269020 13226 269086 13230
rect 273252 13226 273318 13230
rect 86952 13154 87018 13156
rect 91828 13154 91894 13156
rect 86952 13152 91894 13154
rect 86952 13096 86958 13152
rect 87014 13096 91834 13152
rect 91890 13096 91894 13152
rect 86952 13094 91894 13096
rect 86952 13090 87018 13094
rect 91828 13090 91894 13094
rect 225412 13154 225478 13156
rect 227068 13154 227134 13156
rect 225412 13152 227134 13154
rect 225412 13096 225418 13152
rect 225474 13096 227074 13152
rect 227130 13096 227134 13152
rect 225412 13094 227134 13096
rect 225412 13090 225478 13094
rect 227068 13090 227134 13094
rect 77144 13024 77150 13088
rect 77214 13024 77230 13088
rect 77294 13024 77310 13088
rect 77374 13024 77390 13088
rect 77454 13024 77460 13088
rect 77144 13022 77460 13024
rect 153342 13024 153348 13088
rect 153412 13024 153428 13088
rect 153492 13024 153508 13088
rect 153572 13024 153588 13088
rect 153652 13024 153658 13088
rect 153342 13022 153658 13024
rect 229540 13024 229546 13088
rect 229610 13024 229626 13088
rect 229690 13024 229706 13088
rect 229770 13024 229786 13088
rect 229850 13024 229856 13088
rect 229540 13022 229856 13024
rect 256600 13018 256666 13020
rect 257980 13018 258046 13020
rect 256600 13016 258046 13018
rect 256600 12960 256606 13016
rect 256662 12960 257986 13016
rect 258042 12960 258046 13016
rect 256600 12958 258046 12960
rect 256600 12954 256666 12958
rect 257980 12954 258046 12958
rect 155032 12882 155098 12884
rect 194592 12882 194658 12884
rect 195788 12882 195854 12884
rect 155032 12880 195854 12882
rect 155032 12824 155038 12880
rect 155094 12824 194598 12880
rect 194654 12824 195794 12880
rect 195850 12824 195854 12880
rect 155032 12822 195854 12824
rect 155032 12818 155098 12822
rect 194592 12818 194658 12822
rect 195788 12818 195854 12822
rect 197352 12882 197418 12884
rect 299472 12882 299538 12884
rect 197352 12880 299538 12882
rect 197352 12824 197358 12880
rect 197414 12824 299478 12880
rect 299534 12824 299538 12880
rect 197352 12822 299538 12824
rect 197352 12818 197418 12822
rect 299472 12818 299538 12822
rect 87780 12746 87846 12748
rect 90724 12746 90790 12748
rect 87780 12744 90790 12746
rect 87780 12688 87786 12744
rect 87842 12688 90730 12744
rect 90786 12688 90790 12744
rect 87780 12686 90790 12688
rect 87780 12682 87846 12686
rect 90724 12682 90790 12686
rect 195052 12746 195118 12748
rect 207840 12746 207906 12748
rect 195052 12744 207906 12746
rect 195052 12688 195058 12744
rect 195114 12688 207846 12744
rect 207902 12688 207906 12744
rect 195052 12686 207906 12688
rect 195052 12682 195118 12686
rect 207840 12682 207906 12686
rect 238292 12746 238358 12748
rect 242156 12746 242222 12748
rect 238292 12744 242222 12746
rect 238292 12688 238298 12744
rect 238354 12688 242162 12744
rect 242218 12688 242222 12744
rect 238292 12686 242222 12688
rect 238292 12682 238358 12686
rect 242156 12682 242222 12686
rect 262304 12746 262370 12748
rect 263500 12746 263566 12748
rect 262304 12744 263566 12746
rect 262304 12688 262310 12744
rect 262366 12688 263506 12744
rect 263562 12688 263566 12744
rect 262304 12686 263566 12688
rect 262304 12682 262370 12686
rect 263500 12682 263566 12686
rect 264328 12746 264394 12748
rect 267088 12746 267154 12748
rect 264328 12744 267154 12746
rect 264328 12688 264334 12744
rect 264390 12688 267094 12744
rect 267150 12688 267154 12744
rect 264328 12686 267154 12688
rect 264328 12682 264394 12686
rect 267088 12682 267154 12686
rect 267640 12746 267706 12748
rect 268100 12746 268166 12748
rect 267640 12744 268166 12746
rect 267640 12688 267646 12744
rect 267702 12688 268106 12744
rect 268162 12688 268166 12744
rect 267640 12686 268166 12688
rect 267640 12682 267706 12686
rect 268100 12682 268166 12686
rect 157884 12610 157950 12612
rect 160276 12610 160342 12612
rect 157884 12608 160342 12610
rect 157884 12552 157890 12608
rect 157946 12552 160282 12608
rect 160338 12552 160342 12608
rect 157884 12550 160342 12552
rect 157884 12546 157950 12550
rect 160276 12546 160342 12550
rect 191832 12610 191898 12612
rect 192200 12610 192266 12612
rect 191832 12608 192266 12610
rect 191832 12552 191838 12608
rect 191894 12552 192206 12608
rect 192262 12552 192266 12608
rect 191832 12550 192266 12552
rect 191832 12546 191898 12550
rect 192200 12546 192266 12550
rect 200388 12610 200454 12612
rect 205264 12610 205330 12612
rect 200388 12608 205330 12610
rect 200388 12552 200394 12608
rect 200450 12552 205270 12608
rect 205326 12552 205330 12608
rect 200388 12550 205330 12552
rect 200388 12546 200454 12550
rect 205264 12546 205330 12550
rect 251908 12610 251974 12612
rect 257060 12610 257126 12612
rect 251908 12608 257126 12610
rect 251908 12552 251914 12608
rect 251970 12552 257066 12608
rect 257122 12552 257126 12608
rect 251908 12550 257126 12552
rect 251908 12546 251974 12550
rect 257060 12546 257126 12550
rect 39044 12480 39050 12544
rect 39114 12480 39130 12544
rect 39194 12480 39210 12544
rect 39274 12480 39290 12544
rect 39354 12480 39360 12544
rect 39044 12478 39360 12480
rect 115242 12480 115248 12544
rect 115312 12480 115328 12544
rect 115392 12480 115408 12544
rect 115472 12480 115488 12544
rect 115552 12480 115558 12544
rect 115242 12478 115558 12480
rect 191440 12480 191446 12544
rect 191510 12480 191526 12544
rect 191590 12480 191606 12544
rect 191670 12480 191686 12544
rect 191750 12480 191756 12544
rect 191440 12478 191756 12480
rect 267638 12480 267644 12544
rect 267708 12480 267724 12544
rect 267788 12480 267804 12544
rect 267868 12480 267884 12544
rect 267948 12480 267954 12544
rect 267638 12478 267954 12480
rect 251816 12474 251882 12476
rect 257152 12474 257218 12476
rect 251816 12472 257218 12474
rect 251816 12416 251822 12472
rect 251878 12416 257158 12472
rect 257214 12416 257218 12472
rect 251816 12414 257218 12416
rect 251816 12410 251882 12414
rect 257152 12410 257218 12414
rect 88148 12338 88214 12340
rect 89896 12338 89962 12340
rect 88148 12336 89962 12338
rect 88148 12280 88154 12336
rect 88210 12280 89902 12336
rect 89958 12280 89962 12336
rect 88148 12278 89962 12280
rect 88148 12274 88214 12278
rect 89896 12274 89962 12278
rect 163588 12338 163654 12340
rect 193028 12338 193094 12340
rect 163588 12336 193094 12338
rect 163588 12280 163594 12336
rect 163650 12280 193034 12336
rect 193090 12280 193094 12336
rect 163588 12278 193094 12280
rect 163588 12274 163654 12278
rect 193028 12274 193094 12278
rect 29360 12202 29426 12204
rect 30740 12202 30806 12204
rect 31384 12202 31450 12204
rect 29360 12200 31450 12202
rect 29360 12144 29366 12200
rect 29422 12144 30746 12200
rect 30802 12144 31390 12200
rect 31446 12144 31450 12200
rect 29360 12142 31450 12144
rect 29360 12138 29426 12142
rect 30740 12138 30806 12142
rect 31384 12138 31450 12142
rect 40584 12202 40650 12204
rect 42424 12202 42490 12204
rect 40584 12200 42490 12202
rect 40584 12144 40590 12200
rect 40646 12144 42430 12200
rect 42486 12144 42490 12200
rect 40584 12142 42490 12144
rect 40584 12138 40650 12142
rect 42424 12138 42490 12142
rect 77144 11936 77150 12000
rect 77214 11936 77230 12000
rect 77294 11936 77310 12000
rect 77374 11936 77390 12000
rect 77454 11936 77460 12000
rect 77144 11934 77460 11936
rect 153342 11936 153348 12000
rect 153412 11936 153428 12000
rect 153492 11936 153508 12000
rect 153572 11936 153588 12000
rect 153652 11936 153658 12000
rect 153342 11934 153658 11936
rect 229540 11936 229546 12000
rect 229610 11936 229626 12000
rect 229690 11936 229706 12000
rect 229770 11936 229786 12000
rect 229850 11936 229856 12000
rect 229540 11934 229856 11936
rect 189624 11794 189690 11796
rect 193028 11794 193094 11796
rect 189624 11792 193094 11794
rect 189624 11736 189630 11792
rect 189686 11736 193034 11792
rect 193090 11736 193094 11792
rect 189624 11734 193094 11736
rect 189624 11730 189690 11734
rect 193028 11730 193094 11734
rect 39044 11392 39050 11456
rect 39114 11392 39130 11456
rect 39194 11392 39210 11456
rect 39274 11392 39290 11456
rect 39354 11392 39360 11456
rect 39044 11390 39360 11392
rect 115242 11392 115248 11456
rect 115312 11392 115328 11456
rect 115392 11392 115408 11456
rect 115472 11392 115488 11456
rect 115552 11392 115558 11456
rect 115242 11390 115558 11392
rect 191440 11392 191446 11456
rect 191510 11392 191526 11456
rect 191590 11392 191606 11456
rect 191670 11392 191686 11456
rect 191750 11392 191756 11456
rect 191440 11390 191756 11392
rect 267638 11392 267644 11456
rect 267708 11392 267724 11456
rect 267788 11392 267804 11456
rect 267868 11392 267884 11456
rect 267948 11392 267954 11456
rect 267638 11390 267954 11392
rect 77144 10848 77150 10912
rect 77214 10848 77230 10912
rect 77294 10848 77310 10912
rect 77374 10848 77390 10912
rect 77454 10848 77460 10912
rect 77144 10846 77460 10848
rect 153342 10848 153348 10912
rect 153412 10848 153428 10912
rect 153492 10848 153508 10912
rect 153572 10848 153588 10912
rect 153652 10848 153658 10912
rect 153342 10846 153658 10848
rect 229540 10848 229546 10912
rect 229610 10848 229626 10912
rect 229690 10848 229706 10912
rect 229770 10848 229786 10912
rect 229850 10848 229856 10912
rect 229540 10846 229856 10848
rect 39044 10304 39050 10368
rect 39114 10304 39130 10368
rect 39194 10304 39210 10368
rect 39274 10304 39290 10368
rect 39354 10304 39360 10368
rect 39044 10302 39360 10304
rect 115242 10304 115248 10368
rect 115312 10304 115328 10368
rect 115392 10304 115408 10368
rect 115472 10304 115488 10368
rect 115552 10304 115558 10368
rect 115242 10302 115558 10304
rect 191440 10304 191446 10368
rect 191510 10304 191526 10368
rect 191590 10304 191606 10368
rect 191670 10304 191686 10368
rect 191750 10304 191756 10368
rect 191440 10302 191756 10304
rect 267638 10304 267644 10368
rect 267708 10304 267724 10368
rect 267788 10304 267804 10368
rect 267868 10304 267884 10368
rect 267948 10304 267954 10368
rect 267638 10302 267954 10304
rect 304440 10026 304506 10028
rect 306200 10026 307000 10056
rect 304440 10024 307000 10026
rect 304440 9968 304446 10024
rect 304502 9968 307000 10024
rect 304440 9966 307000 9968
rect 304440 9962 304506 9966
rect 306200 9936 307000 9966
rect 77144 9760 77150 9824
rect 77214 9760 77230 9824
rect 77294 9760 77310 9824
rect 77374 9760 77390 9824
rect 77454 9760 77460 9824
rect 77144 9758 77460 9760
rect 153342 9760 153348 9824
rect 153412 9760 153428 9824
rect 153492 9760 153508 9824
rect 153572 9760 153588 9824
rect 153652 9760 153658 9824
rect 153342 9758 153658 9760
rect 229540 9760 229546 9824
rect 229610 9760 229626 9824
rect 229690 9760 229706 9824
rect 229770 9760 229786 9824
rect 229850 9760 229856 9824
rect 229540 9758 229856 9760
rect 39044 9216 39050 9280
rect 39114 9216 39130 9280
rect 39194 9216 39210 9280
rect 39274 9216 39290 9280
rect 39354 9216 39360 9280
rect 39044 9214 39360 9216
rect 115242 9216 115248 9280
rect 115312 9216 115328 9280
rect 115392 9216 115408 9280
rect 115472 9216 115488 9280
rect 115552 9216 115558 9280
rect 115242 9214 115558 9216
rect 191440 9216 191446 9280
rect 191510 9216 191526 9280
rect 191590 9216 191606 9280
rect 191670 9216 191686 9280
rect 191750 9216 191756 9280
rect 191440 9214 191756 9216
rect 267638 9216 267644 9280
rect 267708 9216 267724 9280
rect 267788 9216 267804 9280
rect 267868 9216 267884 9280
rect 267948 9216 267954 9280
rect 267638 9214 267954 9216
rect 77144 8672 77150 8736
rect 77214 8672 77230 8736
rect 77294 8672 77310 8736
rect 77374 8672 77390 8736
rect 77454 8672 77460 8736
rect 77144 8670 77460 8672
rect 153342 8672 153348 8736
rect 153412 8672 153428 8736
rect 153492 8672 153508 8736
rect 153572 8672 153588 8736
rect 153652 8672 153658 8736
rect 153342 8670 153658 8672
rect 229540 8672 229546 8736
rect 229610 8672 229626 8736
rect 229690 8672 229706 8736
rect 229770 8672 229786 8736
rect 229850 8672 229856 8736
rect 229540 8670 229856 8672
rect 0 8122 800 8152
rect 1388 8122 1462 8134
rect 39044 8128 39050 8192
rect 39114 8128 39130 8192
rect 39194 8128 39210 8192
rect 39274 8128 39290 8192
rect 39354 8128 39360 8192
rect 39044 8126 39360 8128
rect 115242 8128 115248 8192
rect 115312 8128 115328 8192
rect 115392 8128 115408 8192
rect 115472 8128 115488 8192
rect 115552 8128 115558 8192
rect 115242 8126 115558 8128
rect 191440 8128 191446 8192
rect 191510 8128 191526 8192
rect 191590 8128 191606 8192
rect 191670 8128 191686 8192
rect 191750 8128 191756 8192
rect 191440 8126 191756 8128
rect 267638 8128 267644 8192
rect 267708 8128 267724 8192
rect 267788 8128 267804 8192
rect 267868 8128 267884 8192
rect 267948 8128 267954 8192
rect 267638 8126 267954 8128
rect 0 8120 1462 8122
rect 0 8064 1398 8120
rect 1454 8064 1462 8120
rect 0 8062 1462 8064
rect 0 8032 800 8062
rect 1388 8044 1462 8062
rect 77144 7584 77150 7648
rect 77214 7584 77230 7648
rect 77294 7584 77310 7648
rect 77374 7584 77390 7648
rect 77454 7584 77460 7648
rect 77144 7582 77460 7584
rect 153342 7584 153348 7648
rect 153412 7584 153428 7648
rect 153492 7584 153508 7648
rect 153572 7584 153588 7648
rect 153652 7584 153658 7648
rect 153342 7582 153658 7584
rect 229540 7584 229546 7648
rect 229610 7584 229626 7648
rect 229690 7584 229706 7648
rect 229770 7584 229786 7648
rect 229850 7584 229856 7648
rect 229540 7582 229856 7584
rect 39044 7040 39050 7104
rect 39114 7040 39130 7104
rect 39194 7040 39210 7104
rect 39274 7040 39290 7104
rect 39354 7040 39360 7104
rect 39044 7038 39360 7040
rect 115242 7040 115248 7104
rect 115312 7040 115328 7104
rect 115392 7040 115408 7104
rect 115472 7040 115488 7104
rect 115552 7040 115558 7104
rect 115242 7038 115558 7040
rect 191440 7040 191446 7104
rect 191510 7040 191526 7104
rect 191590 7040 191606 7104
rect 191670 7040 191686 7104
rect 191750 7040 191756 7104
rect 191440 7038 191756 7040
rect 267638 7040 267644 7104
rect 267708 7040 267724 7104
rect 267788 7040 267804 7104
rect 267868 7040 267884 7104
rect 267948 7040 267954 7104
rect 267638 7038 267954 7040
rect 77144 6496 77150 6560
rect 77214 6496 77230 6560
rect 77294 6496 77310 6560
rect 77374 6496 77390 6560
rect 77454 6496 77460 6560
rect 77144 6494 77460 6496
rect 153342 6496 153348 6560
rect 153412 6496 153428 6560
rect 153492 6496 153508 6560
rect 153572 6496 153588 6560
rect 153652 6496 153658 6560
rect 153342 6494 153658 6496
rect 229540 6496 229546 6560
rect 229610 6496 229626 6560
rect 229690 6496 229706 6560
rect 229770 6496 229786 6560
rect 229850 6496 229856 6560
rect 229540 6494 229856 6496
rect 39044 5952 39050 6016
rect 39114 5952 39130 6016
rect 39194 5952 39210 6016
rect 39274 5952 39290 6016
rect 39354 5952 39360 6016
rect 39044 5950 39360 5952
rect 115242 5952 115248 6016
rect 115312 5952 115328 6016
rect 115392 5952 115408 6016
rect 115472 5952 115488 6016
rect 115552 5952 115558 6016
rect 115242 5950 115558 5952
rect 191440 5952 191446 6016
rect 191510 5952 191526 6016
rect 191590 5952 191606 6016
rect 191670 5952 191686 6016
rect 191750 5952 191756 6016
rect 191440 5950 191756 5952
rect 267638 5952 267644 6016
rect 267708 5952 267724 6016
rect 267788 5952 267804 6016
rect 267868 5952 267884 6016
rect 267948 5952 267954 6016
rect 267638 5950 267954 5952
rect 303980 5946 304046 5948
rect 306200 5946 307000 5976
rect 303980 5944 307000 5946
rect 303980 5888 303986 5944
rect 304042 5888 307000 5944
rect 303980 5886 307000 5888
rect 303980 5882 304046 5886
rect 306200 5856 307000 5886
rect 77144 5408 77150 5472
rect 77214 5408 77230 5472
rect 77294 5408 77310 5472
rect 77374 5408 77390 5472
rect 77454 5408 77460 5472
rect 77144 5406 77460 5408
rect 153342 5408 153348 5472
rect 153412 5408 153428 5472
rect 153492 5408 153508 5472
rect 153572 5408 153588 5472
rect 153652 5408 153658 5472
rect 153342 5406 153658 5408
rect 229540 5408 229546 5472
rect 229610 5408 229626 5472
rect 229690 5408 229706 5472
rect 229770 5408 229786 5472
rect 229850 5408 229856 5472
rect 229540 5406 229856 5408
rect 39044 4864 39050 4928
rect 39114 4864 39130 4928
rect 39194 4864 39210 4928
rect 39274 4864 39290 4928
rect 39354 4864 39360 4928
rect 39044 4862 39360 4864
rect 115242 4864 115248 4928
rect 115312 4864 115328 4928
rect 115392 4864 115408 4928
rect 115472 4864 115488 4928
rect 115552 4864 115558 4928
rect 115242 4862 115558 4864
rect 191440 4864 191446 4928
rect 191510 4864 191526 4928
rect 191590 4864 191606 4928
rect 191670 4864 191686 4928
rect 191750 4864 191756 4928
rect 191440 4862 191756 4864
rect 267638 4864 267644 4928
rect 267708 4864 267724 4928
rect 267788 4864 267804 4928
rect 267868 4864 267884 4928
rect 267948 4864 267954 4928
rect 267638 4862 267954 4864
rect 77144 4320 77150 4384
rect 77214 4320 77230 4384
rect 77294 4320 77310 4384
rect 77374 4320 77390 4384
rect 77454 4320 77460 4384
rect 77144 4318 77460 4320
rect 153342 4320 153348 4384
rect 153412 4320 153428 4384
rect 153492 4320 153508 4384
rect 153572 4320 153588 4384
rect 153652 4320 153658 4384
rect 153342 4318 153658 4320
rect 229540 4320 229546 4384
rect 229610 4320 229626 4384
rect 229690 4320 229706 4384
rect 229770 4320 229786 4384
rect 229850 4320 229856 4384
rect 229540 4318 229856 4320
rect 39044 3776 39050 3840
rect 39114 3776 39130 3840
rect 39194 3776 39210 3840
rect 39274 3776 39290 3840
rect 39354 3776 39360 3840
rect 39044 3774 39360 3776
rect 115242 3776 115248 3840
rect 115312 3776 115328 3840
rect 115392 3776 115408 3840
rect 115472 3776 115488 3840
rect 115552 3776 115558 3840
rect 115242 3774 115558 3776
rect 191440 3776 191446 3840
rect 191510 3776 191526 3840
rect 191590 3776 191606 3840
rect 191670 3776 191686 3840
rect 191750 3776 191756 3840
rect 191440 3774 191756 3776
rect 267638 3776 267644 3840
rect 267708 3776 267724 3840
rect 267788 3776 267804 3840
rect 267868 3776 267884 3840
rect 267948 3776 267954 3840
rect 267638 3774 267954 3776
rect 77144 3232 77150 3296
rect 77214 3232 77230 3296
rect 77294 3232 77310 3296
rect 77374 3232 77390 3296
rect 77454 3232 77460 3296
rect 77144 3230 77460 3232
rect 153342 3232 153348 3296
rect 153412 3232 153428 3296
rect 153492 3232 153508 3296
rect 153572 3232 153588 3296
rect 153652 3232 153658 3296
rect 153342 3230 153658 3232
rect 229540 3232 229546 3296
rect 229610 3232 229626 3296
rect 229690 3232 229706 3296
rect 229770 3232 229786 3296
rect 229850 3232 229856 3296
rect 229540 3230 229856 3232
rect 39044 2688 39050 2752
rect 39114 2688 39130 2752
rect 39194 2688 39210 2752
rect 39274 2688 39290 2752
rect 39354 2688 39360 2752
rect 39044 2686 39360 2688
rect 115242 2688 115248 2752
rect 115312 2688 115328 2752
rect 115392 2688 115408 2752
rect 115472 2688 115488 2752
rect 115552 2688 115558 2752
rect 115242 2686 115558 2688
rect 191440 2688 191446 2752
rect 191510 2688 191526 2752
rect 191590 2688 191606 2752
rect 191670 2688 191686 2752
rect 191750 2688 191756 2752
rect 191440 2686 191756 2688
rect 267638 2688 267644 2752
rect 267708 2688 267724 2752
rect 267788 2688 267804 2752
rect 267868 2688 267884 2752
rect 267948 2688 267954 2752
rect 267638 2686 267954 2688
rect 77144 2144 77150 2208
rect 77214 2144 77230 2208
rect 77294 2144 77310 2208
rect 77374 2144 77390 2208
rect 77454 2144 77460 2208
rect 77144 2142 77460 2144
rect 153342 2144 153348 2208
rect 153412 2144 153428 2208
rect 153492 2144 153508 2208
rect 153572 2144 153588 2208
rect 153652 2144 153658 2208
rect 153342 2142 153658 2144
rect 229540 2144 229546 2208
rect 229610 2144 229626 2208
rect 229690 2144 229706 2208
rect 229770 2144 229786 2208
rect 229850 2144 229856 2208
rect 229540 2142 229856 2144
rect 302232 2002 302298 2004
rect 306200 2002 307000 2032
rect 302232 2000 307000 2002
rect 302232 1944 302238 2000
rect 302294 1944 307000 2000
rect 302232 1942 307000 1944
rect 302232 1938 302298 1942
rect 306200 1912 307000 1942
<< via3 >>
rect 39050 13628 39114 13632
rect 39050 13572 39054 13628
rect 39054 13572 39110 13628
rect 39110 13572 39114 13628
rect 39050 13568 39114 13572
rect 39130 13628 39194 13632
rect 39130 13572 39134 13628
rect 39134 13572 39190 13628
rect 39190 13572 39194 13628
rect 39130 13568 39194 13572
rect 39210 13628 39274 13632
rect 39210 13572 39214 13628
rect 39214 13572 39270 13628
rect 39270 13572 39274 13628
rect 39210 13568 39274 13572
rect 39290 13628 39354 13632
rect 39290 13572 39294 13628
rect 39294 13572 39350 13628
rect 39350 13572 39354 13628
rect 39290 13568 39354 13572
rect 115248 13628 115312 13632
rect 115248 13572 115252 13628
rect 115252 13572 115308 13628
rect 115308 13572 115312 13628
rect 115248 13568 115312 13572
rect 115328 13628 115392 13632
rect 115328 13572 115332 13628
rect 115332 13572 115388 13628
rect 115388 13572 115392 13628
rect 115328 13568 115392 13572
rect 115408 13628 115472 13632
rect 115408 13572 115412 13628
rect 115412 13572 115468 13628
rect 115468 13572 115472 13628
rect 115408 13568 115472 13572
rect 115488 13628 115552 13632
rect 115488 13572 115492 13628
rect 115492 13572 115548 13628
rect 115548 13572 115552 13628
rect 115488 13568 115552 13572
rect 191446 13628 191510 13632
rect 191446 13572 191450 13628
rect 191450 13572 191506 13628
rect 191506 13572 191510 13628
rect 191446 13568 191510 13572
rect 191526 13628 191590 13632
rect 191526 13572 191530 13628
rect 191530 13572 191586 13628
rect 191586 13572 191590 13628
rect 191526 13568 191590 13572
rect 191606 13628 191670 13632
rect 191606 13572 191610 13628
rect 191610 13572 191666 13628
rect 191666 13572 191670 13628
rect 191606 13568 191670 13572
rect 191686 13628 191750 13632
rect 191686 13572 191690 13628
rect 191690 13572 191746 13628
rect 191746 13572 191750 13628
rect 191686 13568 191750 13572
rect 267644 13628 267708 13632
rect 267644 13572 267648 13628
rect 267648 13572 267704 13628
rect 267704 13572 267708 13628
rect 267644 13568 267708 13572
rect 267724 13628 267788 13632
rect 267724 13572 267728 13628
rect 267728 13572 267784 13628
rect 267784 13572 267788 13628
rect 267724 13568 267788 13572
rect 267804 13628 267868 13632
rect 267804 13572 267808 13628
rect 267808 13572 267864 13628
rect 267864 13572 267868 13628
rect 267804 13568 267868 13572
rect 267884 13628 267948 13632
rect 267884 13572 267888 13628
rect 267888 13572 267944 13628
rect 267944 13572 267948 13628
rect 267884 13568 267948 13572
rect 77150 13084 77214 13088
rect 77150 13028 77154 13084
rect 77154 13028 77210 13084
rect 77210 13028 77214 13084
rect 77150 13024 77214 13028
rect 77230 13084 77294 13088
rect 77230 13028 77234 13084
rect 77234 13028 77290 13084
rect 77290 13028 77294 13084
rect 77230 13024 77294 13028
rect 77310 13084 77374 13088
rect 77310 13028 77314 13084
rect 77314 13028 77370 13084
rect 77370 13028 77374 13084
rect 77310 13024 77374 13028
rect 77390 13084 77454 13088
rect 77390 13028 77394 13084
rect 77394 13028 77450 13084
rect 77450 13028 77454 13084
rect 77390 13024 77454 13028
rect 153348 13084 153412 13088
rect 153348 13028 153352 13084
rect 153352 13028 153408 13084
rect 153408 13028 153412 13084
rect 153348 13024 153412 13028
rect 153428 13084 153492 13088
rect 153428 13028 153432 13084
rect 153432 13028 153488 13084
rect 153488 13028 153492 13084
rect 153428 13024 153492 13028
rect 153508 13084 153572 13088
rect 153508 13028 153512 13084
rect 153512 13028 153568 13084
rect 153568 13028 153572 13084
rect 153508 13024 153572 13028
rect 153588 13084 153652 13088
rect 153588 13028 153592 13084
rect 153592 13028 153648 13084
rect 153648 13028 153652 13084
rect 153588 13024 153652 13028
rect 229546 13084 229610 13088
rect 229546 13028 229550 13084
rect 229550 13028 229606 13084
rect 229606 13028 229610 13084
rect 229546 13024 229610 13028
rect 229626 13084 229690 13088
rect 229626 13028 229630 13084
rect 229630 13028 229686 13084
rect 229686 13028 229690 13084
rect 229626 13024 229690 13028
rect 229706 13084 229770 13088
rect 229706 13028 229710 13084
rect 229710 13028 229766 13084
rect 229766 13028 229770 13084
rect 229706 13024 229770 13028
rect 229786 13084 229850 13088
rect 229786 13028 229790 13084
rect 229790 13028 229846 13084
rect 229846 13028 229850 13084
rect 229786 13024 229850 13028
rect 39050 12540 39114 12544
rect 39050 12484 39054 12540
rect 39054 12484 39110 12540
rect 39110 12484 39114 12540
rect 39050 12480 39114 12484
rect 39130 12540 39194 12544
rect 39130 12484 39134 12540
rect 39134 12484 39190 12540
rect 39190 12484 39194 12540
rect 39130 12480 39194 12484
rect 39210 12540 39274 12544
rect 39210 12484 39214 12540
rect 39214 12484 39270 12540
rect 39270 12484 39274 12540
rect 39210 12480 39274 12484
rect 39290 12540 39354 12544
rect 39290 12484 39294 12540
rect 39294 12484 39350 12540
rect 39350 12484 39354 12540
rect 39290 12480 39354 12484
rect 115248 12540 115312 12544
rect 115248 12484 115252 12540
rect 115252 12484 115308 12540
rect 115308 12484 115312 12540
rect 115248 12480 115312 12484
rect 115328 12540 115392 12544
rect 115328 12484 115332 12540
rect 115332 12484 115388 12540
rect 115388 12484 115392 12540
rect 115328 12480 115392 12484
rect 115408 12540 115472 12544
rect 115408 12484 115412 12540
rect 115412 12484 115468 12540
rect 115468 12484 115472 12540
rect 115408 12480 115472 12484
rect 115488 12540 115552 12544
rect 115488 12484 115492 12540
rect 115492 12484 115548 12540
rect 115548 12484 115552 12540
rect 115488 12480 115552 12484
rect 191446 12540 191510 12544
rect 191446 12484 191450 12540
rect 191450 12484 191506 12540
rect 191506 12484 191510 12540
rect 191446 12480 191510 12484
rect 191526 12540 191590 12544
rect 191526 12484 191530 12540
rect 191530 12484 191586 12540
rect 191586 12484 191590 12540
rect 191526 12480 191590 12484
rect 191606 12540 191670 12544
rect 191606 12484 191610 12540
rect 191610 12484 191666 12540
rect 191666 12484 191670 12540
rect 191606 12480 191670 12484
rect 191686 12540 191750 12544
rect 191686 12484 191690 12540
rect 191690 12484 191746 12540
rect 191746 12484 191750 12540
rect 191686 12480 191750 12484
rect 267644 12540 267708 12544
rect 267644 12484 267648 12540
rect 267648 12484 267704 12540
rect 267704 12484 267708 12540
rect 267644 12480 267708 12484
rect 267724 12540 267788 12544
rect 267724 12484 267728 12540
rect 267728 12484 267784 12540
rect 267784 12484 267788 12540
rect 267724 12480 267788 12484
rect 267804 12540 267868 12544
rect 267804 12484 267808 12540
rect 267808 12484 267864 12540
rect 267864 12484 267868 12540
rect 267804 12480 267868 12484
rect 267884 12540 267948 12544
rect 267884 12484 267888 12540
rect 267888 12484 267944 12540
rect 267944 12484 267948 12540
rect 267884 12480 267948 12484
rect 77150 11996 77214 12000
rect 77150 11940 77154 11996
rect 77154 11940 77210 11996
rect 77210 11940 77214 11996
rect 77150 11936 77214 11940
rect 77230 11996 77294 12000
rect 77230 11940 77234 11996
rect 77234 11940 77290 11996
rect 77290 11940 77294 11996
rect 77230 11936 77294 11940
rect 77310 11996 77374 12000
rect 77310 11940 77314 11996
rect 77314 11940 77370 11996
rect 77370 11940 77374 11996
rect 77310 11936 77374 11940
rect 77390 11996 77454 12000
rect 77390 11940 77394 11996
rect 77394 11940 77450 11996
rect 77450 11940 77454 11996
rect 77390 11936 77454 11940
rect 153348 11996 153412 12000
rect 153348 11940 153352 11996
rect 153352 11940 153408 11996
rect 153408 11940 153412 11996
rect 153348 11936 153412 11940
rect 153428 11996 153492 12000
rect 153428 11940 153432 11996
rect 153432 11940 153488 11996
rect 153488 11940 153492 11996
rect 153428 11936 153492 11940
rect 153508 11996 153572 12000
rect 153508 11940 153512 11996
rect 153512 11940 153568 11996
rect 153568 11940 153572 11996
rect 153508 11936 153572 11940
rect 153588 11996 153652 12000
rect 153588 11940 153592 11996
rect 153592 11940 153648 11996
rect 153648 11940 153652 11996
rect 153588 11936 153652 11940
rect 229546 11996 229610 12000
rect 229546 11940 229550 11996
rect 229550 11940 229606 11996
rect 229606 11940 229610 11996
rect 229546 11936 229610 11940
rect 229626 11996 229690 12000
rect 229626 11940 229630 11996
rect 229630 11940 229686 11996
rect 229686 11940 229690 11996
rect 229626 11936 229690 11940
rect 229706 11996 229770 12000
rect 229706 11940 229710 11996
rect 229710 11940 229766 11996
rect 229766 11940 229770 11996
rect 229706 11936 229770 11940
rect 229786 11996 229850 12000
rect 229786 11940 229790 11996
rect 229790 11940 229846 11996
rect 229846 11940 229850 11996
rect 229786 11936 229850 11940
rect 39050 11452 39114 11456
rect 39050 11396 39054 11452
rect 39054 11396 39110 11452
rect 39110 11396 39114 11452
rect 39050 11392 39114 11396
rect 39130 11452 39194 11456
rect 39130 11396 39134 11452
rect 39134 11396 39190 11452
rect 39190 11396 39194 11452
rect 39130 11392 39194 11396
rect 39210 11452 39274 11456
rect 39210 11396 39214 11452
rect 39214 11396 39270 11452
rect 39270 11396 39274 11452
rect 39210 11392 39274 11396
rect 39290 11452 39354 11456
rect 39290 11396 39294 11452
rect 39294 11396 39350 11452
rect 39350 11396 39354 11452
rect 39290 11392 39354 11396
rect 115248 11452 115312 11456
rect 115248 11396 115252 11452
rect 115252 11396 115308 11452
rect 115308 11396 115312 11452
rect 115248 11392 115312 11396
rect 115328 11452 115392 11456
rect 115328 11396 115332 11452
rect 115332 11396 115388 11452
rect 115388 11396 115392 11452
rect 115328 11392 115392 11396
rect 115408 11452 115472 11456
rect 115408 11396 115412 11452
rect 115412 11396 115468 11452
rect 115468 11396 115472 11452
rect 115408 11392 115472 11396
rect 115488 11452 115552 11456
rect 115488 11396 115492 11452
rect 115492 11396 115548 11452
rect 115548 11396 115552 11452
rect 115488 11392 115552 11396
rect 191446 11452 191510 11456
rect 191446 11396 191450 11452
rect 191450 11396 191506 11452
rect 191506 11396 191510 11452
rect 191446 11392 191510 11396
rect 191526 11452 191590 11456
rect 191526 11396 191530 11452
rect 191530 11396 191586 11452
rect 191586 11396 191590 11452
rect 191526 11392 191590 11396
rect 191606 11452 191670 11456
rect 191606 11396 191610 11452
rect 191610 11396 191666 11452
rect 191666 11396 191670 11452
rect 191606 11392 191670 11396
rect 191686 11452 191750 11456
rect 191686 11396 191690 11452
rect 191690 11396 191746 11452
rect 191746 11396 191750 11452
rect 191686 11392 191750 11396
rect 267644 11452 267708 11456
rect 267644 11396 267648 11452
rect 267648 11396 267704 11452
rect 267704 11396 267708 11452
rect 267644 11392 267708 11396
rect 267724 11452 267788 11456
rect 267724 11396 267728 11452
rect 267728 11396 267784 11452
rect 267784 11396 267788 11452
rect 267724 11392 267788 11396
rect 267804 11452 267868 11456
rect 267804 11396 267808 11452
rect 267808 11396 267864 11452
rect 267864 11396 267868 11452
rect 267804 11392 267868 11396
rect 267884 11452 267948 11456
rect 267884 11396 267888 11452
rect 267888 11396 267944 11452
rect 267944 11396 267948 11452
rect 267884 11392 267948 11396
rect 77150 10908 77214 10912
rect 77150 10852 77154 10908
rect 77154 10852 77210 10908
rect 77210 10852 77214 10908
rect 77150 10848 77214 10852
rect 77230 10908 77294 10912
rect 77230 10852 77234 10908
rect 77234 10852 77290 10908
rect 77290 10852 77294 10908
rect 77230 10848 77294 10852
rect 77310 10908 77374 10912
rect 77310 10852 77314 10908
rect 77314 10852 77370 10908
rect 77370 10852 77374 10908
rect 77310 10848 77374 10852
rect 77390 10908 77454 10912
rect 77390 10852 77394 10908
rect 77394 10852 77450 10908
rect 77450 10852 77454 10908
rect 77390 10848 77454 10852
rect 153348 10908 153412 10912
rect 153348 10852 153352 10908
rect 153352 10852 153408 10908
rect 153408 10852 153412 10908
rect 153348 10848 153412 10852
rect 153428 10908 153492 10912
rect 153428 10852 153432 10908
rect 153432 10852 153488 10908
rect 153488 10852 153492 10908
rect 153428 10848 153492 10852
rect 153508 10908 153572 10912
rect 153508 10852 153512 10908
rect 153512 10852 153568 10908
rect 153568 10852 153572 10908
rect 153508 10848 153572 10852
rect 153588 10908 153652 10912
rect 153588 10852 153592 10908
rect 153592 10852 153648 10908
rect 153648 10852 153652 10908
rect 153588 10848 153652 10852
rect 229546 10908 229610 10912
rect 229546 10852 229550 10908
rect 229550 10852 229606 10908
rect 229606 10852 229610 10908
rect 229546 10848 229610 10852
rect 229626 10908 229690 10912
rect 229626 10852 229630 10908
rect 229630 10852 229686 10908
rect 229686 10852 229690 10908
rect 229626 10848 229690 10852
rect 229706 10908 229770 10912
rect 229706 10852 229710 10908
rect 229710 10852 229766 10908
rect 229766 10852 229770 10908
rect 229706 10848 229770 10852
rect 229786 10908 229850 10912
rect 229786 10852 229790 10908
rect 229790 10852 229846 10908
rect 229846 10852 229850 10908
rect 229786 10848 229850 10852
rect 39050 10364 39114 10368
rect 39050 10308 39054 10364
rect 39054 10308 39110 10364
rect 39110 10308 39114 10364
rect 39050 10304 39114 10308
rect 39130 10364 39194 10368
rect 39130 10308 39134 10364
rect 39134 10308 39190 10364
rect 39190 10308 39194 10364
rect 39130 10304 39194 10308
rect 39210 10364 39274 10368
rect 39210 10308 39214 10364
rect 39214 10308 39270 10364
rect 39270 10308 39274 10364
rect 39210 10304 39274 10308
rect 39290 10364 39354 10368
rect 39290 10308 39294 10364
rect 39294 10308 39350 10364
rect 39350 10308 39354 10364
rect 39290 10304 39354 10308
rect 115248 10364 115312 10368
rect 115248 10308 115252 10364
rect 115252 10308 115308 10364
rect 115308 10308 115312 10364
rect 115248 10304 115312 10308
rect 115328 10364 115392 10368
rect 115328 10308 115332 10364
rect 115332 10308 115388 10364
rect 115388 10308 115392 10364
rect 115328 10304 115392 10308
rect 115408 10364 115472 10368
rect 115408 10308 115412 10364
rect 115412 10308 115468 10364
rect 115468 10308 115472 10364
rect 115408 10304 115472 10308
rect 115488 10364 115552 10368
rect 115488 10308 115492 10364
rect 115492 10308 115548 10364
rect 115548 10308 115552 10364
rect 115488 10304 115552 10308
rect 191446 10364 191510 10368
rect 191446 10308 191450 10364
rect 191450 10308 191506 10364
rect 191506 10308 191510 10364
rect 191446 10304 191510 10308
rect 191526 10364 191590 10368
rect 191526 10308 191530 10364
rect 191530 10308 191586 10364
rect 191586 10308 191590 10364
rect 191526 10304 191590 10308
rect 191606 10364 191670 10368
rect 191606 10308 191610 10364
rect 191610 10308 191666 10364
rect 191666 10308 191670 10364
rect 191606 10304 191670 10308
rect 191686 10364 191750 10368
rect 191686 10308 191690 10364
rect 191690 10308 191746 10364
rect 191746 10308 191750 10364
rect 191686 10304 191750 10308
rect 267644 10364 267708 10368
rect 267644 10308 267648 10364
rect 267648 10308 267704 10364
rect 267704 10308 267708 10364
rect 267644 10304 267708 10308
rect 267724 10364 267788 10368
rect 267724 10308 267728 10364
rect 267728 10308 267784 10364
rect 267784 10308 267788 10364
rect 267724 10304 267788 10308
rect 267804 10364 267868 10368
rect 267804 10308 267808 10364
rect 267808 10308 267864 10364
rect 267864 10308 267868 10364
rect 267804 10304 267868 10308
rect 267884 10364 267948 10368
rect 267884 10308 267888 10364
rect 267888 10308 267944 10364
rect 267944 10308 267948 10364
rect 267884 10304 267948 10308
rect 77150 9820 77214 9824
rect 77150 9764 77154 9820
rect 77154 9764 77210 9820
rect 77210 9764 77214 9820
rect 77150 9760 77214 9764
rect 77230 9820 77294 9824
rect 77230 9764 77234 9820
rect 77234 9764 77290 9820
rect 77290 9764 77294 9820
rect 77230 9760 77294 9764
rect 77310 9820 77374 9824
rect 77310 9764 77314 9820
rect 77314 9764 77370 9820
rect 77370 9764 77374 9820
rect 77310 9760 77374 9764
rect 77390 9820 77454 9824
rect 77390 9764 77394 9820
rect 77394 9764 77450 9820
rect 77450 9764 77454 9820
rect 77390 9760 77454 9764
rect 153348 9820 153412 9824
rect 153348 9764 153352 9820
rect 153352 9764 153408 9820
rect 153408 9764 153412 9820
rect 153348 9760 153412 9764
rect 153428 9820 153492 9824
rect 153428 9764 153432 9820
rect 153432 9764 153488 9820
rect 153488 9764 153492 9820
rect 153428 9760 153492 9764
rect 153508 9820 153572 9824
rect 153508 9764 153512 9820
rect 153512 9764 153568 9820
rect 153568 9764 153572 9820
rect 153508 9760 153572 9764
rect 153588 9820 153652 9824
rect 153588 9764 153592 9820
rect 153592 9764 153648 9820
rect 153648 9764 153652 9820
rect 153588 9760 153652 9764
rect 229546 9820 229610 9824
rect 229546 9764 229550 9820
rect 229550 9764 229606 9820
rect 229606 9764 229610 9820
rect 229546 9760 229610 9764
rect 229626 9820 229690 9824
rect 229626 9764 229630 9820
rect 229630 9764 229686 9820
rect 229686 9764 229690 9820
rect 229626 9760 229690 9764
rect 229706 9820 229770 9824
rect 229706 9764 229710 9820
rect 229710 9764 229766 9820
rect 229766 9764 229770 9820
rect 229706 9760 229770 9764
rect 229786 9820 229850 9824
rect 229786 9764 229790 9820
rect 229790 9764 229846 9820
rect 229846 9764 229850 9820
rect 229786 9760 229850 9764
rect 39050 9276 39114 9280
rect 39050 9220 39054 9276
rect 39054 9220 39110 9276
rect 39110 9220 39114 9276
rect 39050 9216 39114 9220
rect 39130 9276 39194 9280
rect 39130 9220 39134 9276
rect 39134 9220 39190 9276
rect 39190 9220 39194 9276
rect 39130 9216 39194 9220
rect 39210 9276 39274 9280
rect 39210 9220 39214 9276
rect 39214 9220 39270 9276
rect 39270 9220 39274 9276
rect 39210 9216 39274 9220
rect 39290 9276 39354 9280
rect 39290 9220 39294 9276
rect 39294 9220 39350 9276
rect 39350 9220 39354 9276
rect 39290 9216 39354 9220
rect 115248 9276 115312 9280
rect 115248 9220 115252 9276
rect 115252 9220 115308 9276
rect 115308 9220 115312 9276
rect 115248 9216 115312 9220
rect 115328 9276 115392 9280
rect 115328 9220 115332 9276
rect 115332 9220 115388 9276
rect 115388 9220 115392 9276
rect 115328 9216 115392 9220
rect 115408 9276 115472 9280
rect 115408 9220 115412 9276
rect 115412 9220 115468 9276
rect 115468 9220 115472 9276
rect 115408 9216 115472 9220
rect 115488 9276 115552 9280
rect 115488 9220 115492 9276
rect 115492 9220 115548 9276
rect 115548 9220 115552 9276
rect 115488 9216 115552 9220
rect 191446 9276 191510 9280
rect 191446 9220 191450 9276
rect 191450 9220 191506 9276
rect 191506 9220 191510 9276
rect 191446 9216 191510 9220
rect 191526 9276 191590 9280
rect 191526 9220 191530 9276
rect 191530 9220 191586 9276
rect 191586 9220 191590 9276
rect 191526 9216 191590 9220
rect 191606 9276 191670 9280
rect 191606 9220 191610 9276
rect 191610 9220 191666 9276
rect 191666 9220 191670 9276
rect 191606 9216 191670 9220
rect 191686 9276 191750 9280
rect 191686 9220 191690 9276
rect 191690 9220 191746 9276
rect 191746 9220 191750 9276
rect 191686 9216 191750 9220
rect 267644 9276 267708 9280
rect 267644 9220 267648 9276
rect 267648 9220 267704 9276
rect 267704 9220 267708 9276
rect 267644 9216 267708 9220
rect 267724 9276 267788 9280
rect 267724 9220 267728 9276
rect 267728 9220 267784 9276
rect 267784 9220 267788 9276
rect 267724 9216 267788 9220
rect 267804 9276 267868 9280
rect 267804 9220 267808 9276
rect 267808 9220 267864 9276
rect 267864 9220 267868 9276
rect 267804 9216 267868 9220
rect 267884 9276 267948 9280
rect 267884 9220 267888 9276
rect 267888 9220 267944 9276
rect 267944 9220 267948 9276
rect 267884 9216 267948 9220
rect 77150 8732 77214 8736
rect 77150 8676 77154 8732
rect 77154 8676 77210 8732
rect 77210 8676 77214 8732
rect 77150 8672 77214 8676
rect 77230 8732 77294 8736
rect 77230 8676 77234 8732
rect 77234 8676 77290 8732
rect 77290 8676 77294 8732
rect 77230 8672 77294 8676
rect 77310 8732 77374 8736
rect 77310 8676 77314 8732
rect 77314 8676 77370 8732
rect 77370 8676 77374 8732
rect 77310 8672 77374 8676
rect 77390 8732 77454 8736
rect 77390 8676 77394 8732
rect 77394 8676 77450 8732
rect 77450 8676 77454 8732
rect 77390 8672 77454 8676
rect 153348 8732 153412 8736
rect 153348 8676 153352 8732
rect 153352 8676 153408 8732
rect 153408 8676 153412 8732
rect 153348 8672 153412 8676
rect 153428 8732 153492 8736
rect 153428 8676 153432 8732
rect 153432 8676 153488 8732
rect 153488 8676 153492 8732
rect 153428 8672 153492 8676
rect 153508 8732 153572 8736
rect 153508 8676 153512 8732
rect 153512 8676 153568 8732
rect 153568 8676 153572 8732
rect 153508 8672 153572 8676
rect 153588 8732 153652 8736
rect 153588 8676 153592 8732
rect 153592 8676 153648 8732
rect 153648 8676 153652 8732
rect 153588 8672 153652 8676
rect 229546 8732 229610 8736
rect 229546 8676 229550 8732
rect 229550 8676 229606 8732
rect 229606 8676 229610 8732
rect 229546 8672 229610 8676
rect 229626 8732 229690 8736
rect 229626 8676 229630 8732
rect 229630 8676 229686 8732
rect 229686 8676 229690 8732
rect 229626 8672 229690 8676
rect 229706 8732 229770 8736
rect 229706 8676 229710 8732
rect 229710 8676 229766 8732
rect 229766 8676 229770 8732
rect 229706 8672 229770 8676
rect 229786 8732 229850 8736
rect 229786 8676 229790 8732
rect 229790 8676 229846 8732
rect 229846 8676 229850 8732
rect 229786 8672 229850 8676
rect 39050 8188 39114 8192
rect 39050 8132 39054 8188
rect 39054 8132 39110 8188
rect 39110 8132 39114 8188
rect 39050 8128 39114 8132
rect 39130 8188 39194 8192
rect 39130 8132 39134 8188
rect 39134 8132 39190 8188
rect 39190 8132 39194 8188
rect 39130 8128 39194 8132
rect 39210 8188 39274 8192
rect 39210 8132 39214 8188
rect 39214 8132 39270 8188
rect 39270 8132 39274 8188
rect 39210 8128 39274 8132
rect 39290 8188 39354 8192
rect 39290 8132 39294 8188
rect 39294 8132 39350 8188
rect 39350 8132 39354 8188
rect 39290 8128 39354 8132
rect 115248 8188 115312 8192
rect 115248 8132 115252 8188
rect 115252 8132 115308 8188
rect 115308 8132 115312 8188
rect 115248 8128 115312 8132
rect 115328 8188 115392 8192
rect 115328 8132 115332 8188
rect 115332 8132 115388 8188
rect 115388 8132 115392 8188
rect 115328 8128 115392 8132
rect 115408 8188 115472 8192
rect 115408 8132 115412 8188
rect 115412 8132 115468 8188
rect 115468 8132 115472 8188
rect 115408 8128 115472 8132
rect 115488 8188 115552 8192
rect 115488 8132 115492 8188
rect 115492 8132 115548 8188
rect 115548 8132 115552 8188
rect 115488 8128 115552 8132
rect 191446 8188 191510 8192
rect 191446 8132 191450 8188
rect 191450 8132 191506 8188
rect 191506 8132 191510 8188
rect 191446 8128 191510 8132
rect 191526 8188 191590 8192
rect 191526 8132 191530 8188
rect 191530 8132 191586 8188
rect 191586 8132 191590 8188
rect 191526 8128 191590 8132
rect 191606 8188 191670 8192
rect 191606 8132 191610 8188
rect 191610 8132 191666 8188
rect 191666 8132 191670 8188
rect 191606 8128 191670 8132
rect 191686 8188 191750 8192
rect 191686 8132 191690 8188
rect 191690 8132 191746 8188
rect 191746 8132 191750 8188
rect 191686 8128 191750 8132
rect 267644 8188 267708 8192
rect 267644 8132 267648 8188
rect 267648 8132 267704 8188
rect 267704 8132 267708 8188
rect 267644 8128 267708 8132
rect 267724 8188 267788 8192
rect 267724 8132 267728 8188
rect 267728 8132 267784 8188
rect 267784 8132 267788 8188
rect 267724 8128 267788 8132
rect 267804 8188 267868 8192
rect 267804 8132 267808 8188
rect 267808 8132 267864 8188
rect 267864 8132 267868 8188
rect 267804 8128 267868 8132
rect 267884 8188 267948 8192
rect 267884 8132 267888 8188
rect 267888 8132 267944 8188
rect 267944 8132 267948 8188
rect 267884 8128 267948 8132
rect 77150 7644 77214 7648
rect 77150 7588 77154 7644
rect 77154 7588 77210 7644
rect 77210 7588 77214 7644
rect 77150 7584 77214 7588
rect 77230 7644 77294 7648
rect 77230 7588 77234 7644
rect 77234 7588 77290 7644
rect 77290 7588 77294 7644
rect 77230 7584 77294 7588
rect 77310 7644 77374 7648
rect 77310 7588 77314 7644
rect 77314 7588 77370 7644
rect 77370 7588 77374 7644
rect 77310 7584 77374 7588
rect 77390 7644 77454 7648
rect 77390 7588 77394 7644
rect 77394 7588 77450 7644
rect 77450 7588 77454 7644
rect 77390 7584 77454 7588
rect 153348 7644 153412 7648
rect 153348 7588 153352 7644
rect 153352 7588 153408 7644
rect 153408 7588 153412 7644
rect 153348 7584 153412 7588
rect 153428 7644 153492 7648
rect 153428 7588 153432 7644
rect 153432 7588 153488 7644
rect 153488 7588 153492 7644
rect 153428 7584 153492 7588
rect 153508 7644 153572 7648
rect 153508 7588 153512 7644
rect 153512 7588 153568 7644
rect 153568 7588 153572 7644
rect 153508 7584 153572 7588
rect 153588 7644 153652 7648
rect 153588 7588 153592 7644
rect 153592 7588 153648 7644
rect 153648 7588 153652 7644
rect 153588 7584 153652 7588
rect 229546 7644 229610 7648
rect 229546 7588 229550 7644
rect 229550 7588 229606 7644
rect 229606 7588 229610 7644
rect 229546 7584 229610 7588
rect 229626 7644 229690 7648
rect 229626 7588 229630 7644
rect 229630 7588 229686 7644
rect 229686 7588 229690 7644
rect 229626 7584 229690 7588
rect 229706 7644 229770 7648
rect 229706 7588 229710 7644
rect 229710 7588 229766 7644
rect 229766 7588 229770 7644
rect 229706 7584 229770 7588
rect 229786 7644 229850 7648
rect 229786 7588 229790 7644
rect 229790 7588 229846 7644
rect 229846 7588 229850 7644
rect 229786 7584 229850 7588
rect 39050 7100 39114 7104
rect 39050 7044 39054 7100
rect 39054 7044 39110 7100
rect 39110 7044 39114 7100
rect 39050 7040 39114 7044
rect 39130 7100 39194 7104
rect 39130 7044 39134 7100
rect 39134 7044 39190 7100
rect 39190 7044 39194 7100
rect 39130 7040 39194 7044
rect 39210 7100 39274 7104
rect 39210 7044 39214 7100
rect 39214 7044 39270 7100
rect 39270 7044 39274 7100
rect 39210 7040 39274 7044
rect 39290 7100 39354 7104
rect 39290 7044 39294 7100
rect 39294 7044 39350 7100
rect 39350 7044 39354 7100
rect 39290 7040 39354 7044
rect 115248 7100 115312 7104
rect 115248 7044 115252 7100
rect 115252 7044 115308 7100
rect 115308 7044 115312 7100
rect 115248 7040 115312 7044
rect 115328 7100 115392 7104
rect 115328 7044 115332 7100
rect 115332 7044 115388 7100
rect 115388 7044 115392 7100
rect 115328 7040 115392 7044
rect 115408 7100 115472 7104
rect 115408 7044 115412 7100
rect 115412 7044 115468 7100
rect 115468 7044 115472 7100
rect 115408 7040 115472 7044
rect 115488 7100 115552 7104
rect 115488 7044 115492 7100
rect 115492 7044 115548 7100
rect 115548 7044 115552 7100
rect 115488 7040 115552 7044
rect 191446 7100 191510 7104
rect 191446 7044 191450 7100
rect 191450 7044 191506 7100
rect 191506 7044 191510 7100
rect 191446 7040 191510 7044
rect 191526 7100 191590 7104
rect 191526 7044 191530 7100
rect 191530 7044 191586 7100
rect 191586 7044 191590 7100
rect 191526 7040 191590 7044
rect 191606 7100 191670 7104
rect 191606 7044 191610 7100
rect 191610 7044 191666 7100
rect 191666 7044 191670 7100
rect 191606 7040 191670 7044
rect 191686 7100 191750 7104
rect 191686 7044 191690 7100
rect 191690 7044 191746 7100
rect 191746 7044 191750 7100
rect 191686 7040 191750 7044
rect 267644 7100 267708 7104
rect 267644 7044 267648 7100
rect 267648 7044 267704 7100
rect 267704 7044 267708 7100
rect 267644 7040 267708 7044
rect 267724 7100 267788 7104
rect 267724 7044 267728 7100
rect 267728 7044 267784 7100
rect 267784 7044 267788 7100
rect 267724 7040 267788 7044
rect 267804 7100 267868 7104
rect 267804 7044 267808 7100
rect 267808 7044 267864 7100
rect 267864 7044 267868 7100
rect 267804 7040 267868 7044
rect 267884 7100 267948 7104
rect 267884 7044 267888 7100
rect 267888 7044 267944 7100
rect 267944 7044 267948 7100
rect 267884 7040 267948 7044
rect 77150 6556 77214 6560
rect 77150 6500 77154 6556
rect 77154 6500 77210 6556
rect 77210 6500 77214 6556
rect 77150 6496 77214 6500
rect 77230 6556 77294 6560
rect 77230 6500 77234 6556
rect 77234 6500 77290 6556
rect 77290 6500 77294 6556
rect 77230 6496 77294 6500
rect 77310 6556 77374 6560
rect 77310 6500 77314 6556
rect 77314 6500 77370 6556
rect 77370 6500 77374 6556
rect 77310 6496 77374 6500
rect 77390 6556 77454 6560
rect 77390 6500 77394 6556
rect 77394 6500 77450 6556
rect 77450 6500 77454 6556
rect 77390 6496 77454 6500
rect 153348 6556 153412 6560
rect 153348 6500 153352 6556
rect 153352 6500 153408 6556
rect 153408 6500 153412 6556
rect 153348 6496 153412 6500
rect 153428 6556 153492 6560
rect 153428 6500 153432 6556
rect 153432 6500 153488 6556
rect 153488 6500 153492 6556
rect 153428 6496 153492 6500
rect 153508 6556 153572 6560
rect 153508 6500 153512 6556
rect 153512 6500 153568 6556
rect 153568 6500 153572 6556
rect 153508 6496 153572 6500
rect 153588 6556 153652 6560
rect 153588 6500 153592 6556
rect 153592 6500 153648 6556
rect 153648 6500 153652 6556
rect 153588 6496 153652 6500
rect 229546 6556 229610 6560
rect 229546 6500 229550 6556
rect 229550 6500 229606 6556
rect 229606 6500 229610 6556
rect 229546 6496 229610 6500
rect 229626 6556 229690 6560
rect 229626 6500 229630 6556
rect 229630 6500 229686 6556
rect 229686 6500 229690 6556
rect 229626 6496 229690 6500
rect 229706 6556 229770 6560
rect 229706 6500 229710 6556
rect 229710 6500 229766 6556
rect 229766 6500 229770 6556
rect 229706 6496 229770 6500
rect 229786 6556 229850 6560
rect 229786 6500 229790 6556
rect 229790 6500 229846 6556
rect 229846 6500 229850 6556
rect 229786 6496 229850 6500
rect 39050 6012 39114 6016
rect 39050 5956 39054 6012
rect 39054 5956 39110 6012
rect 39110 5956 39114 6012
rect 39050 5952 39114 5956
rect 39130 6012 39194 6016
rect 39130 5956 39134 6012
rect 39134 5956 39190 6012
rect 39190 5956 39194 6012
rect 39130 5952 39194 5956
rect 39210 6012 39274 6016
rect 39210 5956 39214 6012
rect 39214 5956 39270 6012
rect 39270 5956 39274 6012
rect 39210 5952 39274 5956
rect 39290 6012 39354 6016
rect 39290 5956 39294 6012
rect 39294 5956 39350 6012
rect 39350 5956 39354 6012
rect 39290 5952 39354 5956
rect 115248 6012 115312 6016
rect 115248 5956 115252 6012
rect 115252 5956 115308 6012
rect 115308 5956 115312 6012
rect 115248 5952 115312 5956
rect 115328 6012 115392 6016
rect 115328 5956 115332 6012
rect 115332 5956 115388 6012
rect 115388 5956 115392 6012
rect 115328 5952 115392 5956
rect 115408 6012 115472 6016
rect 115408 5956 115412 6012
rect 115412 5956 115468 6012
rect 115468 5956 115472 6012
rect 115408 5952 115472 5956
rect 115488 6012 115552 6016
rect 115488 5956 115492 6012
rect 115492 5956 115548 6012
rect 115548 5956 115552 6012
rect 115488 5952 115552 5956
rect 191446 6012 191510 6016
rect 191446 5956 191450 6012
rect 191450 5956 191506 6012
rect 191506 5956 191510 6012
rect 191446 5952 191510 5956
rect 191526 6012 191590 6016
rect 191526 5956 191530 6012
rect 191530 5956 191586 6012
rect 191586 5956 191590 6012
rect 191526 5952 191590 5956
rect 191606 6012 191670 6016
rect 191606 5956 191610 6012
rect 191610 5956 191666 6012
rect 191666 5956 191670 6012
rect 191606 5952 191670 5956
rect 191686 6012 191750 6016
rect 191686 5956 191690 6012
rect 191690 5956 191746 6012
rect 191746 5956 191750 6012
rect 191686 5952 191750 5956
rect 267644 6012 267708 6016
rect 267644 5956 267648 6012
rect 267648 5956 267704 6012
rect 267704 5956 267708 6012
rect 267644 5952 267708 5956
rect 267724 6012 267788 6016
rect 267724 5956 267728 6012
rect 267728 5956 267784 6012
rect 267784 5956 267788 6012
rect 267724 5952 267788 5956
rect 267804 6012 267868 6016
rect 267804 5956 267808 6012
rect 267808 5956 267864 6012
rect 267864 5956 267868 6012
rect 267804 5952 267868 5956
rect 267884 6012 267948 6016
rect 267884 5956 267888 6012
rect 267888 5956 267944 6012
rect 267944 5956 267948 6012
rect 267884 5952 267948 5956
rect 77150 5468 77214 5472
rect 77150 5412 77154 5468
rect 77154 5412 77210 5468
rect 77210 5412 77214 5468
rect 77150 5408 77214 5412
rect 77230 5468 77294 5472
rect 77230 5412 77234 5468
rect 77234 5412 77290 5468
rect 77290 5412 77294 5468
rect 77230 5408 77294 5412
rect 77310 5468 77374 5472
rect 77310 5412 77314 5468
rect 77314 5412 77370 5468
rect 77370 5412 77374 5468
rect 77310 5408 77374 5412
rect 77390 5468 77454 5472
rect 77390 5412 77394 5468
rect 77394 5412 77450 5468
rect 77450 5412 77454 5468
rect 77390 5408 77454 5412
rect 153348 5468 153412 5472
rect 153348 5412 153352 5468
rect 153352 5412 153408 5468
rect 153408 5412 153412 5468
rect 153348 5408 153412 5412
rect 153428 5468 153492 5472
rect 153428 5412 153432 5468
rect 153432 5412 153488 5468
rect 153488 5412 153492 5468
rect 153428 5408 153492 5412
rect 153508 5468 153572 5472
rect 153508 5412 153512 5468
rect 153512 5412 153568 5468
rect 153568 5412 153572 5468
rect 153508 5408 153572 5412
rect 153588 5468 153652 5472
rect 153588 5412 153592 5468
rect 153592 5412 153648 5468
rect 153648 5412 153652 5468
rect 153588 5408 153652 5412
rect 229546 5468 229610 5472
rect 229546 5412 229550 5468
rect 229550 5412 229606 5468
rect 229606 5412 229610 5468
rect 229546 5408 229610 5412
rect 229626 5468 229690 5472
rect 229626 5412 229630 5468
rect 229630 5412 229686 5468
rect 229686 5412 229690 5468
rect 229626 5408 229690 5412
rect 229706 5468 229770 5472
rect 229706 5412 229710 5468
rect 229710 5412 229766 5468
rect 229766 5412 229770 5468
rect 229706 5408 229770 5412
rect 229786 5468 229850 5472
rect 229786 5412 229790 5468
rect 229790 5412 229846 5468
rect 229846 5412 229850 5468
rect 229786 5408 229850 5412
rect 39050 4924 39114 4928
rect 39050 4868 39054 4924
rect 39054 4868 39110 4924
rect 39110 4868 39114 4924
rect 39050 4864 39114 4868
rect 39130 4924 39194 4928
rect 39130 4868 39134 4924
rect 39134 4868 39190 4924
rect 39190 4868 39194 4924
rect 39130 4864 39194 4868
rect 39210 4924 39274 4928
rect 39210 4868 39214 4924
rect 39214 4868 39270 4924
rect 39270 4868 39274 4924
rect 39210 4864 39274 4868
rect 39290 4924 39354 4928
rect 39290 4868 39294 4924
rect 39294 4868 39350 4924
rect 39350 4868 39354 4924
rect 39290 4864 39354 4868
rect 115248 4924 115312 4928
rect 115248 4868 115252 4924
rect 115252 4868 115308 4924
rect 115308 4868 115312 4924
rect 115248 4864 115312 4868
rect 115328 4924 115392 4928
rect 115328 4868 115332 4924
rect 115332 4868 115388 4924
rect 115388 4868 115392 4924
rect 115328 4864 115392 4868
rect 115408 4924 115472 4928
rect 115408 4868 115412 4924
rect 115412 4868 115468 4924
rect 115468 4868 115472 4924
rect 115408 4864 115472 4868
rect 115488 4924 115552 4928
rect 115488 4868 115492 4924
rect 115492 4868 115548 4924
rect 115548 4868 115552 4924
rect 115488 4864 115552 4868
rect 191446 4924 191510 4928
rect 191446 4868 191450 4924
rect 191450 4868 191506 4924
rect 191506 4868 191510 4924
rect 191446 4864 191510 4868
rect 191526 4924 191590 4928
rect 191526 4868 191530 4924
rect 191530 4868 191586 4924
rect 191586 4868 191590 4924
rect 191526 4864 191590 4868
rect 191606 4924 191670 4928
rect 191606 4868 191610 4924
rect 191610 4868 191666 4924
rect 191666 4868 191670 4924
rect 191606 4864 191670 4868
rect 191686 4924 191750 4928
rect 191686 4868 191690 4924
rect 191690 4868 191746 4924
rect 191746 4868 191750 4924
rect 191686 4864 191750 4868
rect 267644 4924 267708 4928
rect 267644 4868 267648 4924
rect 267648 4868 267704 4924
rect 267704 4868 267708 4924
rect 267644 4864 267708 4868
rect 267724 4924 267788 4928
rect 267724 4868 267728 4924
rect 267728 4868 267784 4924
rect 267784 4868 267788 4924
rect 267724 4864 267788 4868
rect 267804 4924 267868 4928
rect 267804 4868 267808 4924
rect 267808 4868 267864 4924
rect 267864 4868 267868 4924
rect 267804 4864 267868 4868
rect 267884 4924 267948 4928
rect 267884 4868 267888 4924
rect 267888 4868 267944 4924
rect 267944 4868 267948 4924
rect 267884 4864 267948 4868
rect 77150 4380 77214 4384
rect 77150 4324 77154 4380
rect 77154 4324 77210 4380
rect 77210 4324 77214 4380
rect 77150 4320 77214 4324
rect 77230 4380 77294 4384
rect 77230 4324 77234 4380
rect 77234 4324 77290 4380
rect 77290 4324 77294 4380
rect 77230 4320 77294 4324
rect 77310 4380 77374 4384
rect 77310 4324 77314 4380
rect 77314 4324 77370 4380
rect 77370 4324 77374 4380
rect 77310 4320 77374 4324
rect 77390 4380 77454 4384
rect 77390 4324 77394 4380
rect 77394 4324 77450 4380
rect 77450 4324 77454 4380
rect 77390 4320 77454 4324
rect 153348 4380 153412 4384
rect 153348 4324 153352 4380
rect 153352 4324 153408 4380
rect 153408 4324 153412 4380
rect 153348 4320 153412 4324
rect 153428 4380 153492 4384
rect 153428 4324 153432 4380
rect 153432 4324 153488 4380
rect 153488 4324 153492 4380
rect 153428 4320 153492 4324
rect 153508 4380 153572 4384
rect 153508 4324 153512 4380
rect 153512 4324 153568 4380
rect 153568 4324 153572 4380
rect 153508 4320 153572 4324
rect 153588 4380 153652 4384
rect 153588 4324 153592 4380
rect 153592 4324 153648 4380
rect 153648 4324 153652 4380
rect 153588 4320 153652 4324
rect 229546 4380 229610 4384
rect 229546 4324 229550 4380
rect 229550 4324 229606 4380
rect 229606 4324 229610 4380
rect 229546 4320 229610 4324
rect 229626 4380 229690 4384
rect 229626 4324 229630 4380
rect 229630 4324 229686 4380
rect 229686 4324 229690 4380
rect 229626 4320 229690 4324
rect 229706 4380 229770 4384
rect 229706 4324 229710 4380
rect 229710 4324 229766 4380
rect 229766 4324 229770 4380
rect 229706 4320 229770 4324
rect 229786 4380 229850 4384
rect 229786 4324 229790 4380
rect 229790 4324 229846 4380
rect 229846 4324 229850 4380
rect 229786 4320 229850 4324
rect 39050 3836 39114 3840
rect 39050 3780 39054 3836
rect 39054 3780 39110 3836
rect 39110 3780 39114 3836
rect 39050 3776 39114 3780
rect 39130 3836 39194 3840
rect 39130 3780 39134 3836
rect 39134 3780 39190 3836
rect 39190 3780 39194 3836
rect 39130 3776 39194 3780
rect 39210 3836 39274 3840
rect 39210 3780 39214 3836
rect 39214 3780 39270 3836
rect 39270 3780 39274 3836
rect 39210 3776 39274 3780
rect 39290 3836 39354 3840
rect 39290 3780 39294 3836
rect 39294 3780 39350 3836
rect 39350 3780 39354 3836
rect 39290 3776 39354 3780
rect 115248 3836 115312 3840
rect 115248 3780 115252 3836
rect 115252 3780 115308 3836
rect 115308 3780 115312 3836
rect 115248 3776 115312 3780
rect 115328 3836 115392 3840
rect 115328 3780 115332 3836
rect 115332 3780 115388 3836
rect 115388 3780 115392 3836
rect 115328 3776 115392 3780
rect 115408 3836 115472 3840
rect 115408 3780 115412 3836
rect 115412 3780 115468 3836
rect 115468 3780 115472 3836
rect 115408 3776 115472 3780
rect 115488 3836 115552 3840
rect 115488 3780 115492 3836
rect 115492 3780 115548 3836
rect 115548 3780 115552 3836
rect 115488 3776 115552 3780
rect 191446 3836 191510 3840
rect 191446 3780 191450 3836
rect 191450 3780 191506 3836
rect 191506 3780 191510 3836
rect 191446 3776 191510 3780
rect 191526 3836 191590 3840
rect 191526 3780 191530 3836
rect 191530 3780 191586 3836
rect 191586 3780 191590 3836
rect 191526 3776 191590 3780
rect 191606 3836 191670 3840
rect 191606 3780 191610 3836
rect 191610 3780 191666 3836
rect 191666 3780 191670 3836
rect 191606 3776 191670 3780
rect 191686 3836 191750 3840
rect 191686 3780 191690 3836
rect 191690 3780 191746 3836
rect 191746 3780 191750 3836
rect 191686 3776 191750 3780
rect 267644 3836 267708 3840
rect 267644 3780 267648 3836
rect 267648 3780 267704 3836
rect 267704 3780 267708 3836
rect 267644 3776 267708 3780
rect 267724 3836 267788 3840
rect 267724 3780 267728 3836
rect 267728 3780 267784 3836
rect 267784 3780 267788 3836
rect 267724 3776 267788 3780
rect 267804 3836 267868 3840
rect 267804 3780 267808 3836
rect 267808 3780 267864 3836
rect 267864 3780 267868 3836
rect 267804 3776 267868 3780
rect 267884 3836 267948 3840
rect 267884 3780 267888 3836
rect 267888 3780 267944 3836
rect 267944 3780 267948 3836
rect 267884 3776 267948 3780
rect 77150 3292 77214 3296
rect 77150 3236 77154 3292
rect 77154 3236 77210 3292
rect 77210 3236 77214 3292
rect 77150 3232 77214 3236
rect 77230 3292 77294 3296
rect 77230 3236 77234 3292
rect 77234 3236 77290 3292
rect 77290 3236 77294 3292
rect 77230 3232 77294 3236
rect 77310 3292 77374 3296
rect 77310 3236 77314 3292
rect 77314 3236 77370 3292
rect 77370 3236 77374 3292
rect 77310 3232 77374 3236
rect 77390 3292 77454 3296
rect 77390 3236 77394 3292
rect 77394 3236 77450 3292
rect 77450 3236 77454 3292
rect 77390 3232 77454 3236
rect 153348 3292 153412 3296
rect 153348 3236 153352 3292
rect 153352 3236 153408 3292
rect 153408 3236 153412 3292
rect 153348 3232 153412 3236
rect 153428 3292 153492 3296
rect 153428 3236 153432 3292
rect 153432 3236 153488 3292
rect 153488 3236 153492 3292
rect 153428 3232 153492 3236
rect 153508 3292 153572 3296
rect 153508 3236 153512 3292
rect 153512 3236 153568 3292
rect 153568 3236 153572 3292
rect 153508 3232 153572 3236
rect 153588 3292 153652 3296
rect 153588 3236 153592 3292
rect 153592 3236 153648 3292
rect 153648 3236 153652 3292
rect 153588 3232 153652 3236
rect 229546 3292 229610 3296
rect 229546 3236 229550 3292
rect 229550 3236 229606 3292
rect 229606 3236 229610 3292
rect 229546 3232 229610 3236
rect 229626 3292 229690 3296
rect 229626 3236 229630 3292
rect 229630 3236 229686 3292
rect 229686 3236 229690 3292
rect 229626 3232 229690 3236
rect 229706 3292 229770 3296
rect 229706 3236 229710 3292
rect 229710 3236 229766 3292
rect 229766 3236 229770 3292
rect 229706 3232 229770 3236
rect 229786 3292 229850 3296
rect 229786 3236 229790 3292
rect 229790 3236 229846 3292
rect 229846 3236 229850 3292
rect 229786 3232 229850 3236
rect 39050 2748 39114 2752
rect 39050 2692 39054 2748
rect 39054 2692 39110 2748
rect 39110 2692 39114 2748
rect 39050 2688 39114 2692
rect 39130 2748 39194 2752
rect 39130 2692 39134 2748
rect 39134 2692 39190 2748
rect 39190 2692 39194 2748
rect 39130 2688 39194 2692
rect 39210 2748 39274 2752
rect 39210 2692 39214 2748
rect 39214 2692 39270 2748
rect 39270 2692 39274 2748
rect 39210 2688 39274 2692
rect 39290 2748 39354 2752
rect 39290 2692 39294 2748
rect 39294 2692 39350 2748
rect 39350 2692 39354 2748
rect 39290 2688 39354 2692
rect 115248 2748 115312 2752
rect 115248 2692 115252 2748
rect 115252 2692 115308 2748
rect 115308 2692 115312 2748
rect 115248 2688 115312 2692
rect 115328 2748 115392 2752
rect 115328 2692 115332 2748
rect 115332 2692 115388 2748
rect 115388 2692 115392 2748
rect 115328 2688 115392 2692
rect 115408 2748 115472 2752
rect 115408 2692 115412 2748
rect 115412 2692 115468 2748
rect 115468 2692 115472 2748
rect 115408 2688 115472 2692
rect 115488 2748 115552 2752
rect 115488 2692 115492 2748
rect 115492 2692 115548 2748
rect 115548 2692 115552 2748
rect 115488 2688 115552 2692
rect 191446 2748 191510 2752
rect 191446 2692 191450 2748
rect 191450 2692 191506 2748
rect 191506 2692 191510 2748
rect 191446 2688 191510 2692
rect 191526 2748 191590 2752
rect 191526 2692 191530 2748
rect 191530 2692 191586 2748
rect 191586 2692 191590 2748
rect 191526 2688 191590 2692
rect 191606 2748 191670 2752
rect 191606 2692 191610 2748
rect 191610 2692 191666 2748
rect 191666 2692 191670 2748
rect 191606 2688 191670 2692
rect 191686 2748 191750 2752
rect 191686 2692 191690 2748
rect 191690 2692 191746 2748
rect 191746 2692 191750 2748
rect 191686 2688 191750 2692
rect 267644 2748 267708 2752
rect 267644 2692 267648 2748
rect 267648 2692 267704 2748
rect 267704 2692 267708 2748
rect 267644 2688 267708 2692
rect 267724 2748 267788 2752
rect 267724 2692 267728 2748
rect 267728 2692 267784 2748
rect 267784 2692 267788 2748
rect 267724 2688 267788 2692
rect 267804 2748 267868 2752
rect 267804 2692 267808 2748
rect 267808 2692 267864 2748
rect 267864 2692 267868 2748
rect 267804 2688 267868 2692
rect 267884 2748 267948 2752
rect 267884 2692 267888 2748
rect 267888 2692 267944 2748
rect 267944 2692 267948 2748
rect 267884 2688 267948 2692
rect 77150 2204 77214 2208
rect 77150 2148 77154 2204
rect 77154 2148 77210 2204
rect 77210 2148 77214 2204
rect 77150 2144 77214 2148
rect 77230 2204 77294 2208
rect 77230 2148 77234 2204
rect 77234 2148 77290 2204
rect 77290 2148 77294 2204
rect 77230 2144 77294 2148
rect 77310 2204 77374 2208
rect 77310 2148 77314 2204
rect 77314 2148 77370 2204
rect 77370 2148 77374 2204
rect 77310 2144 77374 2148
rect 77390 2204 77454 2208
rect 77390 2148 77394 2204
rect 77394 2148 77450 2204
rect 77450 2148 77454 2204
rect 77390 2144 77454 2148
rect 153348 2204 153412 2208
rect 153348 2148 153352 2204
rect 153352 2148 153408 2204
rect 153408 2148 153412 2204
rect 153348 2144 153412 2148
rect 153428 2204 153492 2208
rect 153428 2148 153432 2204
rect 153432 2148 153488 2204
rect 153488 2148 153492 2204
rect 153428 2144 153492 2148
rect 153508 2204 153572 2208
rect 153508 2148 153512 2204
rect 153512 2148 153568 2204
rect 153568 2148 153572 2204
rect 153508 2144 153572 2148
rect 153588 2204 153652 2208
rect 153588 2148 153592 2204
rect 153592 2148 153648 2204
rect 153648 2148 153652 2204
rect 153588 2144 153652 2148
rect 229546 2204 229610 2208
rect 229546 2148 229550 2204
rect 229550 2148 229606 2204
rect 229606 2148 229610 2204
rect 229546 2144 229610 2148
rect 229626 2204 229690 2208
rect 229626 2148 229630 2204
rect 229630 2148 229686 2204
rect 229686 2148 229690 2204
rect 229626 2144 229690 2148
rect 229706 2204 229770 2208
rect 229706 2148 229710 2204
rect 229710 2148 229766 2204
rect 229766 2148 229770 2204
rect 229706 2144 229770 2148
rect 229786 2204 229850 2208
rect 229786 2148 229790 2204
rect 229790 2148 229846 2204
rect 229846 2148 229850 2204
rect 229786 2144 229850 2148
<< metal4 >>
rect -1076 15738 -756 15780
rect -1076 15502 -1034 15738
rect -798 15502 -756 15738
rect -1076 11030 -756 15502
rect -1076 10794 -1034 11030
rect -798 10794 -756 11030
rect -1076 8118 -756 10794
rect -1076 7882 -1034 8118
rect -798 7882 -756 8118
rect -1076 5206 -756 7882
rect -1076 4970 -1034 5206
rect -798 4970 -756 5206
rect -1076 274 -756 4970
rect -416 15078 -96 15120
rect -416 14842 -374 15078
rect -138 14842 -96 15078
rect -416 12486 -96 14842
rect -416 12250 -374 12486
rect -138 12250 -96 12486
rect -416 9574 -96 12250
rect -416 9338 -374 9574
rect -138 9338 -96 9574
rect -416 6662 -96 9338
rect -416 6426 -374 6662
rect -138 6426 -96 6662
rect -416 3750 -96 6426
rect -416 3514 -374 3750
rect -138 3514 -96 3750
rect -416 934 -96 3514
rect -416 698 -374 934
rect -138 698 -96 934
rect -416 656 -96 698
rect 39042 15078 39362 15780
rect 39042 14842 39084 15078
rect 39320 14842 39362 15078
rect 39042 13632 39362 14842
rect 39042 13568 39050 13632
rect 39114 13568 39130 13632
rect 39194 13568 39210 13632
rect 39274 13568 39290 13632
rect 39354 13568 39362 13632
rect 39042 12544 39362 13568
rect 39042 12480 39050 12544
rect 39114 12486 39130 12544
rect 39194 12486 39210 12544
rect 39274 12486 39290 12544
rect 39354 12480 39362 12544
rect 39042 12250 39084 12480
rect 39320 12250 39362 12480
rect 39042 11456 39362 12250
rect 39042 11392 39050 11456
rect 39114 11392 39130 11456
rect 39194 11392 39210 11456
rect 39274 11392 39290 11456
rect 39354 11392 39362 11456
rect 39042 10368 39362 11392
rect 39042 10304 39050 10368
rect 39114 10304 39130 10368
rect 39194 10304 39210 10368
rect 39274 10304 39290 10368
rect 39354 10304 39362 10368
rect 39042 9574 39362 10304
rect 39042 9338 39084 9574
rect 39320 9338 39362 9574
rect 39042 9280 39362 9338
rect 39042 9216 39050 9280
rect 39114 9216 39130 9280
rect 39194 9216 39210 9280
rect 39274 9216 39290 9280
rect 39354 9216 39362 9280
rect 39042 8192 39362 9216
rect 39042 8128 39050 8192
rect 39114 8128 39130 8192
rect 39194 8128 39210 8192
rect 39274 8128 39290 8192
rect 39354 8128 39362 8192
rect 39042 7104 39362 8128
rect 39042 7040 39050 7104
rect 39114 7040 39130 7104
rect 39194 7040 39210 7104
rect 39274 7040 39290 7104
rect 39354 7040 39362 7104
rect 39042 6662 39362 7040
rect 39042 6426 39084 6662
rect 39320 6426 39362 6662
rect 39042 6016 39362 6426
rect 39042 5952 39050 6016
rect 39114 5952 39130 6016
rect 39194 5952 39210 6016
rect 39274 5952 39290 6016
rect 39354 5952 39362 6016
rect 39042 4928 39362 5952
rect 39042 4864 39050 4928
rect 39114 4864 39130 4928
rect 39194 4864 39210 4928
rect 39274 4864 39290 4928
rect 39354 4864 39362 4928
rect 39042 3840 39362 4864
rect 39042 3776 39050 3840
rect 39114 3776 39130 3840
rect 39194 3776 39210 3840
rect 39274 3776 39290 3840
rect 39354 3776 39362 3840
rect 39042 3750 39362 3776
rect 39042 3514 39084 3750
rect 39320 3514 39362 3750
rect 39042 2752 39362 3514
rect 39042 2688 39050 2752
rect 39114 2688 39130 2752
rect 39194 2688 39210 2752
rect 39274 2688 39290 2752
rect 39354 2688 39362 2752
rect 39042 934 39362 2688
rect 39042 698 39084 934
rect 39320 698 39362 934
rect -1076 38 -1034 274
rect -798 38 -756 274
rect -1076 -4 -756 38
rect 39042 -4 39362 698
rect 77142 15738 77462 15780
rect 77142 15502 77184 15738
rect 77420 15502 77462 15738
rect 77142 13088 77462 15502
rect 77142 13024 77150 13088
rect 77214 13024 77230 13088
rect 77294 13024 77310 13088
rect 77374 13024 77390 13088
rect 77454 13024 77462 13088
rect 77142 12000 77462 13024
rect 77142 11936 77150 12000
rect 77214 11936 77230 12000
rect 77294 11936 77310 12000
rect 77374 11936 77390 12000
rect 77454 11936 77462 12000
rect 77142 11030 77462 11936
rect 77142 10912 77184 11030
rect 77420 10912 77462 11030
rect 77142 10848 77150 10912
rect 77454 10848 77462 10912
rect 77142 10794 77184 10848
rect 77420 10794 77462 10848
rect 77142 9824 77462 10794
rect 77142 9760 77150 9824
rect 77214 9760 77230 9824
rect 77294 9760 77310 9824
rect 77374 9760 77390 9824
rect 77454 9760 77462 9824
rect 77142 8736 77462 9760
rect 77142 8672 77150 8736
rect 77214 8672 77230 8736
rect 77294 8672 77310 8736
rect 77374 8672 77390 8736
rect 77454 8672 77462 8736
rect 77142 8118 77462 8672
rect 77142 7882 77184 8118
rect 77420 7882 77462 8118
rect 77142 7648 77462 7882
rect 77142 7584 77150 7648
rect 77214 7584 77230 7648
rect 77294 7584 77310 7648
rect 77374 7584 77390 7648
rect 77454 7584 77462 7648
rect 77142 6560 77462 7584
rect 77142 6496 77150 6560
rect 77214 6496 77230 6560
rect 77294 6496 77310 6560
rect 77374 6496 77390 6560
rect 77454 6496 77462 6560
rect 77142 5472 77462 6496
rect 77142 5408 77150 5472
rect 77214 5408 77230 5472
rect 77294 5408 77310 5472
rect 77374 5408 77390 5472
rect 77454 5408 77462 5472
rect 77142 5206 77462 5408
rect 77142 4970 77184 5206
rect 77420 4970 77462 5206
rect 77142 4384 77462 4970
rect 77142 4320 77150 4384
rect 77214 4320 77230 4384
rect 77294 4320 77310 4384
rect 77374 4320 77390 4384
rect 77454 4320 77462 4384
rect 77142 3296 77462 4320
rect 77142 3232 77150 3296
rect 77214 3232 77230 3296
rect 77294 3232 77310 3296
rect 77374 3232 77390 3296
rect 77454 3232 77462 3296
rect 77142 2208 77462 3232
rect 77142 2144 77150 2208
rect 77214 2144 77230 2208
rect 77294 2144 77310 2208
rect 77374 2144 77390 2208
rect 77454 2144 77462 2208
rect 77142 274 77462 2144
rect 77142 38 77184 274
rect 77420 38 77462 274
rect 77142 -4 77462 38
rect 115240 15078 115560 15780
rect 115240 14842 115282 15078
rect 115518 14842 115560 15078
rect 115240 13632 115560 14842
rect 115240 13568 115248 13632
rect 115312 13568 115328 13632
rect 115392 13568 115408 13632
rect 115472 13568 115488 13632
rect 115552 13568 115560 13632
rect 115240 12544 115560 13568
rect 115240 12480 115248 12544
rect 115312 12486 115328 12544
rect 115392 12486 115408 12544
rect 115472 12486 115488 12544
rect 115552 12480 115560 12544
rect 115240 12250 115282 12480
rect 115518 12250 115560 12480
rect 115240 11456 115560 12250
rect 115240 11392 115248 11456
rect 115312 11392 115328 11456
rect 115392 11392 115408 11456
rect 115472 11392 115488 11456
rect 115552 11392 115560 11456
rect 115240 10368 115560 11392
rect 115240 10304 115248 10368
rect 115312 10304 115328 10368
rect 115392 10304 115408 10368
rect 115472 10304 115488 10368
rect 115552 10304 115560 10368
rect 115240 9574 115560 10304
rect 115240 9338 115282 9574
rect 115518 9338 115560 9574
rect 115240 9280 115560 9338
rect 115240 9216 115248 9280
rect 115312 9216 115328 9280
rect 115392 9216 115408 9280
rect 115472 9216 115488 9280
rect 115552 9216 115560 9280
rect 115240 8192 115560 9216
rect 115240 8128 115248 8192
rect 115312 8128 115328 8192
rect 115392 8128 115408 8192
rect 115472 8128 115488 8192
rect 115552 8128 115560 8192
rect 115240 7104 115560 8128
rect 115240 7040 115248 7104
rect 115312 7040 115328 7104
rect 115392 7040 115408 7104
rect 115472 7040 115488 7104
rect 115552 7040 115560 7104
rect 115240 6662 115560 7040
rect 115240 6426 115282 6662
rect 115518 6426 115560 6662
rect 115240 6016 115560 6426
rect 115240 5952 115248 6016
rect 115312 5952 115328 6016
rect 115392 5952 115408 6016
rect 115472 5952 115488 6016
rect 115552 5952 115560 6016
rect 115240 4928 115560 5952
rect 115240 4864 115248 4928
rect 115312 4864 115328 4928
rect 115392 4864 115408 4928
rect 115472 4864 115488 4928
rect 115552 4864 115560 4928
rect 115240 3840 115560 4864
rect 115240 3776 115248 3840
rect 115312 3776 115328 3840
rect 115392 3776 115408 3840
rect 115472 3776 115488 3840
rect 115552 3776 115560 3840
rect 115240 3750 115560 3776
rect 115240 3514 115282 3750
rect 115518 3514 115560 3750
rect 115240 2752 115560 3514
rect 115240 2688 115248 2752
rect 115312 2688 115328 2752
rect 115392 2688 115408 2752
rect 115472 2688 115488 2752
rect 115552 2688 115560 2752
rect 115240 934 115560 2688
rect 115240 698 115282 934
rect 115518 698 115560 934
rect 115240 -4 115560 698
rect 153340 15738 153660 15780
rect 153340 15502 153382 15738
rect 153618 15502 153660 15738
rect 153340 13088 153660 15502
rect 153340 13024 153348 13088
rect 153412 13024 153428 13088
rect 153492 13024 153508 13088
rect 153572 13024 153588 13088
rect 153652 13024 153660 13088
rect 153340 12000 153660 13024
rect 153340 11936 153348 12000
rect 153412 11936 153428 12000
rect 153492 11936 153508 12000
rect 153572 11936 153588 12000
rect 153652 11936 153660 12000
rect 153340 11030 153660 11936
rect 153340 10912 153382 11030
rect 153618 10912 153660 11030
rect 153340 10848 153348 10912
rect 153652 10848 153660 10912
rect 153340 10794 153382 10848
rect 153618 10794 153660 10848
rect 153340 9824 153660 10794
rect 153340 9760 153348 9824
rect 153412 9760 153428 9824
rect 153492 9760 153508 9824
rect 153572 9760 153588 9824
rect 153652 9760 153660 9824
rect 153340 8736 153660 9760
rect 153340 8672 153348 8736
rect 153412 8672 153428 8736
rect 153492 8672 153508 8736
rect 153572 8672 153588 8736
rect 153652 8672 153660 8736
rect 153340 8118 153660 8672
rect 153340 7882 153382 8118
rect 153618 7882 153660 8118
rect 153340 7648 153660 7882
rect 153340 7584 153348 7648
rect 153412 7584 153428 7648
rect 153492 7584 153508 7648
rect 153572 7584 153588 7648
rect 153652 7584 153660 7648
rect 153340 6560 153660 7584
rect 153340 6496 153348 6560
rect 153412 6496 153428 6560
rect 153492 6496 153508 6560
rect 153572 6496 153588 6560
rect 153652 6496 153660 6560
rect 153340 5472 153660 6496
rect 153340 5408 153348 5472
rect 153412 5408 153428 5472
rect 153492 5408 153508 5472
rect 153572 5408 153588 5472
rect 153652 5408 153660 5472
rect 153340 5206 153660 5408
rect 153340 4970 153382 5206
rect 153618 4970 153660 5206
rect 153340 4384 153660 4970
rect 153340 4320 153348 4384
rect 153412 4320 153428 4384
rect 153492 4320 153508 4384
rect 153572 4320 153588 4384
rect 153652 4320 153660 4384
rect 153340 3296 153660 4320
rect 153340 3232 153348 3296
rect 153412 3232 153428 3296
rect 153492 3232 153508 3296
rect 153572 3232 153588 3296
rect 153652 3232 153660 3296
rect 153340 2208 153660 3232
rect 153340 2144 153348 2208
rect 153412 2144 153428 2208
rect 153492 2144 153508 2208
rect 153572 2144 153588 2208
rect 153652 2144 153660 2208
rect 153340 274 153660 2144
rect 153340 38 153382 274
rect 153618 38 153660 274
rect 153340 -4 153660 38
rect 191438 15078 191758 15780
rect 191438 14842 191480 15078
rect 191716 14842 191758 15078
rect 191438 13632 191758 14842
rect 191438 13568 191446 13632
rect 191510 13568 191526 13632
rect 191590 13568 191606 13632
rect 191670 13568 191686 13632
rect 191750 13568 191758 13632
rect 191438 12544 191758 13568
rect 191438 12480 191446 12544
rect 191510 12486 191526 12544
rect 191590 12486 191606 12544
rect 191670 12486 191686 12544
rect 191750 12480 191758 12544
rect 191438 12250 191480 12480
rect 191716 12250 191758 12480
rect 191438 11456 191758 12250
rect 191438 11392 191446 11456
rect 191510 11392 191526 11456
rect 191590 11392 191606 11456
rect 191670 11392 191686 11456
rect 191750 11392 191758 11456
rect 191438 10368 191758 11392
rect 191438 10304 191446 10368
rect 191510 10304 191526 10368
rect 191590 10304 191606 10368
rect 191670 10304 191686 10368
rect 191750 10304 191758 10368
rect 191438 9574 191758 10304
rect 191438 9338 191480 9574
rect 191716 9338 191758 9574
rect 191438 9280 191758 9338
rect 191438 9216 191446 9280
rect 191510 9216 191526 9280
rect 191590 9216 191606 9280
rect 191670 9216 191686 9280
rect 191750 9216 191758 9280
rect 191438 8192 191758 9216
rect 191438 8128 191446 8192
rect 191510 8128 191526 8192
rect 191590 8128 191606 8192
rect 191670 8128 191686 8192
rect 191750 8128 191758 8192
rect 191438 7104 191758 8128
rect 191438 7040 191446 7104
rect 191510 7040 191526 7104
rect 191590 7040 191606 7104
rect 191670 7040 191686 7104
rect 191750 7040 191758 7104
rect 191438 6662 191758 7040
rect 191438 6426 191480 6662
rect 191716 6426 191758 6662
rect 191438 6016 191758 6426
rect 191438 5952 191446 6016
rect 191510 5952 191526 6016
rect 191590 5952 191606 6016
rect 191670 5952 191686 6016
rect 191750 5952 191758 6016
rect 191438 4928 191758 5952
rect 191438 4864 191446 4928
rect 191510 4864 191526 4928
rect 191590 4864 191606 4928
rect 191670 4864 191686 4928
rect 191750 4864 191758 4928
rect 191438 3840 191758 4864
rect 191438 3776 191446 3840
rect 191510 3776 191526 3840
rect 191590 3776 191606 3840
rect 191670 3776 191686 3840
rect 191750 3776 191758 3840
rect 191438 3750 191758 3776
rect 191438 3514 191480 3750
rect 191716 3514 191758 3750
rect 191438 2752 191758 3514
rect 191438 2688 191446 2752
rect 191510 2688 191526 2752
rect 191590 2688 191606 2752
rect 191670 2688 191686 2752
rect 191750 2688 191758 2752
rect 191438 934 191758 2688
rect 191438 698 191480 934
rect 191716 698 191758 934
rect 191438 -4 191758 698
rect 229538 15738 229858 15780
rect 229538 15502 229580 15738
rect 229816 15502 229858 15738
rect 229538 13088 229858 15502
rect 229538 13024 229546 13088
rect 229610 13024 229626 13088
rect 229690 13024 229706 13088
rect 229770 13024 229786 13088
rect 229850 13024 229858 13088
rect 229538 12000 229858 13024
rect 229538 11936 229546 12000
rect 229610 11936 229626 12000
rect 229690 11936 229706 12000
rect 229770 11936 229786 12000
rect 229850 11936 229858 12000
rect 229538 11030 229858 11936
rect 229538 10912 229580 11030
rect 229816 10912 229858 11030
rect 229538 10848 229546 10912
rect 229850 10848 229858 10912
rect 229538 10794 229580 10848
rect 229816 10794 229858 10848
rect 229538 9824 229858 10794
rect 229538 9760 229546 9824
rect 229610 9760 229626 9824
rect 229690 9760 229706 9824
rect 229770 9760 229786 9824
rect 229850 9760 229858 9824
rect 229538 8736 229858 9760
rect 229538 8672 229546 8736
rect 229610 8672 229626 8736
rect 229690 8672 229706 8736
rect 229770 8672 229786 8736
rect 229850 8672 229858 8736
rect 229538 8118 229858 8672
rect 229538 7882 229580 8118
rect 229816 7882 229858 8118
rect 229538 7648 229858 7882
rect 229538 7584 229546 7648
rect 229610 7584 229626 7648
rect 229690 7584 229706 7648
rect 229770 7584 229786 7648
rect 229850 7584 229858 7648
rect 229538 6560 229858 7584
rect 229538 6496 229546 6560
rect 229610 6496 229626 6560
rect 229690 6496 229706 6560
rect 229770 6496 229786 6560
rect 229850 6496 229858 6560
rect 229538 5472 229858 6496
rect 229538 5408 229546 5472
rect 229610 5408 229626 5472
rect 229690 5408 229706 5472
rect 229770 5408 229786 5472
rect 229850 5408 229858 5472
rect 229538 5206 229858 5408
rect 229538 4970 229580 5206
rect 229816 4970 229858 5206
rect 229538 4384 229858 4970
rect 229538 4320 229546 4384
rect 229610 4320 229626 4384
rect 229690 4320 229706 4384
rect 229770 4320 229786 4384
rect 229850 4320 229858 4384
rect 229538 3296 229858 4320
rect 229538 3232 229546 3296
rect 229610 3232 229626 3296
rect 229690 3232 229706 3296
rect 229770 3232 229786 3296
rect 229850 3232 229858 3296
rect 229538 2208 229858 3232
rect 229538 2144 229546 2208
rect 229610 2144 229626 2208
rect 229690 2144 229706 2208
rect 229770 2144 229786 2208
rect 229850 2144 229858 2208
rect 229538 274 229858 2144
rect 229538 38 229580 274
rect 229816 38 229858 274
rect 229538 -4 229858 38
rect 267636 15078 267956 15780
rect 307668 15738 307988 15780
rect 307668 15502 307710 15738
rect 307946 15502 307988 15738
rect 267636 14842 267678 15078
rect 267914 14842 267956 15078
rect 267636 13632 267956 14842
rect 267636 13568 267644 13632
rect 267708 13568 267724 13632
rect 267788 13568 267804 13632
rect 267868 13568 267884 13632
rect 267948 13568 267956 13632
rect 267636 12544 267956 13568
rect 267636 12480 267644 12544
rect 267708 12486 267724 12544
rect 267788 12486 267804 12544
rect 267868 12486 267884 12544
rect 267948 12480 267956 12544
rect 267636 12250 267678 12480
rect 267914 12250 267956 12480
rect 267636 11456 267956 12250
rect 267636 11392 267644 11456
rect 267708 11392 267724 11456
rect 267788 11392 267804 11456
rect 267868 11392 267884 11456
rect 267948 11392 267956 11456
rect 267636 10368 267956 11392
rect 267636 10304 267644 10368
rect 267708 10304 267724 10368
rect 267788 10304 267804 10368
rect 267868 10304 267884 10368
rect 267948 10304 267956 10368
rect 267636 9574 267956 10304
rect 267636 9338 267678 9574
rect 267914 9338 267956 9574
rect 267636 9280 267956 9338
rect 267636 9216 267644 9280
rect 267708 9216 267724 9280
rect 267788 9216 267804 9280
rect 267868 9216 267884 9280
rect 267948 9216 267956 9280
rect 267636 8192 267956 9216
rect 267636 8128 267644 8192
rect 267708 8128 267724 8192
rect 267788 8128 267804 8192
rect 267868 8128 267884 8192
rect 267948 8128 267956 8192
rect 267636 7104 267956 8128
rect 267636 7040 267644 7104
rect 267708 7040 267724 7104
rect 267788 7040 267804 7104
rect 267868 7040 267884 7104
rect 267948 7040 267956 7104
rect 267636 6662 267956 7040
rect 267636 6426 267678 6662
rect 267914 6426 267956 6662
rect 267636 6016 267956 6426
rect 267636 5952 267644 6016
rect 267708 5952 267724 6016
rect 267788 5952 267804 6016
rect 267868 5952 267884 6016
rect 267948 5952 267956 6016
rect 267636 4928 267956 5952
rect 267636 4864 267644 4928
rect 267708 4864 267724 4928
rect 267788 4864 267804 4928
rect 267868 4864 267884 4928
rect 267948 4864 267956 4928
rect 267636 3840 267956 4864
rect 267636 3776 267644 3840
rect 267708 3776 267724 3840
rect 267788 3776 267804 3840
rect 267868 3776 267884 3840
rect 267948 3776 267956 3840
rect 267636 3750 267956 3776
rect 267636 3514 267678 3750
rect 267914 3514 267956 3750
rect 267636 2752 267956 3514
rect 267636 2688 267644 2752
rect 267708 2688 267724 2752
rect 267788 2688 267804 2752
rect 267868 2688 267884 2752
rect 267948 2688 267956 2752
rect 267636 934 267956 2688
rect 267636 698 267678 934
rect 267914 698 267956 934
rect 267636 -4 267956 698
rect 307008 15078 307328 15120
rect 307008 14842 307050 15078
rect 307286 14842 307328 15078
rect 307008 12486 307328 14842
rect 307008 12250 307050 12486
rect 307286 12250 307328 12486
rect 307008 9574 307328 12250
rect 307008 9338 307050 9574
rect 307286 9338 307328 9574
rect 307008 6662 307328 9338
rect 307008 6426 307050 6662
rect 307286 6426 307328 6662
rect 307008 3750 307328 6426
rect 307008 3514 307050 3750
rect 307286 3514 307328 3750
rect 307008 934 307328 3514
rect 307008 698 307050 934
rect 307286 698 307328 934
rect 307008 656 307328 698
rect 307668 11030 307988 15502
rect 307668 10794 307710 11030
rect 307946 10794 307988 11030
rect 307668 8118 307988 10794
rect 307668 7882 307710 8118
rect 307946 7882 307988 8118
rect 307668 5206 307988 7882
rect 307668 4970 307710 5206
rect 307946 4970 307988 5206
rect 307668 274 307988 4970
rect 307668 38 307710 274
rect 307946 38 307988 274
rect 307668 -4 307988 38
<< via4 >>
rect -1034 15502 -798 15738
rect -1034 10794 -798 11030
rect -1034 7882 -798 8118
rect -1034 4970 -798 5206
rect -374 14842 -138 15078
rect -374 12250 -138 12486
rect -374 9338 -138 9574
rect -374 6426 -138 6662
rect -374 3514 -138 3750
rect -374 698 -138 934
rect 39084 14842 39320 15078
rect 39084 12480 39114 12486
rect 39114 12480 39130 12486
rect 39130 12480 39194 12486
rect 39194 12480 39210 12486
rect 39210 12480 39274 12486
rect 39274 12480 39290 12486
rect 39290 12480 39320 12486
rect 39084 12250 39320 12480
rect 39084 9338 39320 9574
rect 39084 6426 39320 6662
rect 39084 3514 39320 3750
rect 39084 698 39320 934
rect -1034 38 -798 274
rect 77184 15502 77420 15738
rect 77184 10912 77420 11030
rect 77184 10848 77214 10912
rect 77214 10848 77230 10912
rect 77230 10848 77294 10912
rect 77294 10848 77310 10912
rect 77310 10848 77374 10912
rect 77374 10848 77390 10912
rect 77390 10848 77420 10912
rect 77184 10794 77420 10848
rect 77184 7882 77420 8118
rect 77184 4970 77420 5206
rect 77184 38 77420 274
rect 115282 14842 115518 15078
rect 115282 12480 115312 12486
rect 115312 12480 115328 12486
rect 115328 12480 115392 12486
rect 115392 12480 115408 12486
rect 115408 12480 115472 12486
rect 115472 12480 115488 12486
rect 115488 12480 115518 12486
rect 115282 12250 115518 12480
rect 115282 9338 115518 9574
rect 115282 6426 115518 6662
rect 115282 3514 115518 3750
rect 115282 698 115518 934
rect 153382 15502 153618 15738
rect 153382 10912 153618 11030
rect 153382 10848 153412 10912
rect 153412 10848 153428 10912
rect 153428 10848 153492 10912
rect 153492 10848 153508 10912
rect 153508 10848 153572 10912
rect 153572 10848 153588 10912
rect 153588 10848 153618 10912
rect 153382 10794 153618 10848
rect 153382 7882 153618 8118
rect 153382 4970 153618 5206
rect 153382 38 153618 274
rect 191480 14842 191716 15078
rect 191480 12480 191510 12486
rect 191510 12480 191526 12486
rect 191526 12480 191590 12486
rect 191590 12480 191606 12486
rect 191606 12480 191670 12486
rect 191670 12480 191686 12486
rect 191686 12480 191716 12486
rect 191480 12250 191716 12480
rect 191480 9338 191716 9574
rect 191480 6426 191716 6662
rect 191480 3514 191716 3750
rect 191480 698 191716 934
rect 229580 15502 229816 15738
rect 229580 10912 229816 11030
rect 229580 10848 229610 10912
rect 229610 10848 229626 10912
rect 229626 10848 229690 10912
rect 229690 10848 229706 10912
rect 229706 10848 229770 10912
rect 229770 10848 229786 10912
rect 229786 10848 229816 10912
rect 229580 10794 229816 10848
rect 229580 7882 229816 8118
rect 229580 4970 229816 5206
rect 229580 38 229816 274
rect 307710 15502 307946 15738
rect 267678 14842 267914 15078
rect 267678 12480 267708 12486
rect 267708 12480 267724 12486
rect 267724 12480 267788 12486
rect 267788 12480 267804 12486
rect 267804 12480 267868 12486
rect 267868 12480 267884 12486
rect 267884 12480 267914 12486
rect 267678 12250 267914 12480
rect 267678 9338 267914 9574
rect 267678 6426 267914 6662
rect 267678 3514 267914 3750
rect 267678 698 267914 934
rect 307050 14842 307286 15078
rect 307050 12250 307286 12486
rect 307050 9338 307286 9574
rect 307050 6426 307286 6662
rect 307050 3514 307286 3750
rect 307050 698 307286 934
rect 307710 10794 307946 11030
rect 307710 7882 307946 8118
rect 307710 4970 307946 5206
rect 307710 38 307946 274
<< metal5 >>
rect -1076 15738 307988 15780
rect -1076 15502 -1034 15738
rect -798 15502 77184 15738
rect 77420 15502 153382 15738
rect 153618 15502 229580 15738
rect 229816 15502 307710 15738
rect 307946 15502 307988 15738
rect -1076 15460 307988 15502
rect -416 15078 307328 15120
rect -416 14842 -374 15078
rect -138 14842 39084 15078
rect 39320 14842 115282 15078
rect 115518 14842 191480 15078
rect 191716 14842 267678 15078
rect 267914 14842 307050 15078
rect 307286 14842 307328 15078
rect -416 14800 307328 14842
rect -1076 12486 307988 12528
rect -1076 12250 -374 12486
rect -138 12250 39084 12486
rect 39320 12250 115282 12486
rect 115518 12250 191480 12486
rect 191716 12250 267678 12486
rect 267914 12250 307050 12486
rect 307286 12250 307988 12486
rect -1076 12208 307988 12250
rect -1076 11030 307988 11072
rect -1076 10794 -1034 11030
rect -798 10794 77184 11030
rect 77420 10794 153382 11030
rect 153618 10794 229580 11030
rect 229816 10794 307710 11030
rect 307946 10794 307988 11030
rect -1076 10752 307988 10794
rect -1076 9574 307988 9616
rect -1076 9338 -374 9574
rect -138 9338 39084 9574
rect 39320 9338 115282 9574
rect 115518 9338 191480 9574
rect 191716 9338 267678 9574
rect 267914 9338 307050 9574
rect 307286 9338 307988 9574
rect -1076 9296 307988 9338
rect -1076 8118 307988 8160
rect -1076 7882 -1034 8118
rect -798 7882 77184 8118
rect 77420 7882 153382 8118
rect 153618 7882 229580 8118
rect 229816 7882 307710 8118
rect 307946 7882 307988 8118
rect -1076 7840 307988 7882
rect -1076 6662 307988 6704
rect -1076 6426 -374 6662
rect -138 6426 39084 6662
rect 39320 6426 115282 6662
rect 115518 6426 191480 6662
rect 191716 6426 267678 6662
rect 267914 6426 307050 6662
rect 307286 6426 307988 6662
rect -1076 6384 307988 6426
rect -1076 5206 307988 5248
rect -1076 4970 -1034 5206
rect -798 4970 77184 5206
rect 77420 4970 153382 5206
rect 153618 4970 229580 5206
rect 229816 4970 307710 5206
rect 307946 4970 307988 5206
rect -1076 4928 307988 4970
rect -1076 3750 307988 3792
rect -1076 3514 -374 3750
rect -138 3514 39084 3750
rect 39320 3514 115282 3750
rect 115518 3514 191480 3750
rect 191716 3514 267678 3750
rect 267914 3514 307050 3750
rect 307286 3514 307988 3750
rect -1076 3472 307988 3514
rect -416 934 307328 976
rect -416 698 -374 934
rect -138 698 39084 934
rect 39320 698 115282 934
rect 115518 698 191480 934
rect 191716 698 267678 934
rect 267914 698 307050 934
rect 307286 698 307328 934
rect -416 656 307328 698
rect -1076 274 307988 316
rect -1076 38 -1034 274
rect -798 38 77184 274
rect 77420 38 153382 274
rect 153618 38 229580 274
rect 229816 38 307710 274
rect 307946 38 307988 274
rect -1076 -4 307988 38
use sky130_fd_sc_hd__buf_4  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 137724 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _349_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 56948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 58144 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 56212 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1758069660
transform 1 0 56120 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1758069660
transform 1 0 57960 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1758069660
transform 1 0 54924 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp 1758069660
transform 1 0 55292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1758069660
transform 1 0 53544 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _357_
timestamp 1758069660
transform 1 0 51980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1758069660
transform 1 0 50968 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _359_
timestamp 1758069660
transform 1 0 52808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _360_
timestamp 1758069660
transform 1 0 43608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1758069660
transform 1 0 43056 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1758069660
transform 1 0 41676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1758069660
transform 1 0 44988 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1758069660
transform 1 0 41584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _365_
timestamp 1758069660
transform 1 0 40204 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp 1758069660
transform 1 0 40296 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1758069660
transform 1 0 39652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1758069660
transform 1 0 39008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1758069660
transform 1 0 37996 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1758069660
transform 1 0 38456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _371_
timestamp 1758069660
transform 1 0 36984 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1758069660
transform 1 0 34316 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1758069660
transform 1 0 33948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1758069660
transform 1 0 32108 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1758069660
transform 1 0 32752 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1758069660
transform 1 0 31832 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1758069660
transform 1 0 33396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1758069660
transform 1 0 28612 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1758069660
transform 1 0 34960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1758069660
transform 1 0 30268 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _381_
timestamp 1758069660
transform 1 0 32108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _382_
timestamp 1758069660
transform 1 0 36248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1758069660
transform 1 0 28244 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _384_
timestamp 1758069660
transform 1 0 30912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1758069660
transform 1 0 28428 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1758069660
transform 1 0 29624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1758069660
transform 1 0 25668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1758069660
transform 1 0 28796 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1758069660
transform 1 0 27048 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _390_
timestamp 1758069660
transform 1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1758069660
transform 1 0 27416 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _392_
timestamp 1758069660
transform 1 0 31096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 145728 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1758069660
transform 1 0 154468 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _395_
timestamp 1758069660
transform 1 0 150788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1758069660
transform 1 0 195500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _397_
timestamp 1758069660
transform 1 0 188508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1758069660
transform 1 0 194396 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1758069660
transform 1 0 193108 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1758069660
transform 1 0 196972 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _401_
timestamp 1758069660
transform 1 0 192280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1758069660
transform 1 0 198168 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 1758069660
transform 1 0 196236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _404_
timestamp 1758069660
transform 1 0 248952 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _405_
timestamp 1758069660
transform 1 0 262384 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1758069660
transform 1 0 268824 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1758069660
transform 1 0 267720 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1758069660
transform 1 0 272504 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1758069660
transform 1 0 268364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1758069660
transform 1 0 271676 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1758069660
transform 1 0 267076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1758069660
transform 1 0 270020 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1758069660
transform 1 0 267720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1758069660
transform 1 0 271308 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 1758069660
transform 1 0 267996 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _416_
timestamp 1758069660
transform 1 0 261740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 1758069660
transform 1 0 267812 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _418_
timestamp 1758069660
transform 1 0 265788 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp 1758069660
transform 1 0 266800 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 1758069660
transform 1 0 264960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp 1758069660
transform 1 0 267444 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _422_
timestamp 1758069660
transform 1 0 263948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp 1758069660
transform 1 0 265236 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 1758069660
transform 1 0 264592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _425_
timestamp 1758069660
transform 1 0 262660 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1758069660
transform 1 0 264592 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _427_
timestamp 1758069660
transform 1 0 251804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _428_
timestamp 1758069660
transform 1 0 255852 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _429_
timestamp 1758069660
transform 1 0 253644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _430_
timestamp 1758069660
transform 1 0 254748 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _431_
timestamp 1758069660
transform 1 0 253736 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _432_
timestamp 1758069660
transform 1 0 253644 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _433_
timestamp 1758069660
transform 1 0 253092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _434_
timestamp 1758069660
transform 1 0 251988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1758069660
transform 1 0 251804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _436_
timestamp 1758069660
transform 1 0 249504 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _437_
timestamp 1758069660
transform 1 0 251068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _438_
timestamp 1758069660
transform 1 0 243708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _439_
timestamp 1758069660
transform 1 0 242328 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _440_
timestamp 1758069660
transform 1 0 243524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _441_
timestamp 1758069660
transform 1 0 240856 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _442_
timestamp 1758069660
transform 1 0 241408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp 1758069660
transform 1 0 239844 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _444_
timestamp 1758069660
transform 1 0 241040 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _445_
timestamp 1758069660
transform 1 0 238740 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _446_
timestamp 1758069660
transform 1 0 239936 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp 1758069660
transform 1 0 236716 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1758069660
transform 1 0 236808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _449_
timestamp 1758069660
transform 1 0 238556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _450_
timestamp 1758069660
transform 1 0 230920 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _451_
timestamp 1758069660
transform 1 0 231564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp 1758069660
transform 1 0 229080 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _453_
timestamp 1758069660
transform 1 0 229172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp 1758069660
transform 1 0 227884 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _455_
timestamp 1758069660
transform 1 0 230092 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _456_
timestamp 1758069660
transform 1 0 226596 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _457_
timestamp 1758069660
transform 1 0 227148 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _458_
timestamp 1758069660
transform 1 0 223652 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _459_
timestamp 1758069660
transform 1 0 226504 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _460_
timestamp 1758069660
transform 1 0 165784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _461_
timestamp 1758069660
transform 1 0 193384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1758069660
transform 1 0 207276 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _463_
timestamp 1758069660
transform 1 0 202124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _464_
timestamp 1758069660
transform 1 0 204792 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _465_
timestamp 1758069660
transform 1 0 202860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1758069660
transform 1 0 203596 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _467_
timestamp 1758069660
transform 1 0 199824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp 1758069660
transform 1 0 202860 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _469_
timestamp 1758069660
transform 1 0 202860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _470_
timestamp 1758069660
transform 1 0 200468 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _471_
timestamp 1758069660
transform 1 0 201664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _472_
timestamp 1758069660
transform 1 0 189244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _473_
timestamp 1758069660
transform 1 0 196972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _474_
timestamp 1758069660
transform 1 0 192464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp 1758069660
transform 1 0 193016 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _476_
timestamp 1758069660
transform 1 0 189428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _477_
timestamp 1758069660
transform 1 0 190532 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _478_
timestamp 1758069660
transform 1 0 191084 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _479_
timestamp 1758069660
transform 1 0 191820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _480_
timestamp 1758069660
transform 1 0 191820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _481_
timestamp 1758069660
transform 1 0 187956 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _482_
timestamp 1758069660
transform 1 0 190164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _483_
timestamp 1758069660
transform 1 0 175536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _484_
timestamp 1758069660
transform 1 0 181516 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _485_
timestamp 1758069660
transform 1 0 178940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _486_
timestamp 1758069660
transform 1 0 178756 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _487_
timestamp 1758069660
transform 1 0 180780 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _488_
timestamp 1758069660
transform 1 0 177560 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _489_
timestamp 1758069660
transform 1 0 174984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _490_
timestamp 1758069660
transform 1 0 176548 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _491_
timestamp 1758069660
transform 1 0 176456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _492_
timestamp 1758069660
transform 1 0 173788 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _493_
timestamp 1758069660
transform 1 0 175628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _494_
timestamp 1758069660
transform 1 0 167256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _495_
timestamp 1758069660
transform 1 0 166060 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _496_
timestamp 1758069660
transform 1 0 162656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _497_
timestamp 1758069660
transform 1 0 164036 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _498_
timestamp 1758069660
transform 1 0 163484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _499_
timestamp 1758069660
transform 1 0 162012 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _500_
timestamp 1758069660
transform 1 0 162012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _501_
timestamp 1758069660
transform 1 0 160816 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _502_
timestamp 1758069660
transform 1 0 160908 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _503_
timestamp 1758069660
transform 1 0 158792 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp 1758069660
transform 1 0 159988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _505_
timestamp 1758069660
transform 1 0 161092 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _506_
timestamp 1758069660
transform 1 0 153272 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _507_
timestamp 1758069660
transform 1 0 154100 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _508_
timestamp 1758069660
transform 1 0 151064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _509_
timestamp 1758069660
transform 1 0 151064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _510_
timestamp 1758069660
transform 1 0 151616 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _511_
timestamp 1758069660
transform 1 0 148856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _512_
timestamp 1758069660
transform 1 0 148028 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _513_
timestamp 1758069660
transform 1 0 147292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _514_
timestamp 1758069660
transform 1 0 145452 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _515_
timestamp 1758069660
transform 1 0 147568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 131652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _517_
timestamp 1758069660
transform 1 0 125396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _518_
timestamp 1758069660
transform 1 0 133124 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1758069660
transform 1 0 131744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _520_
timestamp 1758069660
transform 1 0 131284 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1758069660
transform 1 0 132388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _522_
timestamp 1758069660
transform 1 0 130456 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1758069660
transform 1 0 128064 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _524_
timestamp 1758069660
transform 1 0 128708 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1758069660
transform 1 0 128432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _526_
timestamp 1758069660
transform 1 0 126132 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _527_
timestamp 1758069660
transform 1 0 127696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _528_
timestamp 1758069660
transform 1 0 113712 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _529_
timestamp 1758069660
transform 1 0 119692 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _530_
timestamp 1758069660
transform 1 0 117116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _531_
timestamp 1758069660
transform 1 0 117116 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _532_
timestamp 1758069660
transform 1 0 116196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _533_
timestamp 1758069660
transform 1 0 115276 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _534_
timestamp 1758069660
transform 1 0 116012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _535_
timestamp 1758069660
transform 1 0 114632 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _536_
timestamp 1758069660
transform 1 0 113804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _537_
timestamp 1758069660
transform 1 0 111872 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _538_
timestamp 1758069660
transform 1 0 113068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _539_
timestamp 1758069660
transform 1 0 102028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _540_
timestamp 1758069660
transform 1 0 104236 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp 1758069660
transform 1 0 102948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _542_
timestamp 1758069660
transform 1 0 102580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1758069660
transform 1 0 103500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _544_
timestamp 1758069660
transform 1 0 101476 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1758069660
transform 1 0 101660 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _546_
timestamp 1758069660
transform 1 0 100372 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1758069660
transform 1 0 100188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _548_
timestamp 1758069660
transform 1 0 97520 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1758069660
transform 1 0 99084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _550_
timestamp 1758069660
transform 1 0 90344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _551_
timestamp 1758069660
transform 1 0 89148 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1758069660
transform 1 0 88228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _553_
timestamp 1758069660
transform 1 0 87584 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1758069660
transform 1 0 87584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _555_
timestamp 1758069660
transform 1 0 86388 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _556_
timestamp 1758069660
transform 1 0 82892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _557_
timestamp 1758069660
transform 1 0 85652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1758069660
transform 1 0 86204 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _559_
timestamp 1758069660
transform 1 0 83996 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1758069660
transform 1 0 85008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _561_
timestamp 1758069660
transform 1 0 87676 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _562_
timestamp 1758069660
transform 1 0 81052 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp 1758069660
transform 1 0 79120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _564_
timestamp 1758069660
transform 1 0 77464 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 1758069660
transform 1 0 78200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _566_
timestamp 1758069660
transform 1 0 76268 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1758069660
transform 1 0 76912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _568_
timestamp 1758069660
transform 1 0 75532 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1758069660
transform 1 0 74888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _570_
timestamp 1758069660
transform 1 0 72036 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1758069660
transform 1 0 76452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _572_
timestamp 1758069660
transform 1 0 135332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _573_
timestamp 1758069660
transform 1 0 86940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 77740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1758069660
transform 1 0 77740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _576_
timestamp 1758069660
transform 1 0 78476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _577_
timestamp 1758069660
transform 1 0 79212 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _578_
timestamp 1758069660
transform 1 0 80132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _579_
timestamp 1758069660
transform 1 0 91724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1758069660
transform 1 0 86848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1758069660
transform 1 0 85468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _582_
timestamp 1758069660
transform 1 0 90068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1758069660
transform 1 0 88780 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1758069660
transform 1 0 88780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _585_
timestamp 1758069660
transform 1 0 101844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _586_
timestamp 1758069660
transform 1 0 99728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _587_
timestamp 1758069660
transform 1 0 100832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _588_
timestamp 1758069660
transform 1 0 105064 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _589_
timestamp 1758069660
transform 1 0 104420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _590_
timestamp 1758069660
transform 1 0 103776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _591_
timestamp 1758069660
transform 1 0 114540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _592_
timestamp 1758069660
transform 1 0 115276 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _593_
timestamp 1758069660
transform 1 0 113068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _594_
timestamp 1758069660
transform 1 0 118312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _595_
timestamp 1758069660
transform 1 0 116840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _596_
timestamp 1758069660
transform 1 0 117484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _597_
timestamp 1758069660
transform 1 0 127328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _598_
timestamp 1758069660
transform 1 0 129260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _599_
timestamp 1758069660
transform 1 0 130364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _600_
timestamp 1758069660
transform 1 0 131100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _601_
timestamp 1758069660
transform 1 0 132572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _602_
timestamp 1758069660
transform 1 0 130180 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _603_
timestamp 1758069660
transform 1 0 165232 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _604_
timestamp 1758069660
transform 1 0 159988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _605_
timestamp 1758069660
transform 1 0 148304 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _606_
timestamp 1758069660
transform 1 0 150604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _607_
timestamp 1758069660
transform 1 0 149868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _608_
timestamp 1758069660
transform 1 0 152444 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _609_
timestamp 1758069660
transform 1 0 152628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _610_
timestamp 1758069660
transform 1 0 166428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _611_
timestamp 1758069660
transform 1 0 162196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _612_
timestamp 1758069660
transform 1 0 162840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _613_
timestamp 1758069660
transform 1 0 163484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _614_
timestamp 1758069660
transform 1 0 164772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _615_
timestamp 1758069660
transform 1 0 164128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _616_
timestamp 1758069660
transform 1 0 177836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _617_
timestamp 1758069660
transform 1 0 177468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _618_
timestamp 1758069660
transform 1 0 178112 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _619_
timestamp 1758069660
transform 1 0 179952 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _620_
timestamp 1758069660
transform 1 0 181516 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _621_
timestamp 1758069660
transform 1 0 182160 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _622_
timestamp 1758069660
transform 1 0 188508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _623_
timestamp 1758069660
transform 1 0 187312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _624_
timestamp 1758069660
transform 1 0 190164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _625_
timestamp 1758069660
transform 1 0 194120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _626_
timestamp 1758069660
transform 1 0 192924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _627_
timestamp 1758069660
transform 1 0 196696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _628_
timestamp 1758069660
transform 1 0 192648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _629_
timestamp 1758069660
transform 1 0 202216 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1758069660
transform 1 0 202768 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _631_
timestamp 1758069660
transform 1 0 203412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _632_
timestamp 1758069660
transform 1 0 201020 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _633_
timestamp 1758069660
transform 1 0 200468 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _634_
timestamp 1758069660
transform 1 0 252632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _635_
timestamp 1758069660
transform 1 0 238004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _636_
timestamp 1758069660
transform 1 0 233036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _637_
timestamp 1758069660
transform 1 0 230276 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _638_
timestamp 1758069660
transform 1 0 230920 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _639_
timestamp 1758069660
transform 1 0 232116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _640_
timestamp 1758069660
transform 1 0 233036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _641_
timestamp 1758069660
transform 1 0 244444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _642_
timestamp 1758069660
transform 1 0 239844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _643_
timestamp 1758069660
transform 1 0 240764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _644_
timestamp 1758069660
transform 1 0 241684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _645_
timestamp 1758069660
transform 1 0 242052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _646_
timestamp 1758069660
transform 1 0 245180 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _647_
timestamp 1758069660
transform 1 0 251252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _648_
timestamp 1758069660
transform 1 0 252448 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _649_
timestamp 1758069660
transform 1 0 254840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _650_
timestamp 1758069660
transform 1 0 255484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _651_
timestamp 1758069660
transform 1 0 257048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _652_
timestamp 1758069660
transform 1 0 256220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _653_
timestamp 1758069660
transform 1 0 261648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _654_
timestamp 1758069660
transform 1 0 263948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _655_
timestamp 1758069660
transform 1 0 266432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _656_
timestamp 1758069660
transform 1 0 264316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _657_
timestamp 1758069660
transform 1 0 264868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _658_
timestamp 1758069660
transform 1 0 267076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _659_
timestamp 1758069660
transform 1 0 263120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _660_
timestamp 1758069660
transform 1 0 270940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _661_
timestamp 1758069660
transform 1 0 268364 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _662_
timestamp 1758069660
transform 1 0 269100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _663_
timestamp 1758069660
transform 1 0 267812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _664_
timestamp 1758069660
transform 1 0 271308 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _665_
timestamp 1758069660
transform 1 0 142968 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _666_
timestamp 1758069660
transform 1 0 149500 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _667_
timestamp 1758069660
transform 1 0 189520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _668_
timestamp 1758069660
transform 1 0 190808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _669_
timestamp 1758069660
transform 1 0 190072 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _670_
timestamp 1758069660
transform 1 0 190716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _671_
timestamp 1758069660
transform 1 0 156400 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _672_
timestamp 1758069660
transform 1 0 36432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _673_
timestamp 1758069660
transform 1 0 31556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _674_
timestamp 1758069660
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _675_
timestamp 1758069660
transform 1 0 33488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _676_
timestamp 1758069660
transform 1 0 32752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _677_
timestamp 1758069660
transform 1 0 32200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _678_
timestamp 1758069660
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _679_
timestamp 1758069660
transform 1 0 33488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _680_
timestamp 1758069660
transform 1 0 35328 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _681_
timestamp 1758069660
transform 1 0 34316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _682_
timestamp 1758069660
transform 1 0 33672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _683_
timestamp 1758069660
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _684_
timestamp 1758069660
transform 1 0 42780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _685_
timestamp 1758069660
transform 1 0 39100 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _686_
timestamp 1758069660
transform 1 0 40940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _687_
timestamp 1758069660
transform 1 0 41032 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _688_
timestamp 1758069660
transform 1 0 41676 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _689_
timestamp 1758069660
transform 1 0 42412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _690_
timestamp 1758069660
transform 1 0 55384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _691_
timestamp 1758069660
transform 1 0 52900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _692_
timestamp 1758069660
transform 1 0 54280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _693_
timestamp 1758069660
transform 1 0 54556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _694_
timestamp 1758069660
transform 1 0 56396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _695_
timestamp 1758069660
transform 1 0 57040 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 73600 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _697_
timestamp 1758069660
transform 1 0 75532 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _698_
timestamp 1758069660
transform 1 0 76176 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _699_
timestamp 1758069660
transform 1 0 78476 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _700_
timestamp 1758069660
transform 1 0 79764 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _701_
timestamp 1758069660
transform 1 0 83996 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _702_
timestamp 1758069660
transform 1 0 83904 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _703_
timestamp 1758069660
transform 1 0 86204 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _704_
timestamp 1758069660
transform 1 0 86480 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _705_
timestamp 1758069660
transform 1 0 88780 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _706_
timestamp 1758069660
transform 1 0 99176 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _707_
timestamp 1758069660
transform 1 0 99360 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _708_
timestamp 1758069660
transform 1 0 101384 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _709_
timestamp 1758069660
transform 1 0 101936 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _710_
timestamp 1758069660
transform 1 0 104236 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _711_
timestamp 1758069660
transform 1 0 112240 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _712_
timestamp 1758069660
transform 1 0 114356 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _713_
timestamp 1758069660
transform 1 0 114816 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _714_
timestamp 1758069660
transform 1 0 116472 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _715_
timestamp 1758069660
transform 1 0 117392 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _716_
timestamp 1758069660
transform 1 0 127512 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _717_
timestamp 1758069660
transform 1 0 129076 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _718_
timestamp 1758069660
transform 1 0 130272 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _719_
timestamp 1758069660
transform 1 0 130824 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _720_
timestamp 1758069660
transform 1 0 132572 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _721_
timestamp 1758069660
transform 1 0 145728 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _722_
timestamp 1758069660
transform 1 0 147476 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _723_
timestamp 1758069660
transform 1 0 148304 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _724_
timestamp 1758069660
transform 1 0 150880 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _725_
timestamp 1758069660
transform 1 0 153456 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _726_
timestamp 1758069660
transform 1 0 158608 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _727_
timestamp 1758069660
transform 1 0 160908 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _728_
timestamp 1758069660
transform 1 0 161828 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _729_
timestamp 1758069660
transform 1 0 163484 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _730_
timestamp 1758069660
transform 1 0 163576 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _731_
timestamp 1758069660
transform 1 0 176364 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _732_
timestamp 1758069660
transform 1 0 176364 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _733_
timestamp 1758069660
transform 1 0 178940 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _734_
timestamp 1758069660
transform 1 0 178572 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _735_
timestamp 1758069660
transform 1 0 179124 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _736_
timestamp 1758069660
transform 1 0 189520 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _737_
timestamp 1758069660
transform 1 0 190808 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _738_
timestamp 1758069660
transform 1 0 191820 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _739_
timestamp 1758069660
transform 1 0 192004 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _740_
timestamp 1758069660
transform 1 0 194028 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _741_
timestamp 1758069660
transform 1 0 202124 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _742_
timestamp 1758069660
transform 1 0 202584 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _743_
timestamp 1758069660
transform 1 0 204700 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _744_
timestamp 1758069660
transform 1 0 204792 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _745_
timestamp 1758069660
transform 1 0 204700 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _746_
timestamp 1758069660
transform 1 0 227884 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _747_
timestamp 1758069660
transform 1 0 227884 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _748_
timestamp 1758069660
transform 1 0 227516 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _749_
timestamp 1758069660
transform 1 0 230460 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _750_
timestamp 1758069660
transform 1 0 230736 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _751_
timestamp 1758069660
transform 1 0 238188 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _752_
timestamp 1758069660
transform 1 0 238464 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _753_
timestamp 1758069660
transform 1 0 240764 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _754_
timestamp 1758069660
transform 1 0 240672 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _755_
timestamp 1758069660
transform 1 0 243340 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _756_
timestamp 1758069660
transform 1 0 251068 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _757_
timestamp 1758069660
transform 1 0 253644 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _758_
timestamp 1758069660
transform 1 0 252540 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _759_
timestamp 1758069660
transform 1 0 253644 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _760_
timestamp 1758069660
transform 1 0 256220 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _761_
timestamp 1758069660
transform 1 0 264224 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _762_
timestamp 1758069660
transform 1 0 265236 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _763_
timestamp 1758069660
transform 1 0 265604 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _764_
timestamp 1758069660
transform 1 0 266524 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _765_
timestamp 1758069660
transform 1 0 269100 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _766_
timestamp 1758069660
transform 1 0 269100 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _767_
timestamp 1758069660
transform 1 0 268732 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _768_
timestamp 1758069660
transform 1 0 271676 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _769_
timestamp 1758069660
transform 1 0 269100 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 266524 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _771_
timestamp 1758069660
transform 1 0 194396 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _772_
timestamp 1758069660
transform 1 0 194396 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _773_
timestamp 1758069660
transform 1 0 191820 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _774_
timestamp 1758069660
transform 1 0 193016 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _775_
timestamp 1758069660
transform 1 0 148028 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _776_
timestamp 1758069660
transform 1 0 29624 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _777_
timestamp 1758069660
transform 1 0 27232 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _778_
timestamp 1758069660
transform 1 0 29624 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _779_
timestamp 1758069660
transform 1 0 29532 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _780_
timestamp 1758069660
transform 1 0 29808 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _781_
timestamp 1758069660
transform 1 0 29808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _782_
timestamp 1758069660
transform 1 0 31740 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _783_
timestamp 1758069660
transform 1 0 32108 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _784_
timestamp 1758069660
transform 1 0 32384 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _785_
timestamp 1758069660
transform 1 0 34684 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _786_
timestamp 1758069660
transform 1 0 37536 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _787_
timestamp 1758069660
transform 1 0 39468 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _788_
timestamp 1758069660
transform 1 0 40112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _789_
timestamp 1758069660
transform 1 0 41400 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _790_
timestamp 1758069660
transform 1 0 42504 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _791_
timestamp 1758069660
transform 1 0 52348 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _792_
timestamp 1758069660
transform 1 0 52992 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _793_
timestamp 1758069660
transform 1 0 54740 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _794_
timestamp 1758069660
transform 1 0 55568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _795_
timestamp 1758069660
transform 1 0 57868 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  _796_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 187128 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform -1 0 43516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1758069660
transform 1 0 55936 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1758069660
transform 1 0 154100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1758069660
transform 1 0 153732 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1758069660
transform 1 0 155940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1758069660
transform 1 0 153364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1758069660
transform 1 0 156308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1758069660
transform 1 0 152996 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1758069660
transform 1 0 156676 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1758069660
transform 1 0 152628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1758069660
transform 1 0 157044 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1758069660
transform 1 0 152260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1758069660
transform -1 0 303508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1758069660
transform -1 0 303140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1758069660
transform -1 0 302312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1758069660
transform -1 0 301944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1758069660
transform -1 0 301576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1758069660
transform 1 0 305348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1758069660
transform 1 0 304888 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1758069660
transform 1 0 305348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1758069660
transform 1 0 304888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1758069660
transform 1 0 305348 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1758069660
transform 1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1758069660
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1758069660
transform 1 0 2576 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1758069660
transform 1 0 2944 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1758069660
transform 1 0 268456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1758069660
transform 1 0 252264 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1758069660
transform 1 0 197984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1758069660
transform 1 0 197800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1758069660
transform 1 0 295872 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 149408 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1758069660
transform 1 0 140668 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1758069660
transform 1 0 140392 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1758069660
transform 1 0 140392 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1758069660
transform 1 0 140668 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1758069660
transform 1 0 156124 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1758069660
transform 1 0 156032 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1758069660
transform 1 0 156032 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1758069660
transform 1 0 156124 0 -1 9792
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1758069660
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1758069660
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1758069660
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1758069660
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1758069660
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1758069660
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1758069660
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1758069660
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1758069660
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1758069660
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1758069660
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1758069660
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1758069660
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1758069660
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1758069660
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1758069660
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1758069660
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1758069660
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1758069660
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1758069660
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1758069660
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1758069660
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1758069660
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1758069660
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1758069660
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1758069660
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1758069660
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1758069660
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1758069660
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1758069660
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1758069660
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1758069660
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1758069660
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1758069660
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1758069660
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1758069660
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1758069660
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1758069660
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1758069660
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1758069660
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1758069660
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1758069660
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1758069660
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1758069660
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1758069660
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1758069660
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1758069660
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1758069660
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1758069660
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1758069660
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1758069660
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1758069660
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1758069660
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1758069660
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1758069660
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1758069660
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1758069660
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1758069660
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1758069660
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1758069660
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1758069660
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1758069660
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1758069660
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1758069660
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1758069660
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1758069660
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1758069660
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1758069660
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1758069660
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1758069660
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1758069660
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1758069660
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1758069660
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1758069660
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1758069660
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1758069660
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1758069660
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1758069660
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1758069660
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1758069660
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1758069660
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1758069660
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1758069660
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1758069660
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1758069660
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1758069660
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1758069660
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1758069660
transform 1 0 78476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1758069660
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1758069660
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1758069660
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1758069660
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1758069660
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1758069660
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1758069660
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1758069660
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1758069660
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1758069660
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1758069660
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1758069660
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1758069660
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1758069660
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1758069660
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1758069660
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1758069660
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1758069660
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1758069660
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1758069660
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1758069660
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1758069660
transform 1 0 97612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1758069660
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1758069660
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1758069660
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1758069660
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1758069660
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1758069660
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1758069660
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1758069660
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1758069660
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1758069660
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1758069660
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1161
timestamp 1758069660
transform 1 0 107916 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1173
timestamp 1758069660
transform 1 0 109020 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1177
timestamp 1758069660
transform 1 0 109388 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1189
timestamp 1758069660
transform 1 0 110492 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1201
timestamp 1758069660
transform 1 0 111596 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1205
timestamp 1758069660
transform 1 0 111964 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1217
timestamp 1758069660
transform 1 0 113068 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1229
timestamp 1758069660
transform 1 0 114172 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1233
timestamp 1758069660
transform 1 0 114540 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1245
timestamp 1758069660
transform 1 0 115644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1257
timestamp 1758069660
transform 1 0 116748 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1261
timestamp 1758069660
transform 1 0 117116 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1273
timestamp 1758069660
transform 1 0 118220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1285
timestamp 1758069660
transform 1 0 119324 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1289
timestamp 1758069660
transform 1 0 119692 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1301
timestamp 1758069660
transform 1 0 120796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1313
timestamp 1758069660
transform 1 0 121900 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1317
timestamp 1758069660
transform 1 0 122268 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1329
timestamp 1758069660
transform 1 0 123372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1341
timestamp 1758069660
transform 1 0 124476 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1345
timestamp 1758069660
transform 1 0 124844 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1357
timestamp 1758069660
transform 1 0 125948 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1369
timestamp 1758069660
transform 1 0 127052 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1373
timestamp 1758069660
transform 1 0 127420 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1385
timestamp 1758069660
transform 1 0 128524 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1397
timestamp 1758069660
transform 1 0 129628 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1401
timestamp 1758069660
transform 1 0 129996 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1413
timestamp 1758069660
transform 1 0 131100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1425
timestamp 1758069660
transform 1 0 132204 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1429
timestamp 1758069660
transform 1 0 132572 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1441
timestamp 1758069660
transform 1 0 133676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1453
timestamp 1758069660
transform 1 0 134780 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1457
timestamp 1758069660
transform 1 0 135148 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1469
timestamp 1758069660
transform 1 0 136252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1481
timestamp 1758069660
transform 1 0 137356 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1485
timestamp 1758069660
transform 1 0 137724 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1497
timestamp 1758069660
transform 1 0 138828 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1509
timestamp 1758069660
transform 1 0 139932 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1513
timestamp 1758069660
transform 1 0 140300 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1525
timestamp 1758069660
transform 1 0 141404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1537
timestamp 1758069660
transform 1 0 142508 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1541
timestamp 1758069660
transform 1 0 142876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1553
timestamp 1758069660
transform 1 0 143980 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1565
timestamp 1758069660
transform 1 0 145084 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1569
timestamp 1758069660
transform 1 0 145452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1581
timestamp 1758069660
transform 1 0 146556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1593
timestamp 1758069660
transform 1 0 147660 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1597
timestamp 1758069660
transform 1 0 148028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1609
timestamp 1758069660
transform 1 0 149132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1621
timestamp 1758069660
transform 1 0 150236 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1625
timestamp 1758069660
transform 1 0 150604 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1637
timestamp 1758069660
transform 1 0 151708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1649
timestamp 1758069660
transform 1 0 152812 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1653
timestamp 1758069660
transform 1 0 153180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1665
timestamp 1758069660
transform 1 0 154284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1677
timestamp 1758069660
transform 1 0 155388 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1681
timestamp 1758069660
transform 1 0 155756 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1693
timestamp 1758069660
transform 1 0 156860 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1705
timestamp 1758069660
transform 1 0 157964 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1709
timestamp 1758069660
transform 1 0 158332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1721
timestamp 1758069660
transform 1 0 159436 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1733
timestamp 1758069660
transform 1 0 160540 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1737
timestamp 1758069660
transform 1 0 160908 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1749
timestamp 1758069660
transform 1 0 162012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1761
timestamp 1758069660
transform 1 0 163116 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1765
timestamp 1758069660
transform 1 0 163484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1777
timestamp 1758069660
transform 1 0 164588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1789
timestamp 1758069660
transform 1 0 165692 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1793
timestamp 1758069660
transform 1 0 166060 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1805
timestamp 1758069660
transform 1 0 167164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1817
timestamp 1758069660
transform 1 0 168268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1821
timestamp 1758069660
transform 1 0 168636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1833
timestamp 1758069660
transform 1 0 169740 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1845
timestamp 1758069660
transform 1 0 170844 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1849
timestamp 1758069660
transform 1 0 171212 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1861
timestamp 1758069660
transform 1 0 172316 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1873
timestamp 1758069660
transform 1 0 173420 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1877
timestamp 1758069660
transform 1 0 173788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1889
timestamp 1758069660
transform 1 0 174892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1901
timestamp 1758069660
transform 1 0 175996 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1905
timestamp 1758069660
transform 1 0 176364 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1917
timestamp 1758069660
transform 1 0 177468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1929
timestamp 1758069660
transform 1 0 178572 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1933
timestamp 1758069660
transform 1 0 178940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1945
timestamp 1758069660
transform 1 0 180044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1957
timestamp 1758069660
transform 1 0 181148 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1961
timestamp 1758069660
transform 1 0 181516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1973
timestamp 1758069660
transform 1 0 182620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1985
timestamp 1758069660
transform 1 0 183724 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1989
timestamp 1758069660
transform 1 0 184092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2001
timestamp 1758069660
transform 1 0 185196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2013
timestamp 1758069660
transform 1 0 186300 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2017
timestamp 1758069660
transform 1 0 186668 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2029
timestamp 1758069660
transform 1 0 187772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2041
timestamp 1758069660
transform 1 0 188876 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2045
timestamp 1758069660
transform 1 0 189244 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2057
timestamp 1758069660
transform 1 0 190348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2069
timestamp 1758069660
transform 1 0 191452 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2073
timestamp 1758069660
transform 1 0 191820 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2085
timestamp 1758069660
transform 1 0 192924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2097
timestamp 1758069660
transform 1 0 194028 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2101
timestamp 1758069660
transform 1 0 194396 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2113
timestamp 1758069660
transform 1 0 195500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2125
timestamp 1758069660
transform 1 0 196604 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2129
timestamp 1758069660
transform 1 0 196972 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2141
timestamp 1758069660
transform 1 0 198076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2153
timestamp 1758069660
transform 1 0 199180 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2157
timestamp 1758069660
transform 1 0 199548 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2169
timestamp 1758069660
transform 1 0 200652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2181
timestamp 1758069660
transform 1 0 201756 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2185
timestamp 1758069660
transform 1 0 202124 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2197
timestamp 1758069660
transform 1 0 203228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2209
timestamp 1758069660
transform 1 0 204332 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2213
timestamp 1758069660
transform 1 0 204700 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2225
timestamp 1758069660
transform 1 0 205804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2237
timestamp 1758069660
transform 1 0 206908 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2241
timestamp 1758069660
transform 1 0 207276 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2253
timestamp 1758069660
transform 1 0 208380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2265
timestamp 1758069660
transform 1 0 209484 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2269
timestamp 1758069660
transform 1 0 209852 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2281
timestamp 1758069660
transform 1 0 210956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2293
timestamp 1758069660
transform 1 0 212060 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2297
timestamp 1758069660
transform 1 0 212428 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2309
timestamp 1758069660
transform 1 0 213532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2321
timestamp 1758069660
transform 1 0 214636 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2325
timestamp 1758069660
transform 1 0 215004 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2337
timestamp 1758069660
transform 1 0 216108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2349
timestamp 1758069660
transform 1 0 217212 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2353
timestamp 1758069660
transform 1 0 217580 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2365
timestamp 1758069660
transform 1 0 218684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2377
timestamp 1758069660
transform 1 0 219788 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2381
timestamp 1758069660
transform 1 0 220156 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2393
timestamp 1758069660
transform 1 0 221260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2405
timestamp 1758069660
transform 1 0 222364 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2409
timestamp 1758069660
transform 1 0 222732 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2421
timestamp 1758069660
transform 1 0 223836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2433
timestamp 1758069660
transform 1 0 224940 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2437
timestamp 1758069660
transform 1 0 225308 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2449
timestamp 1758069660
transform 1 0 226412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2461
timestamp 1758069660
transform 1 0 227516 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2465
timestamp 1758069660
transform 1 0 227884 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2477
timestamp 1758069660
transform 1 0 228988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2489
timestamp 1758069660
transform 1 0 230092 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2493
timestamp 1758069660
transform 1 0 230460 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2505
timestamp 1758069660
transform 1 0 231564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2517
timestamp 1758069660
transform 1 0 232668 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2521
timestamp 1758069660
transform 1 0 233036 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2533
timestamp 1758069660
transform 1 0 234140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2545
timestamp 1758069660
transform 1 0 235244 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2549
timestamp 1758069660
transform 1 0 235612 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2561
timestamp 1758069660
transform 1 0 236716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2573
timestamp 1758069660
transform 1 0 237820 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2577
timestamp 1758069660
transform 1 0 238188 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2589
timestamp 1758069660
transform 1 0 239292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2601
timestamp 1758069660
transform 1 0 240396 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2605
timestamp 1758069660
transform 1 0 240764 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2617
timestamp 1758069660
transform 1 0 241868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2629
timestamp 1758069660
transform 1 0 242972 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2633
timestamp 1758069660
transform 1 0 243340 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2645
timestamp 1758069660
transform 1 0 244444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2657
timestamp 1758069660
transform 1 0 245548 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2661
timestamp 1758069660
transform 1 0 245916 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2673
timestamp 1758069660
transform 1 0 247020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2685
timestamp 1758069660
transform 1 0 248124 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2689
timestamp 1758069660
transform 1 0 248492 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2701
timestamp 1758069660
transform 1 0 249596 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2713
timestamp 1758069660
transform 1 0 250700 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2717
timestamp 1758069660
transform 1 0 251068 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2729
timestamp 1758069660
transform 1 0 252172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2741
timestamp 1758069660
transform 1 0 253276 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2745
timestamp 1758069660
transform 1 0 253644 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2757
timestamp 1758069660
transform 1 0 254748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2769
timestamp 1758069660
transform 1 0 255852 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2773
timestamp 1758069660
transform 1 0 256220 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2785
timestamp 1758069660
transform 1 0 257324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2797
timestamp 1758069660
transform 1 0 258428 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2801
timestamp 1758069660
transform 1 0 258796 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2813
timestamp 1758069660
transform 1 0 259900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2825
timestamp 1758069660
transform 1 0 261004 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2829
timestamp 1758069660
transform 1 0 261372 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2841
timestamp 1758069660
transform 1 0 262476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2853
timestamp 1758069660
transform 1 0 263580 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2857
timestamp 1758069660
transform 1 0 263948 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2869
timestamp 1758069660
transform 1 0 265052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2881
timestamp 1758069660
transform 1 0 266156 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2885
timestamp 1758069660
transform 1 0 266524 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2897
timestamp 1758069660
transform 1 0 267628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2909
timestamp 1758069660
transform 1 0 268732 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2913
timestamp 1758069660
transform 1 0 269100 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2925
timestamp 1758069660
transform 1 0 270204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2937
timestamp 1758069660
transform 1 0 271308 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2941
timestamp 1758069660
transform 1 0 271676 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2953
timestamp 1758069660
transform 1 0 272780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2965
timestamp 1758069660
transform 1 0 273884 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2969
timestamp 1758069660
transform 1 0 274252 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2981
timestamp 1758069660
transform 1 0 275356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2993
timestamp 1758069660
transform 1 0 276460 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2997
timestamp 1758069660
transform 1 0 276828 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3009
timestamp 1758069660
transform 1 0 277932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3021
timestamp 1758069660
transform 1 0 279036 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3025
timestamp 1758069660
transform 1 0 279404 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3037
timestamp 1758069660
transform 1 0 280508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3049
timestamp 1758069660
transform 1 0 281612 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3053
timestamp 1758069660
transform 1 0 281980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3065
timestamp 1758069660
transform 1 0 283084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3077
timestamp 1758069660
transform 1 0 284188 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3081
timestamp 1758069660
transform 1 0 284556 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3093
timestamp 1758069660
transform 1 0 285660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3105
timestamp 1758069660
transform 1 0 286764 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3109
timestamp 1758069660
transform 1 0 287132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3121
timestamp 1758069660
transform 1 0 288236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3133
timestamp 1758069660
transform 1 0 289340 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3137
timestamp 1758069660
transform 1 0 289708 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3149
timestamp 1758069660
transform 1 0 290812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3161
timestamp 1758069660
transform 1 0 291916 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3165
timestamp 1758069660
transform 1 0 292284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3177
timestamp 1758069660
transform 1 0 293388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3189
timestamp 1758069660
transform 1 0 294492 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3193
timestamp 1758069660
transform 1 0 294860 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3205
timestamp 1758069660
transform 1 0 295964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3217
timestamp 1758069660
transform 1 0 297068 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3221
timestamp 1758069660
transform 1 0 297436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3233
timestamp 1758069660
transform 1 0 298540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3245
timestamp 1758069660
transform 1 0 299644 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3249
timestamp 1758069660
transform 1 0 300012 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3261
timestamp 1758069660
transform 1 0 301116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3273
timestamp 1758069660
transform 1 0 302220 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3277
timestamp 1758069660
transform 1 0 302588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3289
timestamp 1758069660
transform 1 0 303692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3301
timestamp 1758069660
transform 1 0 304796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3305 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 305164 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1758069660
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1758069660
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1758069660
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1758069660
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1758069660
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1758069660
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1758069660
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1758069660
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1758069660
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1758069660
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1758069660
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1758069660
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1758069660
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1758069660
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1758069660
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1758069660
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1758069660
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1758069660
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1758069660
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1758069660
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1758069660
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1758069660
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1758069660
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1758069660
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1758069660
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1758069660
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1758069660
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1758069660
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1758069660
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1758069660
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1758069660
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1758069660
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1758069660
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1758069660
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1758069660
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1758069660
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1758069660
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1758069660
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1758069660
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1758069660
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1758069660
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1758069660
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1758069660
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1758069660
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1758069660
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1758069660
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1758069660
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1758069660
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1758069660
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1758069660
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1758069660
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1758069660
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1758069660
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1758069660
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1758069660
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1758069660
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1758069660
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1758069660
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1758069660
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1758069660
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1758069660
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1758069660
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1758069660
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1758069660
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1758069660
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1758069660
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1758069660
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1758069660
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1758069660
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1758069660
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1758069660
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1758069660
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1758069660
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1758069660
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1758069660
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1758069660
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1758069660
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1758069660
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1758069660
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1758069660
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1758069660
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1758069660
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1758069660
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1758069660
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1758069660
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1758069660
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1758069660
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1758069660
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1758069660
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1758069660
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1758069660
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1758069660
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1758069660
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 1758069660
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1758069660
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1758069660
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1758069660
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1758069660
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1758069660
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1758069660
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1758069660
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1758069660
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1758069660
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1758069660
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1758069660
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1758069660
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1758069660
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1758069660
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1758069660
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1758069660
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1758069660
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1758069660
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1758069660
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1758069660
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1758069660
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1758069660
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1758069660
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1758069660
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1758069660
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1758069660
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1758069660
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1758069660
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1157
timestamp 1758069660
transform 1 0 107548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1758069660
transform 1 0 108652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1758069660
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1177
timestamp 1758069660
transform 1 0 109388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1189
timestamp 1758069660
transform 1 0 110492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1201
timestamp 1758069660
transform 1 0 111596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1213
timestamp 1758069660
transform 1 0 112700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1225
timestamp 1758069660
transform 1 0 113804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1758069660
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1233
timestamp 1758069660
transform 1 0 114540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1245
timestamp 1758069660
transform 1 0 115644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1257
timestamp 1758069660
transform 1 0 116748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1269
timestamp 1758069660
transform 1 0 117852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1281
timestamp 1758069660
transform 1 0 118956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1287
timestamp 1758069660
transform 1 0 119508 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1289
timestamp 1758069660
transform 1 0 119692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1301
timestamp 1758069660
transform 1 0 120796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1313
timestamp 1758069660
transform 1 0 121900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1325
timestamp 1758069660
transform 1 0 123004 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1337
timestamp 1758069660
transform 1 0 124108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1343
timestamp 1758069660
transform 1 0 124660 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1345
timestamp 1758069660
transform 1 0 124844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1357
timestamp 1758069660
transform 1 0 125948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1369
timestamp 1758069660
transform 1 0 127052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1381
timestamp 1758069660
transform 1 0 128156 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1393
timestamp 1758069660
transform 1 0 129260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1399
timestamp 1758069660
transform 1 0 129812 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1401
timestamp 1758069660
transform 1 0 129996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1413
timestamp 1758069660
transform 1 0 131100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1425
timestamp 1758069660
transform 1 0 132204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1437
timestamp 1758069660
transform 1 0 133308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1449
timestamp 1758069660
transform 1 0 134412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1455
timestamp 1758069660
transform 1 0 134964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1457
timestamp 1758069660
transform 1 0 135148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1469
timestamp 1758069660
transform 1 0 136252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1481
timestamp 1758069660
transform 1 0 137356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1493
timestamp 1758069660
transform 1 0 138460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1505
timestamp 1758069660
transform 1 0 139564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1511
timestamp 1758069660
transform 1 0 140116 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1513
timestamp 1758069660
transform 1 0 140300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1525
timestamp 1758069660
transform 1 0 141404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1537
timestamp 1758069660
transform 1 0 142508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1549
timestamp 1758069660
transform 1 0 143612 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1561
timestamp 1758069660
transform 1 0 144716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1567
timestamp 1758069660
transform 1 0 145268 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1569
timestamp 1758069660
transform 1 0 145452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1581
timestamp 1758069660
transform 1 0 146556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1593
timestamp 1758069660
transform 1 0 147660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1605
timestamp 1758069660
transform 1 0 148764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1617
timestamp 1758069660
transform 1 0 149868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1623
timestamp 1758069660
transform 1 0 150420 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1625
timestamp 1758069660
transform 1 0 150604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1637
timestamp 1758069660
transform 1 0 151708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1649
timestamp 1758069660
transform 1 0 152812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1661
timestamp 1758069660
transform 1 0 153916 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1673
timestamp 1758069660
transform 1 0 155020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1679
timestamp 1758069660
transform 1 0 155572 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1681
timestamp 1758069660
transform 1 0 155756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1693
timestamp 1758069660
transform 1 0 156860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1705
timestamp 1758069660
transform 1 0 157964 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1717
timestamp 1758069660
transform 1 0 159068 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1729
timestamp 1758069660
transform 1 0 160172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1735
timestamp 1758069660
transform 1 0 160724 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1737
timestamp 1758069660
transform 1 0 160908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1749
timestamp 1758069660
transform 1 0 162012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1761
timestamp 1758069660
transform 1 0 163116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1773
timestamp 1758069660
transform 1 0 164220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1785
timestamp 1758069660
transform 1 0 165324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1791
timestamp 1758069660
transform 1 0 165876 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1793
timestamp 1758069660
transform 1 0 166060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1805
timestamp 1758069660
transform 1 0 167164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1817
timestamp 1758069660
transform 1 0 168268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1829
timestamp 1758069660
transform 1 0 169372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1841
timestamp 1758069660
transform 1 0 170476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1847
timestamp 1758069660
transform 1 0 171028 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1849
timestamp 1758069660
transform 1 0 171212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1861
timestamp 1758069660
transform 1 0 172316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1873
timestamp 1758069660
transform 1 0 173420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1885
timestamp 1758069660
transform 1 0 174524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1897
timestamp 1758069660
transform 1 0 175628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1903
timestamp 1758069660
transform 1 0 176180 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1905
timestamp 1758069660
transform 1 0 176364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1917
timestamp 1758069660
transform 1 0 177468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1929
timestamp 1758069660
transform 1 0 178572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1941
timestamp 1758069660
transform 1 0 179676 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1953
timestamp 1758069660
transform 1 0 180780 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1959
timestamp 1758069660
transform 1 0 181332 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1961
timestamp 1758069660
transform 1 0 181516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1973
timestamp 1758069660
transform 1 0 182620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1985
timestamp 1758069660
transform 1 0 183724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1997
timestamp 1758069660
transform 1 0 184828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2009
timestamp 1758069660
transform 1 0 185932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2015
timestamp 1758069660
transform 1 0 186484 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2017
timestamp 1758069660
transform 1 0 186668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2029
timestamp 1758069660
transform 1 0 187772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2041
timestamp 1758069660
transform 1 0 188876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2053
timestamp 1758069660
transform 1 0 189980 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2065
timestamp 1758069660
transform 1 0 191084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2071
timestamp 1758069660
transform 1 0 191636 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2073
timestamp 1758069660
transform 1 0 191820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2085
timestamp 1758069660
transform 1 0 192924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2097
timestamp 1758069660
transform 1 0 194028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2109
timestamp 1758069660
transform 1 0 195132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2121
timestamp 1758069660
transform 1 0 196236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2127
timestamp 1758069660
transform 1 0 196788 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2129
timestamp 1758069660
transform 1 0 196972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2141
timestamp 1758069660
transform 1 0 198076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2153
timestamp 1758069660
transform 1 0 199180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2165
timestamp 1758069660
transform 1 0 200284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2177
timestamp 1758069660
transform 1 0 201388 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2183
timestamp 1758069660
transform 1 0 201940 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2185
timestamp 1758069660
transform 1 0 202124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2197
timestamp 1758069660
transform 1 0 203228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2209
timestamp 1758069660
transform 1 0 204332 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2221
timestamp 1758069660
transform 1 0 205436 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2233
timestamp 1758069660
transform 1 0 206540 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2239
timestamp 1758069660
transform 1 0 207092 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2241
timestamp 1758069660
transform 1 0 207276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2253
timestamp 1758069660
transform 1 0 208380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2265
timestamp 1758069660
transform 1 0 209484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2277
timestamp 1758069660
transform 1 0 210588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2289
timestamp 1758069660
transform 1 0 211692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2295
timestamp 1758069660
transform 1 0 212244 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2297
timestamp 1758069660
transform 1 0 212428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2309
timestamp 1758069660
transform 1 0 213532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2321
timestamp 1758069660
transform 1 0 214636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2333
timestamp 1758069660
transform 1 0 215740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2345
timestamp 1758069660
transform 1 0 216844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2351
timestamp 1758069660
transform 1 0 217396 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2353
timestamp 1758069660
transform 1 0 217580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2365
timestamp 1758069660
transform 1 0 218684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2377
timestamp 1758069660
transform 1 0 219788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2389
timestamp 1758069660
transform 1 0 220892 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2401
timestamp 1758069660
transform 1 0 221996 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2407
timestamp 1758069660
transform 1 0 222548 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2409
timestamp 1758069660
transform 1 0 222732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2421
timestamp 1758069660
transform 1 0 223836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2433
timestamp 1758069660
transform 1 0 224940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2445
timestamp 1758069660
transform 1 0 226044 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2457
timestamp 1758069660
transform 1 0 227148 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2463
timestamp 1758069660
transform 1 0 227700 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2465
timestamp 1758069660
transform 1 0 227884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2477
timestamp 1758069660
transform 1 0 228988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2489
timestamp 1758069660
transform 1 0 230092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2501
timestamp 1758069660
transform 1 0 231196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2513
timestamp 1758069660
transform 1 0 232300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2519
timestamp 1758069660
transform 1 0 232852 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2521
timestamp 1758069660
transform 1 0 233036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2533
timestamp 1758069660
transform 1 0 234140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2545
timestamp 1758069660
transform 1 0 235244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2557
timestamp 1758069660
transform 1 0 236348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2569
timestamp 1758069660
transform 1 0 237452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2575
timestamp 1758069660
transform 1 0 238004 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2577
timestamp 1758069660
transform 1 0 238188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2589
timestamp 1758069660
transform 1 0 239292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2601
timestamp 1758069660
transform 1 0 240396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2613
timestamp 1758069660
transform 1 0 241500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2625
timestamp 1758069660
transform 1 0 242604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2631
timestamp 1758069660
transform 1 0 243156 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2633
timestamp 1758069660
transform 1 0 243340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2645
timestamp 1758069660
transform 1 0 244444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2657
timestamp 1758069660
transform 1 0 245548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2669
timestamp 1758069660
transform 1 0 246652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2681
timestamp 1758069660
transform 1 0 247756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2687
timestamp 1758069660
transform 1 0 248308 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2689
timestamp 1758069660
transform 1 0 248492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2701
timestamp 1758069660
transform 1 0 249596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2713
timestamp 1758069660
transform 1 0 250700 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2725
timestamp 1758069660
transform 1 0 251804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2737
timestamp 1758069660
transform 1 0 252908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2743
timestamp 1758069660
transform 1 0 253460 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2745
timestamp 1758069660
transform 1 0 253644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2757
timestamp 1758069660
transform 1 0 254748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2769
timestamp 1758069660
transform 1 0 255852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2781
timestamp 1758069660
transform 1 0 256956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2793
timestamp 1758069660
transform 1 0 258060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2799
timestamp 1758069660
transform 1 0 258612 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2801
timestamp 1758069660
transform 1 0 258796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2813
timestamp 1758069660
transform 1 0 259900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2825
timestamp 1758069660
transform 1 0 261004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2837
timestamp 1758069660
transform 1 0 262108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2849
timestamp 1758069660
transform 1 0 263212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2855
timestamp 1758069660
transform 1 0 263764 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2857
timestamp 1758069660
transform 1 0 263948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2869
timestamp 1758069660
transform 1 0 265052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2881
timestamp 1758069660
transform 1 0 266156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2893
timestamp 1758069660
transform 1 0 267260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2905
timestamp 1758069660
transform 1 0 268364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2911
timestamp 1758069660
transform 1 0 268916 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2913
timestamp 1758069660
transform 1 0 269100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2925
timestamp 1758069660
transform 1 0 270204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2937
timestamp 1758069660
transform 1 0 271308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2949
timestamp 1758069660
transform 1 0 272412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2961
timestamp 1758069660
transform 1 0 273516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2967
timestamp 1758069660
transform 1 0 274068 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2969
timestamp 1758069660
transform 1 0 274252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2981
timestamp 1758069660
transform 1 0 275356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2993
timestamp 1758069660
transform 1 0 276460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3005
timestamp 1758069660
transform 1 0 277564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3017
timestamp 1758069660
transform 1 0 278668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3023
timestamp 1758069660
transform 1 0 279220 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3025
timestamp 1758069660
transform 1 0 279404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3037
timestamp 1758069660
transform 1 0 280508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3049
timestamp 1758069660
transform 1 0 281612 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3061
timestamp 1758069660
transform 1 0 282716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3073
timestamp 1758069660
transform 1 0 283820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3079
timestamp 1758069660
transform 1 0 284372 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3081
timestamp 1758069660
transform 1 0 284556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3093
timestamp 1758069660
transform 1 0 285660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3105
timestamp 1758069660
transform 1 0 286764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3117
timestamp 1758069660
transform 1 0 287868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3129
timestamp 1758069660
transform 1 0 288972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3135
timestamp 1758069660
transform 1 0 289524 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3137
timestamp 1758069660
transform 1 0 289708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3149
timestamp 1758069660
transform 1 0 290812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3161
timestamp 1758069660
transform 1 0 291916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3173
timestamp 1758069660
transform 1 0 293020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3185
timestamp 1758069660
transform 1 0 294124 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3191
timestamp 1758069660
transform 1 0 294676 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3193
timestamp 1758069660
transform 1 0 294860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3205
timestamp 1758069660
transform 1 0 295964 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3217
timestamp 1758069660
transform 1 0 297068 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3229
timestamp 1758069660
transform 1 0 298172 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3241
timestamp 1758069660
transform 1 0 299276 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3247
timestamp 1758069660
transform 1 0 299828 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3249
timestamp 1758069660
transform 1 0 300012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3261
timestamp 1758069660
transform 1 0 301116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3273
timestamp 1758069660
transform 1 0 302220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3285
timestamp 1758069660
transform 1 0 303324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3297
timestamp 1758069660
transform 1 0 304428 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3303
timestamp 1758069660
transform 1 0 304980 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3305
timestamp 1758069660
transform 1 0 305164 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1758069660
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1758069660
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1758069660
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1758069660
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1758069660
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1758069660
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1758069660
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1758069660
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1758069660
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1758069660
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1758069660
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1758069660
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1758069660
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1758069660
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1758069660
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1758069660
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1758069660
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1758069660
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1758069660
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1758069660
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1758069660
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1758069660
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1758069660
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1758069660
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1758069660
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1758069660
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1758069660
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1758069660
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1758069660
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1758069660
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1758069660
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1758069660
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1758069660
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1758069660
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1758069660
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1758069660
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1758069660
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1758069660
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1758069660
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1758069660
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1758069660
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1758069660
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1758069660
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1758069660
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1758069660
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1758069660
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1758069660
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1758069660
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1758069660
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1758069660
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1758069660
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1758069660
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1758069660
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1758069660
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1758069660
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1758069660
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1758069660
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1758069660
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1758069660
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1758069660
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1758069660
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1758069660
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1758069660
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1758069660
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1758069660
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1758069660
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1758069660
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1758069660
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1758069660
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1758069660
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1758069660
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1758069660
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1758069660
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1758069660
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1758069660
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1758069660
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1758069660
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1758069660
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1758069660
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1758069660
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1758069660
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1758069660
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1758069660
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1758069660
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1758069660
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1758069660
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1758069660
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1758069660
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1758069660
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1758069660
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1758069660
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1758069660
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1758069660
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1758069660
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1758069660
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1758069660
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1758069660
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1758069660
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1758069660
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1758069660
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1758069660
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1758069660
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1758069660
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1758069660
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1758069660
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1758069660
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1758069660
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1758069660
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1758069660
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1758069660
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1758069660
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1758069660
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1758069660
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1758069660
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1758069660
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1758069660
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1758069660
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1758069660
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1758069660
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1758069660
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1758069660
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1758069660
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1758069660
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1758069660
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1758069660
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1758069660
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1185
timestamp 1758069660
transform 1 0 110124 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1197
timestamp 1758069660
transform 1 0 111228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1758069660
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1758069660
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1217
timestamp 1758069660
transform 1 0 113068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1229
timestamp 1758069660
transform 1 0 114172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1241
timestamp 1758069660
transform 1 0 115276 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1253
timestamp 1758069660
transform 1 0 116380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1259
timestamp 1758069660
transform 1 0 116932 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1261
timestamp 1758069660
transform 1 0 117116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1273
timestamp 1758069660
transform 1 0 118220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1285
timestamp 1758069660
transform 1 0 119324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1297
timestamp 1758069660
transform 1 0 120428 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1309
timestamp 1758069660
transform 1 0 121532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1315
timestamp 1758069660
transform 1 0 122084 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1317
timestamp 1758069660
transform 1 0 122268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1329
timestamp 1758069660
transform 1 0 123372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1341
timestamp 1758069660
transform 1 0 124476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1353
timestamp 1758069660
transform 1 0 125580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1365
timestamp 1758069660
transform 1 0 126684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1371
timestamp 1758069660
transform 1 0 127236 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1373
timestamp 1758069660
transform 1 0 127420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1385
timestamp 1758069660
transform 1 0 128524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1397
timestamp 1758069660
transform 1 0 129628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1409
timestamp 1758069660
transform 1 0 130732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1421
timestamp 1758069660
transform 1 0 131836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1427
timestamp 1758069660
transform 1 0 132388 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1429
timestamp 1758069660
transform 1 0 132572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1441
timestamp 1758069660
transform 1 0 133676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1453
timestamp 1758069660
transform 1 0 134780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1465
timestamp 1758069660
transform 1 0 135884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1477
timestamp 1758069660
transform 1 0 136988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1483
timestamp 1758069660
transform 1 0 137540 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1485
timestamp 1758069660
transform 1 0 137724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1497
timestamp 1758069660
transform 1 0 138828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1509
timestamp 1758069660
transform 1 0 139932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1521
timestamp 1758069660
transform 1 0 141036 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1533
timestamp 1758069660
transform 1 0 142140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1539
timestamp 1758069660
transform 1 0 142692 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1541
timestamp 1758069660
transform 1 0 142876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1553
timestamp 1758069660
transform 1 0 143980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1565
timestamp 1758069660
transform 1 0 145084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1577
timestamp 1758069660
transform 1 0 146188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1589
timestamp 1758069660
transform 1 0 147292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1595
timestamp 1758069660
transform 1 0 147844 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1597
timestamp 1758069660
transform 1 0 148028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1609
timestamp 1758069660
transform 1 0 149132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1621
timestamp 1758069660
transform 1 0 150236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1633
timestamp 1758069660
transform 1 0 151340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1645
timestamp 1758069660
transform 1 0 152444 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1651
timestamp 1758069660
transform 1 0 152996 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1653
timestamp 1758069660
transform 1 0 153180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1665
timestamp 1758069660
transform 1 0 154284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1677
timestamp 1758069660
transform 1 0 155388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1689
timestamp 1758069660
transform 1 0 156492 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1701
timestamp 1758069660
transform 1 0 157596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1707
timestamp 1758069660
transform 1 0 158148 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1709
timestamp 1758069660
transform 1 0 158332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1721
timestamp 1758069660
transform 1 0 159436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1733
timestamp 1758069660
transform 1 0 160540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1745
timestamp 1758069660
transform 1 0 161644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1757
timestamp 1758069660
transform 1 0 162748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1763
timestamp 1758069660
transform 1 0 163300 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1765
timestamp 1758069660
transform 1 0 163484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1777
timestamp 1758069660
transform 1 0 164588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1789
timestamp 1758069660
transform 1 0 165692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1801
timestamp 1758069660
transform 1 0 166796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1813
timestamp 1758069660
transform 1 0 167900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1819
timestamp 1758069660
transform 1 0 168452 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1821
timestamp 1758069660
transform 1 0 168636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1833
timestamp 1758069660
transform 1 0 169740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1845
timestamp 1758069660
transform 1 0 170844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1857
timestamp 1758069660
transform 1 0 171948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1869
timestamp 1758069660
transform 1 0 173052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1875
timestamp 1758069660
transform 1 0 173604 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1877
timestamp 1758069660
transform 1 0 173788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1889
timestamp 1758069660
transform 1 0 174892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1901
timestamp 1758069660
transform 1 0 175996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1913
timestamp 1758069660
transform 1 0 177100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1925
timestamp 1758069660
transform 1 0 178204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1931
timestamp 1758069660
transform 1 0 178756 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1933
timestamp 1758069660
transform 1 0 178940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1945
timestamp 1758069660
transform 1 0 180044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1957
timestamp 1758069660
transform 1 0 181148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1969
timestamp 1758069660
transform 1 0 182252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1981
timestamp 1758069660
transform 1 0 183356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1987
timestamp 1758069660
transform 1 0 183908 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1989
timestamp 1758069660
transform 1 0 184092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2001
timestamp 1758069660
transform 1 0 185196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2013
timestamp 1758069660
transform 1 0 186300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2025
timestamp 1758069660
transform 1 0 187404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2037
timestamp 1758069660
transform 1 0 188508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2043
timestamp 1758069660
transform 1 0 189060 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2045
timestamp 1758069660
transform 1 0 189244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2057
timestamp 1758069660
transform 1 0 190348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2069
timestamp 1758069660
transform 1 0 191452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2081
timestamp 1758069660
transform 1 0 192556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2093
timestamp 1758069660
transform 1 0 193660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2099
timestamp 1758069660
transform 1 0 194212 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2101
timestamp 1758069660
transform 1 0 194396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2113
timestamp 1758069660
transform 1 0 195500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2125
timestamp 1758069660
transform 1 0 196604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2137
timestamp 1758069660
transform 1 0 197708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2149
timestamp 1758069660
transform 1 0 198812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2155
timestamp 1758069660
transform 1 0 199364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2157
timestamp 1758069660
transform 1 0 199548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2169
timestamp 1758069660
transform 1 0 200652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2181
timestamp 1758069660
transform 1 0 201756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2193
timestamp 1758069660
transform 1 0 202860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2205
timestamp 1758069660
transform 1 0 203964 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2211
timestamp 1758069660
transform 1 0 204516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2213
timestamp 1758069660
transform 1 0 204700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2225
timestamp 1758069660
transform 1 0 205804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2237
timestamp 1758069660
transform 1 0 206908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2249
timestamp 1758069660
transform 1 0 208012 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2261
timestamp 1758069660
transform 1 0 209116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2267
timestamp 1758069660
transform 1 0 209668 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2269
timestamp 1758069660
transform 1 0 209852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2281
timestamp 1758069660
transform 1 0 210956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2293
timestamp 1758069660
transform 1 0 212060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2305
timestamp 1758069660
transform 1 0 213164 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2317
timestamp 1758069660
transform 1 0 214268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2323
timestamp 1758069660
transform 1 0 214820 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2325
timestamp 1758069660
transform 1 0 215004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2337
timestamp 1758069660
transform 1 0 216108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2349
timestamp 1758069660
transform 1 0 217212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2361
timestamp 1758069660
transform 1 0 218316 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2373
timestamp 1758069660
transform 1 0 219420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2379
timestamp 1758069660
transform 1 0 219972 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2381
timestamp 1758069660
transform 1 0 220156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2393
timestamp 1758069660
transform 1 0 221260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2405
timestamp 1758069660
transform 1 0 222364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2417
timestamp 1758069660
transform 1 0 223468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2429
timestamp 1758069660
transform 1 0 224572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2435
timestamp 1758069660
transform 1 0 225124 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2437
timestamp 1758069660
transform 1 0 225308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2449
timestamp 1758069660
transform 1 0 226412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2461
timestamp 1758069660
transform 1 0 227516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2473
timestamp 1758069660
transform 1 0 228620 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2485
timestamp 1758069660
transform 1 0 229724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2491
timestamp 1758069660
transform 1 0 230276 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2493
timestamp 1758069660
transform 1 0 230460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2505
timestamp 1758069660
transform 1 0 231564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2517
timestamp 1758069660
transform 1 0 232668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2529
timestamp 1758069660
transform 1 0 233772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2541
timestamp 1758069660
transform 1 0 234876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2547
timestamp 1758069660
transform 1 0 235428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2549
timestamp 1758069660
transform 1 0 235612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2561
timestamp 1758069660
transform 1 0 236716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2573
timestamp 1758069660
transform 1 0 237820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2585
timestamp 1758069660
transform 1 0 238924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2597
timestamp 1758069660
transform 1 0 240028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2603
timestamp 1758069660
transform 1 0 240580 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2605
timestamp 1758069660
transform 1 0 240764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2617
timestamp 1758069660
transform 1 0 241868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2629
timestamp 1758069660
transform 1 0 242972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2641
timestamp 1758069660
transform 1 0 244076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2653
timestamp 1758069660
transform 1 0 245180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2659
timestamp 1758069660
transform 1 0 245732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2661
timestamp 1758069660
transform 1 0 245916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2673
timestamp 1758069660
transform 1 0 247020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2685
timestamp 1758069660
transform 1 0 248124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2697
timestamp 1758069660
transform 1 0 249228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2709
timestamp 1758069660
transform 1 0 250332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2715
timestamp 1758069660
transform 1 0 250884 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2717
timestamp 1758069660
transform 1 0 251068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2729
timestamp 1758069660
transform 1 0 252172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2741
timestamp 1758069660
transform 1 0 253276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2753
timestamp 1758069660
transform 1 0 254380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2765
timestamp 1758069660
transform 1 0 255484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2771
timestamp 1758069660
transform 1 0 256036 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2773
timestamp 1758069660
transform 1 0 256220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2785
timestamp 1758069660
transform 1 0 257324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2797
timestamp 1758069660
transform 1 0 258428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2809
timestamp 1758069660
transform 1 0 259532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2821
timestamp 1758069660
transform 1 0 260636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2827
timestamp 1758069660
transform 1 0 261188 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2829
timestamp 1758069660
transform 1 0 261372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2841
timestamp 1758069660
transform 1 0 262476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2853
timestamp 1758069660
transform 1 0 263580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2865
timestamp 1758069660
transform 1 0 264684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2877
timestamp 1758069660
transform 1 0 265788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2883
timestamp 1758069660
transform 1 0 266340 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2885
timestamp 1758069660
transform 1 0 266524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2897
timestamp 1758069660
transform 1 0 267628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2909
timestamp 1758069660
transform 1 0 268732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2921
timestamp 1758069660
transform 1 0 269836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2933
timestamp 1758069660
transform 1 0 270940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2939
timestamp 1758069660
transform 1 0 271492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2941
timestamp 1758069660
transform 1 0 271676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2953
timestamp 1758069660
transform 1 0 272780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2965
timestamp 1758069660
transform 1 0 273884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2977
timestamp 1758069660
transform 1 0 274988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2989
timestamp 1758069660
transform 1 0 276092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2995
timestamp 1758069660
transform 1 0 276644 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2997
timestamp 1758069660
transform 1 0 276828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3009
timestamp 1758069660
transform 1 0 277932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3021
timestamp 1758069660
transform 1 0 279036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3033
timestamp 1758069660
transform 1 0 280140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3045
timestamp 1758069660
transform 1 0 281244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3051
timestamp 1758069660
transform 1 0 281796 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3053
timestamp 1758069660
transform 1 0 281980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3065
timestamp 1758069660
transform 1 0 283084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3077
timestamp 1758069660
transform 1 0 284188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3089
timestamp 1758069660
transform 1 0 285292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3101
timestamp 1758069660
transform 1 0 286396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3107
timestamp 1758069660
transform 1 0 286948 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3109
timestamp 1758069660
transform 1 0 287132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3121
timestamp 1758069660
transform 1 0 288236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3133
timestamp 1758069660
transform 1 0 289340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3145
timestamp 1758069660
transform 1 0 290444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3157
timestamp 1758069660
transform 1 0 291548 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3163
timestamp 1758069660
transform 1 0 292100 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3165
timestamp 1758069660
transform 1 0 292284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3177
timestamp 1758069660
transform 1 0 293388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3189
timestamp 1758069660
transform 1 0 294492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3201
timestamp 1758069660
transform 1 0 295596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3213
timestamp 1758069660
transform 1 0 296700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3219
timestamp 1758069660
transform 1 0 297252 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3221
timestamp 1758069660
transform 1 0 297436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3233
timestamp 1758069660
transform 1 0 298540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3245
timestamp 1758069660
transform 1 0 299644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3257
timestamp 1758069660
transform 1 0 300748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3269
timestamp 1758069660
transform 1 0 301852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3275
timestamp 1758069660
transform 1 0 302404 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3277
timestamp 1758069660
transform 1 0 302588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3289
timestamp 1758069660
transform 1 0 303692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3301 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 304796 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1758069660
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1758069660
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1758069660
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1758069660
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1758069660
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1758069660
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1758069660
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1758069660
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1758069660
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1758069660
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1758069660
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1758069660
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1758069660
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1758069660
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1758069660
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1758069660
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1758069660
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1758069660
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1758069660
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1758069660
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1758069660
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1758069660
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1758069660
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1758069660
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1758069660
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1758069660
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1758069660
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1758069660
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1758069660
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1758069660
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1758069660
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1758069660
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1758069660
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1758069660
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1758069660
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1758069660
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1758069660
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1758069660
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1758069660
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1758069660
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1758069660
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1758069660
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1758069660
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1758069660
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1758069660
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1758069660
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1758069660
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1758069660
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1758069660
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1758069660
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1758069660
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1758069660
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1758069660
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1758069660
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1758069660
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1758069660
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1758069660
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1758069660
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1758069660
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1758069660
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1758069660
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1758069660
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1758069660
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1758069660
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1758069660
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1758069660
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1758069660
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1758069660
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1758069660
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1758069660
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1758069660
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1758069660
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1758069660
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1758069660
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1758069660
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1758069660
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1758069660
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1758069660
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1758069660
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1758069660
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1758069660
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1758069660
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1758069660
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1758069660
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1758069660
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1758069660
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1758069660
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1758069660
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1758069660
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1758069660
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1758069660
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1758069660
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1758069660
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1758069660
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1758069660
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1758069660
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1758069660
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1758069660
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1758069660
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1758069660
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1758069660
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1758069660
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1758069660
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1758069660
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1758069660
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1758069660
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1758069660
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1758069660
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1758069660
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1758069660
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1758069660
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1758069660
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1758069660
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1758069660
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1758069660
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1758069660
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1758069660
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1758069660
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1758069660
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1758069660
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1758069660
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1758069660
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1758069660
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1758069660
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1758069660
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1758069660
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1758069660
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1758069660
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1758069660
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1758069660
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1758069660
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1758069660
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1758069660
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1758069660
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1257
timestamp 1758069660
transform 1 0 116748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1269
timestamp 1758069660
transform 1 0 117852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1281
timestamp 1758069660
transform 1 0 118956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1287
timestamp 1758069660
transform 1 0 119508 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1289
timestamp 1758069660
transform 1 0 119692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1301
timestamp 1758069660
transform 1 0 120796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1313
timestamp 1758069660
transform 1 0 121900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1325
timestamp 1758069660
transform 1 0 123004 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1337
timestamp 1758069660
transform 1 0 124108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1343
timestamp 1758069660
transform 1 0 124660 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1345
timestamp 1758069660
transform 1 0 124844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1357
timestamp 1758069660
transform 1 0 125948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1369
timestamp 1758069660
transform 1 0 127052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1381
timestamp 1758069660
transform 1 0 128156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1393
timestamp 1758069660
transform 1 0 129260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1399
timestamp 1758069660
transform 1 0 129812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1401
timestamp 1758069660
transform 1 0 129996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1413
timestamp 1758069660
transform 1 0 131100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1425
timestamp 1758069660
transform 1 0 132204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1437
timestamp 1758069660
transform 1 0 133308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1449
timestamp 1758069660
transform 1 0 134412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1455
timestamp 1758069660
transform 1 0 134964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1457
timestamp 1758069660
transform 1 0 135148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1469
timestamp 1758069660
transform 1 0 136252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1481
timestamp 1758069660
transform 1 0 137356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1493
timestamp 1758069660
transform 1 0 138460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1505
timestamp 1758069660
transform 1 0 139564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1511
timestamp 1758069660
transform 1 0 140116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1513
timestamp 1758069660
transform 1 0 140300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1525
timestamp 1758069660
transform 1 0 141404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1537
timestamp 1758069660
transform 1 0 142508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1549
timestamp 1758069660
transform 1 0 143612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1561
timestamp 1758069660
transform 1 0 144716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1567
timestamp 1758069660
transform 1 0 145268 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1569
timestamp 1758069660
transform 1 0 145452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1581
timestamp 1758069660
transform 1 0 146556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1593
timestamp 1758069660
transform 1 0 147660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1605
timestamp 1758069660
transform 1 0 148764 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1617
timestamp 1758069660
transform 1 0 149868 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1623
timestamp 1758069660
transform 1 0 150420 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1625
timestamp 1758069660
transform 1 0 150604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1637
timestamp 1758069660
transform 1 0 151708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1649
timestamp 1758069660
transform 1 0 152812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1661
timestamp 1758069660
transform 1 0 153916 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1673
timestamp 1758069660
transform 1 0 155020 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1679
timestamp 1758069660
transform 1 0 155572 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1681
timestamp 1758069660
transform 1 0 155756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1693
timestamp 1758069660
transform 1 0 156860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1705
timestamp 1758069660
transform 1 0 157964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1717
timestamp 1758069660
transform 1 0 159068 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1729
timestamp 1758069660
transform 1 0 160172 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1735
timestamp 1758069660
transform 1 0 160724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1737
timestamp 1758069660
transform 1 0 160908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1749
timestamp 1758069660
transform 1 0 162012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1761
timestamp 1758069660
transform 1 0 163116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1773
timestamp 1758069660
transform 1 0 164220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1785
timestamp 1758069660
transform 1 0 165324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1791
timestamp 1758069660
transform 1 0 165876 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1793
timestamp 1758069660
transform 1 0 166060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1805
timestamp 1758069660
transform 1 0 167164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1817
timestamp 1758069660
transform 1 0 168268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1829
timestamp 1758069660
transform 1 0 169372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1841
timestamp 1758069660
transform 1 0 170476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1847
timestamp 1758069660
transform 1 0 171028 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1849
timestamp 1758069660
transform 1 0 171212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1861
timestamp 1758069660
transform 1 0 172316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1873
timestamp 1758069660
transform 1 0 173420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1885
timestamp 1758069660
transform 1 0 174524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1897
timestamp 1758069660
transform 1 0 175628 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1903
timestamp 1758069660
transform 1 0 176180 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1905
timestamp 1758069660
transform 1 0 176364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1917
timestamp 1758069660
transform 1 0 177468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1929
timestamp 1758069660
transform 1 0 178572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1941
timestamp 1758069660
transform 1 0 179676 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1953
timestamp 1758069660
transform 1 0 180780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1959
timestamp 1758069660
transform 1 0 181332 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1961
timestamp 1758069660
transform 1 0 181516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1973
timestamp 1758069660
transform 1 0 182620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1985
timestamp 1758069660
transform 1 0 183724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1997
timestamp 1758069660
transform 1 0 184828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2009
timestamp 1758069660
transform 1 0 185932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2015
timestamp 1758069660
transform 1 0 186484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2017
timestamp 1758069660
transform 1 0 186668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2029
timestamp 1758069660
transform 1 0 187772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2041
timestamp 1758069660
transform 1 0 188876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2053
timestamp 1758069660
transform 1 0 189980 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2065
timestamp 1758069660
transform 1 0 191084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2071
timestamp 1758069660
transform 1 0 191636 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2073
timestamp 1758069660
transform 1 0 191820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2085
timestamp 1758069660
transform 1 0 192924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2097
timestamp 1758069660
transform 1 0 194028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2109
timestamp 1758069660
transform 1 0 195132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2121
timestamp 1758069660
transform 1 0 196236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2127
timestamp 1758069660
transform 1 0 196788 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2129
timestamp 1758069660
transform 1 0 196972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2141
timestamp 1758069660
transform 1 0 198076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2153
timestamp 1758069660
transform 1 0 199180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2165
timestamp 1758069660
transform 1 0 200284 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2177
timestamp 1758069660
transform 1 0 201388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2183
timestamp 1758069660
transform 1 0 201940 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2185
timestamp 1758069660
transform 1 0 202124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2197
timestamp 1758069660
transform 1 0 203228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2209
timestamp 1758069660
transform 1 0 204332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2221
timestamp 1758069660
transform 1 0 205436 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2233
timestamp 1758069660
transform 1 0 206540 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2239
timestamp 1758069660
transform 1 0 207092 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2241
timestamp 1758069660
transform 1 0 207276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2253
timestamp 1758069660
transform 1 0 208380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2265
timestamp 1758069660
transform 1 0 209484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2277
timestamp 1758069660
transform 1 0 210588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2289
timestamp 1758069660
transform 1 0 211692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2295
timestamp 1758069660
transform 1 0 212244 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2297
timestamp 1758069660
transform 1 0 212428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2309
timestamp 1758069660
transform 1 0 213532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2321
timestamp 1758069660
transform 1 0 214636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2333
timestamp 1758069660
transform 1 0 215740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2345
timestamp 1758069660
transform 1 0 216844 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2351
timestamp 1758069660
transform 1 0 217396 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2353
timestamp 1758069660
transform 1 0 217580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2365
timestamp 1758069660
transform 1 0 218684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2377
timestamp 1758069660
transform 1 0 219788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2389
timestamp 1758069660
transform 1 0 220892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2401
timestamp 1758069660
transform 1 0 221996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2407
timestamp 1758069660
transform 1 0 222548 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2409
timestamp 1758069660
transform 1 0 222732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2421
timestamp 1758069660
transform 1 0 223836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2433
timestamp 1758069660
transform 1 0 224940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2445
timestamp 1758069660
transform 1 0 226044 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2457
timestamp 1758069660
transform 1 0 227148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2463
timestamp 1758069660
transform 1 0 227700 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2465
timestamp 1758069660
transform 1 0 227884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2477
timestamp 1758069660
transform 1 0 228988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2489
timestamp 1758069660
transform 1 0 230092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2501
timestamp 1758069660
transform 1 0 231196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2513
timestamp 1758069660
transform 1 0 232300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2519
timestamp 1758069660
transform 1 0 232852 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2521
timestamp 1758069660
transform 1 0 233036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2533
timestamp 1758069660
transform 1 0 234140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2545
timestamp 1758069660
transform 1 0 235244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2557
timestamp 1758069660
transform 1 0 236348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2569
timestamp 1758069660
transform 1 0 237452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2575
timestamp 1758069660
transform 1 0 238004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2577
timestamp 1758069660
transform 1 0 238188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2589
timestamp 1758069660
transform 1 0 239292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2601
timestamp 1758069660
transform 1 0 240396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2613
timestamp 1758069660
transform 1 0 241500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2625
timestamp 1758069660
transform 1 0 242604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2631
timestamp 1758069660
transform 1 0 243156 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2633
timestamp 1758069660
transform 1 0 243340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2645
timestamp 1758069660
transform 1 0 244444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2657
timestamp 1758069660
transform 1 0 245548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2669
timestamp 1758069660
transform 1 0 246652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2681
timestamp 1758069660
transform 1 0 247756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2687
timestamp 1758069660
transform 1 0 248308 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2689
timestamp 1758069660
transform 1 0 248492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2701
timestamp 1758069660
transform 1 0 249596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2713
timestamp 1758069660
transform 1 0 250700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2725
timestamp 1758069660
transform 1 0 251804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2737
timestamp 1758069660
transform 1 0 252908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2743
timestamp 1758069660
transform 1 0 253460 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2745
timestamp 1758069660
transform 1 0 253644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2757
timestamp 1758069660
transform 1 0 254748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2769
timestamp 1758069660
transform 1 0 255852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2781
timestamp 1758069660
transform 1 0 256956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2793
timestamp 1758069660
transform 1 0 258060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2799
timestamp 1758069660
transform 1 0 258612 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2801
timestamp 1758069660
transform 1 0 258796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2813
timestamp 1758069660
transform 1 0 259900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2825
timestamp 1758069660
transform 1 0 261004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2837
timestamp 1758069660
transform 1 0 262108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2849
timestamp 1758069660
transform 1 0 263212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2855
timestamp 1758069660
transform 1 0 263764 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2857
timestamp 1758069660
transform 1 0 263948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2869
timestamp 1758069660
transform 1 0 265052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2881
timestamp 1758069660
transform 1 0 266156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2893
timestamp 1758069660
transform 1 0 267260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2905
timestamp 1758069660
transform 1 0 268364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2911
timestamp 1758069660
transform 1 0 268916 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2913
timestamp 1758069660
transform 1 0 269100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2925
timestamp 1758069660
transform 1 0 270204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2937
timestamp 1758069660
transform 1 0 271308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2949
timestamp 1758069660
transform 1 0 272412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2961
timestamp 1758069660
transform 1 0 273516 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2967
timestamp 1758069660
transform 1 0 274068 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2969
timestamp 1758069660
transform 1 0 274252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2981
timestamp 1758069660
transform 1 0 275356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2993
timestamp 1758069660
transform 1 0 276460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3005
timestamp 1758069660
transform 1 0 277564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3017
timestamp 1758069660
transform 1 0 278668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3023
timestamp 1758069660
transform 1 0 279220 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3025
timestamp 1758069660
transform 1 0 279404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3037
timestamp 1758069660
transform 1 0 280508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3049
timestamp 1758069660
transform 1 0 281612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3061
timestamp 1758069660
transform 1 0 282716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3073
timestamp 1758069660
transform 1 0 283820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3079
timestamp 1758069660
transform 1 0 284372 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3081
timestamp 1758069660
transform 1 0 284556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3093
timestamp 1758069660
transform 1 0 285660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3105
timestamp 1758069660
transform 1 0 286764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3117
timestamp 1758069660
transform 1 0 287868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3129
timestamp 1758069660
transform 1 0 288972 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3135
timestamp 1758069660
transform 1 0 289524 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3137
timestamp 1758069660
transform 1 0 289708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3149
timestamp 1758069660
transform 1 0 290812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3161
timestamp 1758069660
transform 1 0 291916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3173
timestamp 1758069660
transform 1 0 293020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3185
timestamp 1758069660
transform 1 0 294124 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3191
timestamp 1758069660
transform 1 0 294676 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3193
timestamp 1758069660
transform 1 0 294860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3205
timestamp 1758069660
transform 1 0 295964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3217
timestamp 1758069660
transform 1 0 297068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3229
timestamp 1758069660
transform 1 0 298172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3241
timestamp 1758069660
transform 1 0 299276 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3247
timestamp 1758069660
transform 1 0 299828 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3249
timestamp 1758069660
transform 1 0 300012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3261
timestamp 1758069660
transform 1 0 301116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3273
timestamp 1758069660
transform 1 0 302220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3285
timestamp 1758069660
transform 1 0 303324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3297
timestamp 1758069660
transform 1 0 304428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3303
timestamp 1758069660
transform 1 0 304980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3305
timestamp 1758069660
transform 1 0 305164 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1758069660
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1758069660
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1758069660
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1758069660
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1758069660
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1758069660
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1758069660
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1758069660
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1758069660
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1758069660
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1758069660
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1758069660
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1758069660
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1758069660
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1758069660
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1758069660
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1758069660
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1758069660
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1758069660
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1758069660
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1758069660
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1758069660
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1758069660
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1758069660
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1758069660
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1758069660
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1758069660
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1758069660
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1758069660
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1758069660
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1758069660
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1758069660
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1758069660
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1758069660
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1758069660
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1758069660
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1758069660
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1758069660
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1758069660
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1758069660
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1758069660
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1758069660
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1758069660
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1758069660
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1758069660
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1758069660
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1758069660
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1758069660
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1758069660
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1758069660
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1758069660
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1758069660
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1758069660
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1758069660
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1758069660
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1758069660
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1758069660
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1758069660
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1758069660
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1758069660
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1758069660
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1758069660
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1758069660
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1758069660
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1758069660
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1758069660
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1758069660
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1758069660
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1758069660
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1758069660
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1758069660
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1758069660
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1758069660
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1758069660
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1758069660
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1758069660
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1758069660
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1758069660
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1758069660
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1758069660
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1758069660
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1758069660
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1758069660
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1758069660
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1758069660
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1758069660
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1758069660
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1758069660
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1758069660
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1758069660
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1758069660
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1758069660
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1758069660
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1758069660
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1758069660
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1758069660
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1758069660
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1758069660
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1758069660
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1758069660
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1758069660
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1758069660
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1758069660
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1758069660
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1758069660
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1758069660
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1758069660
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1758069660
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1758069660
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1758069660
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1758069660
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1758069660
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1758069660
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1758069660
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1758069660
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1758069660
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1758069660
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1758069660
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1758069660
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1758069660
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1758069660
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1758069660
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1758069660
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1758069660
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1758069660
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1758069660
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1758069660
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1758069660
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1758069660
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1758069660
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1217
timestamp 1758069660
transform 1 0 113068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1229
timestamp 1758069660
transform 1 0 114172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1241
timestamp 1758069660
transform 1 0 115276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1253
timestamp 1758069660
transform 1 0 116380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1758069660
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1261
timestamp 1758069660
transform 1 0 117116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1273
timestamp 1758069660
transform 1 0 118220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1285
timestamp 1758069660
transform 1 0 119324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1297
timestamp 1758069660
transform 1 0 120428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1309
timestamp 1758069660
transform 1 0 121532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1315
timestamp 1758069660
transform 1 0 122084 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1317
timestamp 1758069660
transform 1 0 122268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1329
timestamp 1758069660
transform 1 0 123372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1341
timestamp 1758069660
transform 1 0 124476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1353
timestamp 1758069660
transform 1 0 125580 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1365
timestamp 1758069660
transform 1 0 126684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1371
timestamp 1758069660
transform 1 0 127236 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1373
timestamp 1758069660
transform 1 0 127420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1385
timestamp 1758069660
transform 1 0 128524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1397
timestamp 1758069660
transform 1 0 129628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1409
timestamp 1758069660
transform 1 0 130732 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1421
timestamp 1758069660
transform 1 0 131836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1427
timestamp 1758069660
transform 1 0 132388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1429
timestamp 1758069660
transform 1 0 132572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1441
timestamp 1758069660
transform 1 0 133676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1453
timestamp 1758069660
transform 1 0 134780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1465
timestamp 1758069660
transform 1 0 135884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1477
timestamp 1758069660
transform 1 0 136988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1483
timestamp 1758069660
transform 1 0 137540 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1485
timestamp 1758069660
transform 1 0 137724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1497
timestamp 1758069660
transform 1 0 138828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1509
timestamp 1758069660
transform 1 0 139932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1521
timestamp 1758069660
transform 1 0 141036 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1533
timestamp 1758069660
transform 1 0 142140 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1539
timestamp 1758069660
transform 1 0 142692 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1541
timestamp 1758069660
transform 1 0 142876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1553
timestamp 1758069660
transform 1 0 143980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1565
timestamp 1758069660
transform 1 0 145084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1577
timestamp 1758069660
transform 1 0 146188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1589
timestamp 1758069660
transform 1 0 147292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1595
timestamp 1758069660
transform 1 0 147844 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1597
timestamp 1758069660
transform 1 0 148028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1609
timestamp 1758069660
transform 1 0 149132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1621
timestamp 1758069660
transform 1 0 150236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1633
timestamp 1758069660
transform 1 0 151340 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1645
timestamp 1758069660
transform 1 0 152444 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1651
timestamp 1758069660
transform 1 0 152996 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1653
timestamp 1758069660
transform 1 0 153180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1665
timestamp 1758069660
transform 1 0 154284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1677
timestamp 1758069660
transform 1 0 155388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1689
timestamp 1758069660
transform 1 0 156492 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1701
timestamp 1758069660
transform 1 0 157596 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1707
timestamp 1758069660
transform 1 0 158148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1709
timestamp 1758069660
transform 1 0 158332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1721
timestamp 1758069660
transform 1 0 159436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1733
timestamp 1758069660
transform 1 0 160540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1745
timestamp 1758069660
transform 1 0 161644 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1757
timestamp 1758069660
transform 1 0 162748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1763
timestamp 1758069660
transform 1 0 163300 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1765
timestamp 1758069660
transform 1 0 163484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1777
timestamp 1758069660
transform 1 0 164588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1789
timestamp 1758069660
transform 1 0 165692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1801
timestamp 1758069660
transform 1 0 166796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1813
timestamp 1758069660
transform 1 0 167900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1819
timestamp 1758069660
transform 1 0 168452 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1821
timestamp 1758069660
transform 1 0 168636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1833
timestamp 1758069660
transform 1 0 169740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1845
timestamp 1758069660
transform 1 0 170844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1857
timestamp 1758069660
transform 1 0 171948 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1869
timestamp 1758069660
transform 1 0 173052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1875
timestamp 1758069660
transform 1 0 173604 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1877
timestamp 1758069660
transform 1 0 173788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1889
timestamp 1758069660
transform 1 0 174892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1901
timestamp 1758069660
transform 1 0 175996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1913
timestamp 1758069660
transform 1 0 177100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1925
timestamp 1758069660
transform 1 0 178204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1931
timestamp 1758069660
transform 1 0 178756 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1933
timestamp 1758069660
transform 1 0 178940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1945
timestamp 1758069660
transform 1 0 180044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1957
timestamp 1758069660
transform 1 0 181148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1969
timestamp 1758069660
transform 1 0 182252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1981
timestamp 1758069660
transform 1 0 183356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1987
timestamp 1758069660
transform 1 0 183908 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1989
timestamp 1758069660
transform 1 0 184092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2001
timestamp 1758069660
transform 1 0 185196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2013
timestamp 1758069660
transform 1 0 186300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2025
timestamp 1758069660
transform 1 0 187404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2037
timestamp 1758069660
transform 1 0 188508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2043
timestamp 1758069660
transform 1 0 189060 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2045
timestamp 1758069660
transform 1 0 189244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2057
timestamp 1758069660
transform 1 0 190348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2069
timestamp 1758069660
transform 1 0 191452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2081
timestamp 1758069660
transform 1 0 192556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2093
timestamp 1758069660
transform 1 0 193660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2099
timestamp 1758069660
transform 1 0 194212 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2101
timestamp 1758069660
transform 1 0 194396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2113
timestamp 1758069660
transform 1 0 195500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2125
timestamp 1758069660
transform 1 0 196604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2137
timestamp 1758069660
transform 1 0 197708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2149
timestamp 1758069660
transform 1 0 198812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2155
timestamp 1758069660
transform 1 0 199364 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2157
timestamp 1758069660
transform 1 0 199548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2169
timestamp 1758069660
transform 1 0 200652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2181
timestamp 1758069660
transform 1 0 201756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2193
timestamp 1758069660
transform 1 0 202860 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2205
timestamp 1758069660
transform 1 0 203964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2211
timestamp 1758069660
transform 1 0 204516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2213
timestamp 1758069660
transform 1 0 204700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2225
timestamp 1758069660
transform 1 0 205804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2237
timestamp 1758069660
transform 1 0 206908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2249
timestamp 1758069660
transform 1 0 208012 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2261
timestamp 1758069660
transform 1 0 209116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2267
timestamp 1758069660
transform 1 0 209668 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2269
timestamp 1758069660
transform 1 0 209852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2281
timestamp 1758069660
transform 1 0 210956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2293
timestamp 1758069660
transform 1 0 212060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2305
timestamp 1758069660
transform 1 0 213164 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2317
timestamp 1758069660
transform 1 0 214268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2323
timestamp 1758069660
transform 1 0 214820 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2325
timestamp 1758069660
transform 1 0 215004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2337
timestamp 1758069660
transform 1 0 216108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2349
timestamp 1758069660
transform 1 0 217212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2361
timestamp 1758069660
transform 1 0 218316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2373
timestamp 1758069660
transform 1 0 219420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2379
timestamp 1758069660
transform 1 0 219972 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2381
timestamp 1758069660
transform 1 0 220156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2393
timestamp 1758069660
transform 1 0 221260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2405
timestamp 1758069660
transform 1 0 222364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2417
timestamp 1758069660
transform 1 0 223468 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2429
timestamp 1758069660
transform 1 0 224572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2435
timestamp 1758069660
transform 1 0 225124 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2437
timestamp 1758069660
transform 1 0 225308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2449
timestamp 1758069660
transform 1 0 226412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2461
timestamp 1758069660
transform 1 0 227516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2473
timestamp 1758069660
transform 1 0 228620 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2485
timestamp 1758069660
transform 1 0 229724 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2491
timestamp 1758069660
transform 1 0 230276 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2493
timestamp 1758069660
transform 1 0 230460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2505
timestamp 1758069660
transform 1 0 231564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2517
timestamp 1758069660
transform 1 0 232668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2529
timestamp 1758069660
transform 1 0 233772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2541
timestamp 1758069660
transform 1 0 234876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2547
timestamp 1758069660
transform 1 0 235428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2549
timestamp 1758069660
transform 1 0 235612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2561
timestamp 1758069660
transform 1 0 236716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2573
timestamp 1758069660
transform 1 0 237820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2585
timestamp 1758069660
transform 1 0 238924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2597
timestamp 1758069660
transform 1 0 240028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2603
timestamp 1758069660
transform 1 0 240580 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2605
timestamp 1758069660
transform 1 0 240764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2617
timestamp 1758069660
transform 1 0 241868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2629
timestamp 1758069660
transform 1 0 242972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2641
timestamp 1758069660
transform 1 0 244076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2653
timestamp 1758069660
transform 1 0 245180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2659
timestamp 1758069660
transform 1 0 245732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2661
timestamp 1758069660
transform 1 0 245916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2673
timestamp 1758069660
transform 1 0 247020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2685
timestamp 1758069660
transform 1 0 248124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2697
timestamp 1758069660
transform 1 0 249228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2709
timestamp 1758069660
transform 1 0 250332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2715
timestamp 1758069660
transform 1 0 250884 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2717
timestamp 1758069660
transform 1 0 251068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2729
timestamp 1758069660
transform 1 0 252172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2741
timestamp 1758069660
transform 1 0 253276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2753
timestamp 1758069660
transform 1 0 254380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2765
timestamp 1758069660
transform 1 0 255484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2771
timestamp 1758069660
transform 1 0 256036 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2773
timestamp 1758069660
transform 1 0 256220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2785
timestamp 1758069660
transform 1 0 257324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2797
timestamp 1758069660
transform 1 0 258428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2809
timestamp 1758069660
transform 1 0 259532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2821
timestamp 1758069660
transform 1 0 260636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2827
timestamp 1758069660
transform 1 0 261188 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2829
timestamp 1758069660
transform 1 0 261372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2841
timestamp 1758069660
transform 1 0 262476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2853
timestamp 1758069660
transform 1 0 263580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2865
timestamp 1758069660
transform 1 0 264684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2877
timestamp 1758069660
transform 1 0 265788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2883
timestamp 1758069660
transform 1 0 266340 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2885
timestamp 1758069660
transform 1 0 266524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2897
timestamp 1758069660
transform 1 0 267628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2909
timestamp 1758069660
transform 1 0 268732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2921
timestamp 1758069660
transform 1 0 269836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2933
timestamp 1758069660
transform 1 0 270940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2939
timestamp 1758069660
transform 1 0 271492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2941
timestamp 1758069660
transform 1 0 271676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2953
timestamp 1758069660
transform 1 0 272780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2965
timestamp 1758069660
transform 1 0 273884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2977
timestamp 1758069660
transform 1 0 274988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2989
timestamp 1758069660
transform 1 0 276092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2995
timestamp 1758069660
transform 1 0 276644 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2997
timestamp 1758069660
transform 1 0 276828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3009
timestamp 1758069660
transform 1 0 277932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3021
timestamp 1758069660
transform 1 0 279036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3033
timestamp 1758069660
transform 1 0 280140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3045
timestamp 1758069660
transform 1 0 281244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3051
timestamp 1758069660
transform 1 0 281796 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3053
timestamp 1758069660
transform 1 0 281980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3065
timestamp 1758069660
transform 1 0 283084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3077
timestamp 1758069660
transform 1 0 284188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3089
timestamp 1758069660
transform 1 0 285292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3101
timestamp 1758069660
transform 1 0 286396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3107
timestamp 1758069660
transform 1 0 286948 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3109
timestamp 1758069660
transform 1 0 287132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3121
timestamp 1758069660
transform 1 0 288236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3133
timestamp 1758069660
transform 1 0 289340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3145
timestamp 1758069660
transform 1 0 290444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3157
timestamp 1758069660
transform 1 0 291548 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3163
timestamp 1758069660
transform 1 0 292100 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3165
timestamp 1758069660
transform 1 0 292284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3177
timestamp 1758069660
transform 1 0 293388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3189
timestamp 1758069660
transform 1 0 294492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3201
timestamp 1758069660
transform 1 0 295596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3213
timestamp 1758069660
transform 1 0 296700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3219
timestamp 1758069660
transform 1 0 297252 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3221
timestamp 1758069660
transform 1 0 297436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3233
timestamp 1758069660
transform 1 0 298540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3245
timestamp 1758069660
transform 1 0 299644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3257
timestamp 1758069660
transform 1 0 300748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3269
timestamp 1758069660
transform 1 0 301852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3275
timestamp 1758069660
transform 1 0 302404 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3277
timestamp 1758069660
transform 1 0 302588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3289
timestamp 1758069660
transform 1 0 303692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3301
timestamp 1758069660
transform 1 0 304796 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1758069660
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1758069660
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1758069660
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1758069660
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1758069660
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1758069660
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1758069660
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1758069660
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1758069660
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1758069660
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1758069660
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1758069660
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1758069660
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1758069660
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1758069660
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1758069660
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1758069660
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1758069660
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1758069660
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1758069660
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1758069660
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1758069660
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1758069660
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1758069660
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1758069660
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1758069660
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1758069660
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1758069660
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1758069660
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1758069660
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1758069660
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1758069660
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1758069660
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1758069660
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1758069660
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1758069660
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1758069660
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1758069660
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1758069660
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1758069660
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1758069660
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1758069660
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1758069660
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1758069660
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1758069660
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1758069660
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1758069660
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1758069660
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1758069660
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1758069660
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1758069660
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1758069660
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1758069660
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1758069660
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1758069660
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1758069660
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1758069660
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1758069660
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1758069660
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1758069660
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1758069660
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1758069660
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1758069660
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1758069660
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1758069660
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1758069660
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1758069660
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1758069660
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1758069660
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1758069660
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1758069660
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1758069660
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1758069660
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1758069660
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1758069660
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1758069660
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1758069660
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1758069660
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1758069660
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1758069660
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1758069660
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1758069660
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1758069660
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1758069660
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1758069660
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1758069660
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1758069660
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1758069660
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1758069660
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1758069660
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1758069660
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1758069660
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1758069660
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1758069660
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1758069660
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1758069660
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1758069660
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1758069660
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1758069660
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1758069660
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1758069660
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1758069660
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1758069660
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1758069660
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1758069660
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1758069660
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1758069660
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1758069660
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1758069660
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1758069660
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1758069660
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1758069660
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1758069660
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1758069660
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1758069660
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1758069660
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1758069660
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1758069660
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1758069660
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1758069660
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1758069660
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1758069660
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1758069660
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1758069660
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1758069660
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1758069660
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1758069660
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1758069660
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1758069660
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1758069660
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1758069660
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1758069660
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1758069660
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1245
timestamp 1758069660
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1257
timestamp 1758069660
transform 1 0 116748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1269
timestamp 1758069660
transform 1 0 117852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1281
timestamp 1758069660
transform 1 0 118956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1287
timestamp 1758069660
transform 1 0 119508 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1289
timestamp 1758069660
transform 1 0 119692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1301
timestamp 1758069660
transform 1 0 120796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1313
timestamp 1758069660
transform 1 0 121900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1325
timestamp 1758069660
transform 1 0 123004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1337
timestamp 1758069660
transform 1 0 124108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1343
timestamp 1758069660
transform 1 0 124660 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1345
timestamp 1758069660
transform 1 0 124844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1357
timestamp 1758069660
transform 1 0 125948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1369
timestamp 1758069660
transform 1 0 127052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1381
timestamp 1758069660
transform 1 0 128156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1393
timestamp 1758069660
transform 1 0 129260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1399
timestamp 1758069660
transform 1 0 129812 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1401
timestamp 1758069660
transform 1 0 129996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1413
timestamp 1758069660
transform 1 0 131100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1425
timestamp 1758069660
transform 1 0 132204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1437
timestamp 1758069660
transform 1 0 133308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1449
timestamp 1758069660
transform 1 0 134412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1455
timestamp 1758069660
transform 1 0 134964 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1457
timestamp 1758069660
transform 1 0 135148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1469
timestamp 1758069660
transform 1 0 136252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1481
timestamp 1758069660
transform 1 0 137356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1493
timestamp 1758069660
transform 1 0 138460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1505
timestamp 1758069660
transform 1 0 139564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1511
timestamp 1758069660
transform 1 0 140116 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1513
timestamp 1758069660
transform 1 0 140300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1525
timestamp 1758069660
transform 1 0 141404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1537
timestamp 1758069660
transform 1 0 142508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1549
timestamp 1758069660
transform 1 0 143612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1561
timestamp 1758069660
transform 1 0 144716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1567
timestamp 1758069660
transform 1 0 145268 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1569
timestamp 1758069660
transform 1 0 145452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1581
timestamp 1758069660
transform 1 0 146556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1593
timestamp 1758069660
transform 1 0 147660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1605
timestamp 1758069660
transform 1 0 148764 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1617
timestamp 1758069660
transform 1 0 149868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1623
timestamp 1758069660
transform 1 0 150420 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1625
timestamp 1758069660
transform 1 0 150604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1637
timestamp 1758069660
transform 1 0 151708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1649
timestamp 1758069660
transform 1 0 152812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1661
timestamp 1758069660
transform 1 0 153916 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1673
timestamp 1758069660
transform 1 0 155020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1679
timestamp 1758069660
transform 1 0 155572 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1681
timestamp 1758069660
transform 1 0 155756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1693
timestamp 1758069660
transform 1 0 156860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1705
timestamp 1758069660
transform 1 0 157964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1717
timestamp 1758069660
transform 1 0 159068 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1729
timestamp 1758069660
transform 1 0 160172 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1735
timestamp 1758069660
transform 1 0 160724 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1737
timestamp 1758069660
transform 1 0 160908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1749
timestamp 1758069660
transform 1 0 162012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1761
timestamp 1758069660
transform 1 0 163116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1773
timestamp 1758069660
transform 1 0 164220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1785
timestamp 1758069660
transform 1 0 165324 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1791
timestamp 1758069660
transform 1 0 165876 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1793
timestamp 1758069660
transform 1 0 166060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1805
timestamp 1758069660
transform 1 0 167164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1817
timestamp 1758069660
transform 1 0 168268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1829
timestamp 1758069660
transform 1 0 169372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1841
timestamp 1758069660
transform 1 0 170476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1847
timestamp 1758069660
transform 1 0 171028 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1849
timestamp 1758069660
transform 1 0 171212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1861
timestamp 1758069660
transform 1 0 172316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1873
timestamp 1758069660
transform 1 0 173420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1885
timestamp 1758069660
transform 1 0 174524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1897
timestamp 1758069660
transform 1 0 175628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1903
timestamp 1758069660
transform 1 0 176180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1905
timestamp 1758069660
transform 1 0 176364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1917
timestamp 1758069660
transform 1 0 177468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1929
timestamp 1758069660
transform 1 0 178572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1941
timestamp 1758069660
transform 1 0 179676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1953
timestamp 1758069660
transform 1 0 180780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1959
timestamp 1758069660
transform 1 0 181332 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1961
timestamp 1758069660
transform 1 0 181516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1973
timestamp 1758069660
transform 1 0 182620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1985
timestamp 1758069660
transform 1 0 183724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1997
timestamp 1758069660
transform 1 0 184828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2009
timestamp 1758069660
transform 1 0 185932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2015
timestamp 1758069660
transform 1 0 186484 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2017
timestamp 1758069660
transform 1 0 186668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2029
timestamp 1758069660
transform 1 0 187772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2041
timestamp 1758069660
transform 1 0 188876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2053
timestamp 1758069660
transform 1 0 189980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2065
timestamp 1758069660
transform 1 0 191084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2071
timestamp 1758069660
transform 1 0 191636 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2073
timestamp 1758069660
transform 1 0 191820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2085
timestamp 1758069660
transform 1 0 192924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2097
timestamp 1758069660
transform 1 0 194028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2109
timestamp 1758069660
transform 1 0 195132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2121
timestamp 1758069660
transform 1 0 196236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2127
timestamp 1758069660
transform 1 0 196788 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2129
timestamp 1758069660
transform 1 0 196972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2141
timestamp 1758069660
transform 1 0 198076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2153
timestamp 1758069660
transform 1 0 199180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2165
timestamp 1758069660
transform 1 0 200284 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2177
timestamp 1758069660
transform 1 0 201388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2183
timestamp 1758069660
transform 1 0 201940 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2185
timestamp 1758069660
transform 1 0 202124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2197
timestamp 1758069660
transform 1 0 203228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2209
timestamp 1758069660
transform 1 0 204332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2221
timestamp 1758069660
transform 1 0 205436 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2233
timestamp 1758069660
transform 1 0 206540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2239
timestamp 1758069660
transform 1 0 207092 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2241
timestamp 1758069660
transform 1 0 207276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2253
timestamp 1758069660
transform 1 0 208380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2265
timestamp 1758069660
transform 1 0 209484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2277
timestamp 1758069660
transform 1 0 210588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2289
timestamp 1758069660
transform 1 0 211692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2295
timestamp 1758069660
transform 1 0 212244 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2297
timestamp 1758069660
transform 1 0 212428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2309
timestamp 1758069660
transform 1 0 213532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2321
timestamp 1758069660
transform 1 0 214636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2333
timestamp 1758069660
transform 1 0 215740 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2345
timestamp 1758069660
transform 1 0 216844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2351
timestamp 1758069660
transform 1 0 217396 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2353
timestamp 1758069660
transform 1 0 217580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2365
timestamp 1758069660
transform 1 0 218684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2377
timestamp 1758069660
transform 1 0 219788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2389
timestamp 1758069660
transform 1 0 220892 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2401
timestamp 1758069660
transform 1 0 221996 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2407
timestamp 1758069660
transform 1 0 222548 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2409
timestamp 1758069660
transform 1 0 222732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2421
timestamp 1758069660
transform 1 0 223836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2433
timestamp 1758069660
transform 1 0 224940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2445
timestamp 1758069660
transform 1 0 226044 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2457
timestamp 1758069660
transform 1 0 227148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2463
timestamp 1758069660
transform 1 0 227700 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2465
timestamp 1758069660
transform 1 0 227884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2477
timestamp 1758069660
transform 1 0 228988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2489
timestamp 1758069660
transform 1 0 230092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2501
timestamp 1758069660
transform 1 0 231196 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2513
timestamp 1758069660
transform 1 0 232300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2519
timestamp 1758069660
transform 1 0 232852 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2521
timestamp 1758069660
transform 1 0 233036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2533
timestamp 1758069660
transform 1 0 234140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2545
timestamp 1758069660
transform 1 0 235244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2557
timestamp 1758069660
transform 1 0 236348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2569
timestamp 1758069660
transform 1 0 237452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2575
timestamp 1758069660
transform 1 0 238004 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2577
timestamp 1758069660
transform 1 0 238188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2589
timestamp 1758069660
transform 1 0 239292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2601
timestamp 1758069660
transform 1 0 240396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2613
timestamp 1758069660
transform 1 0 241500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2625
timestamp 1758069660
transform 1 0 242604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2631
timestamp 1758069660
transform 1 0 243156 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2633
timestamp 1758069660
transform 1 0 243340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2645
timestamp 1758069660
transform 1 0 244444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2657
timestamp 1758069660
transform 1 0 245548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2669
timestamp 1758069660
transform 1 0 246652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2681
timestamp 1758069660
transform 1 0 247756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2687
timestamp 1758069660
transform 1 0 248308 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2689
timestamp 1758069660
transform 1 0 248492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2701
timestamp 1758069660
transform 1 0 249596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2713
timestamp 1758069660
transform 1 0 250700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2725
timestamp 1758069660
transform 1 0 251804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2737
timestamp 1758069660
transform 1 0 252908 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2743
timestamp 1758069660
transform 1 0 253460 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2745
timestamp 1758069660
transform 1 0 253644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2757
timestamp 1758069660
transform 1 0 254748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2769
timestamp 1758069660
transform 1 0 255852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2781
timestamp 1758069660
transform 1 0 256956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2793
timestamp 1758069660
transform 1 0 258060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2799
timestamp 1758069660
transform 1 0 258612 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2801
timestamp 1758069660
transform 1 0 258796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2813
timestamp 1758069660
transform 1 0 259900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2825
timestamp 1758069660
transform 1 0 261004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2837
timestamp 1758069660
transform 1 0 262108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2849
timestamp 1758069660
transform 1 0 263212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2855
timestamp 1758069660
transform 1 0 263764 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2857
timestamp 1758069660
transform 1 0 263948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2869
timestamp 1758069660
transform 1 0 265052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2881
timestamp 1758069660
transform 1 0 266156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2893
timestamp 1758069660
transform 1 0 267260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2905
timestamp 1758069660
transform 1 0 268364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2911
timestamp 1758069660
transform 1 0 268916 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2913
timestamp 1758069660
transform 1 0 269100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2925
timestamp 1758069660
transform 1 0 270204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2937
timestamp 1758069660
transform 1 0 271308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2949
timestamp 1758069660
transform 1 0 272412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2961
timestamp 1758069660
transform 1 0 273516 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2967
timestamp 1758069660
transform 1 0 274068 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2969
timestamp 1758069660
transform 1 0 274252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2981
timestamp 1758069660
transform 1 0 275356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2993
timestamp 1758069660
transform 1 0 276460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3005
timestamp 1758069660
transform 1 0 277564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3017
timestamp 1758069660
transform 1 0 278668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3023
timestamp 1758069660
transform 1 0 279220 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3025
timestamp 1758069660
transform 1 0 279404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3037
timestamp 1758069660
transform 1 0 280508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3049
timestamp 1758069660
transform 1 0 281612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3061
timestamp 1758069660
transform 1 0 282716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3073
timestamp 1758069660
transform 1 0 283820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3079
timestamp 1758069660
transform 1 0 284372 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3081
timestamp 1758069660
transform 1 0 284556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3093
timestamp 1758069660
transform 1 0 285660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3105
timestamp 1758069660
transform 1 0 286764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3117
timestamp 1758069660
transform 1 0 287868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3129
timestamp 1758069660
transform 1 0 288972 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3135
timestamp 1758069660
transform 1 0 289524 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3137
timestamp 1758069660
transform 1 0 289708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3149
timestamp 1758069660
transform 1 0 290812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3161
timestamp 1758069660
transform 1 0 291916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3173
timestamp 1758069660
transform 1 0 293020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3185
timestamp 1758069660
transform 1 0 294124 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3191
timestamp 1758069660
transform 1 0 294676 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3193
timestamp 1758069660
transform 1 0 294860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3205
timestamp 1758069660
transform 1 0 295964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3217
timestamp 1758069660
transform 1 0 297068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3229
timestamp 1758069660
transform 1 0 298172 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3241
timestamp 1758069660
transform 1 0 299276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3247
timestamp 1758069660
transform 1 0 299828 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3249
timestamp 1758069660
transform 1 0 300012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3261
timestamp 1758069660
transform 1 0 301116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3273
timestamp 1758069660
transform 1 0 302220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3285
timestamp 1758069660
transform 1 0 303324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3297
timestamp 1758069660
transform 1 0 304428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3303
timestamp 1758069660
transform 1 0 304980 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3305
timestamp 1758069660
transform 1 0 305164 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1758069660
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1758069660
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1758069660
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1758069660
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1758069660
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1758069660
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1758069660
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1758069660
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1758069660
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1758069660
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1758069660
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1758069660
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1758069660
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1758069660
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1758069660
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1758069660
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1758069660
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1758069660
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1758069660
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1758069660
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1758069660
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1758069660
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1758069660
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1758069660
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1758069660
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1758069660
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1758069660
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1758069660
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1758069660
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1758069660
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1758069660
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1758069660
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1758069660
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1758069660
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1758069660
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1758069660
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1758069660
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1758069660
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1758069660
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1758069660
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1758069660
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1758069660
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1758069660
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1758069660
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1758069660
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1758069660
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1758069660
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1758069660
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1758069660
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1758069660
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1758069660
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1758069660
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1758069660
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1758069660
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1758069660
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1758069660
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1758069660
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1758069660
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1758069660
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1758069660
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1758069660
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1758069660
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1758069660
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1758069660
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1758069660
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1758069660
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1758069660
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1758069660
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1758069660
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1758069660
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1758069660
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1758069660
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1758069660
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1758069660
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1758069660
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1758069660
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1758069660
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1758069660
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1758069660
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1758069660
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1758069660
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1758069660
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1758069660
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1758069660
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1758069660
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1758069660
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1758069660
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1758069660
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1758069660
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1758069660
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1758069660
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1758069660
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1758069660
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1758069660
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1758069660
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1758069660
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1758069660
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1758069660
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1758069660
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1758069660
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1758069660
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1758069660
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1758069660
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1758069660
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1758069660
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1758069660
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1758069660
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1758069660
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1758069660
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1758069660
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1758069660
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1758069660
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1758069660
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1758069660
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1758069660
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1758069660
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1758069660
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1758069660
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1758069660
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1758069660
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1758069660
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1758069660
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1758069660
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1758069660
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1758069660
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1758069660
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1758069660
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1758069660
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1758069660
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1758069660
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1758069660
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1229
timestamp 1758069660
transform 1 0 114172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1241
timestamp 1758069660
transform 1 0 115276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1758069660
transform 1 0 116380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1758069660
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1261
timestamp 1758069660
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1273
timestamp 1758069660
transform 1 0 118220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1285
timestamp 1758069660
transform 1 0 119324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1297
timestamp 1758069660
transform 1 0 120428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1309
timestamp 1758069660
transform 1 0 121532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1315
timestamp 1758069660
transform 1 0 122084 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1317
timestamp 1758069660
transform 1 0 122268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1329
timestamp 1758069660
transform 1 0 123372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1341
timestamp 1758069660
transform 1 0 124476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1353
timestamp 1758069660
transform 1 0 125580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1365
timestamp 1758069660
transform 1 0 126684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1371
timestamp 1758069660
transform 1 0 127236 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1373
timestamp 1758069660
transform 1 0 127420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1385
timestamp 1758069660
transform 1 0 128524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1397
timestamp 1758069660
transform 1 0 129628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1409
timestamp 1758069660
transform 1 0 130732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1421
timestamp 1758069660
transform 1 0 131836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1427
timestamp 1758069660
transform 1 0 132388 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1429
timestamp 1758069660
transform 1 0 132572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1441
timestamp 1758069660
transform 1 0 133676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1453
timestamp 1758069660
transform 1 0 134780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1465
timestamp 1758069660
transform 1 0 135884 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1477
timestamp 1758069660
transform 1 0 136988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1483
timestamp 1758069660
transform 1 0 137540 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1485
timestamp 1758069660
transform 1 0 137724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1497
timestamp 1758069660
transform 1 0 138828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1509
timestamp 1758069660
transform 1 0 139932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1521
timestamp 1758069660
transform 1 0 141036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1533
timestamp 1758069660
transform 1 0 142140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1539
timestamp 1758069660
transform 1 0 142692 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1541
timestamp 1758069660
transform 1 0 142876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1553
timestamp 1758069660
transform 1 0 143980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1565
timestamp 1758069660
transform 1 0 145084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1577
timestamp 1758069660
transform 1 0 146188 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1589
timestamp 1758069660
transform 1 0 147292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1595
timestamp 1758069660
transform 1 0 147844 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1597
timestamp 1758069660
transform 1 0 148028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1609
timestamp 1758069660
transform 1 0 149132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1621
timestamp 1758069660
transform 1 0 150236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1633
timestamp 1758069660
transform 1 0 151340 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1645
timestamp 1758069660
transform 1 0 152444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1651
timestamp 1758069660
transform 1 0 152996 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1653
timestamp 1758069660
transform 1 0 153180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1665
timestamp 1758069660
transform 1 0 154284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1677
timestamp 1758069660
transform 1 0 155388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1689
timestamp 1758069660
transform 1 0 156492 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1701
timestamp 1758069660
transform 1 0 157596 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1707
timestamp 1758069660
transform 1 0 158148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1709
timestamp 1758069660
transform 1 0 158332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1721
timestamp 1758069660
transform 1 0 159436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1733
timestamp 1758069660
transform 1 0 160540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1745
timestamp 1758069660
transform 1 0 161644 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1757
timestamp 1758069660
transform 1 0 162748 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1763
timestamp 1758069660
transform 1 0 163300 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1765
timestamp 1758069660
transform 1 0 163484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1777
timestamp 1758069660
transform 1 0 164588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1789
timestamp 1758069660
transform 1 0 165692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1801
timestamp 1758069660
transform 1 0 166796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1813
timestamp 1758069660
transform 1 0 167900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1819
timestamp 1758069660
transform 1 0 168452 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1821
timestamp 1758069660
transform 1 0 168636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1833
timestamp 1758069660
transform 1 0 169740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1845
timestamp 1758069660
transform 1 0 170844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1857
timestamp 1758069660
transform 1 0 171948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1869
timestamp 1758069660
transform 1 0 173052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1875
timestamp 1758069660
transform 1 0 173604 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1877
timestamp 1758069660
transform 1 0 173788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1889
timestamp 1758069660
transform 1 0 174892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1901
timestamp 1758069660
transform 1 0 175996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1913
timestamp 1758069660
transform 1 0 177100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1925
timestamp 1758069660
transform 1 0 178204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1931
timestamp 1758069660
transform 1 0 178756 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1933
timestamp 1758069660
transform 1 0 178940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1945
timestamp 1758069660
transform 1 0 180044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1957
timestamp 1758069660
transform 1 0 181148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1969
timestamp 1758069660
transform 1 0 182252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1981
timestamp 1758069660
transform 1 0 183356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1987
timestamp 1758069660
transform 1 0 183908 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1989
timestamp 1758069660
transform 1 0 184092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2001
timestamp 1758069660
transform 1 0 185196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2013
timestamp 1758069660
transform 1 0 186300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2025
timestamp 1758069660
transform 1 0 187404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2037
timestamp 1758069660
transform 1 0 188508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2043
timestamp 1758069660
transform 1 0 189060 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2045
timestamp 1758069660
transform 1 0 189244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2057
timestamp 1758069660
transform 1 0 190348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2069
timestamp 1758069660
transform 1 0 191452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2081
timestamp 1758069660
transform 1 0 192556 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2093
timestamp 1758069660
transform 1 0 193660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2099
timestamp 1758069660
transform 1 0 194212 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2101
timestamp 1758069660
transform 1 0 194396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2113
timestamp 1758069660
transform 1 0 195500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2125
timestamp 1758069660
transform 1 0 196604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2137
timestamp 1758069660
transform 1 0 197708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2149
timestamp 1758069660
transform 1 0 198812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2155
timestamp 1758069660
transform 1 0 199364 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2157
timestamp 1758069660
transform 1 0 199548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2169
timestamp 1758069660
transform 1 0 200652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2181
timestamp 1758069660
transform 1 0 201756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2193
timestamp 1758069660
transform 1 0 202860 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2205
timestamp 1758069660
transform 1 0 203964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2211
timestamp 1758069660
transform 1 0 204516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2213
timestamp 1758069660
transform 1 0 204700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2225
timestamp 1758069660
transform 1 0 205804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2237
timestamp 1758069660
transform 1 0 206908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2249
timestamp 1758069660
transform 1 0 208012 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2261
timestamp 1758069660
transform 1 0 209116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2267
timestamp 1758069660
transform 1 0 209668 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2269
timestamp 1758069660
transform 1 0 209852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2281
timestamp 1758069660
transform 1 0 210956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2293
timestamp 1758069660
transform 1 0 212060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2305
timestamp 1758069660
transform 1 0 213164 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2317
timestamp 1758069660
transform 1 0 214268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2323
timestamp 1758069660
transform 1 0 214820 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2325
timestamp 1758069660
transform 1 0 215004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2337
timestamp 1758069660
transform 1 0 216108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2349
timestamp 1758069660
transform 1 0 217212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2361
timestamp 1758069660
transform 1 0 218316 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2373
timestamp 1758069660
transform 1 0 219420 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2379
timestamp 1758069660
transform 1 0 219972 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2381
timestamp 1758069660
transform 1 0 220156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2393
timestamp 1758069660
transform 1 0 221260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2405
timestamp 1758069660
transform 1 0 222364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2417
timestamp 1758069660
transform 1 0 223468 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2429
timestamp 1758069660
transform 1 0 224572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2435
timestamp 1758069660
transform 1 0 225124 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2437
timestamp 1758069660
transform 1 0 225308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2449
timestamp 1758069660
transform 1 0 226412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2461
timestamp 1758069660
transform 1 0 227516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2473
timestamp 1758069660
transform 1 0 228620 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2485
timestamp 1758069660
transform 1 0 229724 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2491
timestamp 1758069660
transform 1 0 230276 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2493
timestamp 1758069660
transform 1 0 230460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2505
timestamp 1758069660
transform 1 0 231564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2517
timestamp 1758069660
transform 1 0 232668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2529
timestamp 1758069660
transform 1 0 233772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2541
timestamp 1758069660
transform 1 0 234876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2547
timestamp 1758069660
transform 1 0 235428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2549
timestamp 1758069660
transform 1 0 235612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2561
timestamp 1758069660
transform 1 0 236716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2573
timestamp 1758069660
transform 1 0 237820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2585
timestamp 1758069660
transform 1 0 238924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2597
timestamp 1758069660
transform 1 0 240028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2603
timestamp 1758069660
transform 1 0 240580 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2605
timestamp 1758069660
transform 1 0 240764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2617
timestamp 1758069660
transform 1 0 241868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2629
timestamp 1758069660
transform 1 0 242972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2641
timestamp 1758069660
transform 1 0 244076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2653
timestamp 1758069660
transform 1 0 245180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2659
timestamp 1758069660
transform 1 0 245732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2661
timestamp 1758069660
transform 1 0 245916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2673
timestamp 1758069660
transform 1 0 247020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2685
timestamp 1758069660
transform 1 0 248124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2697
timestamp 1758069660
transform 1 0 249228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2709
timestamp 1758069660
transform 1 0 250332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2715
timestamp 1758069660
transform 1 0 250884 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2717
timestamp 1758069660
transform 1 0 251068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2729
timestamp 1758069660
transform 1 0 252172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2741
timestamp 1758069660
transform 1 0 253276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2753
timestamp 1758069660
transform 1 0 254380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2765
timestamp 1758069660
transform 1 0 255484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2771
timestamp 1758069660
transform 1 0 256036 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2773
timestamp 1758069660
transform 1 0 256220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2785
timestamp 1758069660
transform 1 0 257324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2797
timestamp 1758069660
transform 1 0 258428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2809
timestamp 1758069660
transform 1 0 259532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2821
timestamp 1758069660
transform 1 0 260636 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2827
timestamp 1758069660
transform 1 0 261188 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2829
timestamp 1758069660
transform 1 0 261372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2841
timestamp 1758069660
transform 1 0 262476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2853
timestamp 1758069660
transform 1 0 263580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2865
timestamp 1758069660
transform 1 0 264684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2877
timestamp 1758069660
transform 1 0 265788 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2883
timestamp 1758069660
transform 1 0 266340 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2885
timestamp 1758069660
transform 1 0 266524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2897
timestamp 1758069660
transform 1 0 267628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2909
timestamp 1758069660
transform 1 0 268732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2921
timestamp 1758069660
transform 1 0 269836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2933
timestamp 1758069660
transform 1 0 270940 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2939
timestamp 1758069660
transform 1 0 271492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2941
timestamp 1758069660
transform 1 0 271676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2953
timestamp 1758069660
transform 1 0 272780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2965
timestamp 1758069660
transform 1 0 273884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2977
timestamp 1758069660
transform 1 0 274988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2989
timestamp 1758069660
transform 1 0 276092 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2995
timestamp 1758069660
transform 1 0 276644 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2997
timestamp 1758069660
transform 1 0 276828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3009
timestamp 1758069660
transform 1 0 277932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3021
timestamp 1758069660
transform 1 0 279036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3033
timestamp 1758069660
transform 1 0 280140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3045
timestamp 1758069660
transform 1 0 281244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3051
timestamp 1758069660
transform 1 0 281796 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3053
timestamp 1758069660
transform 1 0 281980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3065
timestamp 1758069660
transform 1 0 283084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3077
timestamp 1758069660
transform 1 0 284188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3089
timestamp 1758069660
transform 1 0 285292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3101
timestamp 1758069660
transform 1 0 286396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3107
timestamp 1758069660
transform 1 0 286948 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3109
timestamp 1758069660
transform 1 0 287132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3121
timestamp 1758069660
transform 1 0 288236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3133
timestamp 1758069660
transform 1 0 289340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3145
timestamp 1758069660
transform 1 0 290444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3157
timestamp 1758069660
transform 1 0 291548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3163
timestamp 1758069660
transform 1 0 292100 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3165
timestamp 1758069660
transform 1 0 292284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3177
timestamp 1758069660
transform 1 0 293388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3189
timestamp 1758069660
transform 1 0 294492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3201
timestamp 1758069660
transform 1 0 295596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3213
timestamp 1758069660
transform 1 0 296700 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3219
timestamp 1758069660
transform 1 0 297252 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3221
timestamp 1758069660
transform 1 0 297436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3233
timestamp 1758069660
transform 1 0 298540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3245
timestamp 1758069660
transform 1 0 299644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3257
timestamp 1758069660
transform 1 0 300748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3269
timestamp 1758069660
transform 1 0 301852 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3275
timestamp 1758069660
transform 1 0 302404 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3277
timestamp 1758069660
transform 1 0 302588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3289
timestamp 1758069660
transform 1 0 303692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3301
timestamp 1758069660
transform 1 0 304796 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1758069660
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1758069660
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1758069660
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1758069660
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1758069660
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1758069660
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1758069660
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1758069660
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1758069660
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1758069660
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1758069660
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1758069660
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1758069660
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1758069660
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1758069660
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1758069660
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1758069660
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1758069660
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1758069660
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1758069660
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1758069660
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1758069660
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1758069660
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1758069660
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1758069660
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1758069660
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1758069660
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1758069660
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1758069660
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1758069660
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1758069660
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1758069660
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1758069660
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1758069660
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1758069660
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1758069660
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1758069660
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1758069660
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1758069660
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1758069660
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1758069660
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1758069660
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1758069660
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1758069660
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1758069660
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1758069660
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1758069660
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1758069660
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1758069660
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1758069660
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1758069660
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1758069660
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1758069660
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1758069660
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1758069660
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1758069660
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1758069660
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1758069660
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1758069660
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1758069660
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1758069660
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1758069660
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1758069660
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1758069660
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1758069660
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1758069660
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1758069660
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1758069660
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1758069660
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1758069660
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1758069660
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1758069660
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1758069660
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1758069660
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1758069660
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1758069660
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1758069660
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1758069660
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1758069660
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1758069660
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1758069660
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1758069660
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1758069660
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1758069660
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1758069660
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1758069660
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1758069660
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1758069660
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1758069660
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1758069660
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1758069660
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1758069660
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1758069660
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1758069660
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1758069660
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1758069660
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1758069660
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1758069660
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1758069660
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1758069660
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1758069660
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1758069660
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1758069660
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1758069660
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1758069660
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1758069660
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1758069660
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1758069660
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1758069660
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1758069660
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1758069660
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1758069660
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1758069660
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1758069660
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1758069660
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1758069660
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1758069660
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1758069660
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1758069660
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1758069660
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1758069660
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1758069660
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1758069660
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1758069660
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1758069660
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1758069660
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1758069660
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1189
timestamp 1758069660
transform 1 0 110492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1201
timestamp 1758069660
transform 1 0 111596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1213
timestamp 1758069660
transform 1 0 112700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1758069660
transform 1 0 113804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1758069660
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1233
timestamp 1758069660
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1245
timestamp 1758069660
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1257
timestamp 1758069660
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1269
timestamp 1758069660
transform 1 0 117852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1281
timestamp 1758069660
transform 1 0 118956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1287
timestamp 1758069660
transform 1 0 119508 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1289
timestamp 1758069660
transform 1 0 119692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1301
timestamp 1758069660
transform 1 0 120796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1313
timestamp 1758069660
transform 1 0 121900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1325
timestamp 1758069660
transform 1 0 123004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1337
timestamp 1758069660
transform 1 0 124108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1343
timestamp 1758069660
transform 1 0 124660 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1345
timestamp 1758069660
transform 1 0 124844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1357
timestamp 1758069660
transform 1 0 125948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1369
timestamp 1758069660
transform 1 0 127052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1381
timestamp 1758069660
transform 1 0 128156 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1393
timestamp 1758069660
transform 1 0 129260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1399
timestamp 1758069660
transform 1 0 129812 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1401
timestamp 1758069660
transform 1 0 129996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1413
timestamp 1758069660
transform 1 0 131100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1425
timestamp 1758069660
transform 1 0 132204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1437
timestamp 1758069660
transform 1 0 133308 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1449
timestamp 1758069660
transform 1 0 134412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1455
timestamp 1758069660
transform 1 0 134964 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1457
timestamp 1758069660
transform 1 0 135148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1469
timestamp 1758069660
transform 1 0 136252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1481
timestamp 1758069660
transform 1 0 137356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1493
timestamp 1758069660
transform 1 0 138460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1505
timestamp 1758069660
transform 1 0 139564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1511
timestamp 1758069660
transform 1 0 140116 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1513
timestamp 1758069660
transform 1 0 140300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1525
timestamp 1758069660
transform 1 0 141404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1537
timestamp 1758069660
transform 1 0 142508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1549
timestamp 1758069660
transform 1 0 143612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1561
timestamp 1758069660
transform 1 0 144716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1567
timestamp 1758069660
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1569
timestamp 1758069660
transform 1 0 145452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1581
timestamp 1758069660
transform 1 0 146556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1593
timestamp 1758069660
transform 1 0 147660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1605
timestamp 1758069660
transform 1 0 148764 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1617
timestamp 1758069660
transform 1 0 149868 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1623
timestamp 1758069660
transform 1 0 150420 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1625
timestamp 1758069660
transform 1 0 150604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1637
timestamp 1758069660
transform 1 0 151708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1649
timestamp 1758069660
transform 1 0 152812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1661
timestamp 1758069660
transform 1 0 153916 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1673
timestamp 1758069660
transform 1 0 155020 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1679
timestamp 1758069660
transform 1 0 155572 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1681
timestamp 1758069660
transform 1 0 155756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1693
timestamp 1758069660
transform 1 0 156860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1705
timestamp 1758069660
transform 1 0 157964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1717
timestamp 1758069660
transform 1 0 159068 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1729
timestamp 1758069660
transform 1 0 160172 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1735
timestamp 1758069660
transform 1 0 160724 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1737
timestamp 1758069660
transform 1 0 160908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1749
timestamp 1758069660
transform 1 0 162012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1761
timestamp 1758069660
transform 1 0 163116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1773
timestamp 1758069660
transform 1 0 164220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1785
timestamp 1758069660
transform 1 0 165324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1791
timestamp 1758069660
transform 1 0 165876 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1793
timestamp 1758069660
transform 1 0 166060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1805
timestamp 1758069660
transform 1 0 167164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1817
timestamp 1758069660
transform 1 0 168268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1829
timestamp 1758069660
transform 1 0 169372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1841
timestamp 1758069660
transform 1 0 170476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1847
timestamp 1758069660
transform 1 0 171028 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1849
timestamp 1758069660
transform 1 0 171212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1861
timestamp 1758069660
transform 1 0 172316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1873
timestamp 1758069660
transform 1 0 173420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1885
timestamp 1758069660
transform 1 0 174524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1897
timestamp 1758069660
transform 1 0 175628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1903
timestamp 1758069660
transform 1 0 176180 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1905
timestamp 1758069660
transform 1 0 176364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1917
timestamp 1758069660
transform 1 0 177468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1929
timestamp 1758069660
transform 1 0 178572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1941
timestamp 1758069660
transform 1 0 179676 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1953
timestamp 1758069660
transform 1 0 180780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1959
timestamp 1758069660
transform 1 0 181332 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1961
timestamp 1758069660
transform 1 0 181516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1973
timestamp 1758069660
transform 1 0 182620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1985
timestamp 1758069660
transform 1 0 183724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1997
timestamp 1758069660
transform 1 0 184828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2009
timestamp 1758069660
transform 1 0 185932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2015
timestamp 1758069660
transform 1 0 186484 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2017
timestamp 1758069660
transform 1 0 186668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2029
timestamp 1758069660
transform 1 0 187772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2041
timestamp 1758069660
transform 1 0 188876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2053
timestamp 1758069660
transform 1 0 189980 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2065
timestamp 1758069660
transform 1 0 191084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2071
timestamp 1758069660
transform 1 0 191636 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2073
timestamp 1758069660
transform 1 0 191820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2085
timestamp 1758069660
transform 1 0 192924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2097
timestamp 1758069660
transform 1 0 194028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2109
timestamp 1758069660
transform 1 0 195132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2121
timestamp 1758069660
transform 1 0 196236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2127
timestamp 1758069660
transform 1 0 196788 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2129
timestamp 1758069660
transform 1 0 196972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2141
timestamp 1758069660
transform 1 0 198076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2153
timestamp 1758069660
transform 1 0 199180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2165
timestamp 1758069660
transform 1 0 200284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2177
timestamp 1758069660
transform 1 0 201388 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2183
timestamp 1758069660
transform 1 0 201940 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2185
timestamp 1758069660
transform 1 0 202124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2197
timestamp 1758069660
transform 1 0 203228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2209
timestamp 1758069660
transform 1 0 204332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2221
timestamp 1758069660
transform 1 0 205436 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2233
timestamp 1758069660
transform 1 0 206540 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2239
timestamp 1758069660
transform 1 0 207092 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2241
timestamp 1758069660
transform 1 0 207276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2253
timestamp 1758069660
transform 1 0 208380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2265
timestamp 1758069660
transform 1 0 209484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2277
timestamp 1758069660
transform 1 0 210588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2289
timestamp 1758069660
transform 1 0 211692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2295
timestamp 1758069660
transform 1 0 212244 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2297
timestamp 1758069660
transform 1 0 212428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2309
timestamp 1758069660
transform 1 0 213532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2321
timestamp 1758069660
transform 1 0 214636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2333
timestamp 1758069660
transform 1 0 215740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2345
timestamp 1758069660
transform 1 0 216844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2351
timestamp 1758069660
transform 1 0 217396 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2353
timestamp 1758069660
transform 1 0 217580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2365
timestamp 1758069660
transform 1 0 218684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2377
timestamp 1758069660
transform 1 0 219788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2389
timestamp 1758069660
transform 1 0 220892 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2401
timestamp 1758069660
transform 1 0 221996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2407
timestamp 1758069660
transform 1 0 222548 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2409
timestamp 1758069660
transform 1 0 222732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2421
timestamp 1758069660
transform 1 0 223836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2433
timestamp 1758069660
transform 1 0 224940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2445
timestamp 1758069660
transform 1 0 226044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2457
timestamp 1758069660
transform 1 0 227148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2463
timestamp 1758069660
transform 1 0 227700 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2465
timestamp 1758069660
transform 1 0 227884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2477
timestamp 1758069660
transform 1 0 228988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2489
timestamp 1758069660
transform 1 0 230092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2501
timestamp 1758069660
transform 1 0 231196 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2513
timestamp 1758069660
transform 1 0 232300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2519
timestamp 1758069660
transform 1 0 232852 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2521
timestamp 1758069660
transform 1 0 233036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2533
timestamp 1758069660
transform 1 0 234140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2545
timestamp 1758069660
transform 1 0 235244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2557
timestamp 1758069660
transform 1 0 236348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2569
timestamp 1758069660
transform 1 0 237452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2575
timestamp 1758069660
transform 1 0 238004 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2577
timestamp 1758069660
transform 1 0 238188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2589
timestamp 1758069660
transform 1 0 239292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2601
timestamp 1758069660
transform 1 0 240396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2613
timestamp 1758069660
transform 1 0 241500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2625
timestamp 1758069660
transform 1 0 242604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2631
timestamp 1758069660
transform 1 0 243156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2633
timestamp 1758069660
transform 1 0 243340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2645
timestamp 1758069660
transform 1 0 244444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2657
timestamp 1758069660
transform 1 0 245548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2669
timestamp 1758069660
transform 1 0 246652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2681
timestamp 1758069660
transform 1 0 247756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2687
timestamp 1758069660
transform 1 0 248308 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2689
timestamp 1758069660
transform 1 0 248492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2701
timestamp 1758069660
transform 1 0 249596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2713
timestamp 1758069660
transform 1 0 250700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2725
timestamp 1758069660
transform 1 0 251804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2737
timestamp 1758069660
transform 1 0 252908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2743
timestamp 1758069660
transform 1 0 253460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2745
timestamp 1758069660
transform 1 0 253644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2757
timestamp 1758069660
transform 1 0 254748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2769
timestamp 1758069660
transform 1 0 255852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2781
timestamp 1758069660
transform 1 0 256956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2793
timestamp 1758069660
transform 1 0 258060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2799
timestamp 1758069660
transform 1 0 258612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2801
timestamp 1758069660
transform 1 0 258796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2813
timestamp 1758069660
transform 1 0 259900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2825
timestamp 1758069660
transform 1 0 261004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2837
timestamp 1758069660
transform 1 0 262108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2849
timestamp 1758069660
transform 1 0 263212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2855
timestamp 1758069660
transform 1 0 263764 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2857
timestamp 1758069660
transform 1 0 263948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2869
timestamp 1758069660
transform 1 0 265052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2881
timestamp 1758069660
transform 1 0 266156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2893
timestamp 1758069660
transform 1 0 267260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2905
timestamp 1758069660
transform 1 0 268364 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2911
timestamp 1758069660
transform 1 0 268916 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2913
timestamp 1758069660
transform 1 0 269100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2925
timestamp 1758069660
transform 1 0 270204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2937
timestamp 1758069660
transform 1 0 271308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2949
timestamp 1758069660
transform 1 0 272412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2961
timestamp 1758069660
transform 1 0 273516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2967
timestamp 1758069660
transform 1 0 274068 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2969
timestamp 1758069660
transform 1 0 274252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2981
timestamp 1758069660
transform 1 0 275356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2993
timestamp 1758069660
transform 1 0 276460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3005
timestamp 1758069660
transform 1 0 277564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3017
timestamp 1758069660
transform 1 0 278668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3023
timestamp 1758069660
transform 1 0 279220 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3025
timestamp 1758069660
transform 1 0 279404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3037
timestamp 1758069660
transform 1 0 280508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3049
timestamp 1758069660
transform 1 0 281612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3061
timestamp 1758069660
transform 1 0 282716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3073
timestamp 1758069660
transform 1 0 283820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3079
timestamp 1758069660
transform 1 0 284372 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3081
timestamp 1758069660
transform 1 0 284556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3093
timestamp 1758069660
transform 1 0 285660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3105
timestamp 1758069660
transform 1 0 286764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3117
timestamp 1758069660
transform 1 0 287868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3129
timestamp 1758069660
transform 1 0 288972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3135
timestamp 1758069660
transform 1 0 289524 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3137
timestamp 1758069660
transform 1 0 289708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3149
timestamp 1758069660
transform 1 0 290812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3161
timestamp 1758069660
transform 1 0 291916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3173
timestamp 1758069660
transform 1 0 293020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3185
timestamp 1758069660
transform 1 0 294124 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3191
timestamp 1758069660
transform 1 0 294676 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3193
timestamp 1758069660
transform 1 0 294860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3205
timestamp 1758069660
transform 1 0 295964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3217
timestamp 1758069660
transform 1 0 297068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3229
timestamp 1758069660
transform 1 0 298172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3241
timestamp 1758069660
transform 1 0 299276 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3247
timestamp 1758069660
transform 1 0 299828 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3249
timestamp 1758069660
transform 1 0 300012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3261
timestamp 1758069660
transform 1 0 301116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3273
timestamp 1758069660
transform 1 0 302220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3285
timestamp 1758069660
transform 1 0 303324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3300
timestamp 1758069660
transform 1 0 304704 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3305
timestamp 1758069660
transform 1 0 305164 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1758069660
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1758069660
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1758069660
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1758069660
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1758069660
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1758069660
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1758069660
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1758069660
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1758069660
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1758069660
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1758069660
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1758069660
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1758069660
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1758069660
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1758069660
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1758069660
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1758069660
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1758069660
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1758069660
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1758069660
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1758069660
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1758069660
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1758069660
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1758069660
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1758069660
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1758069660
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1758069660
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1758069660
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1758069660
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1758069660
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1758069660
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1758069660
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1758069660
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1758069660
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1758069660
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1758069660
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1758069660
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1758069660
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1758069660
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1758069660
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1758069660
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1758069660
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1758069660
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1758069660
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1758069660
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1758069660
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1758069660
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1758069660
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1758069660
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1758069660
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1758069660
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1758069660
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1758069660
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1758069660
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1758069660
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1758069660
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1758069660
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1758069660
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1758069660
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1758069660
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1758069660
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1758069660
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1758069660
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1758069660
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1758069660
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1758069660
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1758069660
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1758069660
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1758069660
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1758069660
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1758069660
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1758069660
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1758069660
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1758069660
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1758069660
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1758069660
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1758069660
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1758069660
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1758069660
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1758069660
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1758069660
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1758069660
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1758069660
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1758069660
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1758069660
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1758069660
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1758069660
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1758069660
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1758069660
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1758069660
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1758069660
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1758069660
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1758069660
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1758069660
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1758069660
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1758069660
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1758069660
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1758069660
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1758069660
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1758069660
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1758069660
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1758069660
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1758069660
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1758069660
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1758069660
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1758069660
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1758069660
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1758069660
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1758069660
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1758069660
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1758069660
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1758069660
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1758069660
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1758069660
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1758069660
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1758069660
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1758069660
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1758069660
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1758069660
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1758069660
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1758069660
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1758069660
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1758069660
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1758069660
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1161
timestamp 1758069660
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1758069660
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1185
timestamp 1758069660
transform 1 0 110124 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1758069660
transform 1 0 111228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1758069660
transform 1 0 111780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1205
timestamp 1758069660
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1217
timestamp 1758069660
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1229
timestamp 1758069660
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1241
timestamp 1758069660
transform 1 0 115276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1758069660
transform 1 0 116380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1758069660
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1261
timestamp 1758069660
transform 1 0 117116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1273
timestamp 1758069660
transform 1 0 118220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1285
timestamp 1758069660
transform 1 0 119324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1297
timestamp 1758069660
transform 1 0 120428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1309
timestamp 1758069660
transform 1 0 121532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1315
timestamp 1758069660
transform 1 0 122084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1317
timestamp 1758069660
transform 1 0 122268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1329
timestamp 1758069660
transform 1 0 123372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1341
timestamp 1758069660
transform 1 0 124476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1353
timestamp 1758069660
transform 1 0 125580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1365
timestamp 1758069660
transform 1 0 126684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1371
timestamp 1758069660
transform 1 0 127236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1373
timestamp 1758069660
transform 1 0 127420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1385
timestamp 1758069660
transform 1 0 128524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1397
timestamp 1758069660
transform 1 0 129628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1409
timestamp 1758069660
transform 1 0 130732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1421
timestamp 1758069660
transform 1 0 131836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1427
timestamp 1758069660
transform 1 0 132388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1429
timestamp 1758069660
transform 1 0 132572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1441
timestamp 1758069660
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1453
timestamp 1758069660
transform 1 0 134780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1465
timestamp 1758069660
transform 1 0 135884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1477
timestamp 1758069660
transform 1 0 136988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1483
timestamp 1758069660
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1485
timestamp 1758069660
transform 1 0 137724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1497
timestamp 1758069660
transform 1 0 138828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1509
timestamp 1758069660
transform 1 0 139932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1521
timestamp 1758069660
transform 1 0 141036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1533
timestamp 1758069660
transform 1 0 142140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1539
timestamp 1758069660
transform 1 0 142692 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1541
timestamp 1758069660
transform 1 0 142876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1553
timestamp 1758069660
transform 1 0 143980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1565
timestamp 1758069660
transform 1 0 145084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1577
timestamp 1758069660
transform 1 0 146188 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1589
timestamp 1758069660
transform 1 0 147292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1595
timestamp 1758069660
transform 1 0 147844 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1597
timestamp 1758069660
transform 1 0 148028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1609
timestamp 1758069660
transform 1 0 149132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1621
timestamp 1758069660
transform 1 0 150236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1633
timestamp 1758069660
transform 1 0 151340 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1645
timestamp 1758069660
transform 1 0 152444 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1651
timestamp 1758069660
transform 1 0 152996 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1653
timestamp 1758069660
transform 1 0 153180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1665
timestamp 1758069660
transform 1 0 154284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1677
timestamp 1758069660
transform 1 0 155388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1689
timestamp 1758069660
transform 1 0 156492 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1701
timestamp 1758069660
transform 1 0 157596 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1707
timestamp 1758069660
transform 1 0 158148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1709
timestamp 1758069660
transform 1 0 158332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1721
timestamp 1758069660
transform 1 0 159436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1733
timestamp 1758069660
transform 1 0 160540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1745
timestamp 1758069660
transform 1 0 161644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1757
timestamp 1758069660
transform 1 0 162748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1763
timestamp 1758069660
transform 1 0 163300 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1765
timestamp 1758069660
transform 1 0 163484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1777
timestamp 1758069660
transform 1 0 164588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1789
timestamp 1758069660
transform 1 0 165692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1801
timestamp 1758069660
transform 1 0 166796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1813
timestamp 1758069660
transform 1 0 167900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1819
timestamp 1758069660
transform 1 0 168452 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1821
timestamp 1758069660
transform 1 0 168636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1833
timestamp 1758069660
transform 1 0 169740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1845
timestamp 1758069660
transform 1 0 170844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1857
timestamp 1758069660
transform 1 0 171948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1869
timestamp 1758069660
transform 1 0 173052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1875
timestamp 1758069660
transform 1 0 173604 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1877
timestamp 1758069660
transform 1 0 173788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1889
timestamp 1758069660
transform 1 0 174892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1901
timestamp 1758069660
transform 1 0 175996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1913
timestamp 1758069660
transform 1 0 177100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1925
timestamp 1758069660
transform 1 0 178204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1931
timestamp 1758069660
transform 1 0 178756 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1933
timestamp 1758069660
transform 1 0 178940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1945
timestamp 1758069660
transform 1 0 180044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1957
timestamp 1758069660
transform 1 0 181148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1969
timestamp 1758069660
transform 1 0 182252 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1981
timestamp 1758069660
transform 1 0 183356 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1987
timestamp 1758069660
transform 1 0 183908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1989
timestamp 1758069660
transform 1 0 184092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2001
timestamp 1758069660
transform 1 0 185196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2013
timestamp 1758069660
transform 1 0 186300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2025
timestamp 1758069660
transform 1 0 187404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2037
timestamp 1758069660
transform 1 0 188508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2043
timestamp 1758069660
transform 1 0 189060 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2045
timestamp 1758069660
transform 1 0 189244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2057
timestamp 1758069660
transform 1 0 190348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2069
timestamp 1758069660
transform 1 0 191452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2081
timestamp 1758069660
transform 1 0 192556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2093
timestamp 1758069660
transform 1 0 193660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2099
timestamp 1758069660
transform 1 0 194212 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2101
timestamp 1758069660
transform 1 0 194396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2113
timestamp 1758069660
transform 1 0 195500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2125
timestamp 1758069660
transform 1 0 196604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2137
timestamp 1758069660
transform 1 0 197708 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2149
timestamp 1758069660
transform 1 0 198812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2155
timestamp 1758069660
transform 1 0 199364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2157
timestamp 1758069660
transform 1 0 199548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2169
timestamp 1758069660
transform 1 0 200652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2181
timestamp 1758069660
transform 1 0 201756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2193
timestamp 1758069660
transform 1 0 202860 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2205
timestamp 1758069660
transform 1 0 203964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2211
timestamp 1758069660
transform 1 0 204516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2213
timestamp 1758069660
transform 1 0 204700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2225
timestamp 1758069660
transform 1 0 205804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2237
timestamp 1758069660
transform 1 0 206908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2249
timestamp 1758069660
transform 1 0 208012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2261
timestamp 1758069660
transform 1 0 209116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2267
timestamp 1758069660
transform 1 0 209668 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2269
timestamp 1758069660
transform 1 0 209852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2281
timestamp 1758069660
transform 1 0 210956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2293
timestamp 1758069660
transform 1 0 212060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2305
timestamp 1758069660
transform 1 0 213164 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2317
timestamp 1758069660
transform 1 0 214268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2323
timestamp 1758069660
transform 1 0 214820 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2325
timestamp 1758069660
transform 1 0 215004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2337
timestamp 1758069660
transform 1 0 216108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2349
timestamp 1758069660
transform 1 0 217212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2361
timestamp 1758069660
transform 1 0 218316 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2373
timestamp 1758069660
transform 1 0 219420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2379
timestamp 1758069660
transform 1 0 219972 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2381
timestamp 1758069660
transform 1 0 220156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2393
timestamp 1758069660
transform 1 0 221260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2405
timestamp 1758069660
transform 1 0 222364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2417
timestamp 1758069660
transform 1 0 223468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2429
timestamp 1758069660
transform 1 0 224572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2435
timestamp 1758069660
transform 1 0 225124 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2437
timestamp 1758069660
transform 1 0 225308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2449
timestamp 1758069660
transform 1 0 226412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2461
timestamp 1758069660
transform 1 0 227516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2473
timestamp 1758069660
transform 1 0 228620 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2485
timestamp 1758069660
transform 1 0 229724 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2491
timestamp 1758069660
transform 1 0 230276 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2493
timestamp 1758069660
transform 1 0 230460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2505
timestamp 1758069660
transform 1 0 231564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2517
timestamp 1758069660
transform 1 0 232668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2529
timestamp 1758069660
transform 1 0 233772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2541
timestamp 1758069660
transform 1 0 234876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2547
timestamp 1758069660
transform 1 0 235428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2549
timestamp 1758069660
transform 1 0 235612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2561
timestamp 1758069660
transform 1 0 236716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2573
timestamp 1758069660
transform 1 0 237820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2585
timestamp 1758069660
transform 1 0 238924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2597
timestamp 1758069660
transform 1 0 240028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2603
timestamp 1758069660
transform 1 0 240580 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2605
timestamp 1758069660
transform 1 0 240764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2617
timestamp 1758069660
transform 1 0 241868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2629
timestamp 1758069660
transform 1 0 242972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2641
timestamp 1758069660
transform 1 0 244076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2653
timestamp 1758069660
transform 1 0 245180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2659
timestamp 1758069660
transform 1 0 245732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2661
timestamp 1758069660
transform 1 0 245916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2673
timestamp 1758069660
transform 1 0 247020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2685
timestamp 1758069660
transform 1 0 248124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2697
timestamp 1758069660
transform 1 0 249228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2709
timestamp 1758069660
transform 1 0 250332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2715
timestamp 1758069660
transform 1 0 250884 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2717
timestamp 1758069660
transform 1 0 251068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2729
timestamp 1758069660
transform 1 0 252172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2741
timestamp 1758069660
transform 1 0 253276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2753
timestamp 1758069660
transform 1 0 254380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2765
timestamp 1758069660
transform 1 0 255484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2771
timestamp 1758069660
transform 1 0 256036 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2773
timestamp 1758069660
transform 1 0 256220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2785
timestamp 1758069660
transform 1 0 257324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2797
timestamp 1758069660
transform 1 0 258428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2809
timestamp 1758069660
transform 1 0 259532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2821
timestamp 1758069660
transform 1 0 260636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2827
timestamp 1758069660
transform 1 0 261188 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2829
timestamp 1758069660
transform 1 0 261372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2841
timestamp 1758069660
transform 1 0 262476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2853
timestamp 1758069660
transform 1 0 263580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2865
timestamp 1758069660
transform 1 0 264684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2877
timestamp 1758069660
transform 1 0 265788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2883
timestamp 1758069660
transform 1 0 266340 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2885
timestamp 1758069660
transform 1 0 266524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2897
timestamp 1758069660
transform 1 0 267628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2909
timestamp 1758069660
transform 1 0 268732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2921
timestamp 1758069660
transform 1 0 269836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2933
timestamp 1758069660
transform 1 0 270940 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2939
timestamp 1758069660
transform 1 0 271492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2941
timestamp 1758069660
transform 1 0 271676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2953
timestamp 1758069660
transform 1 0 272780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2965
timestamp 1758069660
transform 1 0 273884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2977
timestamp 1758069660
transform 1 0 274988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2989
timestamp 1758069660
transform 1 0 276092 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2995
timestamp 1758069660
transform 1 0 276644 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2997
timestamp 1758069660
transform 1 0 276828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3009
timestamp 1758069660
transform 1 0 277932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3021
timestamp 1758069660
transform 1 0 279036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3033
timestamp 1758069660
transform 1 0 280140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3045
timestamp 1758069660
transform 1 0 281244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3051
timestamp 1758069660
transform 1 0 281796 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3053
timestamp 1758069660
transform 1 0 281980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3065
timestamp 1758069660
transform 1 0 283084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3077
timestamp 1758069660
transform 1 0 284188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3089
timestamp 1758069660
transform 1 0 285292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3101
timestamp 1758069660
transform 1 0 286396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3107
timestamp 1758069660
transform 1 0 286948 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3109
timestamp 1758069660
transform 1 0 287132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3121
timestamp 1758069660
transform 1 0 288236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3133
timestamp 1758069660
transform 1 0 289340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3145
timestamp 1758069660
transform 1 0 290444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3157
timestamp 1758069660
transform 1 0 291548 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3163
timestamp 1758069660
transform 1 0 292100 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3165
timestamp 1758069660
transform 1 0 292284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3177
timestamp 1758069660
transform 1 0 293388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3189
timestamp 1758069660
transform 1 0 294492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3201
timestamp 1758069660
transform 1 0 295596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3213
timestamp 1758069660
transform 1 0 296700 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3219
timestamp 1758069660
transform 1 0 297252 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3221
timestamp 1758069660
transform 1 0 297436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3233
timestamp 1758069660
transform 1 0 298540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3245
timestamp 1758069660
transform 1 0 299644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3257
timestamp 1758069660
transform 1 0 300748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3269
timestamp 1758069660
transform 1 0 301852 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3275
timestamp 1758069660
transform 1 0 302404 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3277
timestamp 1758069660
transform 1 0 302588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3289
timestamp 1758069660
transform 1 0 303692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3301
timestamp 1758069660
transform 1 0 304796 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1758069660
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1758069660
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1758069660
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1758069660
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1758069660
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1758069660
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1758069660
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1758069660
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1758069660
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1758069660
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1758069660
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1758069660
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1758069660
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1758069660
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1758069660
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1758069660
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1758069660
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1758069660
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1758069660
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1758069660
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1758069660
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1758069660
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1758069660
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1758069660
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1758069660
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1758069660
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1758069660
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1758069660
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1758069660
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1758069660
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1758069660
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1758069660
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1758069660
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1758069660
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1758069660
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1758069660
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1758069660
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1758069660
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1758069660
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1758069660
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1758069660
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1758069660
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1758069660
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1758069660
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1758069660
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1758069660
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1758069660
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1758069660
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1758069660
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1758069660
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1758069660
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1758069660
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1758069660
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1758069660
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1758069660
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1758069660
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1758069660
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1758069660
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1758069660
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1758069660
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1758069660
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1758069660
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1758069660
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1758069660
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1758069660
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1758069660
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1758069660
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1758069660
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1758069660
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1758069660
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1758069660
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1758069660
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1758069660
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1758069660
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1758069660
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1758069660
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1758069660
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1758069660
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1758069660
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1758069660
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1758069660
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1758069660
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1758069660
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1758069660
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1758069660
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1758069660
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1758069660
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_821
timestamp 1758069660
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1758069660
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1758069660
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1758069660
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1758069660
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_865
timestamp 1758069660
transform 1 0 80684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_877
timestamp 1758069660
transform 1 0 81788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_889
timestamp 1758069660
transform 1 0 82892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_895
timestamp 1758069660
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1758069660
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1758069660
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_921
timestamp 1758069660
transform 1 0 85836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_933
timestamp 1758069660
transform 1 0 86940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_945
timestamp 1758069660
transform 1 0 88044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_951
timestamp 1758069660
transform 1 0 88596 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1758069660
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1758069660
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_977
timestamp 1758069660
transform 1 0 90988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_989
timestamp 1758069660
transform 1 0 92092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1001
timestamp 1758069660
transform 1 0 93196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1007
timestamp 1758069660
transform 1 0 93748 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1758069660
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1758069660
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1033
timestamp 1758069660
transform 1 0 96140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1045
timestamp 1758069660
transform 1 0 97244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1057
timestamp 1758069660
transform 1 0 98348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1063
timestamp 1758069660
transform 1 0 98900 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1758069660
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1758069660
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1089
timestamp 1758069660
transform 1 0 101292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1101
timestamp 1758069660
transform 1 0 102396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1113
timestamp 1758069660
transform 1 0 103500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1119
timestamp 1758069660
transform 1 0 104052 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1758069660
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1758069660
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1145
timestamp 1758069660
transform 1 0 106444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1157
timestamp 1758069660
transform 1 0 107548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1169
timestamp 1758069660
transform 1 0 108652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1175
timestamp 1758069660
transform 1 0 109204 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1758069660
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1189
timestamp 1758069660
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1201
timestamp 1758069660
transform 1 0 111596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1213
timestamp 1758069660
transform 1 0 112700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1225
timestamp 1758069660
transform 1 0 113804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1231
timestamp 1758069660
transform 1 0 114356 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1758069660
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1758069660
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1257
timestamp 1758069660
transform 1 0 116748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1269
timestamp 1758069660
transform 1 0 117852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1281
timestamp 1758069660
transform 1 0 118956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1287
timestamp 1758069660
transform 1 0 119508 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1289
timestamp 1758069660
transform 1 0 119692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1301
timestamp 1758069660
transform 1 0 120796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1313
timestamp 1758069660
transform 1 0 121900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1325
timestamp 1758069660
transform 1 0 123004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1337
timestamp 1758069660
transform 1 0 124108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1343
timestamp 1758069660
transform 1 0 124660 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1345
timestamp 1758069660
transform 1 0 124844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1357
timestamp 1758069660
transform 1 0 125948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1369
timestamp 1758069660
transform 1 0 127052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1381
timestamp 1758069660
transform 1 0 128156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1393
timestamp 1758069660
transform 1 0 129260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1399
timestamp 1758069660
transform 1 0 129812 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1401
timestamp 1758069660
transform 1 0 129996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1413
timestamp 1758069660
transform 1 0 131100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1425
timestamp 1758069660
transform 1 0 132204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1437
timestamp 1758069660
transform 1 0 133308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1449
timestamp 1758069660
transform 1 0 134412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1455
timestamp 1758069660
transform 1 0 134964 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1457
timestamp 1758069660
transform 1 0 135148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1469
timestamp 1758069660
transform 1 0 136252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1481
timestamp 1758069660
transform 1 0 137356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1493
timestamp 1758069660
transform 1 0 138460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1505
timestamp 1758069660
transform 1 0 139564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1511
timestamp 1758069660
transform 1 0 140116 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1513
timestamp 1758069660
transform 1 0 140300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1525
timestamp 1758069660
transform 1 0 141404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1537
timestamp 1758069660
transform 1 0 142508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1549
timestamp 1758069660
transform 1 0 143612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1561
timestamp 1758069660
transform 1 0 144716 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1567
timestamp 1758069660
transform 1 0 145268 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1569
timestamp 1758069660
transform 1 0 145452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1581
timestamp 1758069660
transform 1 0 146556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1593
timestamp 1758069660
transform 1 0 147660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1605
timestamp 1758069660
transform 1 0 148764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1617
timestamp 1758069660
transform 1 0 149868 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1623
timestamp 1758069660
transform 1 0 150420 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1625
timestamp 1758069660
transform 1 0 150604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1637
timestamp 1758069660
transform 1 0 151708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1649
timestamp 1758069660
transform 1 0 152812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1661
timestamp 1758069660
transform 1 0 153916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1673
timestamp 1758069660
transform 1 0 155020 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1679
timestamp 1758069660
transform 1 0 155572 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1681
timestamp 1758069660
transform 1 0 155756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1693
timestamp 1758069660
transform 1 0 156860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1705
timestamp 1758069660
transform 1 0 157964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1717
timestamp 1758069660
transform 1 0 159068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1729
timestamp 1758069660
transform 1 0 160172 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1735
timestamp 1758069660
transform 1 0 160724 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1737
timestamp 1758069660
transform 1 0 160908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1749
timestamp 1758069660
transform 1 0 162012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1761
timestamp 1758069660
transform 1 0 163116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1773
timestamp 1758069660
transform 1 0 164220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1785
timestamp 1758069660
transform 1 0 165324 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1791
timestamp 1758069660
transform 1 0 165876 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1793
timestamp 1758069660
transform 1 0 166060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1805
timestamp 1758069660
transform 1 0 167164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1817
timestamp 1758069660
transform 1 0 168268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1829
timestamp 1758069660
transform 1 0 169372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1841
timestamp 1758069660
transform 1 0 170476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1847
timestamp 1758069660
transform 1 0 171028 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1849
timestamp 1758069660
transform 1 0 171212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1861
timestamp 1758069660
transform 1 0 172316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1873
timestamp 1758069660
transform 1 0 173420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1885
timestamp 1758069660
transform 1 0 174524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1897
timestamp 1758069660
transform 1 0 175628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1903
timestamp 1758069660
transform 1 0 176180 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1905
timestamp 1758069660
transform 1 0 176364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1917
timestamp 1758069660
transform 1 0 177468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1929
timestamp 1758069660
transform 1 0 178572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1941
timestamp 1758069660
transform 1 0 179676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1953
timestamp 1758069660
transform 1 0 180780 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1959
timestamp 1758069660
transform 1 0 181332 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1961
timestamp 1758069660
transform 1 0 181516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1973
timestamp 1758069660
transform 1 0 182620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1985
timestamp 1758069660
transform 1 0 183724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1997
timestamp 1758069660
transform 1 0 184828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2009
timestamp 1758069660
transform 1 0 185932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2015
timestamp 1758069660
transform 1 0 186484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2017
timestamp 1758069660
transform 1 0 186668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2029
timestamp 1758069660
transform 1 0 187772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2041
timestamp 1758069660
transform 1 0 188876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2053
timestamp 1758069660
transform 1 0 189980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2065
timestamp 1758069660
transform 1 0 191084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2071
timestamp 1758069660
transform 1 0 191636 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2073
timestamp 1758069660
transform 1 0 191820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2085
timestamp 1758069660
transform 1 0 192924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2097
timestamp 1758069660
transform 1 0 194028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2109
timestamp 1758069660
transform 1 0 195132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2121
timestamp 1758069660
transform 1 0 196236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2127
timestamp 1758069660
transform 1 0 196788 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2129
timestamp 1758069660
transform 1 0 196972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2141
timestamp 1758069660
transform 1 0 198076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2153
timestamp 1758069660
transform 1 0 199180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2165
timestamp 1758069660
transform 1 0 200284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2177
timestamp 1758069660
transform 1 0 201388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2183
timestamp 1758069660
transform 1 0 201940 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2185
timestamp 1758069660
transform 1 0 202124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2197
timestamp 1758069660
transform 1 0 203228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2209
timestamp 1758069660
transform 1 0 204332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2221
timestamp 1758069660
transform 1 0 205436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2233
timestamp 1758069660
transform 1 0 206540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2239
timestamp 1758069660
transform 1 0 207092 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2241
timestamp 1758069660
transform 1 0 207276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2253
timestamp 1758069660
transform 1 0 208380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2265
timestamp 1758069660
transform 1 0 209484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2277
timestamp 1758069660
transform 1 0 210588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2289
timestamp 1758069660
transform 1 0 211692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2295
timestamp 1758069660
transform 1 0 212244 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2297
timestamp 1758069660
transform 1 0 212428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2309
timestamp 1758069660
transform 1 0 213532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2321
timestamp 1758069660
transform 1 0 214636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2333
timestamp 1758069660
transform 1 0 215740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2345
timestamp 1758069660
transform 1 0 216844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2351
timestamp 1758069660
transform 1 0 217396 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2353
timestamp 1758069660
transform 1 0 217580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2365
timestamp 1758069660
transform 1 0 218684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2377
timestamp 1758069660
transform 1 0 219788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2389
timestamp 1758069660
transform 1 0 220892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2401
timestamp 1758069660
transform 1 0 221996 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2407
timestamp 1758069660
transform 1 0 222548 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2409
timestamp 1758069660
transform 1 0 222732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2421
timestamp 1758069660
transform 1 0 223836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2433
timestamp 1758069660
transform 1 0 224940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2445
timestamp 1758069660
transform 1 0 226044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2457
timestamp 1758069660
transform 1 0 227148 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2463
timestamp 1758069660
transform 1 0 227700 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2465
timestamp 1758069660
transform 1 0 227884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2477
timestamp 1758069660
transform 1 0 228988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2489
timestamp 1758069660
transform 1 0 230092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2501
timestamp 1758069660
transform 1 0 231196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2513
timestamp 1758069660
transform 1 0 232300 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2519
timestamp 1758069660
transform 1 0 232852 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2521
timestamp 1758069660
transform 1 0 233036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2533
timestamp 1758069660
transform 1 0 234140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2545
timestamp 1758069660
transform 1 0 235244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2557
timestamp 1758069660
transform 1 0 236348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2569
timestamp 1758069660
transform 1 0 237452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2575
timestamp 1758069660
transform 1 0 238004 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2577
timestamp 1758069660
transform 1 0 238188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2589
timestamp 1758069660
transform 1 0 239292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2601
timestamp 1758069660
transform 1 0 240396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2613
timestamp 1758069660
transform 1 0 241500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2625
timestamp 1758069660
transform 1 0 242604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2631
timestamp 1758069660
transform 1 0 243156 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2633
timestamp 1758069660
transform 1 0 243340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2645
timestamp 1758069660
transform 1 0 244444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2657
timestamp 1758069660
transform 1 0 245548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2669
timestamp 1758069660
transform 1 0 246652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2681
timestamp 1758069660
transform 1 0 247756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2687
timestamp 1758069660
transform 1 0 248308 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2689
timestamp 1758069660
transform 1 0 248492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2701
timestamp 1758069660
transform 1 0 249596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2713
timestamp 1758069660
transform 1 0 250700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2725
timestamp 1758069660
transform 1 0 251804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2737
timestamp 1758069660
transform 1 0 252908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2743
timestamp 1758069660
transform 1 0 253460 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2745
timestamp 1758069660
transform 1 0 253644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2757
timestamp 1758069660
transform 1 0 254748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2769
timestamp 1758069660
transform 1 0 255852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2781
timestamp 1758069660
transform 1 0 256956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2793
timestamp 1758069660
transform 1 0 258060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2799
timestamp 1758069660
transform 1 0 258612 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2801
timestamp 1758069660
transform 1 0 258796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2813
timestamp 1758069660
transform 1 0 259900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2825
timestamp 1758069660
transform 1 0 261004 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2837
timestamp 1758069660
transform 1 0 262108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2849
timestamp 1758069660
transform 1 0 263212 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2855
timestamp 1758069660
transform 1 0 263764 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2857
timestamp 1758069660
transform 1 0 263948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2869
timestamp 1758069660
transform 1 0 265052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2881
timestamp 1758069660
transform 1 0 266156 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2893
timestamp 1758069660
transform 1 0 267260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2905
timestamp 1758069660
transform 1 0 268364 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2911
timestamp 1758069660
transform 1 0 268916 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2913
timestamp 1758069660
transform 1 0 269100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2925
timestamp 1758069660
transform 1 0 270204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2937
timestamp 1758069660
transform 1 0 271308 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2949
timestamp 1758069660
transform 1 0 272412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2961
timestamp 1758069660
transform 1 0 273516 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2967
timestamp 1758069660
transform 1 0 274068 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2969
timestamp 1758069660
transform 1 0 274252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2981
timestamp 1758069660
transform 1 0 275356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2993
timestamp 1758069660
transform 1 0 276460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3005
timestamp 1758069660
transform 1 0 277564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3017
timestamp 1758069660
transform 1 0 278668 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3023
timestamp 1758069660
transform 1 0 279220 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3025
timestamp 1758069660
transform 1 0 279404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3037
timestamp 1758069660
transform 1 0 280508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3049
timestamp 1758069660
transform 1 0 281612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3061
timestamp 1758069660
transform 1 0 282716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3073
timestamp 1758069660
transform 1 0 283820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3079
timestamp 1758069660
transform 1 0 284372 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3081
timestamp 1758069660
transform 1 0 284556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3093
timestamp 1758069660
transform 1 0 285660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3105
timestamp 1758069660
transform 1 0 286764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3117
timestamp 1758069660
transform 1 0 287868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3129
timestamp 1758069660
transform 1 0 288972 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3135
timestamp 1758069660
transform 1 0 289524 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3137
timestamp 1758069660
transform 1 0 289708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3149
timestamp 1758069660
transform 1 0 290812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3161
timestamp 1758069660
transform 1 0 291916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3173
timestamp 1758069660
transform 1 0 293020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3185
timestamp 1758069660
transform 1 0 294124 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3191
timestamp 1758069660
transform 1 0 294676 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3193
timestamp 1758069660
transform 1 0 294860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3205
timestamp 1758069660
transform 1 0 295964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3217
timestamp 1758069660
transform 1 0 297068 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3229
timestamp 1758069660
transform 1 0 298172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3241
timestamp 1758069660
transform 1 0 299276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3247
timestamp 1758069660
transform 1 0 299828 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3249
timestamp 1758069660
transform 1 0 300012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3261
timestamp 1758069660
transform 1 0 301116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3273
timestamp 1758069660
transform 1 0 302220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3285
timestamp 1758069660
transform 1 0 303324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3297
timestamp 1758069660
transform 1 0 304428 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3303
timestamp 1758069660
transform 1 0 304980 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3305
timestamp 1758069660
transform 1 0 305164 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1758069660
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1758069660
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1758069660
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1758069660
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1758069660
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1758069660
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1758069660
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1758069660
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1758069660
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1758069660
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1758069660
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1758069660
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1758069660
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1758069660
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1758069660
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1758069660
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1758069660
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1758069660
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1758069660
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1758069660
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1758069660
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1758069660
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1758069660
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1758069660
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1758069660
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1758069660
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1758069660
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1758069660
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1758069660
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1758069660
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1758069660
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1758069660
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1758069660
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1758069660
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1758069660
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1758069660
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1758069660
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1758069660
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1758069660
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1758069660
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1758069660
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1758069660
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1758069660
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1758069660
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1758069660
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1758069660
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1758069660
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1758069660
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1758069660
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1758069660
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1758069660
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1758069660
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1758069660
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1758069660
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1758069660
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1758069660
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1758069660
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1758069660
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1758069660
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1758069660
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1758069660
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1758069660
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1758069660
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1758069660
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1758069660
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1758069660
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1758069660
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1758069660
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1758069660
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1758069660
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1758069660
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1758069660
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1758069660
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1758069660
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1758069660
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1758069660
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1758069660
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1758069660
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1758069660
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1758069660
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1758069660
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1758069660
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1758069660
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1758069660
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1758069660
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1758069660
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1758069660
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_813
timestamp 1758069660
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_825
timestamp 1758069660
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_837
timestamp 1758069660
transform 1 0 78108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_849
timestamp 1758069660
transform 1 0 79212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_861
timestamp 1758069660
transform 1 0 80316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_867
timestamp 1758069660
transform 1 0 80868 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_869
timestamp 1758069660
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_881
timestamp 1758069660
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_893
timestamp 1758069660
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_905
timestamp 1758069660
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_917
timestamp 1758069660
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_923
timestamp 1758069660
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_925
timestamp 1758069660
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_937
timestamp 1758069660
transform 1 0 87308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_949
timestamp 1758069660
transform 1 0 88412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_961
timestamp 1758069660
transform 1 0 89516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_973
timestamp 1758069660
transform 1 0 90620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_979
timestamp 1758069660
transform 1 0 91172 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_981
timestamp 1758069660
transform 1 0 91356 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_993
timestamp 1758069660
transform 1 0 92460 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1005
timestamp 1758069660
transform 1 0 93564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1017
timestamp 1758069660
transform 1 0 94668 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1029
timestamp 1758069660
transform 1 0 95772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1035
timestamp 1758069660
transform 1 0 96324 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1037
timestamp 1758069660
transform 1 0 96508 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1049
timestamp 1758069660
transform 1 0 97612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1061
timestamp 1758069660
transform 1 0 98716 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1073
timestamp 1758069660
transform 1 0 99820 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1085
timestamp 1758069660
transform 1 0 100924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1091
timestamp 1758069660
transform 1 0 101476 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1093
timestamp 1758069660
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1105
timestamp 1758069660
transform 1 0 102764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1117
timestamp 1758069660
transform 1 0 103868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1129
timestamp 1758069660
transform 1 0 104972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1141
timestamp 1758069660
transform 1 0 106076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1147
timestamp 1758069660
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1149
timestamp 1758069660
transform 1 0 106812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1161
timestamp 1758069660
transform 1 0 107916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1173
timestamp 1758069660
transform 1 0 109020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1185
timestamp 1758069660
transform 1 0 110124 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1197
timestamp 1758069660
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1203
timestamp 1758069660
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1205
timestamp 1758069660
transform 1 0 111964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1217
timestamp 1758069660
transform 1 0 113068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1229
timestamp 1758069660
transform 1 0 114172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1241
timestamp 1758069660
transform 1 0 115276 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1253
timestamp 1758069660
transform 1 0 116380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1259
timestamp 1758069660
transform 1 0 116932 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1261
timestamp 1758069660
transform 1 0 117116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1273
timestamp 1758069660
transform 1 0 118220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1285
timestamp 1758069660
transform 1 0 119324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1297
timestamp 1758069660
transform 1 0 120428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1309
timestamp 1758069660
transform 1 0 121532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1315
timestamp 1758069660
transform 1 0 122084 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1317
timestamp 1758069660
transform 1 0 122268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1329
timestamp 1758069660
transform 1 0 123372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1341
timestamp 1758069660
transform 1 0 124476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1353
timestamp 1758069660
transform 1 0 125580 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1365
timestamp 1758069660
transform 1 0 126684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1371
timestamp 1758069660
transform 1 0 127236 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1373
timestamp 1758069660
transform 1 0 127420 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1385
timestamp 1758069660
transform 1 0 128524 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1397
timestamp 1758069660
transform 1 0 129628 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1409
timestamp 1758069660
transform 1 0 130732 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1421
timestamp 1758069660
transform 1 0 131836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1427
timestamp 1758069660
transform 1 0 132388 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1429
timestamp 1758069660
transform 1 0 132572 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1441
timestamp 1758069660
transform 1 0 133676 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1453
timestamp 1758069660
transform 1 0 134780 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1465
timestamp 1758069660
transform 1 0 135884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1477
timestamp 1758069660
transform 1 0 136988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1483
timestamp 1758069660
transform 1 0 137540 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1485
timestamp 1758069660
transform 1 0 137724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1497
timestamp 1758069660
transform 1 0 138828 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1509
timestamp 1758069660
transform 1 0 139932 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1521
timestamp 1758069660
transform 1 0 141036 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1533
timestamp 1758069660
transform 1 0 142140 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1539
timestamp 1758069660
transform 1 0 142692 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1541
timestamp 1758069660
transform 1 0 142876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1553
timestamp 1758069660
transform 1 0 143980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1565
timestamp 1758069660
transform 1 0 145084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1577
timestamp 1758069660
transform 1 0 146188 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1589
timestamp 1758069660
transform 1 0 147292 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1595
timestamp 1758069660
transform 1 0 147844 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1597
timestamp 1758069660
transform 1 0 148028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1609
timestamp 1758069660
transform 1 0 149132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1621
timestamp 1758069660
transform 1 0 150236 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1633
timestamp 1758069660
transform 1 0 151340 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1645
timestamp 1758069660
transform 1 0 152444 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1651
timestamp 1758069660
transform 1 0 152996 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1653
timestamp 1758069660
transform 1 0 153180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1665
timestamp 1758069660
transform 1 0 154284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1677
timestamp 1758069660
transform 1 0 155388 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1689
timestamp 1758069660
transform 1 0 156492 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1701
timestamp 1758069660
transform 1 0 157596 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1707
timestamp 1758069660
transform 1 0 158148 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1709
timestamp 1758069660
transform 1 0 158332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1721
timestamp 1758069660
transform 1 0 159436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1733
timestamp 1758069660
transform 1 0 160540 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1745
timestamp 1758069660
transform 1 0 161644 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1757
timestamp 1758069660
transform 1 0 162748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1763
timestamp 1758069660
transform 1 0 163300 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1765
timestamp 1758069660
transform 1 0 163484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1777
timestamp 1758069660
transform 1 0 164588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1789
timestamp 1758069660
transform 1 0 165692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1801
timestamp 1758069660
transform 1 0 166796 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1813
timestamp 1758069660
transform 1 0 167900 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1819
timestamp 1758069660
transform 1 0 168452 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1821
timestamp 1758069660
transform 1 0 168636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1833
timestamp 1758069660
transform 1 0 169740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1845
timestamp 1758069660
transform 1 0 170844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1857
timestamp 1758069660
transform 1 0 171948 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1869
timestamp 1758069660
transform 1 0 173052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1875
timestamp 1758069660
transform 1 0 173604 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1877
timestamp 1758069660
transform 1 0 173788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1889
timestamp 1758069660
transform 1 0 174892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1901
timestamp 1758069660
transform 1 0 175996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1913
timestamp 1758069660
transform 1 0 177100 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1925
timestamp 1758069660
transform 1 0 178204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1931
timestamp 1758069660
transform 1 0 178756 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1933
timestamp 1758069660
transform 1 0 178940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1945
timestamp 1758069660
transform 1 0 180044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1957
timestamp 1758069660
transform 1 0 181148 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1969
timestamp 1758069660
transform 1 0 182252 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1981
timestamp 1758069660
transform 1 0 183356 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1987
timestamp 1758069660
transform 1 0 183908 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1989
timestamp 1758069660
transform 1 0 184092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2001
timestamp 1758069660
transform 1 0 185196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2013
timestamp 1758069660
transform 1 0 186300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2025
timestamp 1758069660
transform 1 0 187404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2037
timestamp 1758069660
transform 1 0 188508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2043
timestamp 1758069660
transform 1 0 189060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2045
timestamp 1758069660
transform 1 0 189244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2057
timestamp 1758069660
transform 1 0 190348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2069
timestamp 1758069660
transform 1 0 191452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2081
timestamp 1758069660
transform 1 0 192556 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2093
timestamp 1758069660
transform 1 0 193660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2099
timestamp 1758069660
transform 1 0 194212 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2101
timestamp 1758069660
transform 1 0 194396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2113
timestamp 1758069660
transform 1 0 195500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2125
timestamp 1758069660
transform 1 0 196604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2137
timestamp 1758069660
transform 1 0 197708 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2149
timestamp 1758069660
transform 1 0 198812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2155
timestamp 1758069660
transform 1 0 199364 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2157
timestamp 1758069660
transform 1 0 199548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2169
timestamp 1758069660
transform 1 0 200652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2181
timestamp 1758069660
transform 1 0 201756 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2193
timestamp 1758069660
transform 1 0 202860 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2205
timestamp 1758069660
transform 1 0 203964 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2211
timestamp 1758069660
transform 1 0 204516 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2213
timestamp 1758069660
transform 1 0 204700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2225
timestamp 1758069660
transform 1 0 205804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2237
timestamp 1758069660
transform 1 0 206908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2249
timestamp 1758069660
transform 1 0 208012 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2261
timestamp 1758069660
transform 1 0 209116 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2267
timestamp 1758069660
transform 1 0 209668 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2269
timestamp 1758069660
transform 1 0 209852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2281
timestamp 1758069660
transform 1 0 210956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2293
timestamp 1758069660
transform 1 0 212060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2305
timestamp 1758069660
transform 1 0 213164 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2317
timestamp 1758069660
transform 1 0 214268 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2323
timestamp 1758069660
transform 1 0 214820 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2325
timestamp 1758069660
transform 1 0 215004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2337
timestamp 1758069660
transform 1 0 216108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2349
timestamp 1758069660
transform 1 0 217212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2361
timestamp 1758069660
transform 1 0 218316 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2373
timestamp 1758069660
transform 1 0 219420 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2379
timestamp 1758069660
transform 1 0 219972 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2381
timestamp 1758069660
transform 1 0 220156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2393
timestamp 1758069660
transform 1 0 221260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2405
timestamp 1758069660
transform 1 0 222364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2417
timestamp 1758069660
transform 1 0 223468 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2429
timestamp 1758069660
transform 1 0 224572 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2435
timestamp 1758069660
transform 1 0 225124 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2437
timestamp 1758069660
transform 1 0 225308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2449
timestamp 1758069660
transform 1 0 226412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2461
timestamp 1758069660
transform 1 0 227516 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2473
timestamp 1758069660
transform 1 0 228620 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2485
timestamp 1758069660
transform 1 0 229724 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2491
timestamp 1758069660
transform 1 0 230276 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2493
timestamp 1758069660
transform 1 0 230460 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2505
timestamp 1758069660
transform 1 0 231564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2517
timestamp 1758069660
transform 1 0 232668 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2529
timestamp 1758069660
transform 1 0 233772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2541
timestamp 1758069660
transform 1 0 234876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2547
timestamp 1758069660
transform 1 0 235428 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2549
timestamp 1758069660
transform 1 0 235612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2561
timestamp 1758069660
transform 1 0 236716 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2573
timestamp 1758069660
transform 1 0 237820 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2585
timestamp 1758069660
transform 1 0 238924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2597
timestamp 1758069660
transform 1 0 240028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2603
timestamp 1758069660
transform 1 0 240580 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2605
timestamp 1758069660
transform 1 0 240764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2617
timestamp 1758069660
transform 1 0 241868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2629
timestamp 1758069660
transform 1 0 242972 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2641
timestamp 1758069660
transform 1 0 244076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2653
timestamp 1758069660
transform 1 0 245180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2659
timestamp 1758069660
transform 1 0 245732 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2661
timestamp 1758069660
transform 1 0 245916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2673
timestamp 1758069660
transform 1 0 247020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2685
timestamp 1758069660
transform 1 0 248124 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2697
timestamp 1758069660
transform 1 0 249228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2709
timestamp 1758069660
transform 1 0 250332 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2715
timestamp 1758069660
transform 1 0 250884 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2717
timestamp 1758069660
transform 1 0 251068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2729
timestamp 1758069660
transform 1 0 252172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2741
timestamp 1758069660
transform 1 0 253276 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2753
timestamp 1758069660
transform 1 0 254380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2765
timestamp 1758069660
transform 1 0 255484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2771
timestamp 1758069660
transform 1 0 256036 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2773
timestamp 1758069660
transform 1 0 256220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2785
timestamp 1758069660
transform 1 0 257324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2797
timestamp 1758069660
transform 1 0 258428 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2809
timestamp 1758069660
transform 1 0 259532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2821
timestamp 1758069660
transform 1 0 260636 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2827
timestamp 1758069660
transform 1 0 261188 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2829
timestamp 1758069660
transform 1 0 261372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2841
timestamp 1758069660
transform 1 0 262476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2853
timestamp 1758069660
transform 1 0 263580 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2865
timestamp 1758069660
transform 1 0 264684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2877
timestamp 1758069660
transform 1 0 265788 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2883
timestamp 1758069660
transform 1 0 266340 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2885
timestamp 1758069660
transform 1 0 266524 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2897
timestamp 1758069660
transform 1 0 267628 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2909
timestamp 1758069660
transform 1 0 268732 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2921
timestamp 1758069660
transform 1 0 269836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2933
timestamp 1758069660
transform 1 0 270940 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2939
timestamp 1758069660
transform 1 0 271492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2941
timestamp 1758069660
transform 1 0 271676 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2953
timestamp 1758069660
transform 1 0 272780 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2965
timestamp 1758069660
transform 1 0 273884 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2977
timestamp 1758069660
transform 1 0 274988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2989
timestamp 1758069660
transform 1 0 276092 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2995
timestamp 1758069660
transform 1 0 276644 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2997
timestamp 1758069660
transform 1 0 276828 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3009
timestamp 1758069660
transform 1 0 277932 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3021
timestamp 1758069660
transform 1 0 279036 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3033
timestamp 1758069660
transform 1 0 280140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3045
timestamp 1758069660
transform 1 0 281244 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3051
timestamp 1758069660
transform 1 0 281796 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3053
timestamp 1758069660
transform 1 0 281980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3065
timestamp 1758069660
transform 1 0 283084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3077
timestamp 1758069660
transform 1 0 284188 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3089
timestamp 1758069660
transform 1 0 285292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3101
timestamp 1758069660
transform 1 0 286396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3107
timestamp 1758069660
transform 1 0 286948 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3109
timestamp 1758069660
transform 1 0 287132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3121
timestamp 1758069660
transform 1 0 288236 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3133
timestamp 1758069660
transform 1 0 289340 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3145
timestamp 1758069660
transform 1 0 290444 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3157
timestamp 1758069660
transform 1 0 291548 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3163
timestamp 1758069660
transform 1 0 292100 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3165
timestamp 1758069660
transform 1 0 292284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3177
timestamp 1758069660
transform 1 0 293388 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3189
timestamp 1758069660
transform 1 0 294492 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3201
timestamp 1758069660
transform 1 0 295596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3213
timestamp 1758069660
transform 1 0 296700 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3219
timestamp 1758069660
transform 1 0 297252 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3221
timestamp 1758069660
transform 1 0 297436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3233
timestamp 1758069660
transform 1 0 298540 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3245
timestamp 1758069660
transform 1 0 299644 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3257
timestamp 1758069660
transform 1 0 300748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3269
timestamp 1758069660
transform 1 0 301852 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3275
timestamp 1758069660
transform 1 0 302404 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3277
timestamp 1758069660
transform 1 0 302588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3289
timestamp 1758069660
transform 1 0 303692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3301
timestamp 1758069660
transform 1 0 304796 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_10
timestamp 1758069660
transform 1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_14
timestamp 1758069660
transform 1 0 2392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_18
timestamp 1758069660
transform 1 0 2760 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_22
timestamp 1758069660
transform 1 0 3128 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 1758069660
transform 1 0 4232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp 1758069660
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1758069660
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1758069660
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1758069660
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1758069660
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1758069660
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1758069660
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1758069660
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1758069660
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1758069660
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1758069660
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1758069660
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1758069660
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1758069660
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1758069660
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1758069660
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1758069660
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1758069660
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1758069660
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1758069660
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1758069660
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1758069660
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1758069660
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1758069660
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1758069660
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1758069660
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1758069660
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1758069660
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1758069660
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1758069660
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1758069660
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1758069660
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1758069660
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1758069660
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1758069660
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1758069660
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1758069660
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1758069660
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1758069660
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1758069660
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1758069660
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1758069660
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1758069660
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1758069660
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1758069660
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1758069660
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1758069660
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1758069660
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1758069660
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1758069660
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1758069660
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1758069660
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1758069660
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1758069660
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1758069660
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1758069660
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1758069660
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1758069660
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1758069660
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1758069660
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1758069660
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1758069660
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1758069660
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1758069660
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1758069660
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1758069660
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1758069660
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1758069660
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1758069660
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1758069660
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1758069660
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1758069660
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1758069660
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1758069660
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1758069660
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1758069660
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1758069660
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1758069660
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1758069660
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1758069660
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1758069660
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1758069660
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1758069660
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_821
timestamp 1758069660
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1758069660
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1758069660
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_841
timestamp 1758069660
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_853
timestamp 1758069660
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_865
timestamp 1758069660
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_877
timestamp 1758069660
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1758069660
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1758069660
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_897
timestamp 1758069660
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_909
timestamp 1758069660
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_921
timestamp 1758069660
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_933
timestamp 1758069660
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_945
timestamp 1758069660
transform 1 0 88044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1758069660
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_953
timestamp 1758069660
transform 1 0 88780 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_965
timestamp 1758069660
transform 1 0 89884 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_977
timestamp 1758069660
transform 1 0 90988 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_989
timestamp 1758069660
transform 1 0 92092 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1001
timestamp 1758069660
transform 1 0 93196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1007
timestamp 1758069660
transform 1 0 93748 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1009
timestamp 1758069660
transform 1 0 93932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1021
timestamp 1758069660
transform 1 0 95036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1033
timestamp 1758069660
transform 1 0 96140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1045
timestamp 1758069660
transform 1 0 97244 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1057
timestamp 1758069660
transform 1 0 98348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1063
timestamp 1758069660
transform 1 0 98900 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1065
timestamp 1758069660
transform 1 0 99084 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1077
timestamp 1758069660
transform 1 0 100188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1089
timestamp 1758069660
transform 1 0 101292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1101
timestamp 1758069660
transform 1 0 102396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1113
timestamp 1758069660
transform 1 0 103500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1119
timestamp 1758069660
transform 1 0 104052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1121
timestamp 1758069660
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1133
timestamp 1758069660
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1145
timestamp 1758069660
transform 1 0 106444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1157
timestamp 1758069660
transform 1 0 107548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1169
timestamp 1758069660
transform 1 0 108652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1175
timestamp 1758069660
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1177
timestamp 1758069660
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1189
timestamp 1758069660
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1201
timestamp 1758069660
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1213
timestamp 1758069660
transform 1 0 112700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1225
timestamp 1758069660
transform 1 0 113804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1231
timestamp 1758069660
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1233
timestamp 1758069660
transform 1 0 114540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1245
timestamp 1758069660
transform 1 0 115644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1257
timestamp 1758069660
transform 1 0 116748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1269
timestamp 1758069660
transform 1 0 117852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1281
timestamp 1758069660
transform 1 0 118956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1287
timestamp 1758069660
transform 1 0 119508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1289
timestamp 1758069660
transform 1 0 119692 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1301
timestamp 1758069660
transform 1 0 120796 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1313
timestamp 1758069660
transform 1 0 121900 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1325
timestamp 1758069660
transform 1 0 123004 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1337
timestamp 1758069660
transform 1 0 124108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1343
timestamp 1758069660
transform 1 0 124660 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1345
timestamp 1758069660
transform 1 0 124844 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1357
timestamp 1758069660
transform 1 0 125948 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1369
timestamp 1758069660
transform 1 0 127052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1381
timestamp 1758069660
transform 1 0 128156 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1393
timestamp 1758069660
transform 1 0 129260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1399
timestamp 1758069660
transform 1 0 129812 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1401
timestamp 1758069660
transform 1 0 129996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1413
timestamp 1758069660
transform 1 0 131100 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1425
timestamp 1758069660
transform 1 0 132204 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1437
timestamp 1758069660
transform 1 0 133308 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1449
timestamp 1758069660
transform 1 0 134412 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1455
timestamp 1758069660
transform 1 0 134964 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1457
timestamp 1758069660
transform 1 0 135148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1469
timestamp 1758069660
transform 1 0 136252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1481
timestamp 1758069660
transform 1 0 137356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1493
timestamp 1758069660
transform 1 0 138460 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1505
timestamp 1758069660
transform 1 0 139564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1511
timestamp 1758069660
transform 1 0 140116 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1513
timestamp 1758069660
transform 1 0 140300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1525
timestamp 1758069660
transform 1 0 141404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1537
timestamp 1758069660
transform 1 0 142508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1549
timestamp 1758069660
transform 1 0 143612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1561
timestamp 1758069660
transform 1 0 144716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1567
timestamp 1758069660
transform 1 0 145268 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1569
timestamp 1758069660
transform 1 0 145452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1581
timestamp 1758069660
transform 1 0 146556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1593
timestamp 1758069660
transform 1 0 147660 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1605
timestamp 1758069660
transform 1 0 148764 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1617
timestamp 1758069660
transform 1 0 149868 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1623
timestamp 1758069660
transform 1 0 150420 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1625
timestamp 1758069660
transform 1 0 150604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1637
timestamp 1758069660
transform 1 0 151708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1649
timestamp 1758069660
transform 1 0 152812 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1661
timestamp 1758069660
transform 1 0 153916 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1673
timestamp 1758069660
transform 1 0 155020 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1679
timestamp 1758069660
transform 1 0 155572 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1681
timestamp 1758069660
transform 1 0 155756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1693
timestamp 1758069660
transform 1 0 156860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1705
timestamp 1758069660
transform 1 0 157964 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1717
timestamp 1758069660
transform 1 0 159068 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1729
timestamp 1758069660
transform 1 0 160172 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1735
timestamp 1758069660
transform 1 0 160724 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1737
timestamp 1758069660
transform 1 0 160908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1749
timestamp 1758069660
transform 1 0 162012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1761
timestamp 1758069660
transform 1 0 163116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1773
timestamp 1758069660
transform 1 0 164220 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1785
timestamp 1758069660
transform 1 0 165324 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1791
timestamp 1758069660
transform 1 0 165876 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1793
timestamp 1758069660
transform 1 0 166060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1805
timestamp 1758069660
transform 1 0 167164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1817
timestamp 1758069660
transform 1 0 168268 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1829
timestamp 1758069660
transform 1 0 169372 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1841
timestamp 1758069660
transform 1 0 170476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1847
timestamp 1758069660
transform 1 0 171028 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1849
timestamp 1758069660
transform 1 0 171212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1861
timestamp 1758069660
transform 1 0 172316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1873
timestamp 1758069660
transform 1 0 173420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1885
timestamp 1758069660
transform 1 0 174524 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1897
timestamp 1758069660
transform 1 0 175628 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1903
timestamp 1758069660
transform 1 0 176180 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1905
timestamp 1758069660
transform 1 0 176364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1917
timestamp 1758069660
transform 1 0 177468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1929
timestamp 1758069660
transform 1 0 178572 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1941
timestamp 1758069660
transform 1 0 179676 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1953
timestamp 1758069660
transform 1 0 180780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1959
timestamp 1758069660
transform 1 0 181332 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1961
timestamp 1758069660
transform 1 0 181516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1973
timestamp 1758069660
transform 1 0 182620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1985
timestamp 1758069660
transform 1 0 183724 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1997
timestamp 1758069660
transform 1 0 184828 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2009
timestamp 1758069660
transform 1 0 185932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2015
timestamp 1758069660
transform 1 0 186484 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2017
timestamp 1758069660
transform 1 0 186668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2029
timestamp 1758069660
transform 1 0 187772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2041
timestamp 1758069660
transform 1 0 188876 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2053
timestamp 1758069660
transform 1 0 189980 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2065
timestamp 1758069660
transform 1 0 191084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2071
timestamp 1758069660
transform 1 0 191636 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2073
timestamp 1758069660
transform 1 0 191820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2085
timestamp 1758069660
transform 1 0 192924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2097
timestamp 1758069660
transform 1 0 194028 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2109
timestamp 1758069660
transform 1 0 195132 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2121
timestamp 1758069660
transform 1 0 196236 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2127
timestamp 1758069660
transform 1 0 196788 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2129
timestamp 1758069660
transform 1 0 196972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2141
timestamp 1758069660
transform 1 0 198076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2153
timestamp 1758069660
transform 1 0 199180 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2165
timestamp 1758069660
transform 1 0 200284 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2177
timestamp 1758069660
transform 1 0 201388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2183
timestamp 1758069660
transform 1 0 201940 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2185
timestamp 1758069660
transform 1 0 202124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2197
timestamp 1758069660
transform 1 0 203228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2209
timestamp 1758069660
transform 1 0 204332 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2221
timestamp 1758069660
transform 1 0 205436 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2233
timestamp 1758069660
transform 1 0 206540 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2239
timestamp 1758069660
transform 1 0 207092 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2241
timestamp 1758069660
transform 1 0 207276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2253
timestamp 1758069660
transform 1 0 208380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2265
timestamp 1758069660
transform 1 0 209484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2277
timestamp 1758069660
transform 1 0 210588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2289
timestamp 1758069660
transform 1 0 211692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2295
timestamp 1758069660
transform 1 0 212244 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2297
timestamp 1758069660
transform 1 0 212428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2309
timestamp 1758069660
transform 1 0 213532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2321
timestamp 1758069660
transform 1 0 214636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2333
timestamp 1758069660
transform 1 0 215740 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2345
timestamp 1758069660
transform 1 0 216844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2351
timestamp 1758069660
transform 1 0 217396 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2353
timestamp 1758069660
transform 1 0 217580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2365
timestamp 1758069660
transform 1 0 218684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2377
timestamp 1758069660
transform 1 0 219788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2389
timestamp 1758069660
transform 1 0 220892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2401
timestamp 1758069660
transform 1 0 221996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2407
timestamp 1758069660
transform 1 0 222548 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2409
timestamp 1758069660
transform 1 0 222732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2421
timestamp 1758069660
transform 1 0 223836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2433
timestamp 1758069660
transform 1 0 224940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2445
timestamp 1758069660
transform 1 0 226044 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2457
timestamp 1758069660
transform 1 0 227148 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2463
timestamp 1758069660
transform 1 0 227700 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2465
timestamp 1758069660
transform 1 0 227884 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2477
timestamp 1758069660
transform 1 0 228988 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2489
timestamp 1758069660
transform 1 0 230092 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2501
timestamp 1758069660
transform 1 0 231196 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2513
timestamp 1758069660
transform 1 0 232300 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2519
timestamp 1758069660
transform 1 0 232852 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2521
timestamp 1758069660
transform 1 0 233036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2533
timestamp 1758069660
transform 1 0 234140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2545
timestamp 1758069660
transform 1 0 235244 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2557
timestamp 1758069660
transform 1 0 236348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2569
timestamp 1758069660
transform 1 0 237452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2575
timestamp 1758069660
transform 1 0 238004 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2577
timestamp 1758069660
transform 1 0 238188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2589
timestamp 1758069660
transform 1 0 239292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2601
timestamp 1758069660
transform 1 0 240396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2613
timestamp 1758069660
transform 1 0 241500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2625
timestamp 1758069660
transform 1 0 242604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2631
timestamp 1758069660
transform 1 0 243156 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2633
timestamp 1758069660
transform 1 0 243340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2645
timestamp 1758069660
transform 1 0 244444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2657
timestamp 1758069660
transform 1 0 245548 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2669
timestamp 1758069660
transform 1 0 246652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2681
timestamp 1758069660
transform 1 0 247756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2687
timestamp 1758069660
transform 1 0 248308 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2689
timestamp 1758069660
transform 1 0 248492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2701
timestamp 1758069660
transform 1 0 249596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2713
timestamp 1758069660
transform 1 0 250700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2725
timestamp 1758069660
transform 1 0 251804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2737
timestamp 1758069660
transform 1 0 252908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2743
timestamp 1758069660
transform 1 0 253460 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2745
timestamp 1758069660
transform 1 0 253644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2757
timestamp 1758069660
transform 1 0 254748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2769
timestamp 1758069660
transform 1 0 255852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2781
timestamp 1758069660
transform 1 0 256956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2793
timestamp 1758069660
transform 1 0 258060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2799
timestamp 1758069660
transform 1 0 258612 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2801
timestamp 1758069660
transform 1 0 258796 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2813
timestamp 1758069660
transform 1 0 259900 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2825
timestamp 1758069660
transform 1 0 261004 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2837
timestamp 1758069660
transform 1 0 262108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2849
timestamp 1758069660
transform 1 0 263212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2855
timestamp 1758069660
transform 1 0 263764 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2857
timestamp 1758069660
transform 1 0 263948 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2869
timestamp 1758069660
transform 1 0 265052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2881
timestamp 1758069660
transform 1 0 266156 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2893
timestamp 1758069660
transform 1 0 267260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2905
timestamp 1758069660
transform 1 0 268364 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2911
timestamp 1758069660
transform 1 0 268916 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2913
timestamp 1758069660
transform 1 0 269100 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2925
timestamp 1758069660
transform 1 0 270204 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2937
timestamp 1758069660
transform 1 0 271308 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2949
timestamp 1758069660
transform 1 0 272412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2961
timestamp 1758069660
transform 1 0 273516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2967
timestamp 1758069660
transform 1 0 274068 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2969
timestamp 1758069660
transform 1 0 274252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2981
timestamp 1758069660
transform 1 0 275356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2993
timestamp 1758069660
transform 1 0 276460 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3005
timestamp 1758069660
transform 1 0 277564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3017
timestamp 1758069660
transform 1 0 278668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3023
timestamp 1758069660
transform 1 0 279220 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3025
timestamp 1758069660
transform 1 0 279404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3037
timestamp 1758069660
transform 1 0 280508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3049
timestamp 1758069660
transform 1 0 281612 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3061
timestamp 1758069660
transform 1 0 282716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3073
timestamp 1758069660
transform 1 0 283820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3079
timestamp 1758069660
transform 1 0 284372 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3081
timestamp 1758069660
transform 1 0 284556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3093
timestamp 1758069660
transform 1 0 285660 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3105
timestamp 1758069660
transform 1 0 286764 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3117
timestamp 1758069660
transform 1 0 287868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3129
timestamp 1758069660
transform 1 0 288972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3135
timestamp 1758069660
transform 1 0 289524 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3137
timestamp 1758069660
transform 1 0 289708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3149
timestamp 1758069660
transform 1 0 290812 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3161
timestamp 1758069660
transform 1 0 291916 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3173
timestamp 1758069660
transform 1 0 293020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3185
timestamp 1758069660
transform 1 0 294124 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3191
timestamp 1758069660
transform 1 0 294676 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3193
timestamp 1758069660
transform 1 0 294860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3205
timestamp 1758069660
transform 1 0 295964 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3217
timestamp 1758069660
transform 1 0 297068 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3229
timestamp 1758069660
transform 1 0 298172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3241
timestamp 1758069660
transform 1 0 299276 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3247
timestamp 1758069660
transform 1 0 299828 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3249
timestamp 1758069660
transform 1 0 300012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3261
timestamp 1758069660
transform 1 0 301116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3273
timestamp 1758069660
transform 1 0 302220 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3285
timestamp 1758069660
transform 1 0 303324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3297
timestamp 1758069660
transform 1 0 304428 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3303
timestamp 1758069660
transform 1 0 304980 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3305
timestamp 1758069660
transform 1 0 305164 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1758069660
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1758069660
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1758069660
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1758069660
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1758069660
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1758069660
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1758069660
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1758069660
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1758069660
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1758069660
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1758069660
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1758069660
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1758069660
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1758069660
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1758069660
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1758069660
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1758069660
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1758069660
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1758069660
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1758069660
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1758069660
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1758069660
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1758069660
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1758069660
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1758069660
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1758069660
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1758069660
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1758069660
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1758069660
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1758069660
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1758069660
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1758069660
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1758069660
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1758069660
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1758069660
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1758069660
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1758069660
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1758069660
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1758069660
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1758069660
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1758069660
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1758069660
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1758069660
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1758069660
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1758069660
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1758069660
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1758069660
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1758069660
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1758069660
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1758069660
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1758069660
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1758069660
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1758069660
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1758069660
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1758069660
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1758069660
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1758069660
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1758069660
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1758069660
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1758069660
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1758069660
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1758069660
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1758069660
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1758069660
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1758069660
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1758069660
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1758069660
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1758069660
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1758069660
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1758069660
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1758069660
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1758069660
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1758069660
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1758069660
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1758069660
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1758069660
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1758069660
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1758069660
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1758069660
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1758069660
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1758069660
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1758069660
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1758069660
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1758069660
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1758069660
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1758069660
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1758069660
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_813
timestamp 1758069660
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_825
timestamp 1758069660
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_837
timestamp 1758069660
transform 1 0 78108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_849
timestamp 1758069660
transform 1 0 79212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_861
timestamp 1758069660
transform 1 0 80316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_867
timestamp 1758069660
transform 1 0 80868 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_869
timestamp 1758069660
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_881
timestamp 1758069660
transform 1 0 82156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_893
timestamp 1758069660
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_905
timestamp 1758069660
transform 1 0 84364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1758069660
transform 1 0 85468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1758069660
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_925
timestamp 1758069660
transform 1 0 86204 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_937
timestamp 1758069660
transform 1 0 87308 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_949
timestamp 1758069660
transform 1 0 88412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_961
timestamp 1758069660
transform 1 0 89516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_973
timestamp 1758069660
transform 1 0 90620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_979
timestamp 1758069660
transform 1 0 91172 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_981
timestamp 1758069660
transform 1 0 91356 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_993
timestamp 1758069660
transform 1 0 92460 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1005
timestamp 1758069660
transform 1 0 93564 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1017
timestamp 1758069660
transform 1 0 94668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1029
timestamp 1758069660
transform 1 0 95772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1035
timestamp 1758069660
transform 1 0 96324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1037
timestamp 1758069660
transform 1 0 96508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1049
timestamp 1758069660
transform 1 0 97612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1061
timestamp 1758069660
transform 1 0 98716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1073
timestamp 1758069660
transform 1 0 99820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1085
timestamp 1758069660
transform 1 0 100924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1091
timestamp 1758069660
transform 1 0 101476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1093
timestamp 1758069660
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1105
timestamp 1758069660
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1117
timestamp 1758069660
transform 1 0 103868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1129
timestamp 1758069660
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1141
timestamp 1758069660
transform 1 0 106076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1147
timestamp 1758069660
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1149
timestamp 1758069660
transform 1 0 106812 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1161
timestamp 1758069660
transform 1 0 107916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1173
timestamp 1758069660
transform 1 0 109020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1185
timestamp 1758069660
transform 1 0 110124 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1197
timestamp 1758069660
transform 1 0 111228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1203
timestamp 1758069660
transform 1 0 111780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1205
timestamp 1758069660
transform 1 0 111964 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1217
timestamp 1758069660
transform 1 0 113068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1229
timestamp 1758069660
transform 1 0 114172 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1241
timestamp 1758069660
transform 1 0 115276 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1253
timestamp 1758069660
transform 1 0 116380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1259
timestamp 1758069660
transform 1 0 116932 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1261
timestamp 1758069660
transform 1 0 117116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1273
timestamp 1758069660
transform 1 0 118220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1285
timestamp 1758069660
transform 1 0 119324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1297
timestamp 1758069660
transform 1 0 120428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1309
timestamp 1758069660
transform 1 0 121532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1315
timestamp 1758069660
transform 1 0 122084 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1317
timestamp 1758069660
transform 1 0 122268 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1329
timestamp 1758069660
transform 1 0 123372 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1341
timestamp 1758069660
transform 1 0 124476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1353
timestamp 1758069660
transform 1 0 125580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1365
timestamp 1758069660
transform 1 0 126684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1371
timestamp 1758069660
transform 1 0 127236 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1373
timestamp 1758069660
transform 1 0 127420 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1385
timestamp 1758069660
transform 1 0 128524 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1397
timestamp 1758069660
transform 1 0 129628 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1409
timestamp 1758069660
transform 1 0 130732 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1421
timestamp 1758069660
transform 1 0 131836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1427
timestamp 1758069660
transform 1 0 132388 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1429
timestamp 1758069660
transform 1 0 132572 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1441
timestamp 1758069660
transform 1 0 133676 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1453
timestamp 1758069660
transform 1 0 134780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1465
timestamp 1758069660
transform 1 0 135884 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1477
timestamp 1758069660
transform 1 0 136988 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1483
timestamp 1758069660
transform 1 0 137540 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1485
timestamp 1758069660
transform 1 0 137724 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1497
timestamp 1758069660
transform 1 0 138828 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1509
timestamp 1758069660
transform 1 0 139932 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1521
timestamp 1758069660
transform 1 0 141036 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1533
timestamp 1758069660
transform 1 0 142140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1539
timestamp 1758069660
transform 1 0 142692 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1541
timestamp 1758069660
transform 1 0 142876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1553
timestamp 1758069660
transform 1 0 143980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1565
timestamp 1758069660
transform 1 0 145084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1577
timestamp 1758069660
transform 1 0 146188 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1589
timestamp 1758069660
transform 1 0 147292 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1595
timestamp 1758069660
transform 1 0 147844 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1597
timestamp 1758069660
transform 1 0 148028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1609
timestamp 1758069660
transform 1 0 149132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1621
timestamp 1758069660
transform 1 0 150236 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1633
timestamp 1758069660
transform 1 0 151340 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1645
timestamp 1758069660
transform 1 0 152444 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1651
timestamp 1758069660
transform 1 0 152996 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1653
timestamp 1758069660
transform 1 0 153180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1665
timestamp 1758069660
transform 1 0 154284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1677
timestamp 1758069660
transform 1 0 155388 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1689
timestamp 1758069660
transform 1 0 156492 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1701
timestamp 1758069660
transform 1 0 157596 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1707
timestamp 1758069660
transform 1 0 158148 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1709
timestamp 1758069660
transform 1 0 158332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1721
timestamp 1758069660
transform 1 0 159436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1733
timestamp 1758069660
transform 1 0 160540 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1745
timestamp 1758069660
transform 1 0 161644 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1757
timestamp 1758069660
transform 1 0 162748 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1763
timestamp 1758069660
transform 1 0 163300 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1765
timestamp 1758069660
transform 1 0 163484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1777
timestamp 1758069660
transform 1 0 164588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1789
timestamp 1758069660
transform 1 0 165692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1801
timestamp 1758069660
transform 1 0 166796 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1813
timestamp 1758069660
transform 1 0 167900 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1819
timestamp 1758069660
transform 1 0 168452 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1821
timestamp 1758069660
transform 1 0 168636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1833
timestamp 1758069660
transform 1 0 169740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1845
timestamp 1758069660
transform 1 0 170844 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1857
timestamp 1758069660
transform 1 0 171948 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1869
timestamp 1758069660
transform 1 0 173052 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1875
timestamp 1758069660
transform 1 0 173604 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1877
timestamp 1758069660
transform 1 0 173788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1889
timestamp 1758069660
transform 1 0 174892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1901
timestamp 1758069660
transform 1 0 175996 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1913
timestamp 1758069660
transform 1 0 177100 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1925
timestamp 1758069660
transform 1 0 178204 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1931
timestamp 1758069660
transform 1 0 178756 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1933
timestamp 1758069660
transform 1 0 178940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1945
timestamp 1758069660
transform 1 0 180044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1957
timestamp 1758069660
transform 1 0 181148 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1969
timestamp 1758069660
transform 1 0 182252 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1981
timestamp 1758069660
transform 1 0 183356 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1987
timestamp 1758069660
transform 1 0 183908 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1989
timestamp 1758069660
transform 1 0 184092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2001
timestamp 1758069660
transform 1 0 185196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2013
timestamp 1758069660
transform 1 0 186300 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2025
timestamp 1758069660
transform 1 0 187404 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2037
timestamp 1758069660
transform 1 0 188508 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2043
timestamp 1758069660
transform 1 0 189060 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2045
timestamp 1758069660
transform 1 0 189244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2057
timestamp 1758069660
transform 1 0 190348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2069
timestamp 1758069660
transform 1 0 191452 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2081
timestamp 1758069660
transform 1 0 192556 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2093
timestamp 1758069660
transform 1 0 193660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2099
timestamp 1758069660
transform 1 0 194212 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2101
timestamp 1758069660
transform 1 0 194396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2113
timestamp 1758069660
transform 1 0 195500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2125
timestamp 1758069660
transform 1 0 196604 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2137
timestamp 1758069660
transform 1 0 197708 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2149
timestamp 1758069660
transform 1 0 198812 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2155
timestamp 1758069660
transform 1 0 199364 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2157
timestamp 1758069660
transform 1 0 199548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2169
timestamp 1758069660
transform 1 0 200652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2181
timestamp 1758069660
transform 1 0 201756 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2193
timestamp 1758069660
transform 1 0 202860 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2205
timestamp 1758069660
transform 1 0 203964 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2211
timestamp 1758069660
transform 1 0 204516 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2213
timestamp 1758069660
transform 1 0 204700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2225
timestamp 1758069660
transform 1 0 205804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2237
timestamp 1758069660
transform 1 0 206908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2249
timestamp 1758069660
transform 1 0 208012 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2261
timestamp 1758069660
transform 1 0 209116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2267
timestamp 1758069660
transform 1 0 209668 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2269
timestamp 1758069660
transform 1 0 209852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2281
timestamp 1758069660
transform 1 0 210956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2293
timestamp 1758069660
transform 1 0 212060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2305
timestamp 1758069660
transform 1 0 213164 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2317
timestamp 1758069660
transform 1 0 214268 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2323
timestamp 1758069660
transform 1 0 214820 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2325
timestamp 1758069660
transform 1 0 215004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2337
timestamp 1758069660
transform 1 0 216108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2349
timestamp 1758069660
transform 1 0 217212 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2361
timestamp 1758069660
transform 1 0 218316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2373
timestamp 1758069660
transform 1 0 219420 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2379
timestamp 1758069660
transform 1 0 219972 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2381
timestamp 1758069660
transform 1 0 220156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2393
timestamp 1758069660
transform 1 0 221260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2405
timestamp 1758069660
transform 1 0 222364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2417
timestamp 1758069660
transform 1 0 223468 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2429
timestamp 1758069660
transform 1 0 224572 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2435
timestamp 1758069660
transform 1 0 225124 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2437
timestamp 1758069660
transform 1 0 225308 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2449
timestamp 1758069660
transform 1 0 226412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2461
timestamp 1758069660
transform 1 0 227516 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2473
timestamp 1758069660
transform 1 0 228620 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2485
timestamp 1758069660
transform 1 0 229724 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2491
timestamp 1758069660
transform 1 0 230276 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2493
timestamp 1758069660
transform 1 0 230460 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2505
timestamp 1758069660
transform 1 0 231564 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2517
timestamp 1758069660
transform 1 0 232668 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2529
timestamp 1758069660
transform 1 0 233772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2541
timestamp 1758069660
transform 1 0 234876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2547
timestamp 1758069660
transform 1 0 235428 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2549
timestamp 1758069660
transform 1 0 235612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2561
timestamp 1758069660
transform 1 0 236716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2573
timestamp 1758069660
transform 1 0 237820 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2585
timestamp 1758069660
transform 1 0 238924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2597
timestamp 1758069660
transform 1 0 240028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2603
timestamp 1758069660
transform 1 0 240580 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2605
timestamp 1758069660
transform 1 0 240764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2617
timestamp 1758069660
transform 1 0 241868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2629
timestamp 1758069660
transform 1 0 242972 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2641
timestamp 1758069660
transform 1 0 244076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2653
timestamp 1758069660
transform 1 0 245180 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2659
timestamp 1758069660
transform 1 0 245732 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2661
timestamp 1758069660
transform 1 0 245916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2673
timestamp 1758069660
transform 1 0 247020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2685
timestamp 1758069660
transform 1 0 248124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2697
timestamp 1758069660
transform 1 0 249228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2709
timestamp 1758069660
transform 1 0 250332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2715
timestamp 1758069660
transform 1 0 250884 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2717
timestamp 1758069660
transform 1 0 251068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2729
timestamp 1758069660
transform 1 0 252172 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2741
timestamp 1758069660
transform 1 0 253276 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2753
timestamp 1758069660
transform 1 0 254380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2765
timestamp 1758069660
transform 1 0 255484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2771
timestamp 1758069660
transform 1 0 256036 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2773
timestamp 1758069660
transform 1 0 256220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2785
timestamp 1758069660
transform 1 0 257324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2797
timestamp 1758069660
transform 1 0 258428 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2809
timestamp 1758069660
transform 1 0 259532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2821
timestamp 1758069660
transform 1 0 260636 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2827
timestamp 1758069660
transform 1 0 261188 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2829
timestamp 1758069660
transform 1 0 261372 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2841
timestamp 1758069660
transform 1 0 262476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2853
timestamp 1758069660
transform 1 0 263580 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2865
timestamp 1758069660
transform 1 0 264684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2877
timestamp 1758069660
transform 1 0 265788 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2883
timestamp 1758069660
transform 1 0 266340 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2885
timestamp 1758069660
transform 1 0 266524 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2897
timestamp 1758069660
transform 1 0 267628 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2909
timestamp 1758069660
transform 1 0 268732 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2921
timestamp 1758069660
transform 1 0 269836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2933
timestamp 1758069660
transform 1 0 270940 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2939
timestamp 1758069660
transform 1 0 271492 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2941
timestamp 1758069660
transform 1 0 271676 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2953
timestamp 1758069660
transform 1 0 272780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2965
timestamp 1758069660
transform 1 0 273884 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2977
timestamp 1758069660
transform 1 0 274988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2989
timestamp 1758069660
transform 1 0 276092 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2995
timestamp 1758069660
transform 1 0 276644 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2997
timestamp 1758069660
transform 1 0 276828 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3009
timestamp 1758069660
transform 1 0 277932 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3021
timestamp 1758069660
transform 1 0 279036 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3033
timestamp 1758069660
transform 1 0 280140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3045
timestamp 1758069660
transform 1 0 281244 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3051
timestamp 1758069660
transform 1 0 281796 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3053
timestamp 1758069660
transform 1 0 281980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3065
timestamp 1758069660
transform 1 0 283084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3077
timestamp 1758069660
transform 1 0 284188 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3089
timestamp 1758069660
transform 1 0 285292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3101
timestamp 1758069660
transform 1 0 286396 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3107
timestamp 1758069660
transform 1 0 286948 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3109
timestamp 1758069660
transform 1 0 287132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3121
timestamp 1758069660
transform 1 0 288236 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3133
timestamp 1758069660
transform 1 0 289340 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3145
timestamp 1758069660
transform 1 0 290444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3157
timestamp 1758069660
transform 1 0 291548 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3163
timestamp 1758069660
transform 1 0 292100 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3165
timestamp 1758069660
transform 1 0 292284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3177
timestamp 1758069660
transform 1 0 293388 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3189
timestamp 1758069660
transform 1 0 294492 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3201
timestamp 1758069660
transform 1 0 295596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3213
timestamp 1758069660
transform 1 0 296700 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3219
timestamp 1758069660
transform 1 0 297252 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3221
timestamp 1758069660
transform 1 0 297436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3233
timestamp 1758069660
transform 1 0 298540 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3245
timestamp 1758069660
transform 1 0 299644 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3257
timestamp 1758069660
transform 1 0 300748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3269
timestamp 1758069660
transform 1 0 301852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3275
timestamp 1758069660
transform 1 0 302404 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3277
timestamp 1758069660
transform 1 0 302588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3289
timestamp 1758069660
transform 1 0 303692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3301
timestamp 1758069660
transform 1 0 304796 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1758069660
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1758069660
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1758069660
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1758069660
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1758069660
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1758069660
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1758069660
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1758069660
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1758069660
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1758069660
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1758069660
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1758069660
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1758069660
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1758069660
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1758069660
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1758069660
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1758069660
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1758069660
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1758069660
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1758069660
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1758069660
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1758069660
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1758069660
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1758069660
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1758069660
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1758069660
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1758069660
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1758069660
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1758069660
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1758069660
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1758069660
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1758069660
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1758069660
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_317
timestamp 1758069660
transform 1 0 30268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_325
timestamp 1758069660
transform 1 0 31004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1758069660
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1758069660
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_340
timestamp 1758069660
transform 1 0 32384 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_347
timestamp 1758069660
transform 1 0 33028 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_359
timestamp 1758069660
transform 1 0 34132 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_371
timestamp 1758069660
transform 1 0 35236 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_383
timestamp 1758069660
transform 1 0 36340 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1758069660
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1758069660
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1758069660
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1758069660
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1758069660
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1758069660
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1758069660
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1758069660
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1758069660
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1758069660
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1758069660
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1758069660
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1758069660
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1758069660
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1758069660
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1758069660
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1758069660
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1758069660
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1758069660
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1758069660
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1758069660
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1758069660
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1758069660
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1758069660
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1758069660
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1758069660
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1758069660
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1758069660
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1758069660
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1758069660
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1758069660
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1758069660
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1758069660
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1758069660
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1758069660
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1758069660
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1758069660
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1758069660
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1758069660
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1758069660
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1758069660
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1758069660
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1758069660
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1758069660
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1758069660
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1758069660
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_821
timestamp 1758069660
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1758069660
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1758069660
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_841
timestamp 1758069660
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_853
timestamp 1758069660
transform 1 0 79580 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_865
timestamp 1758069660
transform 1 0 80684 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_877
timestamp 1758069660
transform 1 0 81788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_889
timestamp 1758069660
transform 1 0 82892 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_895
timestamp 1758069660
transform 1 0 83444 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_897
timestamp 1758069660
transform 1 0 83628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_909
timestamp 1758069660
transform 1 0 84732 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_921
timestamp 1758069660
transform 1 0 85836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_933
timestamp 1758069660
transform 1 0 86940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_945
timestamp 1758069660
transform 1 0 88044 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_951
timestamp 1758069660
transform 1 0 88596 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_953
timestamp 1758069660
transform 1 0 88780 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_965
timestamp 1758069660
transform 1 0 89884 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_977
timestamp 1758069660
transform 1 0 90988 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_989
timestamp 1758069660
transform 1 0 92092 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1001
timestamp 1758069660
transform 1 0 93196 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1007
timestamp 1758069660
transform 1 0 93748 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1009
timestamp 1758069660
transform 1 0 93932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1021
timestamp 1758069660
transform 1 0 95036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1033
timestamp 1758069660
transform 1 0 96140 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1045
timestamp 1758069660
transform 1 0 97244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1057
timestamp 1758069660
transform 1 0 98348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1063
timestamp 1758069660
transform 1 0 98900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1065
timestamp 1758069660
transform 1 0 99084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1077
timestamp 1758069660
transform 1 0 100188 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1089
timestamp 1758069660
transform 1 0 101292 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1101
timestamp 1758069660
transform 1 0 102396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1113
timestamp 1758069660
transform 1 0 103500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1119
timestamp 1758069660
transform 1 0 104052 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1121
timestamp 1758069660
transform 1 0 104236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1133
timestamp 1758069660
transform 1 0 105340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1145
timestamp 1758069660
transform 1 0 106444 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1157
timestamp 1758069660
transform 1 0 107548 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1169
timestamp 1758069660
transform 1 0 108652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1175
timestamp 1758069660
transform 1 0 109204 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1177
timestamp 1758069660
transform 1 0 109388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1189
timestamp 1758069660
transform 1 0 110492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1201
timestamp 1758069660
transform 1 0 111596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1213
timestamp 1758069660
transform 1 0 112700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1225
timestamp 1758069660
transform 1 0 113804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1231
timestamp 1758069660
transform 1 0 114356 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1233
timestamp 1758069660
transform 1 0 114540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1245
timestamp 1758069660
transform 1 0 115644 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1257
timestamp 1758069660
transform 1 0 116748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1269
timestamp 1758069660
transform 1 0 117852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1281
timestamp 1758069660
transform 1 0 118956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1287
timestamp 1758069660
transform 1 0 119508 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1289
timestamp 1758069660
transform 1 0 119692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1301
timestamp 1758069660
transform 1 0 120796 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1313
timestamp 1758069660
transform 1 0 121900 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1325
timestamp 1758069660
transform 1 0 123004 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1337
timestamp 1758069660
transform 1 0 124108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1343
timestamp 1758069660
transform 1 0 124660 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1345
timestamp 1758069660
transform 1 0 124844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1357
timestamp 1758069660
transform 1 0 125948 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1369
timestamp 1758069660
transform 1 0 127052 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1381
timestamp 1758069660
transform 1 0 128156 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1393
timestamp 1758069660
transform 1 0 129260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1399
timestamp 1758069660
transform 1 0 129812 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1401
timestamp 1758069660
transform 1 0 129996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1413
timestamp 1758069660
transform 1 0 131100 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1425
timestamp 1758069660
transform 1 0 132204 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1437
timestamp 1758069660
transform 1 0 133308 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1449
timestamp 1758069660
transform 1 0 134412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1455
timestamp 1758069660
transform 1 0 134964 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1457
timestamp 1758069660
transform 1 0 135148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1469
timestamp 1758069660
transform 1 0 136252 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1481
timestamp 1758069660
transform 1 0 137356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1493
timestamp 1758069660
transform 1 0 138460 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1505
timestamp 1758069660
transform 1 0 139564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1511
timestamp 1758069660
transform 1 0 140116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1513
timestamp 1758069660
transform 1 0 140300 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1537
timestamp 1758069660
transform 1 0 142508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1549
timestamp 1758069660
transform 1 0 143612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1561
timestamp 1758069660
transform 1 0 144716 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1567
timestamp 1758069660
transform 1 0 145268 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1569
timestamp 1758069660
transform 1 0 145452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1581
timestamp 1758069660
transform 1 0 146556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1593
timestamp 1758069660
transform 1 0 147660 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1605
timestamp 1758069660
transform 1 0 148764 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1617
timestamp 1758069660
transform 1 0 149868 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1623
timestamp 1758069660
transform 1 0 150420 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1625
timestamp 1758069660
transform 1 0 150604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1637
timestamp 1758069660
transform 1 0 151708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1649
timestamp 1758069660
transform 1 0 152812 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1661
timestamp 1758069660
transform 1 0 153916 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1673
timestamp 1758069660
transform 1 0 155020 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1679
timestamp 1758069660
transform 1 0 155572 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1681
timestamp 1758069660
transform 1 0 155756 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1705
timestamp 1758069660
transform 1 0 157964 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1717
timestamp 1758069660
transform 1 0 159068 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1729
timestamp 1758069660
transform 1 0 160172 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1735
timestamp 1758069660
transform 1 0 160724 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1737
timestamp 1758069660
transform 1 0 160908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1749
timestamp 1758069660
transform 1 0 162012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1761
timestamp 1758069660
transform 1 0 163116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1773
timestamp 1758069660
transform 1 0 164220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1785
timestamp 1758069660
transform 1 0 165324 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1791
timestamp 1758069660
transform 1 0 165876 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1793
timestamp 1758069660
transform 1 0 166060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1805
timestamp 1758069660
transform 1 0 167164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1817
timestamp 1758069660
transform 1 0 168268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1829
timestamp 1758069660
transform 1 0 169372 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1841
timestamp 1758069660
transform 1 0 170476 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1847
timestamp 1758069660
transform 1 0 171028 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1849
timestamp 1758069660
transform 1 0 171212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1861
timestamp 1758069660
transform 1 0 172316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1873
timestamp 1758069660
transform 1 0 173420 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1885
timestamp 1758069660
transform 1 0 174524 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1897
timestamp 1758069660
transform 1 0 175628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1903
timestamp 1758069660
transform 1 0 176180 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1905
timestamp 1758069660
transform 1 0 176364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1917
timestamp 1758069660
transform 1 0 177468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1929
timestamp 1758069660
transform 1 0 178572 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1941
timestamp 1758069660
transform 1 0 179676 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1953
timestamp 1758069660
transform 1 0 180780 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1959
timestamp 1758069660
transform 1 0 181332 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1961
timestamp 1758069660
transform 1 0 181516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1973
timestamp 1758069660
transform 1 0 182620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1985
timestamp 1758069660
transform 1 0 183724 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1997
timestamp 1758069660
transform 1 0 184828 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2009
timestamp 1758069660
transform 1 0 185932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2015
timestamp 1758069660
transform 1 0 186484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2017
timestamp 1758069660
transform 1 0 186668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2029
timestamp 1758069660
transform 1 0 187772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2041
timestamp 1758069660
transform 1 0 188876 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2053
timestamp 1758069660
transform 1 0 189980 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2065
timestamp 1758069660
transform 1 0 191084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2071
timestamp 1758069660
transform 1 0 191636 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2073
timestamp 1758069660
transform 1 0 191820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2077
timestamp 1758069660
transform 1 0 192188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2081
timestamp 1758069660
transform 1 0 192556 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2088
timestamp 1758069660
transform 1 0 193200 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2100
timestamp 1758069660
transform 1 0 194304 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2112
timestamp 1758069660
transform 1 0 195408 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2124
timestamp 1758069660
transform 1 0 196512 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2129
timestamp 1758069660
transform 1 0 196972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2141
timestamp 1758069660
transform 1 0 198076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2153
timestamp 1758069660
transform 1 0 199180 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2165
timestamp 1758069660
transform 1 0 200284 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2177
timestamp 1758069660
transform 1 0 201388 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2183
timestamp 1758069660
transform 1 0 201940 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2185
timestamp 1758069660
transform 1 0 202124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2197
timestamp 1758069660
transform 1 0 203228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2209
timestamp 1758069660
transform 1 0 204332 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2221
timestamp 1758069660
transform 1 0 205436 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2233
timestamp 1758069660
transform 1 0 206540 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2239
timestamp 1758069660
transform 1 0 207092 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2241
timestamp 1758069660
transform 1 0 207276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2253
timestamp 1758069660
transform 1 0 208380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2265
timestamp 1758069660
transform 1 0 209484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2277
timestamp 1758069660
transform 1 0 210588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2289
timestamp 1758069660
transform 1 0 211692 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2295
timestamp 1758069660
transform 1 0 212244 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2297
timestamp 1758069660
transform 1 0 212428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2309
timestamp 1758069660
transform 1 0 213532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2321
timestamp 1758069660
transform 1 0 214636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2333
timestamp 1758069660
transform 1 0 215740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2345
timestamp 1758069660
transform 1 0 216844 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2351
timestamp 1758069660
transform 1 0 217396 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2353
timestamp 1758069660
transform 1 0 217580 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2365
timestamp 1758069660
transform 1 0 218684 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2377
timestamp 1758069660
transform 1 0 219788 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2389
timestamp 1758069660
transform 1 0 220892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2401
timestamp 1758069660
transform 1 0 221996 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2407
timestamp 1758069660
transform 1 0 222548 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2409
timestamp 1758069660
transform 1 0 222732 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2421
timestamp 1758069660
transform 1 0 223836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2433
timestamp 1758069660
transform 1 0 224940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2445
timestamp 1758069660
transform 1 0 226044 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2457
timestamp 1758069660
transform 1 0 227148 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2463
timestamp 1758069660
transform 1 0 227700 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2465
timestamp 1758069660
transform 1 0 227884 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2477
timestamp 1758069660
transform 1 0 228988 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2489
timestamp 1758069660
transform 1 0 230092 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2501
timestamp 1758069660
transform 1 0 231196 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2513
timestamp 1758069660
transform 1 0 232300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2519
timestamp 1758069660
transform 1 0 232852 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2521
timestamp 1758069660
transform 1 0 233036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2533
timestamp 1758069660
transform 1 0 234140 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2545
timestamp 1758069660
transform 1 0 235244 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2557
timestamp 1758069660
transform 1 0 236348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2569
timestamp 1758069660
transform 1 0 237452 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2575
timestamp 1758069660
transform 1 0 238004 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2577
timestamp 1758069660
transform 1 0 238188 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2589
timestamp 1758069660
transform 1 0 239292 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2601
timestamp 1758069660
transform 1 0 240396 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2613
timestamp 1758069660
transform 1 0 241500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2625
timestamp 1758069660
transform 1 0 242604 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2631
timestamp 1758069660
transform 1 0 243156 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2633
timestamp 1758069660
transform 1 0 243340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2645
timestamp 1758069660
transform 1 0 244444 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2657
timestamp 1758069660
transform 1 0 245548 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2669
timestamp 1758069660
transform 1 0 246652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2681
timestamp 1758069660
transform 1 0 247756 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2687
timestamp 1758069660
transform 1 0 248308 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2689
timestamp 1758069660
transform 1 0 248492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2701
timestamp 1758069660
transform 1 0 249596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2713
timestamp 1758069660
transform 1 0 250700 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2725
timestamp 1758069660
transform 1 0 251804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2737
timestamp 1758069660
transform 1 0 252908 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2743
timestamp 1758069660
transform 1 0 253460 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2745
timestamp 1758069660
transform 1 0 253644 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2757
timestamp 1758069660
transform 1 0 254748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2769
timestamp 1758069660
transform 1 0 255852 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2781
timestamp 1758069660
transform 1 0 256956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2793
timestamp 1758069660
transform 1 0 258060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2799
timestamp 1758069660
transform 1 0 258612 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2801
timestamp 1758069660
transform 1 0 258796 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2813
timestamp 1758069660
transform 1 0 259900 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2825
timestamp 1758069660
transform 1 0 261004 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2837
timestamp 1758069660
transform 1 0 262108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2849
timestamp 1758069660
transform 1 0 263212 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2855
timestamp 1758069660
transform 1 0 263764 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2857
timestamp 1758069660
transform 1 0 263948 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2869
timestamp 1758069660
transform 1 0 265052 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2881
timestamp 1758069660
transform 1 0 266156 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2893
timestamp 1758069660
transform 1 0 267260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2902
timestamp 1758069660
transform 1 0 268088 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2910
timestamp 1758069660
transform 1 0 268824 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2913
timestamp 1758069660
transform 1 0 269100 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2925
timestamp 1758069660
transform 1 0 270204 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2937
timestamp 1758069660
transform 1 0 271308 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2949
timestamp 1758069660
transform 1 0 272412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2961
timestamp 1758069660
transform 1 0 273516 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2967
timestamp 1758069660
transform 1 0 274068 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2969
timestamp 1758069660
transform 1 0 274252 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2981
timestamp 1758069660
transform 1 0 275356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2993
timestamp 1758069660
transform 1 0 276460 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3005
timestamp 1758069660
transform 1 0 277564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3017
timestamp 1758069660
transform 1 0 278668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3023
timestamp 1758069660
transform 1 0 279220 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3025
timestamp 1758069660
transform 1 0 279404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3037
timestamp 1758069660
transform 1 0 280508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3049
timestamp 1758069660
transform 1 0 281612 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3061
timestamp 1758069660
transform 1 0 282716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3073
timestamp 1758069660
transform 1 0 283820 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3079
timestamp 1758069660
transform 1 0 284372 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3081
timestamp 1758069660
transform 1 0 284556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3093
timestamp 1758069660
transform 1 0 285660 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3105
timestamp 1758069660
transform 1 0 286764 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3117
timestamp 1758069660
transform 1 0 287868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3129
timestamp 1758069660
transform 1 0 288972 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3135
timestamp 1758069660
transform 1 0 289524 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3137
timestamp 1758069660
transform 1 0 289708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3149
timestamp 1758069660
transform 1 0 290812 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3161
timestamp 1758069660
transform 1 0 291916 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3173
timestamp 1758069660
transform 1 0 293020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3185
timestamp 1758069660
transform 1 0 294124 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3191
timestamp 1758069660
transform 1 0 294676 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3193
timestamp 1758069660
transform 1 0 294860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3205
timestamp 1758069660
transform 1 0 295964 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3217
timestamp 1758069660
transform 1 0 297068 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3229
timestamp 1758069660
transform 1 0 298172 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3241
timestamp 1758069660
transform 1 0 299276 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3247
timestamp 1758069660
transform 1 0 299828 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3249
timestamp 1758069660
transform 1 0 300012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3261
timestamp 1758069660
transform 1 0 301116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3273
timestamp 1758069660
transform 1 0 302220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3285
timestamp 1758069660
transform 1 0 303324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3297
timestamp 1758069660
transform 1 0 304428 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3303
timestamp 1758069660
transform 1 0 304980 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3305
timestamp 1758069660
transform 1 0 305164 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1758069660
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1758069660
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1758069660
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1758069660
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1758069660
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1758069660
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1758069660
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1758069660
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1758069660
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1758069660
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1758069660
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1758069660
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1758069660
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1758069660
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1758069660
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1758069660
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1758069660
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1758069660
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1758069660
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1758069660
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1758069660
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1758069660
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1758069660
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1758069660
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1758069660
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1758069660
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1758069660
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1758069660
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1758069660
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1758069660
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1758069660
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1758069660
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1758069660
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_309
timestamp 1758069660
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_320
timestamp 1758069660
transform 1 0 30544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_327
timestamp 1758069660
transform 1 0 31188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_334
timestamp 1758069660
transform 1 0 31832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_341
timestamp 1758069660
transform 1 0 32476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_348
timestamp 1758069660
transform 1 0 33120 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_355
timestamp 1758069660
transform 1 0 33764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1758069660
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1758069660
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1758069660
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1758069660
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1758069660
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1758069660
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1758069660
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1758069660
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1758069660
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1758069660
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1758069660
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1758069660
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1758069660
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1758069660
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1758069660
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1758069660
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1758069660
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1758069660
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1758069660
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1758069660
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1758069660
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1758069660
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1758069660
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1758069660
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1758069660
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1758069660
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1758069660
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1758069660
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1758069660
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1758069660
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1758069660
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1758069660
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1758069660
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1758069660
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1758069660
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1758069660
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1758069660
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1758069660
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1758069660
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1758069660
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1758069660
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1758069660
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1758069660
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1758069660
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1758069660
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1758069660
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1758069660
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1758069660
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1758069660
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_813
timestamp 1758069660
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_825
timestamp 1758069660
transform 1 0 77004 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_837
timestamp 1758069660
transform 1 0 78108 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_849
timestamp 1758069660
transform 1 0 79212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_861
timestamp 1758069660
transform 1 0 80316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_867
timestamp 1758069660
transform 1 0 80868 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_869
timestamp 1758069660
transform 1 0 81052 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_881
timestamp 1758069660
transform 1 0 82156 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_893
timestamp 1758069660
transform 1 0 83260 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_905
timestamp 1758069660
transform 1 0 84364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_917
timestamp 1758069660
transform 1 0 85468 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_923
timestamp 1758069660
transform 1 0 86020 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_925
timestamp 1758069660
transform 1 0 86204 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_937
timestamp 1758069660
transform 1 0 87308 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_949
timestamp 1758069660
transform 1 0 88412 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_961
timestamp 1758069660
transform 1 0 89516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_973
timestamp 1758069660
transform 1 0 90620 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_979
timestamp 1758069660
transform 1 0 91172 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_981
timestamp 1758069660
transform 1 0 91356 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_993
timestamp 1758069660
transform 1 0 92460 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1005
timestamp 1758069660
transform 1 0 93564 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1017
timestamp 1758069660
transform 1 0 94668 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1029
timestamp 1758069660
transform 1 0 95772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1035
timestamp 1758069660
transform 1 0 96324 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1037
timestamp 1758069660
transform 1 0 96508 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1049
timestamp 1758069660
transform 1 0 97612 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1061
timestamp 1758069660
transform 1 0 98716 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1073
timestamp 1758069660
transform 1 0 99820 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1085
timestamp 1758069660
transform 1 0 100924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1091
timestamp 1758069660
transform 1 0 101476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1093
timestamp 1758069660
transform 1 0 101660 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1105
timestamp 1758069660
transform 1 0 102764 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1117
timestamp 1758069660
transform 1 0 103868 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1129
timestamp 1758069660
transform 1 0 104972 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1141
timestamp 1758069660
transform 1 0 106076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1147
timestamp 1758069660
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1149
timestamp 1758069660
transform 1 0 106812 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1161
timestamp 1758069660
transform 1 0 107916 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1173
timestamp 1758069660
transform 1 0 109020 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1185
timestamp 1758069660
transform 1 0 110124 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1197
timestamp 1758069660
transform 1 0 111228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1203
timestamp 1758069660
transform 1 0 111780 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1205
timestamp 1758069660
transform 1 0 111964 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1217
timestamp 1758069660
transform 1 0 113068 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1229
timestamp 1758069660
transform 1 0 114172 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1241
timestamp 1758069660
transform 1 0 115276 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1253
timestamp 1758069660
transform 1 0 116380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1259
timestamp 1758069660
transform 1 0 116932 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1261
timestamp 1758069660
transform 1 0 117116 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1273
timestamp 1758069660
transform 1 0 118220 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1285
timestamp 1758069660
transform 1 0 119324 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1297
timestamp 1758069660
transform 1 0 120428 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1309
timestamp 1758069660
transform 1 0 121532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1315
timestamp 1758069660
transform 1 0 122084 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1317
timestamp 1758069660
transform 1 0 122268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1329
timestamp 1758069660
transform 1 0 123372 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1341
timestamp 1758069660
transform 1 0 124476 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1353
timestamp 1758069660
transform 1 0 125580 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1365
timestamp 1758069660
transform 1 0 126684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1371
timestamp 1758069660
transform 1 0 127236 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1373
timestamp 1758069660
transform 1 0 127420 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1385
timestamp 1758069660
transform 1 0 128524 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1397
timestamp 1758069660
transform 1 0 129628 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1409
timestamp 1758069660
transform 1 0 130732 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1421
timestamp 1758069660
transform 1 0 131836 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1427
timestamp 1758069660
transform 1 0 132388 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1429
timestamp 1758069660
transform 1 0 132572 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1441
timestamp 1758069660
transform 1 0 133676 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1453
timestamp 1758069660
transform 1 0 134780 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1465
timestamp 1758069660
transform 1 0 135884 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1477
timestamp 1758069660
transform 1 0 136988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1483
timestamp 1758069660
transform 1 0 137540 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1485
timestamp 1758069660
transform 1 0 137724 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1497
timestamp 1758069660
transform 1 0 138828 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1509
timestamp 1758069660
transform 1 0 139932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1513
timestamp 1758069660
transform 1 0 140300 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1534
timestamp 1758069660
transform 1 0 142232 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1541
timestamp 1758069660
transform 1 0 142876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1553
timestamp 1758069660
transform 1 0 143980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1565
timestamp 1758069660
transform 1 0 145084 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1577
timestamp 1758069660
transform 1 0 146188 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1589
timestamp 1758069660
transform 1 0 147292 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1595
timestamp 1758069660
transform 1 0 147844 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1597
timestamp 1758069660
transform 1 0 148028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1609
timestamp 1758069660
transform 1 0 149132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1621
timestamp 1758069660
transform 1 0 150236 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1633
timestamp 1758069660
transform 1 0 151340 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1645
timestamp 1758069660
transform 1 0 152444 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1651
timestamp 1758069660
transform 1 0 152996 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1653
timestamp 1758069660
transform 1 0 153180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1665
timestamp 1758069660
transform 1 0 154284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1677
timestamp 1758069660
transform 1 0 155388 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1683
timestamp 1758069660
transform 1 0 155940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1704
timestamp 1758069660
transform 1 0 157872 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1709
timestamp 1758069660
transform 1 0 158332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1721
timestamp 1758069660
transform 1 0 159436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1733
timestamp 1758069660
transform 1 0 160540 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1745
timestamp 1758069660
transform 1 0 161644 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1757
timestamp 1758069660
transform 1 0 162748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1763
timestamp 1758069660
transform 1 0 163300 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1765
timestamp 1758069660
transform 1 0 163484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1777
timestamp 1758069660
transform 1 0 164588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1789
timestamp 1758069660
transform 1 0 165692 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1801
timestamp 1758069660
transform 1 0 166796 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1813
timestamp 1758069660
transform 1 0 167900 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1819
timestamp 1758069660
transform 1 0 168452 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1821
timestamp 1758069660
transform 1 0 168636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1833
timestamp 1758069660
transform 1 0 169740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1845
timestamp 1758069660
transform 1 0 170844 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1857
timestamp 1758069660
transform 1 0 171948 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1869
timestamp 1758069660
transform 1 0 173052 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1875
timestamp 1758069660
transform 1 0 173604 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1877
timestamp 1758069660
transform 1 0 173788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1889
timestamp 1758069660
transform 1 0 174892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1901
timestamp 1758069660
transform 1 0 175996 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1913
timestamp 1758069660
transform 1 0 177100 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1925
timestamp 1758069660
transform 1 0 178204 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1931
timestamp 1758069660
transform 1 0 178756 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1933
timestamp 1758069660
transform 1 0 178940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1945
timestamp 1758069660
transform 1 0 180044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1957
timestamp 1758069660
transform 1 0 181148 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1969
timestamp 1758069660
transform 1 0 182252 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1981
timestamp 1758069660
transform 1 0 183356 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1987
timestamp 1758069660
transform 1 0 183908 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1989
timestamp 1758069660
transform 1 0 184092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2001
timestamp 1758069660
transform 1 0 185196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2013
timestamp 1758069660
transform 1 0 186300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2025
timestamp 1758069660
transform 1 0 187404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2037
timestamp 1758069660
transform 1 0 188508 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2043
timestamp 1758069660
transform 1 0 189060 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2045
timestamp 1758069660
transform 1 0 189244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2057
timestamp 1758069660
transform 1 0 190348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2069
timestamp 1758069660
transform 1 0 191452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2076
timestamp 1758069660
transform 1 0 192096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2083
timestamp 1758069660
transform 1 0 192740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_2090
timestamp 1758069660
transform 1 0 193384 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_2098
timestamp 1758069660
transform 1 0 194120 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2101
timestamp 1758069660
transform 1 0 194396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2113
timestamp 1758069660
transform 1 0 195500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2125
timestamp 1758069660
transform 1 0 196604 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2137
timestamp 1758069660
transform 1 0 197708 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2149
timestamp 1758069660
transform 1 0 198812 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2155
timestamp 1758069660
transform 1 0 199364 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2157
timestamp 1758069660
transform 1 0 199548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2169
timestamp 1758069660
transform 1 0 200652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2181
timestamp 1758069660
transform 1 0 201756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2193
timestamp 1758069660
transform 1 0 202860 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2205
timestamp 1758069660
transform 1 0 203964 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2211
timestamp 1758069660
transform 1 0 204516 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2213
timestamp 1758069660
transform 1 0 204700 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2225
timestamp 1758069660
transform 1 0 205804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2237
timestamp 1758069660
transform 1 0 206908 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2249
timestamp 1758069660
transform 1 0 208012 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2261
timestamp 1758069660
transform 1 0 209116 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2267
timestamp 1758069660
transform 1 0 209668 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2269
timestamp 1758069660
transform 1 0 209852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2281
timestamp 1758069660
transform 1 0 210956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2293
timestamp 1758069660
transform 1 0 212060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2305
timestamp 1758069660
transform 1 0 213164 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2317
timestamp 1758069660
transform 1 0 214268 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2323
timestamp 1758069660
transform 1 0 214820 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2325
timestamp 1758069660
transform 1 0 215004 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2337
timestamp 1758069660
transform 1 0 216108 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2349
timestamp 1758069660
transform 1 0 217212 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2361
timestamp 1758069660
transform 1 0 218316 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2373
timestamp 1758069660
transform 1 0 219420 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2379
timestamp 1758069660
transform 1 0 219972 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2381
timestamp 1758069660
transform 1 0 220156 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2393
timestamp 1758069660
transform 1 0 221260 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2405
timestamp 1758069660
transform 1 0 222364 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2417
timestamp 1758069660
transform 1 0 223468 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2429
timestamp 1758069660
transform 1 0 224572 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2435
timestamp 1758069660
transform 1 0 225124 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2437
timestamp 1758069660
transform 1 0 225308 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2449
timestamp 1758069660
transform 1 0 226412 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2461
timestamp 1758069660
transform 1 0 227516 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2473
timestamp 1758069660
transform 1 0 228620 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2485
timestamp 1758069660
transform 1 0 229724 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2491
timestamp 1758069660
transform 1 0 230276 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2493
timestamp 1758069660
transform 1 0 230460 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2505
timestamp 1758069660
transform 1 0 231564 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2517
timestamp 1758069660
transform 1 0 232668 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2529
timestamp 1758069660
transform 1 0 233772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2541
timestamp 1758069660
transform 1 0 234876 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2547
timestamp 1758069660
transform 1 0 235428 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2549
timestamp 1758069660
transform 1 0 235612 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2561
timestamp 1758069660
transform 1 0 236716 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2573
timestamp 1758069660
transform 1 0 237820 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2585
timestamp 1758069660
transform 1 0 238924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2597
timestamp 1758069660
transform 1 0 240028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2603
timestamp 1758069660
transform 1 0 240580 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2605
timestamp 1758069660
transform 1 0 240764 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2617
timestamp 1758069660
transform 1 0 241868 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2629
timestamp 1758069660
transform 1 0 242972 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2641
timestamp 1758069660
transform 1 0 244076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2653
timestamp 1758069660
transform 1 0 245180 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2659
timestamp 1758069660
transform 1 0 245732 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2661
timestamp 1758069660
transform 1 0 245916 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2673
timestamp 1758069660
transform 1 0 247020 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2685
timestamp 1758069660
transform 1 0 248124 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2697
timestamp 1758069660
transform 1 0 249228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2709
timestamp 1758069660
transform 1 0 250332 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2715
timestamp 1758069660
transform 1 0 250884 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2717
timestamp 1758069660
transform 1 0 251068 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2729
timestamp 1758069660
transform 1 0 252172 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2741
timestamp 1758069660
transform 1 0 253276 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2753
timestamp 1758069660
transform 1 0 254380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2765
timestamp 1758069660
transform 1 0 255484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2771
timestamp 1758069660
transform 1 0 256036 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2773
timestamp 1758069660
transform 1 0 256220 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2785
timestamp 1758069660
transform 1 0 257324 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2797
timestamp 1758069660
transform 1 0 258428 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2809
timestamp 1758069660
transform 1 0 259532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2821
timestamp 1758069660
transform 1 0 260636 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2827
timestamp 1758069660
transform 1 0 261188 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2829
timestamp 1758069660
transform 1 0 261372 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2841
timestamp 1758069660
transform 1 0 262476 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2853
timestamp 1758069660
transform 1 0 263580 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2865
timestamp 1758069660
transform 1 0 264684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2877
timestamp 1758069660
transform 1 0 265788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2883
timestamp 1758069660
transform 1 0 266340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2885
timestamp 1758069660
transform 1 0 266524 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2894
timestamp 1758069660
transform 1 0 267352 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2901
timestamp 1758069660
transform 1 0 267996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2908
timestamp 1758069660
transform 1 0 268640 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2915
timestamp 1758069660
transform 1 0 269284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2927
timestamp 1758069660
transform 1 0 270388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2939
timestamp 1758069660
transform 1 0 271492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2941
timestamp 1758069660
transform 1 0 271676 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2953
timestamp 1758069660
transform 1 0 272780 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2965
timestamp 1758069660
transform 1 0 273884 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2977
timestamp 1758069660
transform 1 0 274988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2989
timestamp 1758069660
transform 1 0 276092 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2995
timestamp 1758069660
transform 1 0 276644 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2997
timestamp 1758069660
transform 1 0 276828 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3009
timestamp 1758069660
transform 1 0 277932 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3021
timestamp 1758069660
transform 1 0 279036 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3033
timestamp 1758069660
transform 1 0 280140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3045
timestamp 1758069660
transform 1 0 281244 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3051
timestamp 1758069660
transform 1 0 281796 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3053
timestamp 1758069660
transform 1 0 281980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3065
timestamp 1758069660
transform 1 0 283084 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3077
timestamp 1758069660
transform 1 0 284188 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3089
timestamp 1758069660
transform 1 0 285292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3101
timestamp 1758069660
transform 1 0 286396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3107
timestamp 1758069660
transform 1 0 286948 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3109
timestamp 1758069660
transform 1 0 287132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3121
timestamp 1758069660
transform 1 0 288236 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3133
timestamp 1758069660
transform 1 0 289340 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3145
timestamp 1758069660
transform 1 0 290444 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3157
timestamp 1758069660
transform 1 0 291548 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3163
timestamp 1758069660
transform 1 0 292100 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3165
timestamp 1758069660
transform 1 0 292284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3177
timestamp 1758069660
transform 1 0 293388 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3189
timestamp 1758069660
transform 1 0 294492 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3201
timestamp 1758069660
transform 1 0 295596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3213
timestamp 1758069660
transform 1 0 296700 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3219
timestamp 1758069660
transform 1 0 297252 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3221
timestamp 1758069660
transform 1 0 297436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3233
timestamp 1758069660
transform 1 0 298540 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3245
timestamp 1758069660
transform 1 0 299644 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3257
timestamp 1758069660
transform 1 0 300748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3269
timestamp 1758069660
transform 1 0 301852 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3275
timestamp 1758069660
transform 1 0 302404 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3277
timestamp 1758069660
transform 1 0 302588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3289
timestamp 1758069660
transform 1 0 303692 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3295
timestamp 1758069660
transform 1 0 304244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3305
timestamp 1758069660
transform 1 0 305164 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1758069660
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1758069660
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1758069660
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1758069660
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1758069660
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1758069660
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1758069660
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1758069660
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1758069660
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1758069660
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1758069660
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1758069660
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1758069660
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1758069660
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1758069660
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1758069660
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1758069660
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1758069660
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1758069660
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1758069660
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1758069660
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1758069660
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1758069660
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1758069660
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1758069660
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1758069660
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1758069660
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1758069660
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1758069660
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1758069660
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1758069660
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1758069660
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_305
timestamp 1758069660
transform 1 0 29164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_309
timestamp 1758069660
transform 1 0 29532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_313
timestamp 1758069660
transform 1 0 29900 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1758069660
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1758069660
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_340
timestamp 1758069660
transform 1 0 32384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_347
timestamp 1758069660
transform 1 0 33028 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_354
timestamp 1758069660
transform 1 0 33672 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_366
timestamp 1758069660
transform 1 0 34776 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_378
timestamp 1758069660
transform 1 0 35880 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1758069660
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1758069660
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1758069660
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1758069660
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1758069660
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1758069660
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1758069660
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1758069660
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1758069660
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1758069660
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1758069660
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1758069660
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1758069660
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1758069660
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1758069660
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1758069660
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1758069660
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1758069660
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1758069660
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1758069660
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1758069660
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1758069660
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1758069660
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1758069660
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1758069660
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1758069660
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1758069660
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1758069660
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1758069660
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1758069660
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1758069660
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1758069660
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1758069660
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1758069660
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1758069660
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1758069660
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1758069660
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1758069660
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1758069660
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1758069660
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1758069660
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1758069660
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1758069660
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1758069660
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1758069660
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1758069660
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_821
timestamp 1758069660
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1758069660
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1758069660
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_841
timestamp 1758069660
transform 1 0 78476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_853
timestamp 1758069660
transform 1 0 79580 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_865
timestamp 1758069660
transform 1 0 80684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_877
timestamp 1758069660
transform 1 0 81788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_889
timestamp 1758069660
transform 1 0 82892 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_895
timestamp 1758069660
transform 1 0 83444 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_897
timestamp 1758069660
transform 1 0 83628 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_909
timestamp 1758069660
transform 1 0 84732 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_921
timestamp 1758069660
transform 1 0 85836 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_933
timestamp 1758069660
transform 1 0 86940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_945
timestamp 1758069660
transform 1 0 88044 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_951
timestamp 1758069660
transform 1 0 88596 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_953
timestamp 1758069660
transform 1 0 88780 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_965
timestamp 1758069660
transform 1 0 89884 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_977
timestamp 1758069660
transform 1 0 90988 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_989
timestamp 1758069660
transform 1 0 92092 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1001
timestamp 1758069660
transform 1 0 93196 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1007
timestamp 1758069660
transform 1 0 93748 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1009
timestamp 1758069660
transform 1 0 93932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1021
timestamp 1758069660
transform 1 0 95036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1033
timestamp 1758069660
transform 1 0 96140 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1045
timestamp 1758069660
transform 1 0 97244 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1057
timestamp 1758069660
transform 1 0 98348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1063
timestamp 1758069660
transform 1 0 98900 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1065
timestamp 1758069660
transform 1 0 99084 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1077
timestamp 1758069660
transform 1 0 100188 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1089
timestamp 1758069660
transform 1 0 101292 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1096
timestamp 1758069660
transform 1 0 101936 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1108
timestamp 1758069660
transform 1 0 103040 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1121
timestamp 1758069660
transform 1 0 104236 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1133
timestamp 1758069660
transform 1 0 105340 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1145
timestamp 1758069660
transform 1 0 106444 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1157
timestamp 1758069660
transform 1 0 107548 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1169
timestamp 1758069660
transform 1 0 108652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1175
timestamp 1758069660
transform 1 0 109204 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1177
timestamp 1758069660
transform 1 0 109388 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1189
timestamp 1758069660
transform 1 0 110492 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1201
timestamp 1758069660
transform 1 0 111596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1213
timestamp 1758069660
transform 1 0 112700 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1225
timestamp 1758069660
transform 1 0 113804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1231
timestamp 1758069660
transform 1 0 114356 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1233
timestamp 1758069660
transform 1 0 114540 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1245
timestamp 1758069660
transform 1 0 115644 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1257
timestamp 1758069660
transform 1 0 116748 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1269
timestamp 1758069660
transform 1 0 117852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1281
timestamp 1758069660
transform 1 0 118956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1287
timestamp 1758069660
transform 1 0 119508 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1289
timestamp 1758069660
transform 1 0 119692 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1301
timestamp 1758069660
transform 1 0 120796 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1313
timestamp 1758069660
transform 1 0 121900 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1325
timestamp 1758069660
transform 1 0 123004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1337
timestamp 1758069660
transform 1 0 124108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1343
timestamp 1758069660
transform 1 0 124660 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1345
timestamp 1758069660
transform 1 0 124844 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1357
timestamp 1758069660
transform 1 0 125948 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1369
timestamp 1758069660
transform 1 0 127052 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1381
timestamp 1758069660
transform 1 0 128156 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1393
timestamp 1758069660
transform 1 0 129260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1399
timestamp 1758069660
transform 1 0 129812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1401
timestamp 1758069660
transform 1 0 129996 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1408
timestamp 1758069660
transform 1 0 130640 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1420
timestamp 1758069660
transform 1 0 131744 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1432
timestamp 1758069660
transform 1 0 132848 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1444
timestamp 1758069660
transform 1 0 133952 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1457
timestamp 1758069660
transform 1 0 135148 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1469
timestamp 1758069660
transform 1 0 136252 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1481
timestamp 1758069660
transform 1 0 137356 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1493
timestamp 1758069660
transform 1 0 138460 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1505
timestamp 1758069660
transform 1 0 139564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1511
timestamp 1758069660
transform 1 0 140116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1513
timestamp 1758069660
transform 1 0 140300 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1537
timestamp 1758069660
transform 1 0 142508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1549
timestamp 1758069660
transform 1 0 143612 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1561
timestamp 1758069660
transform 1 0 144716 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1567
timestamp 1758069660
transform 1 0 145268 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1569
timestamp 1758069660
transform 1 0 145452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1581
timestamp 1758069660
transform 1 0 146556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1593
timestamp 1758069660
transform 1 0 147660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1605
timestamp 1758069660
transform 1 0 148764 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1609
timestamp 1758069660
transform 1 0 149132 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_1621
timestamp 1758069660
transform 1 0 150236 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1628
timestamp 1758069660
transform 1 0 150880 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1640
timestamp 1758069660
transform 1 0 151984 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1652
timestamp 1758069660
transform 1 0 153088 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1664
timestamp 1758069660
transform 1 0 154192 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1676
timestamp 1758069660
transform 1 0 155296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1681
timestamp 1758069660
transform 1 0 155756 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1705
timestamp 1758069660
transform 1 0 157964 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1717
timestamp 1758069660
transform 1 0 159068 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1729
timestamp 1758069660
transform 1 0 160172 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1735
timestamp 1758069660
transform 1 0 160724 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1737
timestamp 1758069660
transform 1 0 160908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1749
timestamp 1758069660
transform 1 0 162012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1761
timestamp 1758069660
transform 1 0 163116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1773
timestamp 1758069660
transform 1 0 164220 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1785
timestamp 1758069660
transform 1 0 165324 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1791
timestamp 1758069660
transform 1 0 165876 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1793
timestamp 1758069660
transform 1 0 166060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1805
timestamp 1758069660
transform 1 0 167164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1817
timestamp 1758069660
transform 1 0 168268 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1829
timestamp 1758069660
transform 1 0 169372 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1841
timestamp 1758069660
transform 1 0 170476 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1847
timestamp 1758069660
transform 1 0 171028 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1849
timestamp 1758069660
transform 1 0 171212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1861
timestamp 1758069660
transform 1 0 172316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1873
timestamp 1758069660
transform 1 0 173420 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1885
timestamp 1758069660
transform 1 0 174524 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1897
timestamp 1758069660
transform 1 0 175628 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1903
timestamp 1758069660
transform 1 0 176180 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1905
timestamp 1758069660
transform 1 0 176364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1917
timestamp 1758069660
transform 1 0 177468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1929
timestamp 1758069660
transform 1 0 178572 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1941
timestamp 1758069660
transform 1 0 179676 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1953
timestamp 1758069660
transform 1 0 180780 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1959
timestamp 1758069660
transform 1 0 181332 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1961
timestamp 1758069660
transform 1 0 181516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1973
timestamp 1758069660
transform 1 0 182620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1985
timestamp 1758069660
transform 1 0 183724 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1997
timestamp 1758069660
transform 1 0 184828 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2009
timestamp 1758069660
transform 1 0 185932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2015
timestamp 1758069660
transform 1 0 186484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2017
timestamp 1758069660
transform 1 0 186668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2021
timestamp 1758069660
transform 1 0 187036 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2031
timestamp 1758069660
transform 1 0 187956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2043
timestamp 1758069660
transform 1 0 189060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2055
timestamp 1758069660
transform 1 0 190164 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_2063
timestamp 1758069660
transform 1 0 190900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2068
timestamp 1758069660
transform 1 0 191360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2076
timestamp 1758069660
transform 1 0 192096 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2086
timestamp 1758069660
transform 1 0 193016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2094
timestamp 1758069660
transform 1 0 193752 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2101
timestamp 1758069660
transform 1 0 194396 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2113
timestamp 1758069660
transform 1 0 195500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_2125
timestamp 1758069660
transform 1 0 196604 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2129
timestamp 1758069660
transform 1 0 196972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2141
timestamp 1758069660
transform 1 0 198076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2153
timestamp 1758069660
transform 1 0 199180 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2165
timestamp 1758069660
transform 1 0 200284 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2177
timestamp 1758069660
transform 1 0 201388 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2183
timestamp 1758069660
transform 1 0 201940 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2185
timestamp 1758069660
transform 1 0 202124 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2196
timestamp 1758069660
transform 1 0 203136 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2208
timestamp 1758069660
transform 1 0 204240 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2220
timestamp 1758069660
transform 1 0 205344 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2232
timestamp 1758069660
transform 1 0 206448 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2241
timestamp 1758069660
transform 1 0 207276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2253
timestamp 1758069660
transform 1 0 208380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2265
timestamp 1758069660
transform 1 0 209484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2277
timestamp 1758069660
transform 1 0 210588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2289
timestamp 1758069660
transform 1 0 211692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2295
timestamp 1758069660
transform 1 0 212244 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2297
timestamp 1758069660
transform 1 0 212428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2309
timestamp 1758069660
transform 1 0 213532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2321
timestamp 1758069660
transform 1 0 214636 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2333
timestamp 1758069660
transform 1 0 215740 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2345
timestamp 1758069660
transform 1 0 216844 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2351
timestamp 1758069660
transform 1 0 217396 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2353
timestamp 1758069660
transform 1 0 217580 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2365
timestamp 1758069660
transform 1 0 218684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2377
timestamp 1758069660
transform 1 0 219788 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2389
timestamp 1758069660
transform 1 0 220892 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2401
timestamp 1758069660
transform 1 0 221996 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2407
timestamp 1758069660
transform 1 0 222548 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2409
timestamp 1758069660
transform 1 0 222732 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2421
timestamp 1758069660
transform 1 0 223836 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2433
timestamp 1758069660
transform 1 0 224940 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2445
timestamp 1758069660
transform 1 0 226044 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2457
timestamp 1758069660
transform 1 0 227148 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2463
timestamp 1758069660
transform 1 0 227700 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2465
timestamp 1758069660
transform 1 0 227884 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2477
timestamp 1758069660
transform 1 0 228988 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2489
timestamp 1758069660
transform 1 0 230092 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2501
timestamp 1758069660
transform 1 0 231196 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2513
timestamp 1758069660
transform 1 0 232300 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2519
timestamp 1758069660
transform 1 0 232852 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2521
timestamp 1758069660
transform 1 0 233036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2533
timestamp 1758069660
transform 1 0 234140 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2545
timestamp 1758069660
transform 1 0 235244 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2557
timestamp 1758069660
transform 1 0 236348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2569
timestamp 1758069660
transform 1 0 237452 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2575
timestamp 1758069660
transform 1 0 238004 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2577
timestamp 1758069660
transform 1 0 238188 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2589
timestamp 1758069660
transform 1 0 239292 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2601
timestamp 1758069660
transform 1 0 240396 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2613
timestamp 1758069660
transform 1 0 241500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2625
timestamp 1758069660
transform 1 0 242604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2631
timestamp 1758069660
transform 1 0 243156 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2633
timestamp 1758069660
transform 1 0 243340 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2645
timestamp 1758069660
transform 1 0 244444 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2657
timestamp 1758069660
transform 1 0 245548 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2669
timestamp 1758069660
transform 1 0 246652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2681
timestamp 1758069660
transform 1 0 247756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2687
timestamp 1758069660
transform 1 0 248308 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2689
timestamp 1758069660
transform 1 0 248492 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2701
timestamp 1758069660
transform 1 0 249596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2713
timestamp 1758069660
transform 1 0 250700 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2725
timestamp 1758069660
transform 1 0 251804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2737
timestamp 1758069660
transform 1 0 252908 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2743
timestamp 1758069660
transform 1 0 253460 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2748
timestamp 1758069660
transform 1 0 253920 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2760
timestamp 1758069660
transform 1 0 255024 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2772
timestamp 1758069660
transform 1 0 256128 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2784
timestamp 1758069660
transform 1 0 257232 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2796
timestamp 1758069660
transform 1 0 258336 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2801
timestamp 1758069660
transform 1 0 258796 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2813
timestamp 1758069660
transform 1 0 259900 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2825
timestamp 1758069660
transform 1 0 261004 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2837
timestamp 1758069660
transform 1 0 262108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2849
timestamp 1758069660
transform 1 0 263212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2855
timestamp 1758069660
transform 1 0 263764 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2857
timestamp 1758069660
transform 1 0 263948 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2869
timestamp 1758069660
transform 1 0 265052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2880
timestamp 1758069660
transform 1 0 266064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2887
timestamp 1758069660
transform 1 0 266708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2894
timestamp 1758069660
transform 1 0 267352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2901
timestamp 1758069660
transform 1 0 267996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2908
timestamp 1758069660
transform 1 0 268640 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2916
timestamp 1758069660
transform 1 0 269376 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2928
timestamp 1758069660
transform 1 0 270480 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2940
timestamp 1758069660
transform 1 0 271584 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2952
timestamp 1758069660
transform 1 0 272688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2964
timestamp 1758069660
transform 1 0 273792 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2969
timestamp 1758069660
transform 1 0 274252 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2981
timestamp 1758069660
transform 1 0 275356 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2993
timestamp 1758069660
transform 1 0 276460 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3005
timestamp 1758069660
transform 1 0 277564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3017
timestamp 1758069660
transform 1 0 278668 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3023
timestamp 1758069660
transform 1 0 279220 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3025
timestamp 1758069660
transform 1 0 279404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3037
timestamp 1758069660
transform 1 0 280508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3049
timestamp 1758069660
transform 1 0 281612 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3061
timestamp 1758069660
transform 1 0 282716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3073
timestamp 1758069660
transform 1 0 283820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3079
timestamp 1758069660
transform 1 0 284372 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3081
timestamp 1758069660
transform 1 0 284556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3093
timestamp 1758069660
transform 1 0 285660 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3105
timestamp 1758069660
transform 1 0 286764 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3117
timestamp 1758069660
transform 1 0 287868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3129
timestamp 1758069660
transform 1 0 288972 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3135
timestamp 1758069660
transform 1 0 289524 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3137
timestamp 1758069660
transform 1 0 289708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3149
timestamp 1758069660
transform 1 0 290812 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3161
timestamp 1758069660
transform 1 0 291916 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3173
timestamp 1758069660
transform 1 0 293020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3185
timestamp 1758069660
transform 1 0 294124 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3191
timestamp 1758069660
transform 1 0 294676 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3193
timestamp 1758069660
transform 1 0 294860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3205
timestamp 1758069660
transform 1 0 295964 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3217
timestamp 1758069660
transform 1 0 297068 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3229
timestamp 1758069660
transform 1 0 298172 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3241
timestamp 1758069660
transform 1 0 299276 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3247
timestamp 1758069660
transform 1 0 299828 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3249
timestamp 1758069660
transform 1 0 300012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3261
timestamp 1758069660
transform 1 0 301116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3273
timestamp 1758069660
transform 1 0 302220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3285
timestamp 1758069660
transform 1 0 303324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3297
timestamp 1758069660
transform 1 0 304428 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3303
timestamp 1758069660
transform 1 0 304980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3305
timestamp 1758069660
transform 1 0 305164 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1758069660
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1758069660
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1758069660
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1758069660
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1758069660
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1758069660
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1758069660
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1758069660
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1758069660
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1758069660
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1758069660
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1758069660
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1758069660
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1758069660
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1758069660
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1758069660
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1758069660
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1758069660
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1758069660
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1758069660
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1758069660
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1758069660
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1758069660
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1758069660
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1758069660
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1758069660
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1758069660
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1758069660
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1758069660
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1758069660
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1758069660
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1758069660
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_309
timestamp 1758069660
transform 1 0 29532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_330
timestamp 1758069660
transform 1 0 31464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_343
timestamp 1758069660
transform 1 0 32660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_351
timestamp 1758069660
transform 1 0 33396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_355
timestamp 1758069660
transform 1 0 33764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1758069660
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1758069660
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1758069660
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1758069660
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1758069660
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1758069660
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1758069660
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_421
timestamp 1758069660
transform 1 0 39836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_425
timestamp 1758069660
transform 1 0 40204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_429
timestamp 1758069660
transform 1 0 40572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_436
timestamp 1758069660
transform 1 0 41216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_443
timestamp 1758069660
transform 1 0 41860 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_450
timestamp 1758069660
transform 1 0 42504 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_462
timestamp 1758069660
transform 1 0 43608 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1758069660
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1758069660
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1758069660
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1758069660
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1758069660
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1758069660
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1758069660
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1758069660
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1758069660
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1758069660
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1758069660
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1758069660
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1758069660
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_592
timestamp 1758069660
transform 1 0 55568 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_598
timestamp 1758069660
transform 1 0 56120 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_602
timestamp 1758069660
transform 1 0 56488 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_614
timestamp 1758069660
transform 1 0 57592 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_626
timestamp 1758069660
transform 1 0 58696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_638
timestamp 1758069660
transform 1 0 59800 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1758069660
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1758069660
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1758069660
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1758069660
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1758069660
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1758069660
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1758069660
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1758069660
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_725
timestamp 1758069660
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_737
timestamp 1758069660
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1758069660
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1758069660
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1758069660
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1758069660
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1758069660
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1758069660
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1758069660
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1758069660
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_813
timestamp 1758069660
transform 1 0 75900 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_822
timestamp 1758069660
transform 1 0 76728 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_834
timestamp 1758069660
transform 1 0 77832 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_841
timestamp 1758069660
transform 1 0 78476 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_853
timestamp 1758069660
transform 1 0 79580 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_865
timestamp 1758069660
transform 1 0 80684 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_869
timestamp 1758069660
transform 1 0 81052 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_881
timestamp 1758069660
transform 1 0 82156 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_893
timestamp 1758069660
transform 1 0 83260 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_905
timestamp 1758069660
transform 1 0 84364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_917
timestamp 1758069660
transform 1 0 85468 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_923
timestamp 1758069660
transform 1 0 86020 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_928
timestamp 1758069660
transform 1 0 86480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_935
timestamp 1758069660
transform 1 0 87124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_939
timestamp 1758069660
transform 1 0 87492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_943
timestamp 1758069660
transform 1 0 87860 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_950
timestamp 1758069660
transform 1 0 88504 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_962
timestamp 1758069660
transform 1 0 89608 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_974
timestamp 1758069660
transform 1 0 90712 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_981
timestamp 1758069660
transform 1 0 91356 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_993
timestamp 1758069660
transform 1 0 92460 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1005
timestamp 1758069660
transform 1 0 93564 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1017
timestamp 1758069660
transform 1 0 94668 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1029
timestamp 1758069660
transform 1 0 95772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1035
timestamp 1758069660
transform 1 0 96324 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1037
timestamp 1758069660
transform 1 0 96508 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1049
timestamp 1758069660
transform 1 0 97612 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1061
timestamp 1758069660
transform 1 0 98716 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1073
timestamp 1758069660
transform 1 0 99820 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1085
timestamp 1758069660
transform 1 0 100924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1091
timestamp 1758069660
transform 1 0 101476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1093
timestamp 1758069660
transform 1 0 101660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1101
timestamp 1758069660
transform 1 0 102396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1105
timestamp 1758069660
transform 1 0 102764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1109
timestamp 1758069660
transform 1 0 103132 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1116
timestamp 1758069660
transform 1 0 103776 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1128
timestamp 1758069660
transform 1 0 104880 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1140
timestamp 1758069660
transform 1 0 105984 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1149
timestamp 1758069660
transform 1 0 106812 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1161
timestamp 1758069660
transform 1 0 107916 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1173
timestamp 1758069660
transform 1 0 109020 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1185
timestamp 1758069660
transform 1 0 110124 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1197
timestamp 1758069660
transform 1 0 111228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1203
timestamp 1758069660
transform 1 0 111780 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1205
timestamp 1758069660
transform 1 0 111964 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1217
timestamp 1758069660
transform 1 0 113068 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1229
timestamp 1758069660
transform 1 0 114172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1244
timestamp 1758069660
transform 1 0 115552 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1248
timestamp 1758069660
transform 1 0 115920 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1252
timestamp 1758069660
transform 1 0 116288 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1264
timestamp 1758069660
transform 1 0 117392 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1276
timestamp 1758069660
transform 1 0 118496 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1288
timestamp 1758069660
transform 1 0 119600 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1300
timestamp 1758069660
transform 1 0 120704 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1312
timestamp 1758069660
transform 1 0 121808 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1317
timestamp 1758069660
transform 1 0 122268 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1329
timestamp 1758069660
transform 1 0 123372 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1341
timestamp 1758069660
transform 1 0 124476 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1353
timestamp 1758069660
transform 1 0 125580 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1365
timestamp 1758069660
transform 1 0 126684 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1371
timestamp 1758069660
transform 1 0 127236 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1373
timestamp 1758069660
transform 1 0 127420 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1385
timestamp 1758069660
transform 1 0 128524 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1397
timestamp 1758069660
transform 1 0 129628 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1405
timestamp 1758069660
transform 1 0 130364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1409
timestamp 1758069660
transform 1 0 130732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1416
timestamp 1758069660
transform 1 0 131376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1423
timestamp 1758069660
transform 1 0 132020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1427
timestamp 1758069660
transform 1 0 132388 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1429
timestamp 1758069660
transform 1 0 132572 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1441
timestamp 1758069660
transform 1 0 133676 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1453
timestamp 1758069660
transform 1 0 134780 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1465
timestamp 1758069660
transform 1 0 135884 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1477
timestamp 1758069660
transform 1 0 136988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1483
timestamp 1758069660
transform 1 0 137540 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1485
timestamp 1758069660
transform 1 0 137724 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1497
timestamp 1758069660
transform 1 0 138828 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1509
timestamp 1758069660
transform 1 0 139932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1513
timestamp 1758069660
transform 1 0 140300 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1534
timestamp 1758069660
transform 1 0 142232 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1541
timestamp 1758069660
transform 1 0 142876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1553
timestamp 1758069660
transform 1 0 143980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1565
timestamp 1758069660
transform 1 0 145084 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1577
timestamp 1758069660
transform 1 0 146188 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1589
timestamp 1758069660
transform 1 0 147292 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1595
timestamp 1758069660
transform 1 0 147844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1606
timestamp 1758069660
transform 1 0 148856 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1612
timestamp 1758069660
transform 1 0 149408 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1619
timestamp 1758069660
transform 1 0 150052 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1630
timestamp 1758069660
transform 1 0 151064 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1642
timestamp 1758069660
transform 1 0 152168 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1650
timestamp 1758069660
transform 1 0 152904 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1653
timestamp 1758069660
transform 1 0 153180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1665
timestamp 1758069660
transform 1 0 154284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1677
timestamp 1758069660
transform 1 0 155388 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1683
timestamp 1758069660
transform 1 0 155940 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1704
timestamp 1758069660
transform 1 0 157872 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1709
timestamp 1758069660
transform 1 0 158332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1721
timestamp 1758069660
transform 1 0 159436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1733
timestamp 1758069660
transform 1 0 160540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1745
timestamp 1758069660
transform 1 0 161644 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1752
timestamp 1758069660
transform 1 0 162288 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1759
timestamp 1758069660
transform 1 0 162932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1763
timestamp 1758069660
transform 1 0 163300 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1768
timestamp 1758069660
transform 1 0 163760 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1780
timestamp 1758069660
transform 1 0 164864 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1792
timestamp 1758069660
transform 1 0 165968 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1804
timestamp 1758069660
transform 1 0 167072 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1816
timestamp 1758069660
transform 1 0 168176 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1821
timestamp 1758069660
transform 1 0 168636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1833
timestamp 1758069660
transform 1 0 169740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1845
timestamp 1758069660
transform 1 0 170844 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1857
timestamp 1758069660
transform 1 0 171948 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1869
timestamp 1758069660
transform 1 0 173052 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1875
timestamp 1758069660
transform 1 0 173604 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1877
timestamp 1758069660
transform 1 0 173788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1889
timestamp 1758069660
transform 1 0 174892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1901
timestamp 1758069660
transform 1 0 175996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1913
timestamp 1758069660
transform 1 0 177100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1920
timestamp 1758069660
transform 1 0 177744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1927
timestamp 1758069660
transform 1 0 178388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1931
timestamp 1758069660
transform 1 0 178756 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1936
timestamp 1758069660
transform 1 0 179216 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1948
timestamp 1758069660
transform 1 0 180320 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1960
timestamp 1758069660
transform 1 0 181424 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1972
timestamp 1758069660
transform 1 0 182528 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1984
timestamp 1758069660
transform 1 0 183632 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1989
timestamp 1758069660
transform 1 0 184092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2001
timestamp 1758069660
transform 1 0 185196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2013
timestamp 1758069660
transform 1 0 186300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2025
timestamp 1758069660
transform 1 0 187404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2037
timestamp 1758069660
transform 1 0 188508 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2043
timestamp 1758069660
transform 1 0 189060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2045
timestamp 1758069660
transform 1 0 189244 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2053
timestamp 1758069660
transform 1 0 189980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2058
timestamp 1758069660
transform 1 0 190440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2065
timestamp 1758069660
transform 1 0 191084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2073
timestamp 1758069660
transform 1 0 191820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2095
timestamp 1758069660
transform 1 0 193844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2099
timestamp 1758069660
transform 1 0 194212 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2110
timestamp 1758069660
transform 1 0 195224 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2117
timestamp 1758069660
transform 1 0 195868 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2129
timestamp 1758069660
transform 1 0 196972 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2141
timestamp 1758069660
transform 1 0 198076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_2153
timestamp 1758069660
transform 1 0 199180 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2157
timestamp 1758069660
transform 1 0 199548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2169
timestamp 1758069660
transform 1 0 200652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2181
timestamp 1758069660
transform 1 0 201756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2188
timestamp 1758069660
transform 1 0 202400 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2195
timestamp 1758069660
transform 1 0 203044 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2202
timestamp 1758069660
transform 1 0 203688 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2210
timestamp 1758069660
transform 1 0 204424 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2216
timestamp 1758069660
transform 1 0 204976 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2228
timestamp 1758069660
transform 1 0 206080 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2240
timestamp 1758069660
transform 1 0 207184 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2252
timestamp 1758069660
transform 1 0 208288 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2264
timestamp 1758069660
transform 1 0 209392 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2269
timestamp 1758069660
transform 1 0 209852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2281
timestamp 1758069660
transform 1 0 210956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2293
timestamp 1758069660
transform 1 0 212060 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2305
timestamp 1758069660
transform 1 0 213164 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2317
timestamp 1758069660
transform 1 0 214268 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2323
timestamp 1758069660
transform 1 0 214820 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2325
timestamp 1758069660
transform 1 0 215004 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2337
timestamp 1758069660
transform 1 0 216108 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2349
timestamp 1758069660
transform 1 0 217212 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2361
timestamp 1758069660
transform 1 0 218316 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2373
timestamp 1758069660
transform 1 0 219420 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2379
timestamp 1758069660
transform 1 0 219972 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2381
timestamp 1758069660
transform 1 0 220156 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2393
timestamp 1758069660
transform 1 0 221260 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2405
timestamp 1758069660
transform 1 0 222364 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2417
timestamp 1758069660
transform 1 0 223468 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2429
timestamp 1758069660
transform 1 0 224572 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2435
timestamp 1758069660
transform 1 0 225124 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2437
timestamp 1758069660
transform 1 0 225308 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2449
timestamp 1758069660
transform 1 0 226412 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2461
timestamp 1758069660
transform 1 0 227516 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2473
timestamp 1758069660
transform 1 0 228620 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2482
timestamp 1758069660
transform 1 0 229448 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2490
timestamp 1758069660
transform 1 0 230184 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2493
timestamp 1758069660
transform 1 0 230460 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2505
timestamp 1758069660
transform 1 0 231564 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2517
timestamp 1758069660
transform 1 0 232668 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2529
timestamp 1758069660
transform 1 0 233772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2541
timestamp 1758069660
transform 1 0 234876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2547
timestamp 1758069660
transform 1 0 235428 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2549
timestamp 1758069660
transform 1 0 235612 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2561
timestamp 1758069660
transform 1 0 236716 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2573
timestamp 1758069660
transform 1 0 237820 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2585
timestamp 1758069660
transform 1 0 238924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2593
timestamp 1758069660
transform 1 0 239660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2598
timestamp 1758069660
transform 1 0 240120 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2608
timestamp 1758069660
transform 1 0 241040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2615
timestamp 1758069660
transform 1 0 241684 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2622
timestamp 1758069660
transform 1 0 242328 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2634
timestamp 1758069660
transform 1 0 243432 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2646
timestamp 1758069660
transform 1 0 244536 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2658
timestamp 1758069660
transform 1 0 245640 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2661
timestamp 1758069660
transform 1 0 245916 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2673
timestamp 1758069660
transform 1 0 247020 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2685
timestamp 1758069660
transform 1 0 248124 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2697
timestamp 1758069660
transform 1 0 249228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2709
timestamp 1758069660
transform 1 0 250332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2715
timestamp 1758069660
transform 1 0 250884 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2717
timestamp 1758069660
transform 1 0 251068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_2729
timestamp 1758069660
transform 1 0 252172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2735
timestamp 1758069660
transform 1 0 252724 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2742
timestamp 1758069660
transform 1 0 253368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2749
timestamp 1758069660
transform 1 0 254012 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2756
timestamp 1758069660
transform 1 0 254656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2768
timestamp 1758069660
transform 1 0 255760 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2773
timestamp 1758069660
transform 1 0 256220 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2785
timestamp 1758069660
transform 1 0 257324 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2797
timestamp 1758069660
transform 1 0 258428 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2809
timestamp 1758069660
transform 1 0 259532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2821
timestamp 1758069660
transform 1 0 260636 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2827
timestamp 1758069660
transform 1 0 261188 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2829
timestamp 1758069660
transform 1 0 261372 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2841
timestamp 1758069660
transform 1 0 262476 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2853
timestamp 1758069660
transform 1 0 263580 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2865
timestamp 1758069660
transform 1 0 264684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2870
timestamp 1758069660
transform 1 0 265144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2877
timestamp 1758069660
transform 1 0 265788 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2883
timestamp 1758069660
transform 1 0 266340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_2885
timestamp 1758069660
transform 1 0 266524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2897
timestamp 1758069660
transform 1 0 267628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2904
timestamp 1758069660
transform 1 0 268272 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2908
timestamp 1758069660
transform 1 0 268640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2919
timestamp 1758069660
transform 1 0 269652 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2932
timestamp 1758069660
transform 1 0 270848 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2941
timestamp 1758069660
transform 1 0 271676 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2953
timestamp 1758069660
transform 1 0 272780 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2965
timestamp 1758069660
transform 1 0 273884 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2977
timestamp 1758069660
transform 1 0 274988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2989
timestamp 1758069660
transform 1 0 276092 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2995
timestamp 1758069660
transform 1 0 276644 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2997
timestamp 1758069660
transform 1 0 276828 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3009
timestamp 1758069660
transform 1 0 277932 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3021
timestamp 1758069660
transform 1 0 279036 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3033
timestamp 1758069660
transform 1 0 280140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3045
timestamp 1758069660
transform 1 0 281244 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3051
timestamp 1758069660
transform 1 0 281796 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3053
timestamp 1758069660
transform 1 0 281980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3065
timestamp 1758069660
transform 1 0 283084 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3077
timestamp 1758069660
transform 1 0 284188 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3089
timestamp 1758069660
transform 1 0 285292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3101
timestamp 1758069660
transform 1 0 286396 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3107
timestamp 1758069660
transform 1 0 286948 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3109
timestamp 1758069660
transform 1 0 287132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3121
timestamp 1758069660
transform 1 0 288236 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3133
timestamp 1758069660
transform 1 0 289340 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3145
timestamp 1758069660
transform 1 0 290444 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3157
timestamp 1758069660
transform 1 0 291548 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3163
timestamp 1758069660
transform 1 0 292100 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3165
timestamp 1758069660
transform 1 0 292284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3177
timestamp 1758069660
transform 1 0 293388 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3189
timestamp 1758069660
transform 1 0 294492 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3201
timestamp 1758069660
transform 1 0 295596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3213
timestamp 1758069660
transform 1 0 296700 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3219
timestamp 1758069660
transform 1 0 297252 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3221
timestamp 1758069660
transform 1 0 297436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3233
timestamp 1758069660
transform 1 0 298540 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3245
timestamp 1758069660
transform 1 0 299644 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3257
timestamp 1758069660
transform 1 0 300748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3269
timestamp 1758069660
transform 1 0 301852 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3275
timestamp 1758069660
transform 1 0 302404 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3277
timestamp 1758069660
transform 1 0 302588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3289
timestamp 1758069660
transform 1 0 303692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3301
timestamp 1758069660
transform 1 0 304796 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1758069660
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1758069660
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1758069660
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1758069660
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1758069660
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1758069660
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1758069660
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1758069660
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1758069660
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1758069660
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1758069660
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1758069660
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1758069660
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1758069660
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1758069660
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1758069660
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1758069660
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1758069660
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1758069660
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1758069660
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1758069660
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1758069660
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1758069660
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1758069660
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1758069660
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1758069660
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1758069660
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1758069660
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1758069660
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1758069660
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_281
timestamp 1758069660
transform 1 0 26956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_289
timestamp 1758069660
transform 1 0 27692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1758069660
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1758069660
transform 1 0 29256 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_330
timestamp 1758069660
transform 1 0 31464 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_346
timestamp 1758069660
transform 1 0 32936 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_357
timestamp 1758069660
transform 1 0 33948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_364
timestamp 1758069660
transform 1 0 34592 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_371
timestamp 1758069660
transform 1 0 35236 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_383
timestamp 1758069660
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1758069660
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1758069660
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_408
timestamp 1758069660
transform 1 0 38640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_415
timestamp 1758069660
transform 1 0 39284 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_428
timestamp 1758069660
transform 1 0 40480 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_437
timestamp 1758069660
transform 1 0 41308 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_444
timestamp 1758069660
transform 1 0 41952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_449
timestamp 1758069660
transform 1 0 42412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_457
timestamp 1758069660
transform 1 0 43148 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1758069660
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1758069660
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1758069660
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1758069660
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1758069660
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1758069660
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1758069660
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1758069660
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1758069660
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1758069660
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1758069660
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_561
timestamp 1758069660
transform 1 0 52716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_565
timestamp 1758069660
transform 1 0 53084 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_574
timestamp 1758069660
transform 1 0 53912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_581
timestamp 1758069660
transform 1 0 54556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_594
timestamp 1758069660
transform 1 0 55752 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_600
timestamp 1758069660
transform 1 0 56304 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_604
timestamp 1758069660
transform 1 0 56672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_611
timestamp 1758069660
transform 1 0 57316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1758069660
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1758069660
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1758069660
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1758069660
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1758069660
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1758069660
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1758069660
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1758069660
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1758069660
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1758069660
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1758069660
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1758069660
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1758069660
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_729
timestamp 1758069660
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_741
timestamp 1758069660
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_753
timestamp 1758069660
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_765
timestamp 1758069660
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1758069660
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1758069660
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1758069660
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1758069660
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_818
timestamp 1758069660
transform 1 0 76360 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_827
timestamp 1758069660
transform 1 0 77188 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_836
timestamp 1758069660
transform 1 0 78016 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_844
timestamp 1758069660
transform 1 0 78752 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_856
timestamp 1758069660
transform 1 0 79856 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_868
timestamp 1758069660
transform 1 0 80960 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_880
timestamp 1758069660
transform 1 0 82064 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_892
timestamp 1758069660
transform 1 0 83168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_897
timestamp 1758069660
transform 1 0 83628 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_908
timestamp 1758069660
transform 1 0 84640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_915
timestamp 1758069660
transform 1 0 85284 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_928
timestamp 1758069660
transform 1 0 86480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_932
timestamp 1758069660
transform 1 0 86848 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_937
timestamp 1758069660
transform 1 0 87308 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_945
timestamp 1758069660
transform 1 0 88044 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_951
timestamp 1758069660
transform 1 0 88596 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_956
timestamp 1758069660
transform 1 0 89056 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_968
timestamp 1758069660
transform 1 0 90160 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_980
timestamp 1758069660
transform 1 0 91264 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_992
timestamp 1758069660
transform 1 0 92368 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1004
timestamp 1758069660
transform 1 0 93472 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1009
timestamp 1758069660
transform 1 0 93932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1021
timestamp 1758069660
transform 1 0 95036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1033
timestamp 1758069660
transform 1 0 96140 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1045
timestamp 1758069660
transform 1 0 97244 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1057
timestamp 1758069660
transform 1 0 98348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1063
timestamp 1758069660
transform 1 0 98900 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1065
timestamp 1758069660
transform 1 0 99084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1080
timestamp 1758069660
transform 1 0 100464 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1087
timestamp 1758069660
transform 1 0 101108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1100
timestamp 1758069660
transform 1 0 102304 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1106
timestamp 1758069660
transform 1 0 102856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1110
timestamp 1758069660
transform 1 0 103224 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1118
timestamp 1758069660
transform 1 0 103960 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1121
timestamp 1758069660
transform 1 0 104236 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1133
timestamp 1758069660
transform 1 0 105340 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1145
timestamp 1758069660
transform 1 0 106444 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1157
timestamp 1758069660
transform 1 0 107548 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1169
timestamp 1758069660
transform 1 0 108652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1175
timestamp 1758069660
transform 1 0 109204 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1177
timestamp 1758069660
transform 1 0 109388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1189
timestamp 1758069660
transform 1 0 110492 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1201
timestamp 1758069660
transform 1 0 111596 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1213
timestamp 1758069660
transform 1 0 112700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1228
timestamp 1758069660
transform 1 0 114080 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1233
timestamp 1758069660
transform 1 0 114540 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1243
timestamp 1758069660
transform 1 0 115460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1254
timestamp 1758069660
transform 1 0 116472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1261
timestamp 1758069660
transform 1 0 117116 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1268
timestamp 1758069660
transform 1 0 117760 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1280
timestamp 1758069660
transform 1 0 118864 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1289
timestamp 1758069660
transform 1 0 119692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1301
timestamp 1758069660
transform 1 0 120796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1313
timestamp 1758069660
transform 1 0 121900 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1325
timestamp 1758069660
transform 1 0 123004 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1337
timestamp 1758069660
transform 1 0 124108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1343
timestamp 1758069660
transform 1 0 124660 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1345
timestamp 1758069660
transform 1 0 124844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1357
timestamp 1758069660
transform 1 0 125948 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1369
timestamp 1758069660
transform 1 0 127052 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1381
timestamp 1758069660
transform 1 0 128156 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1396
timestamp 1758069660
transform 1 0 129536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1401
timestamp 1758069660
transform 1 0 129996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1405
timestamp 1758069660
transform 1 0 130364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1415
timestamp 1758069660
transform 1 0 131284 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1423
timestamp 1758069660
transform 1 0 132020 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1430
timestamp 1758069660
transform 1 0 132664 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1442
timestamp 1758069660
transform 1 0 133768 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1454
timestamp 1758069660
transform 1 0 134872 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1457
timestamp 1758069660
transform 1 0 135148 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1469
timestamp 1758069660
transform 1 0 136252 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1481
timestamp 1758069660
transform 1 0 137356 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1493
timestamp 1758069660
transform 1 0 138460 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1505
timestamp 1758069660
transform 1 0 139564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1511
timestamp 1758069660
transform 1 0 140116 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1513
timestamp 1758069660
transform 1 0 140300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1525
timestamp 1758069660
transform 1 0 141404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1537
timestamp 1758069660
transform 1 0 142508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1549
timestamp 1758069660
transform 1 0 143612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1561
timestamp 1758069660
transform 1 0 144716 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1567
timestamp 1758069660
transform 1 0 145268 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1569
timestamp 1758069660
transform 1 0 145452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1581
timestamp 1758069660
transform 1 0 146556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_1589
timestamp 1758069660
transform 1 0 147292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1595
timestamp 1758069660
transform 1 0 147844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1599
timestamp 1758069660
transform 1 0 148212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1620
timestamp 1758069660
transform 1 0 150144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1625
timestamp 1758069660
transform 1 0 150604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1629
timestamp 1758069660
transform 1 0 150972 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1633
timestamp 1758069660
transform 1 0 151340 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1639
timestamp 1758069660
transform 1 0 151892 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1643
timestamp 1758069660
transform 1 0 152260 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1650
timestamp 1758069660
transform 1 0 152904 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1662
timestamp 1758069660
transform 1 0 154008 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1674
timestamp 1758069660
transform 1 0 155112 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1681
timestamp 1758069660
transform 1 0 155756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1693
timestamp 1758069660
transform 1 0 156860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1705
timestamp 1758069660
transform 1 0 157964 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1717
timestamp 1758069660
transform 1 0 159068 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1729
timestamp 1758069660
transform 1 0 160172 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1735
timestamp 1758069660
transform 1 0 160724 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1740
timestamp 1758069660
transform 1 0 161184 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1747
timestamp 1758069660
transform 1 0 161828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1754
timestamp 1758069660
transform 1 0 162472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1761
timestamp 1758069660
transform 1 0 163116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1768
timestamp 1758069660
transform 1 0 163760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1775
timestamp 1758069660
transform 1 0 164404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1782
timestamp 1758069660
transform 1 0 165048 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1790
timestamp 1758069660
transform 1 0 165784 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1793
timestamp 1758069660
transform 1 0 166060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1805
timestamp 1758069660
transform 1 0 167164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1817
timestamp 1758069660
transform 1 0 168268 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1829
timestamp 1758069660
transform 1 0 169372 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1841
timestamp 1758069660
transform 1 0 170476 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1847
timestamp 1758069660
transform 1 0 171028 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1849
timestamp 1758069660
transform 1 0 171212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1861
timestamp 1758069660
transform 1 0 172316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1873
timestamp 1758069660
transform 1 0 173420 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1885
timestamp 1758069660
transform 1 0 174524 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1897
timestamp 1758069660
transform 1 0 175628 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1903
timestamp 1758069660
transform 1 0 176180 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1905
timestamp 1758069660
transform 1 0 176364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1909
timestamp 1758069660
transform 1 0 176732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1917
timestamp 1758069660
transform 1 0 177468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1927
timestamp 1758069660
transform 1 0 178388 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1940
timestamp 1758069660
transform 1 0 179584 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1947
timestamp 1758069660
transform 1 0 180228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1959
timestamp 1758069660
transform 1 0 181332 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1961
timestamp 1758069660
transform 1 0 181516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1973
timestamp 1758069660
transform 1 0 182620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1985
timestamp 1758069660
transform 1 0 183724 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1997
timestamp 1758069660
transform 1 0 184828 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2009
timestamp 1758069660
transform 1 0 185932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2015
timestamp 1758069660
transform 1 0 186484 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2017
timestamp 1758069660
transform 1 0 186668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2029
timestamp 1758069660
transform 1 0 187772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2041
timestamp 1758069660
transform 1 0 188876 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2050
timestamp 1758069660
transform 1 0 189704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2057
timestamp 1758069660
transform 1 0 190348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_2064
timestamp 1758069660
transform 1 0 190992 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2093
timestamp 1758069660
transform 1 0 193660 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2117
timestamp 1758069660
transform 1 0 195868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2124
timestamp 1758069660
transform 1 0 196512 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2129
timestamp 1758069660
transform 1 0 196972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2141
timestamp 1758069660
transform 1 0 198076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2153
timestamp 1758069660
transform 1 0 199180 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2165
timestamp 1758069660
transform 1 0 200284 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2177
timestamp 1758069660
transform 1 0 201388 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2183
timestamp 1758069660
transform 1 0 201940 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2185
timestamp 1758069660
transform 1 0 202124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2189
timestamp 1758069660
transform 1 0 202492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2196
timestamp 1758069660
transform 1 0 203136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2200
timestamp 1758069660
transform 1 0 203504 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2210
timestamp 1758069660
transform 1 0 204424 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2223
timestamp 1758069660
transform 1 0 205620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2235
timestamp 1758069660
transform 1 0 206724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2239
timestamp 1758069660
transform 1 0 207092 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2241
timestamp 1758069660
transform 1 0 207276 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2253
timestamp 1758069660
transform 1 0 208380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2265
timestamp 1758069660
transform 1 0 209484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2277
timestamp 1758069660
transform 1 0 210588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2289
timestamp 1758069660
transform 1 0 211692 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2295
timestamp 1758069660
transform 1 0 212244 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2297
timestamp 1758069660
transform 1 0 212428 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2309
timestamp 1758069660
transform 1 0 213532 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2321
timestamp 1758069660
transform 1 0 214636 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2333
timestamp 1758069660
transform 1 0 215740 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2345
timestamp 1758069660
transform 1 0 216844 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2351
timestamp 1758069660
transform 1 0 217396 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2353
timestamp 1758069660
transform 1 0 217580 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2365
timestamp 1758069660
transform 1 0 218684 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2377
timestamp 1758069660
transform 1 0 219788 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2389
timestamp 1758069660
transform 1 0 220892 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2401
timestamp 1758069660
transform 1 0 221996 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2407
timestamp 1758069660
transform 1 0 222548 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2409
timestamp 1758069660
transform 1 0 222732 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2421
timestamp 1758069660
transform 1 0 223836 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2433
timestamp 1758069660
transform 1 0 224940 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2445
timestamp 1758069660
transform 1 0 226044 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2457
timestamp 1758069660
transform 1 0 227148 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2463
timestamp 1758069660
transform 1 0 227700 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2474
timestamp 1758069660
transform 1 0 228712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2487
timestamp 1758069660
transform 1 0 229908 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2494
timestamp 1758069660
transform 1 0 230552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2501
timestamp 1758069660
transform 1 0 231196 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2508
timestamp 1758069660
transform 1 0 231840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2521
timestamp 1758069660
transform 1 0 233036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2533
timestamp 1758069660
transform 1 0 234140 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2545
timestamp 1758069660
transform 1 0 235244 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2557
timestamp 1758069660
transform 1 0 236348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2569
timestamp 1758069660
transform 1 0 237452 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2575
timestamp 1758069660
transform 1 0 238004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2577
timestamp 1758069660
transform 1 0 238188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_2585
timestamp 1758069660
transform 1 0 238924 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_2593
timestamp 1758069660
transform 1 0 239660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2604
timestamp 1758069660
transform 1 0 240672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2611
timestamp 1758069660
transform 1 0 241316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2618
timestamp 1758069660
transform 1 0 241960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2625
timestamp 1758069660
transform 1 0 242604 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2631
timestamp 1758069660
transform 1 0 243156 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2633
timestamp 1758069660
transform 1 0 243340 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2645
timestamp 1758069660
transform 1 0 244444 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2657
timestamp 1758069660
transform 1 0 245548 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2669
timestamp 1758069660
transform 1 0 246652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2681
timestamp 1758069660
transform 1 0 247756 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2687
timestamp 1758069660
transform 1 0 248308 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2689
timestamp 1758069660
transform 1 0 248492 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2701
timestamp 1758069660
transform 1 0 249596 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2713
timestamp 1758069660
transform 1 0 250700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_2728
timestamp 1758069660
transform 1 0 252080 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_2732
timestamp 1758069660
transform 1 0 252448 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2738
timestamp 1758069660
transform 1 0 253000 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2754
timestamp 1758069660
transform 1 0 254472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2761
timestamp 1758069660
transform 1 0 255116 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2768
timestamp 1758069660
transform 1 0 255760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2780
timestamp 1758069660
transform 1 0 256864 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_2792
timestamp 1758069660
transform 1 0 257968 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2801
timestamp 1758069660
transform 1 0 258796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2813
timestamp 1758069660
transform 1 0 259900 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2825
timestamp 1758069660
transform 1 0 261004 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2837
timestamp 1758069660
transform 1 0 262108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2849
timestamp 1758069660
transform 1 0 263212 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2855
timestamp 1758069660
transform 1 0 263764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2857
timestamp 1758069660
transform 1 0 263948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2864
timestamp 1758069660
transform 1 0 264592 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2871
timestamp 1758069660
transform 1 0 265236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2895
timestamp 1758069660
transform 1 0 267444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2908
timestamp 1758069660
transform 1 0 268640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2933
timestamp 1758069660
transform 1 0 270940 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2940
timestamp 1758069660
transform 1 0 271584 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2952
timestamp 1758069660
transform 1 0 272688 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2964
timestamp 1758069660
transform 1 0 273792 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2969
timestamp 1758069660
transform 1 0 274252 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2981
timestamp 1758069660
transform 1 0 275356 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2993
timestamp 1758069660
transform 1 0 276460 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3005
timestamp 1758069660
transform 1 0 277564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3017
timestamp 1758069660
transform 1 0 278668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3023
timestamp 1758069660
transform 1 0 279220 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3025
timestamp 1758069660
transform 1 0 279404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3037
timestamp 1758069660
transform 1 0 280508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3049
timestamp 1758069660
transform 1 0 281612 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3061
timestamp 1758069660
transform 1 0 282716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3073
timestamp 1758069660
transform 1 0 283820 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3079
timestamp 1758069660
transform 1 0 284372 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3081
timestamp 1758069660
transform 1 0 284556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3093
timestamp 1758069660
transform 1 0 285660 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3105
timestamp 1758069660
transform 1 0 286764 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3117
timestamp 1758069660
transform 1 0 287868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3129
timestamp 1758069660
transform 1 0 288972 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3135
timestamp 1758069660
transform 1 0 289524 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3137
timestamp 1758069660
transform 1 0 289708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3149
timestamp 1758069660
transform 1 0 290812 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3161
timestamp 1758069660
transform 1 0 291916 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3173
timestamp 1758069660
transform 1 0 293020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3185
timestamp 1758069660
transform 1 0 294124 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3191
timestamp 1758069660
transform 1 0 294676 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3193
timestamp 1758069660
transform 1 0 294860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3205
timestamp 1758069660
transform 1 0 295964 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3217
timestamp 1758069660
transform 1 0 297068 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3229
timestamp 1758069660
transform 1 0 298172 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3241
timestamp 1758069660
transform 1 0 299276 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3247
timestamp 1758069660
transform 1 0 299828 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3249
timestamp 1758069660
transform 1 0 300012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3261
timestamp 1758069660
transform 1 0 301116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3273
timestamp 1758069660
transform 1 0 302220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3285
timestamp 1758069660
transform 1 0 303324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3297
timestamp 1758069660
transform 1 0 304428 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3303
timestamp 1758069660
transform 1 0 304980 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3305
timestamp 1758069660
transform 1 0 305164 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1758069660
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1758069660
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1758069660
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1758069660
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1758069660
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1758069660
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1758069660
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1758069660
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1758069660
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1758069660
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1758069660
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1758069660
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1758069660
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1758069660
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1758069660
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1758069660
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1758069660
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1758069660
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1758069660
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1758069660
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1758069660
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1758069660
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1758069660
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1758069660
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1758069660
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1758069660
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1758069660
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1758069660
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1758069660
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_277
timestamp 1758069660
transform 1 0 26588 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_281
timestamp 1758069660
transform 1 0 26956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_291
timestamp 1758069660
transform 1 0 27876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1758069660
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_329
timestamp 1758069660
transform 1 0 31372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_353
timestamp 1758069660
transform 1 0 33580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1758069660
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_368
timestamp 1758069660
transform 1 0 34960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_375
timestamp 1758069660
transform 1 0 35604 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_381
timestamp 1758069660
transform 1 0 36156 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_386
timestamp 1758069660
transform 1 0 36616 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_394
timestamp 1758069660
transform 1 0 37352 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_409
timestamp 1758069660
transform 1 0 38732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1758069660
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1758069660
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_434
timestamp 1758069660
transform 1 0 41032 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_458
timestamp 1758069660
transform 1 0 43240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_466
timestamp 1758069660
transform 1 0 43976 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_474
timestamp 1758069660
transform 1 0 44712 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1758069660
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1758069660
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1758069660
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1758069660
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1758069660
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1758069660
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1758069660
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1758069660
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_577
timestamp 1758069660
transform 1 0 54188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_584
timestamp 1758069660
transform 1 0 54832 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_589
timestamp 1758069660
transform 1 0 55292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_594
timestamp 1758069660
transform 1 0 55752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_607
timestamp 1758069660
transform 1 0 56948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_614
timestamp 1758069660
transform 1 0 57592 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_621
timestamp 1758069660
transform 1 0 58236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_633
timestamp 1758069660
transform 1 0 59340 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_641
timestamp 1758069660
transform 1 0 60076 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1758069660
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1758069660
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1758069660
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1758069660
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1758069660
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1758069660
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1758069660
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1758069660
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_725
timestamp 1758069660
transform 1 0 67804 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_737
timestamp 1758069660
transform 1 0 68908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1758069660
transform 1 0 70012 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1758069660
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_757
timestamp 1758069660
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_769
timestamp 1758069660
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_781
timestamp 1758069660
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_793
timestamp 1758069660
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_808
timestamp 1758069660
transform 1 0 75440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_813
timestamp 1758069660
transform 1 0 75900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_826
timestamp 1758069660
transform 1 0 77096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_839
timestamp 1758069660
transform 1 0 78292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_847
timestamp 1758069660
transform 1 0 79028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_852
timestamp 1758069660
transform 1 0 79488 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_858
timestamp 1758069660
transform 1 0 80040 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_862
timestamp 1758069660
transform 1 0 80408 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_869
timestamp 1758069660
transform 1 0 81052 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_881
timestamp 1758069660
transform 1 0 82156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_893
timestamp 1758069660
transform 1 0 83260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_910
timestamp 1758069660
transform 1 0 84824 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_916
timestamp 1758069660
transform 1 0 85376 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_920
timestamp 1758069660
transform 1 0 85744 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_925
timestamp 1758069660
transform 1 0 86204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_936
timestamp 1758069660
transform 1 0 87216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_949
timestamp 1758069660
transform 1 0 88412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_956
timestamp 1758069660
transform 1 0 89056 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_963
timestamp 1758069660
transform 1 0 89700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_970
timestamp 1758069660
transform 1 0 90344 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_978
timestamp 1758069660
transform 1 0 91080 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_981
timestamp 1758069660
transform 1 0 91356 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_993
timestamp 1758069660
transform 1 0 92460 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1005
timestamp 1758069660
transform 1 0 93564 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1017
timestamp 1758069660
transform 1 0 94668 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1029
timestamp 1758069660
transform 1 0 95772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1035
timestamp 1758069660
transform 1 0 96324 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1037
timestamp 1758069660
transform 1 0 96508 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1049
timestamp 1758069660
transform 1 0 97612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1061
timestamp 1758069660
transform 1 0 98716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1068
timestamp 1758069660
transform 1 0 99360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1075
timestamp 1758069660
transform 1 0 100004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1088
timestamp 1758069660
transform 1 0 101200 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1093
timestamp 1758069660
transform 1 0 101660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1099
timestamp 1758069660
transform 1 0 102212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1112
timestamp 1758069660
transform 1 0 103408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1119
timestamp 1758069660
transform 1 0 104052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1126
timestamp 1758069660
transform 1 0 104696 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1133
timestamp 1758069660
transform 1 0 105340 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1145
timestamp 1758069660
transform 1 0 106444 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1149
timestamp 1758069660
transform 1 0 106812 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1161
timestamp 1758069660
transform 1 0 107916 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1173
timestamp 1758069660
transform 1 0 109020 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1185
timestamp 1758069660
transform 1 0 110124 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1197
timestamp 1758069660
transform 1 0 111228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1203
timestamp 1758069660
transform 1 0 111780 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1205
timestamp 1758069660
transform 1 0 111964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1220
timestamp 1758069660
transform 1 0 113344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1227
timestamp 1758069660
transform 1 0 113988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1251
timestamp 1758069660
transform 1 0 116196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1259
timestamp 1758069660
transform 1 0 116932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1270
timestamp 1758069660
transform 1 0 117944 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1277
timestamp 1758069660
transform 1 0 118588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1289
timestamp 1758069660
transform 1 0 119692 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1301
timestamp 1758069660
transform 1 0 120796 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1313
timestamp 1758069660
transform 1 0 121900 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1317
timestamp 1758069660
transform 1 0 122268 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1329
timestamp 1758069660
transform 1 0 123372 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1341
timestamp 1758069660
transform 1 0 124476 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1353
timestamp 1758069660
transform 1 0 125580 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1365
timestamp 1758069660
transform 1 0 126684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1371
timestamp 1758069660
transform 1 0 127236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1373
timestamp 1758069660
transform 1 0 127420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1379
timestamp 1758069660
transform 1 0 127972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1383
timestamp 1758069660
transform 1 0 128340 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1387
timestamp 1758069660
transform 1 0 128708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1411
timestamp 1758069660
transform 1 0 130916 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1424
timestamp 1758069660
transform 1 0 132112 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1432
timestamp 1758069660
transform 1 0 132848 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1444
timestamp 1758069660
transform 1 0 133952 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1456
timestamp 1758069660
transform 1 0 135056 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1468
timestamp 1758069660
transform 1 0 136160 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1480
timestamp 1758069660
transform 1 0 137264 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1491
timestamp 1758069660
transform 1 0 138276 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1503
timestamp 1758069660
transform 1 0 139380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1515
timestamp 1758069660
transform 1 0 140484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1527
timestamp 1758069660
transform 1 0 141588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1539
timestamp 1758069660
transform 1 0 142692 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1541
timestamp 1758069660
transform 1 0 142876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1553
timestamp 1758069660
transform 1 0 143980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1565
timestamp 1758069660
transform 1 0 145084 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1571
timestamp 1758069660
transform 1 0 145636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1578
timestamp 1758069660
transform 1 0 146280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1586
timestamp 1758069660
transform 1 0 147016 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1592
timestamp 1758069660
transform 1 0 147568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1597
timestamp 1758069660
transform 1 0 148028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1603
timestamp 1758069660
transform 1 0 148580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1611
timestamp 1758069660
transform 1 0 149316 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1632
timestamp 1758069660
transform 1 0 151248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1648
timestamp 1758069660
transform 1 0 152720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1653
timestamp 1758069660
transform 1 0 153180 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1666
timestamp 1758069660
transform 1 0 154376 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1678
timestamp 1758069660
transform 1 0 155480 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1690
timestamp 1758069660
transform 1 0 156584 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1702
timestamp 1758069660
transform 1 0 157688 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1709
timestamp 1758069660
transform 1 0 158332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1721
timestamp 1758069660
transform 1 0 159436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1730
timestamp 1758069660
transform 1 0 160264 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1745
timestamp 1758069660
transform 1 0 161644 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1758
timestamp 1758069660
transform 1 0 162840 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1765
timestamp 1758069660
transform 1 0 163484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1786
timestamp 1758069660
transform 1 0 165416 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1794
timestamp 1758069660
transform 1 0 166152 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1806
timestamp 1758069660
transform 1 0 167256 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1818
timestamp 1758069660
transform 1 0 168360 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1821
timestamp 1758069660
transform 1 0 168636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1833
timestamp 1758069660
transform 1 0 169740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1845
timestamp 1758069660
transform 1 0 170844 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1857
timestamp 1758069660
transform 1 0 171948 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1869
timestamp 1758069660
transform 1 0 173052 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1875
timestamp 1758069660
transform 1 0 173604 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1877
timestamp 1758069660
transform 1 0 173788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1889
timestamp 1758069660
transform 1 0 174892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1897
timestamp 1758069660
transform 1 0 175628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1903
timestamp 1758069660
transform 1 0 176180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1916
timestamp 1758069660
transform 1 0 177376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1920
timestamp 1758069660
transform 1 0 177744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1925
timestamp 1758069660
transform 1 0 178204 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1931
timestamp 1758069660
transform 1 0 178756 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1933
timestamp 1758069660
transform 1 0 178940 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1955
timestamp 1758069660
transform 1 0 180964 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1962
timestamp 1758069660
transform 1 0 181608 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1974
timestamp 1758069660
transform 1 0 182712 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1986
timestamp 1758069660
transform 1 0 183816 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1989
timestamp 1758069660
transform 1 0 184092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2001
timestamp 1758069660
transform 1 0 185196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2013
timestamp 1758069660
transform 1 0 186300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2025
timestamp 1758069660
transform 1 0 187404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2040
timestamp 1758069660
transform 1 0 188784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_2045
timestamp 1758069660
transform 1 0 189244 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2051
timestamp 1758069660
transform 1 0 189796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2058
timestamp 1758069660
transform 1 0 190440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2082
timestamp 1758069660
transform 1 0 192648 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2095
timestamp 1758069660
transform 1 0 193844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2099
timestamp 1758069660
transform 1 0 194212 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2124
timestamp 1758069660
transform 1 0 196512 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2138
timestamp 1758069660
transform 1 0 197800 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2150
timestamp 1758069660
transform 1 0 198904 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2157
timestamp 1758069660
transform 1 0 199548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2169
timestamp 1758069660
transform 1 0 200652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2176
timestamp 1758069660
transform 1 0 201296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2183
timestamp 1758069660
transform 1 0 201940 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2191
timestamp 1758069660
transform 1 0 202676 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2202
timestamp 1758069660
transform 1 0 203688 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2210
timestamp 1758069660
transform 1 0 204424 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2233
timestamp 1758069660
transform 1 0 206540 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2245
timestamp 1758069660
transform 1 0 207644 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2257
timestamp 1758069660
transform 1 0 208748 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_2265
timestamp 1758069660
transform 1 0 209484 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2269
timestamp 1758069660
transform 1 0 209852 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2281
timestamp 1758069660
transform 1 0 210956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2293
timestamp 1758069660
transform 1 0 212060 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2305
timestamp 1758069660
transform 1 0 213164 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2317
timestamp 1758069660
transform 1 0 214268 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2323
timestamp 1758069660
transform 1 0 214820 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2325
timestamp 1758069660
transform 1 0 215004 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2337
timestamp 1758069660
transform 1 0 216108 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2349
timestamp 1758069660
transform 1 0 217212 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2361
timestamp 1758069660
transform 1 0 218316 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2373
timestamp 1758069660
transform 1 0 219420 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2379
timestamp 1758069660
transform 1 0 219972 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2381
timestamp 1758069660
transform 1 0 220156 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2393
timestamp 1758069660
transform 1 0 221260 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2405
timestamp 1758069660
transform 1 0 222364 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2417
timestamp 1758069660
transform 1 0 223468 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2429
timestamp 1758069660
transform 1 0 224572 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2435
timestamp 1758069660
transform 1 0 225124 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2437
timestamp 1758069660
transform 1 0 225308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2449
timestamp 1758069660
transform 1 0 226412 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2481
timestamp 1758069660
transform 1 0 229356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2488
timestamp 1758069660
transform 1 0 230000 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2493
timestamp 1758069660
transform 1 0 230460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2497
timestamp 1758069660
transform 1 0 230828 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2507
timestamp 1758069660
transform 1 0 231748 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2514
timestamp 1758069660
transform 1 0 232392 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2526
timestamp 1758069660
transform 1 0 233496 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2538
timestamp 1758069660
transform 1 0 234600 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2546
timestamp 1758069660
transform 1 0 235336 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2549
timestamp 1758069660
transform 1 0 235612 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2561
timestamp 1758069660
transform 1 0 236716 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2573
timestamp 1758069660
transform 1 0 237820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2579
timestamp 1758069660
transform 1 0 238372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2592
timestamp 1758069660
transform 1 0 239568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2599
timestamp 1758069660
transform 1 0 240212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2603
timestamp 1758069660
transform 1 0 240580 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2605
timestamp 1758069660
transform 1 0 240764 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2615
timestamp 1758069660
transform 1 0 241684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2621
timestamp 1758069660
transform 1 0 242236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2631
timestamp 1758069660
transform 1 0 243156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2638
timestamp 1758069660
transform 1 0 243800 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2645
timestamp 1758069660
transform 1 0 244444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_2657
timestamp 1758069660
transform 1 0 245548 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2661
timestamp 1758069660
transform 1 0 245916 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2673
timestamp 1758069660
transform 1 0 247020 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2685
timestamp 1758069660
transform 1 0 248124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2693
timestamp 1758069660
transform 1 0 248860 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2698
timestamp 1758069660
transform 1 0 249320 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2710
timestamp 1758069660
transform 1 0 250424 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2720
timestamp 1758069660
transform 1 0 251344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2724
timestamp 1758069660
transform 1 0 251712 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2729
timestamp 1758069660
transform 1 0 252172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2753
timestamp 1758069660
transform 1 0 254380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2766
timestamp 1758069660
transform 1 0 255576 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2776
timestamp 1758069660
transform 1 0 256496 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2783
timestamp 1758069660
transform 1 0 257140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2795
timestamp 1758069660
transform 1 0 258244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2807
timestamp 1758069660
transform 1 0 259348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2819
timestamp 1758069660
transform 1 0 260452 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2827
timestamp 1758069660
transform 1 0 261188 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2829
timestamp 1758069660
transform 1 0 261372 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2844
timestamp 1758069660
transform 1 0 262752 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2856
timestamp 1758069660
transform 1 0 263856 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2860
timestamp 1758069660
transform 1 0 264224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2867
timestamp 1758069660
transform 1 0 264868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2880
timestamp 1758069660
transform 1 0 266064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2905
timestamp 1758069660
transform 1 0 268364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2929
timestamp 1758069660
transform 1 0 270572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2936
timestamp 1758069660
transform 1 0 271216 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2950
timestamp 1758069660
transform 1 0 272504 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2962
timestamp 1758069660
transform 1 0 273608 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2974
timestamp 1758069660
transform 1 0 274712 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2986
timestamp 1758069660
transform 1 0 275816 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2994
timestamp 1758069660
transform 1 0 276552 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2997
timestamp 1758069660
transform 1 0 276828 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3009
timestamp 1758069660
transform 1 0 277932 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3021
timestamp 1758069660
transform 1 0 279036 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3033
timestamp 1758069660
transform 1 0 280140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3045
timestamp 1758069660
transform 1 0 281244 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3051
timestamp 1758069660
transform 1 0 281796 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3053
timestamp 1758069660
transform 1 0 281980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3065
timestamp 1758069660
transform 1 0 283084 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3077
timestamp 1758069660
transform 1 0 284188 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3089
timestamp 1758069660
transform 1 0 285292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3101
timestamp 1758069660
transform 1 0 286396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3107
timestamp 1758069660
transform 1 0 286948 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3109
timestamp 1758069660
transform 1 0 287132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3121
timestamp 1758069660
transform 1 0 288236 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3133
timestamp 1758069660
transform 1 0 289340 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3145
timestamp 1758069660
transform 1 0 290444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3157
timestamp 1758069660
transform 1 0 291548 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3163
timestamp 1758069660
transform 1 0 292100 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3165
timestamp 1758069660
transform 1 0 292284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3177
timestamp 1758069660
transform 1 0 293388 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3189
timestamp 1758069660
transform 1 0 294492 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3201
timestamp 1758069660
transform 1 0 295596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3213
timestamp 1758069660
transform 1 0 296700 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3219
timestamp 1758069660
transform 1 0 297252 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3221
timestamp 1758069660
transform 1 0 297436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3233
timestamp 1758069660
transform 1 0 298540 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3245
timestamp 1758069660
transform 1 0 299644 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3257
timestamp 1758069660
transform 1 0 300748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3269
timestamp 1758069660
transform 1 0 301852 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3275
timestamp 1758069660
transform 1 0 302404 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3277
timestamp 1758069660
transform 1 0 302588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3289
timestamp 1758069660
transform 1 0 303692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3301
timestamp 1758069660
transform 1 0 304796 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1758069660
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1758069660
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1758069660
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1758069660
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1758069660
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1758069660
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1758069660
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1758069660
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1758069660
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1758069660
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1758069660
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1758069660
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1758069660
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1758069660
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1758069660
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1758069660
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1758069660
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1758069660
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1758069660
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1758069660
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1758069660
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1758069660
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1758069660
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1758069660
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1758069660
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1758069660
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1758069660
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_261
timestamp 1758069660
transform 1 0 25116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_269
timestamp 1758069660
transform 1 0 25852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1758069660
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1758069660
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1758069660
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1758069660
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_308
timestamp 1758069660
transform 1 0 29440 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1758069660
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_357
timestamp 1758069660
transform 1 0 33948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_370
timestamp 1758069660
transform 1 0 35144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_377
timestamp 1758069660
transform 1 0 35788 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_383
timestamp 1758069660
transform 1 0 36340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1758069660
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_397
timestamp 1758069660
transform 1 0 37628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_410
timestamp 1758069660
transform 1 0 38824 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_416
timestamp 1758069660
transform 1 0 39376 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_437
timestamp 1758069660
transform 1 0 41308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1758069660
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_452
timestamp 1758069660
transform 1 0 42688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_465
timestamp 1758069660
transform 1 0 43884 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_471
timestamp 1758069660
transform 1 0 44436 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_475
timestamp 1758069660
transform 1 0 44804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_487
timestamp 1758069660
transform 1 0 45908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_499
timestamp 1758069660
transform 1 0 47012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1758069660
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1758069660
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1758069660
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1758069660
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1758069660
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_556
timestamp 1758069660
transform 1 0 52256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_561
timestamp 1758069660
transform 1 0 52716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_566
timestamp 1758069660
transform 1 0 53176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_579
timestamp 1758069660
transform 1 0 54372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_603
timestamp 1758069660
transform 1 0 56580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_611
timestamp 1758069660
transform 1 0 57316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1758069660
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_617
timestamp 1758069660
transform 1 0 57868 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1758069660
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1758069660
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1758069660
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1758069660
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1758069660
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1758069660
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1758069660
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1758069660
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1758069660
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1758069660
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1758069660
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_729
timestamp 1758069660
transform 1 0 68172 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_741
timestamp 1758069660
transform 1 0 69276 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_753
timestamp 1758069660
transform 1 0 70380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_765
timestamp 1758069660
transform 1 0 71484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_771
timestamp 1758069660
transform 1 0 72036 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_775
timestamp 1758069660
transform 1 0 72404 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1758069660
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1758069660
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_797
timestamp 1758069660
transform 1 0 74428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_801
timestamp 1758069660
transform 1 0 74796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_805
timestamp 1758069660
transform 1 0 75164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_829
timestamp 1758069660
transform 1 0 77372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_836
timestamp 1758069660
transform 1 0 78016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_844
timestamp 1758069660
transform 1 0 78752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_851
timestamp 1758069660
transform 1 0 79396 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_875
timestamp 1758069660
transform 1 0 81604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_887
timestamp 1758069660
transform 1 0 82708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_895
timestamp 1758069660
transform 1 0 83444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_897
timestamp 1758069660
transform 1 0 83628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_921
timestamp 1758069660
transform 1 0 85836 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_945
timestamp 1758069660
transform 1 0 88044 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_951
timestamp 1758069660
transform 1 0 88596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_953
timestamp 1758069660
transform 1 0 88780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_966
timestamp 1758069660
transform 1 0 89976 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_974
timestamp 1758069660
transform 1 0 90712 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_981
timestamp 1758069660
transform 1 0 91356 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_993
timestamp 1758069660
transform 1 0 92460 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1005
timestamp 1758069660
transform 1 0 93564 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1009
timestamp 1758069660
transform 1 0 93932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1021
timestamp 1758069660
transform 1 0 95036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1033
timestamp 1758069660
transform 1 0 96140 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1045
timestamp 1758069660
transform 1 0 97244 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1060
timestamp 1758069660
transform 1 0 98624 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1065
timestamp 1758069660
transform 1 0 99084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1086
timestamp 1758069660
transform 1 0 101016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1110
timestamp 1758069660
transform 1 0 103224 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1118
timestamp 1758069660
transform 1 0 103960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1130
timestamp 1758069660
transform 1 0 105064 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1138
timestamp 1758069660
transform 1 0 105800 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1142
timestamp 1758069660
transform 1 0 106168 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1154
timestamp 1758069660
transform 1 0 107272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1166
timestamp 1758069660
transform 1 0 108376 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1174
timestamp 1758069660
transform 1 0 109112 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1177
timestamp 1758069660
transform 1 0 109388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1189
timestamp 1758069660
transform 1 0 110492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1201
timestamp 1758069660
transform 1 0 111596 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1213
timestamp 1758069660
transform 1 0 112700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1220
timestamp 1758069660
transform 1 0 113344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1228
timestamp 1758069660
transform 1 0 114080 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1237
timestamp 1758069660
transform 1 0 114908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1250
timestamp 1758069660
transform 1 0 116104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1274
timestamp 1758069660
transform 1 0 118312 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1281
timestamp 1758069660
transform 1 0 118956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1287
timestamp 1758069660
transform 1 0 119508 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1289
timestamp 1758069660
transform 1 0 119692 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1301
timestamp 1758069660
transform 1 0 120796 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1313
timestamp 1758069660
transform 1 0 121900 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1325
timestamp 1758069660
transform 1 0 123004 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1337
timestamp 1758069660
transform 1 0 124108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1343
timestamp 1758069660
transform 1 0 124660 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1345
timestamp 1758069660
transform 1 0 124844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1357
timestamp 1758069660
transform 1 0 125948 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1368
timestamp 1758069660
transform 1 0 126960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1376
timestamp 1758069660
transform 1 0 127696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1383
timestamp 1758069660
transform 1 0 128340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1396
timestamp 1758069660
transform 1 0 129536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1401
timestamp 1758069660
transform 1 0 129996 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1406
timestamp 1758069660
transform 1 0 130456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1430
timestamp 1758069660
transform 1 0 132664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1434
timestamp 1758069660
transform 1 0 133032 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1444
timestamp 1758069660
transform 1 0 133952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1451
timestamp 1758069660
transform 1 0 134596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1455
timestamp 1758069660
transform 1 0 134964 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1457
timestamp 1758069660
transform 1 0 135148 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1463
timestamp 1758069660
transform 1 0 135700 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1475
timestamp 1758069660
transform 1 0 136804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1487
timestamp 1758069660
transform 1 0 137908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1499
timestamp 1758069660
transform 1 0 139012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1511
timestamp 1758069660
transform 1 0 140116 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1513
timestamp 1758069660
transform 1 0 140300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1525
timestamp 1758069660
transform 1 0 141404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1537
timestamp 1758069660
transform 1 0 142508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1541
timestamp 1758069660
transform 1 0 142876 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1548
timestamp 1758069660
transform 1 0 143520 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1560
timestamp 1758069660
transform 1 0 144624 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1578
timestamp 1758069660
transform 1 0 146280 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1587
timestamp 1758069660
transform 1 0 147108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1611
timestamp 1758069660
transform 1 0 149316 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1620
timestamp 1758069660
transform 1 0 150144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1625
timestamp 1758069660
transform 1 0 150604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1629
timestamp 1758069660
transform 1 0 150972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1639
timestamp 1758069660
transform 1 0 151892 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1645
timestamp 1758069660
transform 1 0 152444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1649
timestamp 1758069660
transform 1 0 152812 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1653
timestamp 1758069660
transform 1 0 153180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1657
timestamp 1758069660
transform 1 0 153548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1661
timestamp 1758069660
transform 1 0 153916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1665
timestamp 1758069660
transform 1 0 154284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1676
timestamp 1758069660
transform 1 0 155296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1681
timestamp 1758069660
transform 1 0 155756 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1685
timestamp 1758069660
transform 1 0 156124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1689
timestamp 1758069660
transform 1 0 156492 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1693
timestamp 1758069660
transform 1 0 156860 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1697
timestamp 1758069660
transform 1 0 157228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1709
timestamp 1758069660
transform 1 0 158332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1713
timestamp 1758069660
transform 1 0 158700 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1723
timestamp 1758069660
transform 1 0 159620 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1731
timestamp 1758069660
transform 1 0 160356 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1735
timestamp 1758069660
transform 1 0 160724 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1737
timestamp 1758069660
transform 1 0 160908 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1743
timestamp 1758069660
transform 1 0 161460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1767
timestamp 1758069660
transform 1 0 163668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1780
timestamp 1758069660
transform 1 0 164864 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1788
timestamp 1758069660
transform 1 0 165600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1793
timestamp 1758069660
transform 1 0 166060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1801
timestamp 1758069660
transform 1 0 166796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1808
timestamp 1758069660
transform 1 0 167440 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1815
timestamp 1758069660
transform 1 0 168084 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1827
timestamp 1758069660
transform 1 0 169188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1839
timestamp 1758069660
transform 1 0 170292 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1847
timestamp 1758069660
transform 1 0 171028 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1849
timestamp 1758069660
transform 1 0 171212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1861
timestamp 1758069660
transform 1 0 172316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1873
timestamp 1758069660
transform 1 0 173420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1885
timestamp 1758069660
transform 1 0 174524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1889
timestamp 1758069660
transform 1 0 174892 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1893
timestamp 1758069660
transform 1 0 175260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1900
timestamp 1758069660
transform 1 0 175904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1925
timestamp 1758069660
transform 1 0 178204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1949
timestamp 1758069660
transform 1 0 180412 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1956
timestamp 1758069660
transform 1 0 181056 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1964
timestamp 1758069660
transform 1 0 181792 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1971
timestamp 1758069660
transform 1 0 182436 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1983
timestamp 1758069660
transform 1 0 183540 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1995
timestamp 1758069660
transform 1 0 184644 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2007
timestamp 1758069660
transform 1 0 185748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2015
timestamp 1758069660
transform 1 0 186484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2017
timestamp 1758069660
transform 1 0 186668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2029
timestamp 1758069660
transform 1 0 187772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2033
timestamp 1758069660
transform 1 0 188140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2041
timestamp 1758069660
transform 1 0 188876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2049
timestamp 1758069660
transform 1 0 189612 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_2057
timestamp 1758069660
transform 1 0 190348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2068
timestamp 1758069660
transform 1 0 191360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2082
timestamp 1758069660
transform 1 0 192648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2109
timestamp 1758069660
transform 1 0 195132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2122
timestamp 1758069660
transform 1 0 196328 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_2138
timestamp 1758069660
transform 1 0 197800 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2145
timestamp 1758069660
transform 1 0 198444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2157
timestamp 1758069660
transform 1 0 199548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_2165
timestamp 1758069660
transform 1 0 200284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2170
timestamp 1758069660
transform 1 0 200744 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2177
timestamp 1758069660
transform 1 0 201388 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2183
timestamp 1758069660
transform 1 0 201940 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2185
timestamp 1758069660
transform 1 0 202124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2189
timestamp 1758069660
transform 1 0 202492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2210
timestamp 1758069660
transform 1 0 204424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2234
timestamp 1758069660
transform 1 0 206632 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2244
timestamp 1758069660
transform 1 0 207552 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2256
timestamp 1758069660
transform 1 0 208656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2268
timestamp 1758069660
transform 1 0 209760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2280
timestamp 1758069660
transform 1 0 210864 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2292
timestamp 1758069660
transform 1 0 211968 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2297
timestamp 1758069660
transform 1 0 212428 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2309
timestamp 1758069660
transform 1 0 213532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2321
timestamp 1758069660
transform 1 0 214636 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2333
timestamp 1758069660
transform 1 0 215740 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2345
timestamp 1758069660
transform 1 0 216844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2351
timestamp 1758069660
transform 1 0 217396 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2353
timestamp 1758069660
transform 1 0 217580 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2365
timestamp 1758069660
transform 1 0 218684 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2377
timestamp 1758069660
transform 1 0 219788 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2389
timestamp 1758069660
transform 1 0 220892 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2401
timestamp 1758069660
transform 1 0 221996 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2407
timestamp 1758069660
transform 1 0 222548 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2409
timestamp 1758069660
transform 1 0 222732 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2421
timestamp 1758069660
transform 1 0 223836 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2433
timestamp 1758069660
transform 1 0 224940 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2445
timestamp 1758069660
transform 1 0 226044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2449
timestamp 1758069660
transform 1 0 226412 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2453
timestamp 1758069660
transform 1 0 226780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2460
timestamp 1758069660
transform 1 0 227424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2485
timestamp 1758069660
transform 1 0 229724 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2492
timestamp 1758069660
transform 1 0 230368 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2516
timestamp 1758069660
transform 1 0 232576 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2524
timestamp 1758069660
transform 1 0 233312 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2536
timestamp 1758069660
transform 1 0 234416 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2548
timestamp 1758069660
transform 1 0 235520 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_2560
timestamp 1758069660
transform 1 0 236624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2565
timestamp 1758069660
transform 1 0 237084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2572
timestamp 1758069660
transform 1 0 237728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_2577
timestamp 1758069660
transform 1 0 238188 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2600
timestamp 1758069660
transform 1 0 240304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2624
timestamp 1758069660
transform 1 0 242512 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2633
timestamp 1758069660
transform 1 0 243340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2641
timestamp 1758069660
transform 1 0 244076 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2649
timestamp 1758069660
transform 1 0 244812 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2656
timestamp 1758069660
transform 1 0 245456 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2668
timestamp 1758069660
transform 1 0 246560 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2680
timestamp 1758069660
transform 1 0 247664 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2689
timestamp 1758069660
transform 1 0 248492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2701
timestamp 1758069660
transform 1 0 249596 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2710
timestamp 1758069660
transform 1 0 250424 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2718
timestamp 1758069660
transform 1 0 251160 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2723
timestamp 1758069660
transform 1 0 251620 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2736
timestamp 1758069660
transform 1 0 252816 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2765
timestamp 1758069660
transform 1 0 255484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2778
timestamp 1758069660
transform 1 0 256680 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2785
timestamp 1758069660
transform 1 0 257324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_2797
timestamp 1758069660
transform 1 0 258428 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2801
timestamp 1758069660
transform 1 0 258796 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2813
timestamp 1758069660
transform 1 0 259900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2825
timestamp 1758069660
transform 1 0 261004 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2831
timestamp 1758069660
transform 1 0 261556 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2836
timestamp 1758069660
transform 1 0 262016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2844
timestamp 1758069660
transform 1 0 262752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2852
timestamp 1758069660
transform 1 0 263488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2860
timestamp 1758069660
transform 1 0 264224 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2867
timestamp 1758069660
transform 1 0 264868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2891
timestamp 1758069660
transform 1 0 267076 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2904
timestamp 1758069660
transform 1 0 268272 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2933
timestamp 1758069660
transform 1 0 270940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2946
timestamp 1758069660
transform 1 0 272136 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2959
timestamp 1758069660
transform 1 0 273332 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2967
timestamp 1758069660
transform 1 0 274068 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2969
timestamp 1758069660
transform 1 0 274252 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2981
timestamp 1758069660
transform 1 0 275356 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2993
timestamp 1758069660
transform 1 0 276460 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3005
timestamp 1758069660
transform 1 0 277564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3017
timestamp 1758069660
transform 1 0 278668 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3023
timestamp 1758069660
transform 1 0 279220 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3025
timestamp 1758069660
transform 1 0 279404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3037
timestamp 1758069660
transform 1 0 280508 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3049
timestamp 1758069660
transform 1 0 281612 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3061
timestamp 1758069660
transform 1 0 282716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3073
timestamp 1758069660
transform 1 0 283820 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3079
timestamp 1758069660
transform 1 0 284372 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3081
timestamp 1758069660
transform 1 0 284556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3093
timestamp 1758069660
transform 1 0 285660 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3105
timestamp 1758069660
transform 1 0 286764 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3117
timestamp 1758069660
transform 1 0 287868 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3129
timestamp 1758069660
transform 1 0 288972 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3135
timestamp 1758069660
transform 1 0 289524 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3137
timestamp 1758069660
transform 1 0 289708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3149
timestamp 1758069660
transform 1 0 290812 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3161
timestamp 1758069660
transform 1 0 291916 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3173
timestamp 1758069660
transform 1 0 293020 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3185
timestamp 1758069660
transform 1 0 294124 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3191
timestamp 1758069660
transform 1 0 294676 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3193
timestamp 1758069660
transform 1 0 294860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3205
timestamp 1758069660
transform 1 0 295964 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3217
timestamp 1758069660
transform 1 0 297068 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3229
timestamp 1758069660
transform 1 0 298172 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3241
timestamp 1758069660
transform 1 0 299276 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3247
timestamp 1758069660
transform 1 0 299828 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3249
timestamp 1758069660
transform 1 0 300012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3261
timestamp 1758069660
transform 1 0 301116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3273
timestamp 1758069660
transform 1 0 302220 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3280
timestamp 1758069660
transform 1 0 302864 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3292
timestamp 1758069660
transform 1 0 303968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3296
timestamp 1758069660
transform 1 0 304336 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3300
timestamp 1758069660
transform 1 0 304704 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3305
timestamp 1758069660
transform 1 0 305164 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1758069660
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1758069660
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1758069660
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1758069660
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_37
timestamp 1758069660
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1758069660
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_53
timestamp 1758069660
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_57
timestamp 1758069660
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_69
timestamp 1758069660
transform 1 0 7452 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_74
timestamp 1758069660
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1758069660
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1758069660
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_97
timestamp 1758069660
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1758069660
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_113
timestamp 1758069660
transform 1 0 11500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_125
timestamp 1758069660
transform 1 0 12604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1758069660
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_144
timestamp 1758069660
transform 1 0 14352 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_156
timestamp 1758069660
transform 1 0 15456 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_169
timestamp 1758069660
transform 1 0 16652 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_174
timestamp 1758069660
transform 1 0 17112 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1758069660
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1758069660
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1758069660
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_208
timestamp 1758069660
transform 1 0 20240 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1758069660
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_225
timestamp 1758069660
transform 1 0 21804 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_237
timestamp 1758069660
transform 1 0 22908 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_241
timestamp 1758069660
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1758069660
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1758069660
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_265
timestamp 1758069660
transform 1 0 25484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp 1758069660
transform 1 0 26496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_281
timestamp 1758069660
transform 1 0 26956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1758069660
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1758069660
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_332
timestamp 1758069660
transform 1 0 31648 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_337
timestamp 1758069660
transform 1 0 32108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1758069660
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_385
timestamp 1758069660
transform 1 0 36524 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_391
timestamp 1758069660
transform 1 0 37076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_393
timestamp 1758069660
transform 1 0 37260 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1758069660
transform 1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_421
timestamp 1758069660
transform 1 0 39836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_444
timestamp 1758069660
transform 1 0 41952 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_449
timestamp 1758069660
transform 1 0 42412 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_470
timestamp 1758069660
transform 1 0 44344 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_486
timestamp 1758069660
transform 1 0 45816 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_498
timestamp 1758069660
transform 1 0 46920 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_508
timestamp 1758069660
transform 1 0 47840 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_520
timestamp 1758069660
transform 1 0 48944 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_533
timestamp 1758069660
transform 1 0 50140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_538
timestamp 1758069660
transform 1 0 50600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_551
timestamp 1758069660
transform 1 0 51796 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_559
timestamp 1758069660
transform 1 0 52532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_561
timestamp 1758069660
transform 1 0 52716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_584
timestamp 1758069660
transform 1 0 54832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_589
timestamp 1758069660
transform 1 0 55292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_612
timestamp 1758069660
transform 1 0 57408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1758069660
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1758069660
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_648
timestamp 1758069660
transform 1 0 60720 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_660
timestamp 1758069660
transform 1 0 61824 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_676
timestamp 1758069660
transform 1 0 63296 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_688
timestamp 1758069660
transform 1 0 64400 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_701
timestamp 1758069660
transform 1 0 65596 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_708
timestamp 1758069660
transform 1 0 66240 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_720
timestamp 1758069660
transform 1 0 67344 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_729
timestamp 1758069660
transform 1 0 68172 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_737
timestamp 1758069660
transform 1 0 68908 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_742
timestamp 1758069660
transform 1 0 69368 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_754
timestamp 1758069660
transform 1 0 70472 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_757
timestamp 1758069660
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_769
timestamp 1758069660
transform 1 0 71852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_780
timestamp 1758069660
transform 1 0 72864 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_785
timestamp 1758069660
transform 1 0 73324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_808
timestamp 1758069660
transform 1 0 75440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_813
timestamp 1758069660
transform 1 0 75900 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_836
timestamp 1758069660
transform 1 0 78016 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_861
timestamp 1758069660
transform 1 0 80316 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_867
timestamp 1758069660
transform 1 0 80868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_878
timestamp 1758069660
transform 1 0 81880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_885
timestamp 1758069660
transform 1 0 82524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_892
timestamp 1758069660
transform 1 0 83168 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_897
timestamp 1758069660
transform 1 0 83628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_920
timestamp 1758069660
transform 1 0 85744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_925
timestamp 1758069660
transform 1 0 86204 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_948
timestamp 1758069660
transform 1 0 88320 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_973
timestamp 1758069660
transform 1 0 90620 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_979
timestamp 1758069660
transform 1 0 91172 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_981
timestamp 1758069660
transform 1 0 91356 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_989
timestamp 1758069660
transform 1 0 92092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1001
timestamp 1758069660
transform 1 0 93196 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1007
timestamp 1758069660
transform 1 0 93748 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1012
timestamp 1758069660
transform 1 0 94208 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1024
timestamp 1758069660
transform 1 0 95312 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1037
timestamp 1758069660
transform 1 0 96508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1042
timestamp 1758069660
transform 1 0 96968 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1057
timestamp 1758069660
transform 1 0 98348 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1063
timestamp 1758069660
transform 1 0 98900 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1065
timestamp 1758069660
transform 1 0 99084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1088
timestamp 1758069660
transform 1 0 101200 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1093
timestamp 1758069660
transform 1 0 101660 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1116
timestamp 1758069660
transform 1 0 103776 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1141
timestamp 1758069660
transform 1 0 106076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1147
timestamp 1758069660
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1149
timestamp 1758069660
transform 1 0 106812 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1161
timestamp 1758069660
transform 1 0 107916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1173
timestamp 1758069660
transform 1 0 109020 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1180
timestamp 1758069660
transform 1 0 109664 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1192
timestamp 1758069660
transform 1 0 110768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1196
timestamp 1758069660
transform 1 0 111136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1200
timestamp 1758069660
transform 1 0 111504 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1205
timestamp 1758069660
transform 1 0 111964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1228
timestamp 1758069660
transform 1 0 114080 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1233
timestamp 1758069660
transform 1 0 114540 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1256
timestamp 1758069660
transform 1 0 116656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1261
timestamp 1758069660
transform 1 0 117116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1284
timestamp 1758069660
transform 1 0 119232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1298
timestamp 1758069660
transform 1 0 120520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1309
timestamp 1758069660
transform 1 0 121532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1315
timestamp 1758069660
transform 1 0 122084 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1317
timestamp 1758069660
transform 1 0 122268 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1329
timestamp 1758069660
transform 1 0 123372 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1340
timestamp 1758069660
transform 1 0 124384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1345
timestamp 1758069660
transform 1 0 124844 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1355
timestamp 1758069660
transform 1 0 125764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1368
timestamp 1758069660
transform 1 0 126960 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1373
timestamp 1758069660
transform 1 0 127420 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1394
timestamp 1758069660
transform 1 0 129352 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1401
timestamp 1758069660
transform 1 0 129996 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1424
timestamp 1758069660
transform 1 0 132112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1449
timestamp 1758069660
transform 1 0 134412 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1455
timestamp 1758069660
transform 1 0 134964 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1457
timestamp 1758069660
transform 1 0 135148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1469
timestamp 1758069660
transform 1 0 136252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1476
timestamp 1758069660
transform 1 0 136896 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1485
timestamp 1758069660
transform 1 0 137724 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1497
timestamp 1758069660
transform 1 0 138828 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1509
timestamp 1758069660
transform 1 0 139932 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1516
timestamp 1758069660
transform 1 0 140576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1528
timestamp 1758069660
transform 1 0 141680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1544
timestamp 1758069660
transform 1 0 143152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1556
timestamp 1758069660
transform 1 0 144256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1560
timestamp 1758069660
transform 1 0 144624 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1564
timestamp 1758069660
transform 1 0 144992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1569
timestamp 1758069660
transform 1 0 145452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1592
timestamp 1758069660
transform 1 0 147568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1620
timestamp 1758069660
transform 1 0 150144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1625
timestamp 1758069660
transform 1 0 150604 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1648
timestamp 1758069660
transform 1 0 152720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1653
timestamp 1758069660
transform 1 0 153180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1676
timestamp 1758069660
transform 1 0 155296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1684
timestamp 1758069660
transform 1 0 156032 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1691
timestamp 1758069660
transform 1 0 156676 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1699
timestamp 1758069660
transform 1 0 157412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1704
timestamp 1758069660
transform 1 0 157872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1709
timestamp 1758069660
transform 1 0 158332 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1732
timestamp 1758069660
transform 1 0 160448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1757
timestamp 1758069660
transform 1 0 162748 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1763
timestamp 1758069660
transform 1 0 163300 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1785
timestamp 1758069660
transform 1 0 165324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1791
timestamp 1758069660
transform 1 0 165876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1802
timestamp 1758069660
transform 1 0 166888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1810
timestamp 1758069660
transform 1 0 167624 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1818
timestamp 1758069660
transform 1 0 168360 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1821
timestamp 1758069660
transform 1 0 168636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1833
timestamp 1758069660
transform 1 0 169740 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1839
timestamp 1758069660
transform 1 0 170292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1843
timestamp 1758069660
transform 1 0 170660 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1847
timestamp 1758069660
transform 1 0 171028 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1849
timestamp 1758069660
transform 1 0 171212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1861
timestamp 1758069660
transform 1 0 172316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1872
timestamp 1758069660
transform 1 0 173328 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1886
timestamp 1758069660
transform 1 0 174616 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1894
timestamp 1758069660
transform 1 0 175352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1900
timestamp 1758069660
transform 1 0 175904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1925
timestamp 1758069660
transform 1 0 178204 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1931
timestamp 1758069660
transform 1 0 178756 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1953
timestamp 1758069660
transform 1 0 180780 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1959
timestamp 1758069660
transform 1 0 181332 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1970
timestamp 1758069660
transform 1 0 182344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1977
timestamp 1758069660
transform 1 0 182988 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1985
timestamp 1758069660
transform 1 0 183724 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1989
timestamp 1758069660
transform 1 0 184092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2001
timestamp 1758069660
transform 1 0 185196 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2010
timestamp 1758069660
transform 1 0 186024 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2017
timestamp 1758069660
transform 1 0 186668 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2023
timestamp 1758069660
transform 1 0 187220 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2027
timestamp 1758069660
transform 1 0 187588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2040
timestamp 1758069660
transform 1 0 188784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2045
timestamp 1758069660
transform 1 0 189244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2068
timestamp 1758069660
transform 1 0 191360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2096
timestamp 1758069660
transform 1 0 193936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2124
timestamp 1758069660
transform 1 0 196512 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2129
timestamp 1758069660
transform 1 0 196972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2137
timestamp 1758069660
transform 1 0 197708 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_2140
timestamp 1758069660
transform 1 0 197984 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2151
timestamp 1758069660
transform 1 0 198996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2155
timestamp 1758069660
transform 1 0 199364 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2157
timestamp 1758069660
transform 1 0 199548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2163
timestamp 1758069660
transform 1 0 200100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2176
timestamp 1758069660
transform 1 0 201296 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2205
timestamp 1758069660
transform 1 0 203964 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2211
timestamp 1758069660
transform 1 0 204516 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2233
timestamp 1758069660
transform 1 0 206540 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2239
timestamp 1758069660
transform 1 0 207092 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2250
timestamp 1758069660
transform 1 0 208104 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2262
timestamp 1758069660
transform 1 0 209208 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2269
timestamp 1758069660
transform 1 0 209852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2273
timestamp 1758069660
transform 1 0 210220 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2277
timestamp 1758069660
transform 1 0 210588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2289
timestamp 1758069660
transform 1 0 211692 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2295
timestamp 1758069660
transform 1 0 212244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2297
timestamp 1758069660
transform 1 0 212428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_2305
timestamp 1758069660
transform 1 0 213164 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2310
timestamp 1758069660
transform 1 0 213624 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_2322
timestamp 1758069660
transform 1 0 214728 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2325
timestamp 1758069660
transform 1 0 215004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2337
timestamp 1758069660
transform 1 0 216108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2343
timestamp 1758069660
transform 1 0 216660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2351
timestamp 1758069660
transform 1 0 217396 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2353
timestamp 1758069660
transform 1 0 217580 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2365
timestamp 1758069660
transform 1 0 218684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2377
timestamp 1758069660
transform 1 0 219788 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2384
timestamp 1758069660
transform 1 0 220432 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2396
timestamp 1758069660
transform 1 0 221536 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2412
timestamp 1758069660
transform 1 0 223008 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2418
timestamp 1758069660
transform 1 0 223560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2428
timestamp 1758069660
transform 1 0 224480 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2437
timestamp 1758069660
transform 1 0 225308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2444
timestamp 1758069660
transform 1 0 225952 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2450
timestamp 1758069660
transform 1 0 226504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2460
timestamp 1758069660
transform 1 0 227424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2485
timestamp 1758069660
transform 1 0 229724 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2491
timestamp 1758069660
transform 1 0 230276 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2513
timestamp 1758069660
transform 1 0 232300 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2519
timestamp 1758069660
transform 1 0 232852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2524
timestamp 1758069660
transform 1 0 233312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2531
timestamp 1758069660
transform 1 0 233956 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_2539
timestamp 1758069660
transform 1 0 234692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2544
timestamp 1758069660
transform 1 0 235152 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2549
timestamp 1758069660
transform 1 0 235612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2570
timestamp 1758069660
transform 1 0 237544 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2597
timestamp 1758069660
transform 1 0 240028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2603
timestamp 1758069660
transform 1 0 240580 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2625
timestamp 1758069660
transform 1 0 242604 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2631
timestamp 1758069660
transform 1 0 243156 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2653
timestamp 1758069660
transform 1 0 245180 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2659
timestamp 1758069660
transform 1 0 245732 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2661
timestamp 1758069660
transform 1 0 245916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2673
timestamp 1758069660
transform 1 0 247020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2677
timestamp 1758069660
transform 1 0 247388 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2685
timestamp 1758069660
transform 1 0 248124 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2689
timestamp 1758069660
transform 1 0 248492 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2697
timestamp 1758069660
transform 1 0 249228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2709
timestamp 1758069660
transform 1 0 250332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2715
timestamp 1758069660
transform 1 0 250884 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2737
timestamp 1758069660
transform 1 0 252908 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2743
timestamp 1758069660
transform 1 0 253460 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2765
timestamp 1758069660
transform 1 0 255484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2771
timestamp 1758069660
transform 1 0 256036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2793
timestamp 1758069660
transform 1 0 258060 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2799
timestamp 1758069660
transform 1 0 258612 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2801
timestamp 1758069660
transform 1 0 258796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2807
timestamp 1758069660
transform 1 0 259348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2811
timestamp 1758069660
transform 1 0 259716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2823
timestamp 1758069660
transform 1 0 260820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2827
timestamp 1758069660
transform 1 0 261188 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2829
timestamp 1758069660
transform 1 0 261372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2837
timestamp 1758069660
transform 1 0 262108 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2852
timestamp 1758069660
transform 1 0 263488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2857
timestamp 1758069660
transform 1 0 263948 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2880
timestamp 1758069660
transform 1 0 266064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2908
timestamp 1758069660
transform 1 0 268640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2933
timestamp 1758069660
transform 1 0 270940 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2939
timestamp 1758069660
transform 1 0 271492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2961
timestamp 1758069660
transform 1 0 273516 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2967
timestamp 1758069660
transform 1 0 274068 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2972
timestamp 1758069660
transform 1 0 274528 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2979
timestamp 1758069660
transform 1 0 275172 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2991
timestamp 1758069660
transform 1 0 276276 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2995
timestamp 1758069660
transform 1 0 276644 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2997
timestamp 1758069660
transform 1 0 276828 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3005
timestamp 1758069660
transform 1 0 277564 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3011
timestamp 1758069660
transform 1 0 278116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3023
timestamp 1758069660
transform 1 0 279220 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3025
timestamp 1758069660
transform 1 0 279404 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3037
timestamp 1758069660
transform 1 0 280508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3044
timestamp 1758069660
transform 1 0 281152 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3053
timestamp 1758069660
transform 1 0 281980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3065
timestamp 1758069660
transform 1 0 283084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3077
timestamp 1758069660
transform 1 0 284188 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3084
timestamp 1758069660
transform 1 0 284832 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3096
timestamp 1758069660
transform 1 0 285936 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3112
timestamp 1758069660
transform 1 0 287408 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3124
timestamp 1758069660
transform 1 0 288512 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3137
timestamp 1758069660
transform 1 0 289708 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3144
timestamp 1758069660
transform 1 0 290352 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3156
timestamp 1758069660
transform 1 0 291456 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3165
timestamp 1758069660
transform 1 0 292284 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3173
timestamp 1758069660
transform 1 0 293020 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3178
timestamp 1758069660
transform 1 0 293480 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3190
timestamp 1758069660
transform 1 0 294584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3193
timestamp 1758069660
transform 1 0 294860 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3201
timestamp 1758069660
transform 1 0 295596 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3206
timestamp 1758069660
transform 1 0 296056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3211
timestamp 1758069660
transform 1 0 296516 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3219
timestamp 1758069660
transform 1 0 297252 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3221
timestamp 1758069660
transform 1 0 297436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3233
timestamp 1758069660
transform 1 0 298540 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3244
timestamp 1758069660
transform 1 0 299552 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3249
timestamp 1758069660
transform 1 0 300012 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3261
timestamp 1758069660
transform 1 0 301116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3266
timestamp 1758069660
transform 1 0 301576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3270
timestamp 1758069660
transform 1 0 301944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3274
timestamp 1758069660
transform 1 0 302312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3277
timestamp 1758069660
transform 1 0 302588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3283
timestamp 1758069660
transform 1 0 303140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3287
timestamp 1758069660
transform 1 0 303508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3300
timestamp 1758069660
transform 1 0 304704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3305
timestamp 1758069660
transform 1 0 305164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_8  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 303692 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 1758069660
transform 1 0 303876 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input3
timestamp 1758069660
transform 1 0 304336 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  output4
timestamp 1758069660
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output5
timestamp 1758069660
transform 1 0 32844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output6
timestamp 1758069660
transform 1 0 35512 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output7
timestamp 1758069660
transform 1 0 38364 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output8
timestamp 1758069660
transform 1 0 42228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output9
timestamp 1758069660
transform 1 0 44528 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1758069660
transform 1 0 47564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1758069660
transform 1 0 50324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1758069660
transform 1 0 53636 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 1758069660
transform 1 0 57316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output14
timestamp 1758069660
transform 1 0 60444 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output15
timestamp 1758069660
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output16
timestamp 1758069660
transform 1 0 63020 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1758069660
transform 1 0 65964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output18
timestamp 1758069660
transform 1 0 69092 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output19
timestamp 1758069660
transform 1 0 72128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output20
timestamp 1758069660
transform 1 0 75164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output21
timestamp 1758069660
transform 1 0 78476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output22
timestamp 1758069660
transform 1 0 82248 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output23
timestamp 1758069660
transform 1 0 84364 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output24
timestamp 1758069660
transform 1 0 89424 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output25
timestamp 1758069660
transform 1 0 91080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output26
timestamp 1758069660
transform 1 0 7636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output27
timestamp 1758069660
transform 1 0 93932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output28
timestamp 1758069660
transform 1 0 96692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output29
timestamp 1758069660
transform 1 0 98348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output30
timestamp 1758069660
transform 1 0 102856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output31
timestamp 1758069660
transform 1 0 105892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output32
timestamp 1758069660
transform 1 0 109388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output33
timestamp 1758069660
transform 1 0 111228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output34
timestamp 1758069660
transform 1 0 113712 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output35
timestamp 1758069660
transform 1 0 118680 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output36
timestamp 1758069660
transform 1 0 121256 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1758069660
transform 1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output38
timestamp 1758069660
transform 1 0 124108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output39
timestamp 1758069660
transform 1 0 126684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output40
timestamp 1758069660
transform 1 0 130456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output41
timestamp 1758069660
transform 1 0 134320 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output42
timestamp 1758069660
transform 1 0 136620 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output43
timestamp 1758069660
transform 1 0 140300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output44
timestamp 1758069660
transform 1 0 142876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output45
timestamp 1758069660
transform 1 0 144716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output46
timestamp 1758069660
transform 1 0 146832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output47
timestamp 1758069660
transform 1 0 151984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output48
timestamp 1758069660
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output49
timestamp 1758069660
transform 1 0 155756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output50
timestamp 1758069660
transform 1 0 157596 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output51
timestamp 1758069660
transform 1 0 161552 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output52
timestamp 1758069660
transform 1 0 167164 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output53
timestamp 1758069660
transform 1 0 167808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output54
timestamp 1758069660
transform 1 0 170384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output55
timestamp 1758069660
transform 1 0 173052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output56
timestamp 1758069660
transform 1 0 175904 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output57
timestamp 1758069660
transform 1 0 181332 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output58
timestamp 1758069660
transform 1 0 182712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output59
timestamp 1758069660
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output60
timestamp 1758069660
transform 1 0 185748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output61
timestamp 1758069660
transform 1 0 187864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output62
timestamp 1758069660
transform 1 0 191820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output63
timestamp 1758069660
transform 1 0 195592 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output64
timestamp 1758069660
transform 1 0 198168 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output65
timestamp 1758069660
transform 1 0 201112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output66
timestamp 1758069660
transform 1 0 204700 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output67
timestamp 1758069660
transform 1 0 207276 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output68
timestamp 1758069660
transform 1 0 210312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output69
timestamp 1758069660
transform 1 0 213348 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output70
timestamp 1758069660
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output71
timestamp 1758069660
transform 1 0 216384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output72
timestamp 1758069660
transform 1 0 220156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output73
timestamp 1758069660
transform 1 0 222732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output74
timestamp 1758069660
transform 1 0 225676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output75
timestamp 1758069660
transform 1 0 229724 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output76
timestamp 1758069660
transform 1 0 233680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output77
timestamp 1758069660
transform 1 0 234876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output78
timestamp 1758069660
transform 1 0 237452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output79
timestamp 1758069660
transform 1 0 242328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output80
timestamp 1758069660
transform 1 0 244168 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output81
timestamp 1758069660
transform 1 0 23000 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output82
timestamp 1758069660
transform 1 0 247112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output83
timestamp 1758069660
transform 1 0 250148 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output84
timestamp 1758069660
transform 1 0 254380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output85
timestamp 1758069660
transform 1 0 256864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output86
timestamp 1758069660
transform 1 0 259440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output87
timestamp 1758069660
transform 1 0 262476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output88
timestamp 1758069660
transform 1 0 265512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output89
timestamp 1758069660
transform 1 0 269008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output90
timestamp 1758069660
transform 1 0 274252 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output91
timestamp 1758069660
transform 1 0 274896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output92
timestamp 1758069660
transform 1 0 26036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output93
timestamp 1758069660
transform 1 0 277840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output94
timestamp 1758069660
transform 1 0 280876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output95
timestamp 1758069660
transform 1 0 284556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output96
timestamp 1758069660
transform 1 0 287132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output97
timestamp 1758069660
transform 1 0 290076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output98
timestamp 1758069660
transform 1 0 293204 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output99
timestamp 1758069660
transform 1 0 296240 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output100
timestamp 1758069660
transform 1 0 299276 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output101
timestamp 1758069660
transform 1 0 302588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output102
timestamp 1758069660
transform 1 0 304428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output103
timestamp 1758069660
transform 1 0 27784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output104
timestamp 1758069660
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1758069660
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1758069660
transform -1 0 305808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1758069660
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1758069660
transform -1 0 305808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1758069660
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1758069660
transform -1 0 305808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1758069660
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1758069660
transform -1 0 305808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1758069660
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1758069660
transform -1 0 305808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1758069660
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1758069660
transform -1 0 305808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1758069660
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1758069660
transform -1 0 305808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1758069660
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1758069660
transform -1 0 305808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1758069660
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1758069660
transform -1 0 305808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1758069660
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1758069660
transform -1 0 305808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1758069660
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1758069660
transform -1 0 305808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1758069660
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1758069660
transform -1 0 305808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1758069660
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1758069660
transform -1 0 305808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1758069660
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1758069660
transform -1 0 305808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1758069660
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1758069660
transform -1 0 305808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1758069660
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1758069660
transform -1 0 305808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1758069660
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1758069660
transform -1 0 305808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1758069660
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1758069660
transform -1 0 305808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1758069660
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1758069660
transform -1 0 305808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1758069660
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1758069660
transform -1 0 305808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1758069660
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1758069660
transform -1 0 305808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1758069660
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1758069660
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1758069660
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1758069660
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1758069660
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1758069660
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1758069660
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1758069660
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1758069660
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1758069660
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1758069660
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1758069660
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1758069660
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1758069660
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1758069660
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1758069660
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1758069660
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1758069660
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1758069660
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1758069660
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1758069660
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1758069660
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1758069660
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1758069660
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1758069660
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1758069660
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1758069660
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1758069660
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1758069660
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1758069660
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1758069660
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1758069660
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1758069660
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1758069660
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1758069660
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1758069660
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1758069660
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1758069660
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1758069660
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1758069660
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1758069660
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1758069660
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1758069660
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1758069660
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1758069660
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1758069660
transform 1 0 119600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1758069660
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1758069660
transform 1 0 124752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1758069660
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1758069660
transform 1 0 129904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1758069660
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1758069660
transform 1 0 135056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1758069660
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1758069660
transform 1 0 140208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1758069660
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1758069660
transform 1 0 145360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1758069660
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1758069660
transform 1 0 150512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1758069660
transform 1 0 153088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1758069660
transform 1 0 155664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1758069660
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1758069660
transform 1 0 160816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1758069660
transform 1 0 163392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1758069660
transform 1 0 165968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1758069660
transform 1 0 168544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1758069660
transform 1 0 171120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1758069660
transform 1 0 173696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1758069660
transform 1 0 176272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1758069660
transform 1 0 178848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1758069660
transform 1 0 181424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1758069660
transform 1 0 184000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1758069660
transform 1 0 186576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1758069660
transform 1 0 189152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1758069660
transform 1 0 191728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1758069660
transform 1 0 194304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1758069660
transform 1 0 196880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1758069660
transform 1 0 199456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1758069660
transform 1 0 202032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1758069660
transform 1 0 204608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1758069660
transform 1 0 207184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1758069660
transform 1 0 209760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1758069660
transform 1 0 212336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1758069660
transform 1 0 214912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1758069660
transform 1 0 217488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1758069660
transform 1 0 220064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1758069660
transform 1 0 222640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1758069660
transform 1 0 225216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1758069660
transform 1 0 227792 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1758069660
transform 1 0 230368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1758069660
transform 1 0 232944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1758069660
transform 1 0 235520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1758069660
transform 1 0 238096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1758069660
transform 1 0 240672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1758069660
transform 1 0 243248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1758069660
transform 1 0 245824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1758069660
transform 1 0 248400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1758069660
transform 1 0 250976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1758069660
transform 1 0 253552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1758069660
transform 1 0 256128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1758069660
transform 1 0 258704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1758069660
transform 1 0 261280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1758069660
transform 1 0 263856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1758069660
transform 1 0 266432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1758069660
transform 1 0 269008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1758069660
transform 1 0 271584 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1758069660
transform 1 0 274160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1758069660
transform 1 0 276736 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1758069660
transform 1 0 279312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1758069660
transform 1 0 281888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1758069660
transform 1 0 284464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1758069660
transform 1 0 287040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1758069660
transform 1 0 289616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1758069660
transform 1 0 292192 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1758069660
transform 1 0 294768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1758069660
transform 1 0 297344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1758069660
transform 1 0 299920 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1758069660
transform 1 0 302496 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1758069660
transform 1 0 305072 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1758069660
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1758069660
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1758069660
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1758069660
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1758069660
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1758069660
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1758069660
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1758069660
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1758069660
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1758069660
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1758069660
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1758069660
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1758069660
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1758069660
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1758069660
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1758069660
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1758069660
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1758069660
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1758069660
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1758069660
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1758069660
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1758069660
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1758069660
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1758069660
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1758069660
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1758069660
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1758069660
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1758069660
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1758069660
transform 1 0 150512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1758069660
transform 1 0 155664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1758069660
transform 1 0 160816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1758069660
transform 1 0 165968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1758069660
transform 1 0 171120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1758069660
transform 1 0 176272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1758069660
transform 1 0 181424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1758069660
transform 1 0 186576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1758069660
transform 1 0 191728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1758069660
transform 1 0 196880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1758069660
transform 1 0 202032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1758069660
transform 1 0 207184 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1758069660
transform 1 0 212336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1758069660
transform 1 0 217488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1758069660
transform 1 0 222640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1758069660
transform 1 0 227792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1758069660
transform 1 0 232944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1758069660
transform 1 0 238096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1758069660
transform 1 0 243248 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1758069660
transform 1 0 248400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1758069660
transform 1 0 253552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1758069660
transform 1 0 258704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1758069660
transform 1 0 263856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1758069660
transform 1 0 269008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1758069660
transform 1 0 274160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1758069660
transform 1 0 279312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1758069660
transform 1 0 284464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1758069660
transform 1 0 289616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1758069660
transform 1 0 294768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1758069660
transform 1 0 299920 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1758069660
transform 1 0 305072 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1758069660
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1758069660
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1758069660
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1758069660
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1758069660
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1758069660
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1758069660
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1758069660
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1758069660
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1758069660
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1758069660
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1758069660
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1758069660
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1758069660
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1758069660
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1758069660
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1758069660
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1758069660
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1758069660
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1758069660
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1758069660
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1758069660
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1758069660
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1758069660
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1758069660
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1758069660
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1758069660
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1758069660
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1758069660
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1758069660
transform 1 0 153088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1758069660
transform 1 0 158240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1758069660
transform 1 0 163392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1758069660
transform 1 0 168544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1758069660
transform 1 0 173696 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1758069660
transform 1 0 178848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1758069660
transform 1 0 184000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1758069660
transform 1 0 189152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1758069660
transform 1 0 194304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1758069660
transform 1 0 199456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1758069660
transform 1 0 204608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1758069660
transform 1 0 209760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1758069660
transform 1 0 214912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1758069660
transform 1 0 220064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1758069660
transform 1 0 225216 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1758069660
transform 1 0 230368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1758069660
transform 1 0 235520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1758069660
transform 1 0 240672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1758069660
transform 1 0 245824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1758069660
transform 1 0 250976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1758069660
transform 1 0 256128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1758069660
transform 1 0 261280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1758069660
transform 1 0 266432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1758069660
transform 1 0 271584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1758069660
transform 1 0 276736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1758069660
transform 1 0 281888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1758069660
transform 1 0 287040 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1758069660
transform 1 0 292192 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1758069660
transform 1 0 297344 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1758069660
transform 1 0 302496 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1758069660
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1758069660
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1758069660
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1758069660
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1758069660
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1758069660
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1758069660
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1758069660
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1758069660
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1758069660
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1758069660
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1758069660
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1758069660
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1758069660
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1758069660
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1758069660
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1758069660
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1758069660
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1758069660
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1758069660
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1758069660
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1758069660
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1758069660
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1758069660
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1758069660
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1758069660
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1758069660
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1758069660
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1758069660
transform 1 0 150512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1758069660
transform 1 0 155664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1758069660
transform 1 0 160816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1758069660
transform 1 0 165968 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1758069660
transform 1 0 171120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1758069660
transform 1 0 176272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1758069660
transform 1 0 181424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1758069660
transform 1 0 186576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1758069660
transform 1 0 191728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1758069660
transform 1 0 196880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1758069660
transform 1 0 202032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1758069660
transform 1 0 207184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1758069660
transform 1 0 212336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1758069660
transform 1 0 217488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1758069660
transform 1 0 222640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1758069660
transform 1 0 227792 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1758069660
transform 1 0 232944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1758069660
transform 1 0 238096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1758069660
transform 1 0 243248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1758069660
transform 1 0 248400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1758069660
transform 1 0 253552 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1758069660
transform 1 0 258704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1758069660
transform 1 0 263856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1758069660
transform 1 0 269008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1758069660
transform 1 0 274160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1758069660
transform 1 0 279312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1758069660
transform 1 0 284464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1758069660
transform 1 0 289616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1758069660
transform 1 0 294768 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1758069660
transform 1 0 299920 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1758069660
transform 1 0 305072 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1758069660
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1758069660
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1758069660
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1758069660
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1758069660
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1758069660
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1758069660
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1758069660
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1758069660
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1758069660
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1758069660
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1758069660
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1758069660
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1758069660
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1758069660
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1758069660
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1758069660
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1758069660
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1758069660
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1758069660
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1758069660
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1758069660
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1758069660
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1758069660
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1758069660
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1758069660
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1758069660
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1758069660
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1758069660
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1758069660
transform 1 0 153088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1758069660
transform 1 0 158240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1758069660
transform 1 0 163392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1758069660
transform 1 0 168544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1758069660
transform 1 0 173696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1758069660
transform 1 0 178848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1758069660
transform 1 0 184000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1758069660
transform 1 0 189152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1758069660
transform 1 0 194304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1758069660
transform 1 0 199456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1758069660
transform 1 0 204608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1758069660
transform 1 0 209760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1758069660
transform 1 0 214912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1758069660
transform 1 0 220064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1758069660
transform 1 0 225216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1758069660
transform 1 0 230368 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1758069660
transform 1 0 235520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1758069660
transform 1 0 240672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1758069660
transform 1 0 245824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1758069660
transform 1 0 250976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1758069660
transform 1 0 256128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1758069660
transform 1 0 261280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1758069660
transform 1 0 266432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1758069660
transform 1 0 271584 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1758069660
transform 1 0 276736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1758069660
transform 1 0 281888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1758069660
transform 1 0 287040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1758069660
transform 1 0 292192 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1758069660
transform 1 0 297344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1758069660
transform 1 0 302496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1758069660
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1758069660
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1758069660
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1758069660
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1758069660
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1758069660
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1758069660
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1758069660
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1758069660
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1758069660
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1758069660
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1758069660
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1758069660
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1758069660
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1758069660
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1758069660
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1758069660
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1758069660
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1758069660
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1758069660
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1758069660
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1758069660
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1758069660
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1758069660
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1758069660
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1758069660
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1758069660
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1758069660
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1758069660
transform 1 0 150512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1758069660
transform 1 0 155664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1758069660
transform 1 0 160816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1758069660
transform 1 0 165968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1758069660
transform 1 0 171120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1758069660
transform 1 0 176272 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1758069660
transform 1 0 181424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1758069660
transform 1 0 186576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1758069660
transform 1 0 191728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1758069660
transform 1 0 196880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1758069660
transform 1 0 202032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1758069660
transform 1 0 207184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1758069660
transform 1 0 212336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1758069660
transform 1 0 217488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1758069660
transform 1 0 222640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1758069660
transform 1 0 227792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1758069660
transform 1 0 232944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1758069660
transform 1 0 238096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1758069660
transform 1 0 243248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1758069660
transform 1 0 248400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1758069660
transform 1 0 253552 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1758069660
transform 1 0 258704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1758069660
transform 1 0 263856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1758069660
transform 1 0 269008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1758069660
transform 1 0 274160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1758069660
transform 1 0 279312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1758069660
transform 1 0 284464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1758069660
transform 1 0 289616 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1758069660
transform 1 0 294768 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1758069660
transform 1 0 299920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1758069660
transform 1 0 305072 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1758069660
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1758069660
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1758069660
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1758069660
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1758069660
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1758069660
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1758069660
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1758069660
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1758069660
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1758069660
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1758069660
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1758069660
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1758069660
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1758069660
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1758069660
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1758069660
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1758069660
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1758069660
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1758069660
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1758069660
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1758069660
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1758069660
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1758069660
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1758069660
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1758069660
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1758069660
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1758069660
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1758069660
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1758069660
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1758069660
transform 1 0 153088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1758069660
transform 1 0 158240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1758069660
transform 1 0 163392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1758069660
transform 1 0 168544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1758069660
transform 1 0 173696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1758069660
transform 1 0 178848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1758069660
transform 1 0 184000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1758069660
transform 1 0 189152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1758069660
transform 1 0 194304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1758069660
transform 1 0 199456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1758069660
transform 1 0 204608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1758069660
transform 1 0 209760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1758069660
transform 1 0 214912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1758069660
transform 1 0 220064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1758069660
transform 1 0 225216 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1758069660
transform 1 0 230368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1758069660
transform 1 0 235520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1758069660
transform 1 0 240672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1758069660
transform 1 0 245824 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1758069660
transform 1 0 250976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1758069660
transform 1 0 256128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1758069660
transform 1 0 261280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1758069660
transform 1 0 266432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1758069660
transform 1 0 271584 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1758069660
transform 1 0 276736 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1758069660
transform 1 0 281888 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1758069660
transform 1 0 287040 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1758069660
transform 1 0 292192 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1758069660
transform 1 0 297344 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1758069660
transform 1 0 302496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1758069660
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1758069660
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1758069660
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1758069660
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1758069660
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1758069660
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1758069660
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1758069660
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1758069660
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1758069660
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1758069660
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1758069660
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1758069660
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1758069660
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1758069660
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1758069660
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1758069660
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1758069660
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1758069660
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1758069660
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1758069660
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1758069660
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1758069660
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1758069660
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1758069660
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1758069660
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1758069660
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1758069660
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1758069660
transform 1 0 150512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1758069660
transform 1 0 155664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1758069660
transform 1 0 160816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1758069660
transform 1 0 165968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1758069660
transform 1 0 171120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1758069660
transform 1 0 176272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1758069660
transform 1 0 181424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1758069660
transform 1 0 186576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1758069660
transform 1 0 191728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1758069660
transform 1 0 196880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1758069660
transform 1 0 202032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1758069660
transform 1 0 207184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1758069660
transform 1 0 212336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1758069660
transform 1 0 217488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1758069660
transform 1 0 222640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1758069660
transform 1 0 227792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1758069660
transform 1 0 232944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1758069660
transform 1 0 238096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1758069660
transform 1 0 243248 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1758069660
transform 1 0 248400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1758069660
transform 1 0 253552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1758069660
transform 1 0 258704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1758069660
transform 1 0 263856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1758069660
transform 1 0 269008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1758069660
transform 1 0 274160 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1758069660
transform 1 0 279312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1758069660
transform 1 0 284464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1758069660
transform 1 0 289616 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1758069660
transform 1 0 294768 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1758069660
transform 1 0 299920 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1758069660
transform 1 0 305072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1758069660
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1758069660
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1758069660
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1758069660
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1758069660
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1758069660
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1758069660
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1758069660
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1758069660
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1758069660
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1758069660
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1758069660
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1758069660
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1758069660
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1758069660
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1758069660
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1758069660
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1758069660
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1758069660
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1758069660
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1758069660
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1758069660
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1758069660
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1758069660
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1758069660
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1758069660
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1758069660
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1758069660
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1758069660
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1758069660
transform 1 0 153088 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1758069660
transform 1 0 158240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1758069660
transform 1 0 163392 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1758069660
transform 1 0 168544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1758069660
transform 1 0 173696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1758069660
transform 1 0 178848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1758069660
transform 1 0 184000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1758069660
transform 1 0 189152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1758069660
transform 1 0 194304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1758069660
transform 1 0 199456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1758069660
transform 1 0 204608 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1758069660
transform 1 0 209760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1758069660
transform 1 0 214912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1758069660
transform 1 0 220064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1758069660
transform 1 0 225216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1758069660
transform 1 0 230368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1758069660
transform 1 0 235520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1758069660
transform 1 0 240672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1758069660
transform 1 0 245824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1758069660
transform 1 0 250976 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1758069660
transform 1 0 256128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1758069660
transform 1 0 261280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1758069660
transform 1 0 266432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1758069660
transform 1 0 271584 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1758069660
transform 1 0 276736 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1758069660
transform 1 0 281888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1758069660
transform 1 0 287040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1758069660
transform 1 0 292192 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1758069660
transform 1 0 297344 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1758069660
transform 1 0 302496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1758069660
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1758069660
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1758069660
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1758069660
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1758069660
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1758069660
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1758069660
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1758069660
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1758069660
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1758069660
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1758069660
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1758069660
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1758069660
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1758069660
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1758069660
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1758069660
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1758069660
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1758069660
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1758069660
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1758069660
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1758069660
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1758069660
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1758069660
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1758069660
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1758069660
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1758069660
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1758069660
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1758069660
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1758069660
transform 1 0 150512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1758069660
transform 1 0 155664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1758069660
transform 1 0 160816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1758069660
transform 1 0 165968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1758069660
transform 1 0 171120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1758069660
transform 1 0 176272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1758069660
transform 1 0 181424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1758069660
transform 1 0 186576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1758069660
transform 1 0 191728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1758069660
transform 1 0 196880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1758069660
transform 1 0 202032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1758069660
transform 1 0 207184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1758069660
transform 1 0 212336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1758069660
transform 1 0 217488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1758069660
transform 1 0 222640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1758069660
transform 1 0 227792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1758069660
transform 1 0 232944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1758069660
transform 1 0 238096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1758069660
transform 1 0 243248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1758069660
transform 1 0 248400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1758069660
transform 1 0 253552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1758069660
transform 1 0 258704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1758069660
transform 1 0 263856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1758069660
transform 1 0 269008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1758069660
transform 1 0 274160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1758069660
transform 1 0 279312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1758069660
transform 1 0 284464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1758069660
transform 1 0 289616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1758069660
transform 1 0 294768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1758069660
transform 1 0 299920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1758069660
transform 1 0 305072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1758069660
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1758069660
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1758069660
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1758069660
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1758069660
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1758069660
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1758069660
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1758069660
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1758069660
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1758069660
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1758069660
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1758069660
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1758069660
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1758069660
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1758069660
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1758069660
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1758069660
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1758069660
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1758069660
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1758069660
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1758069660
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1758069660
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1758069660
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1758069660
transform 1 0 122176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1758069660
transform 1 0 127328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1758069660
transform 1 0 132480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1758069660
transform 1 0 137632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1758069660
transform 1 0 142784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1758069660
transform 1 0 147936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1758069660
transform 1 0 153088 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1758069660
transform 1 0 158240 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1758069660
transform 1 0 163392 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1758069660
transform 1 0 168544 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1758069660
transform 1 0 173696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1758069660
transform 1 0 178848 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1758069660
transform 1 0 184000 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1758069660
transform 1 0 189152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1758069660
transform 1 0 194304 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1758069660
transform 1 0 199456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1758069660
transform 1 0 204608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1758069660
transform 1 0 209760 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1758069660
transform 1 0 214912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1758069660
transform 1 0 220064 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1758069660
transform 1 0 225216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1758069660
transform 1 0 230368 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1758069660
transform 1 0 235520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1758069660
transform 1 0 240672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1758069660
transform 1 0 245824 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1758069660
transform 1 0 250976 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1758069660
transform 1 0 256128 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1758069660
transform 1 0 261280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1758069660
transform 1 0 266432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1758069660
transform 1 0 271584 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1758069660
transform 1 0 276736 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1758069660
transform 1 0 281888 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1758069660
transform 1 0 287040 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1758069660
transform 1 0 292192 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1758069660
transform 1 0 297344 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1758069660
transform 1 0 302496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1758069660
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1758069660
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1758069660
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1758069660
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1758069660
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1758069660
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1758069660
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1758069660
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1758069660
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1758069660
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1758069660
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1758069660
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1758069660
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1758069660
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1758069660
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1758069660
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1758069660
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1758069660
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1758069660
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1758069660
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1758069660
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1758069660
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1758069660
transform 1 0 119600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1758069660
transform 1 0 124752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1758069660
transform 1 0 129904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1758069660
transform 1 0 135056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1758069660
transform 1 0 140208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1758069660
transform 1 0 145360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1758069660
transform 1 0 150512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1758069660
transform 1 0 155664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1758069660
transform 1 0 160816 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1758069660
transform 1 0 165968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1758069660
transform 1 0 171120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1758069660
transform 1 0 176272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1758069660
transform 1 0 181424 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1758069660
transform 1 0 186576 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1758069660
transform 1 0 191728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1758069660
transform 1 0 196880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1758069660
transform 1 0 202032 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1758069660
transform 1 0 207184 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1758069660
transform 1 0 212336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1758069660
transform 1 0 217488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1758069660
transform 1 0 222640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1758069660
transform 1 0 227792 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1758069660
transform 1 0 232944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1758069660
transform 1 0 238096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1758069660
transform 1 0 243248 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1758069660
transform 1 0 248400 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1758069660
transform 1 0 253552 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1758069660
transform 1 0 258704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1758069660
transform 1 0 263856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1758069660
transform 1 0 269008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1758069660
transform 1 0 274160 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1758069660
transform 1 0 279312 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1758069660
transform 1 0 284464 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1758069660
transform 1 0 289616 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1758069660
transform 1 0 294768 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1758069660
transform 1 0 299920 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1758069660
transform 1 0 305072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1758069660
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1758069660
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1758069660
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1758069660
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1758069660
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1758069660
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1758069660
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1758069660
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1758069660
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1758069660
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1758069660
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1758069660
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1758069660
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1758069660
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1758069660
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1758069660
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1758069660
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1758069660
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1758069660
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1758069660
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1758069660
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1758069660
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1758069660
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1758069660
transform 1 0 122176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1758069660
transform 1 0 127328 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1758069660
transform 1 0 132480 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1758069660
transform 1 0 137632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1758069660
transform 1 0 142784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1758069660
transform 1 0 147936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1758069660
transform 1 0 153088 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1758069660
transform 1 0 158240 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1758069660
transform 1 0 163392 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1758069660
transform 1 0 168544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1758069660
transform 1 0 173696 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1758069660
transform 1 0 178848 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1758069660
transform 1 0 184000 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1758069660
transform 1 0 189152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1758069660
transform 1 0 194304 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1758069660
transform 1 0 199456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1758069660
transform 1 0 204608 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1758069660
transform 1 0 209760 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1758069660
transform 1 0 214912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1758069660
transform 1 0 220064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1758069660
transform 1 0 225216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1758069660
transform 1 0 230368 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1758069660
transform 1 0 235520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1758069660
transform 1 0 240672 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1758069660
transform 1 0 245824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1758069660
transform 1 0 250976 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1758069660
transform 1 0 256128 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1758069660
transform 1 0 261280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1758069660
transform 1 0 266432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1758069660
transform 1 0 271584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1758069660
transform 1 0 276736 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1758069660
transform 1 0 281888 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1758069660
transform 1 0 287040 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1758069660
transform 1 0 292192 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1758069660
transform 1 0 297344 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1758069660
transform 1 0 302496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1758069660
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1758069660
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1758069660
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1758069660
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1758069660
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1758069660
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1758069660
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1758069660
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1758069660
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1758069660
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1758069660
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1758069660
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1758069660
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1758069660
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1758069660
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1758069660
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1758069660
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1758069660
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1758069660
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1758069660
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1758069660
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1758069660
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1758069660
transform 1 0 119600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1758069660
transform 1 0 124752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1758069660
transform 1 0 129904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1758069660
transform 1 0 135056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1758069660
transform 1 0 140208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1758069660
transform 1 0 145360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1758069660
transform 1 0 150512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1758069660
transform 1 0 155664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1758069660
transform 1 0 160816 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1758069660
transform 1 0 165968 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1758069660
transform 1 0 171120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1758069660
transform 1 0 176272 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1758069660
transform 1 0 181424 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1758069660
transform 1 0 186576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1758069660
transform 1 0 191728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1758069660
transform 1 0 196880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1758069660
transform 1 0 202032 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1758069660
transform 1 0 207184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1758069660
transform 1 0 212336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1758069660
transform 1 0 217488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1758069660
transform 1 0 222640 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1758069660
transform 1 0 227792 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1758069660
transform 1 0 232944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1758069660
transform 1 0 238096 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1758069660
transform 1 0 243248 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1758069660
transform 1 0 248400 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1758069660
transform 1 0 253552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1758069660
transform 1 0 258704 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1758069660
transform 1 0 263856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1758069660
transform 1 0 269008 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1758069660
transform 1 0 274160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1758069660
transform 1 0 279312 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1758069660
transform 1 0 284464 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1758069660
transform 1 0 289616 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1758069660
transform 1 0 294768 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1758069660
transform 1 0 299920 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1758069660
transform 1 0 305072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1758069660
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1758069660
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1758069660
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1758069660
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1758069660
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1758069660
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1758069660
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1758069660
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1758069660
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1758069660
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1758069660
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1758069660
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1758069660
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1758069660
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1758069660
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1758069660
transform 1 0 80960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1758069660
transform 1 0 86112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1758069660
transform 1 0 91264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1758069660
transform 1 0 96416 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1758069660
transform 1 0 101568 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1758069660
transform 1 0 106720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1758069660
transform 1 0 111872 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1758069660
transform 1 0 117024 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1758069660
transform 1 0 122176 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1758069660
transform 1 0 127328 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1758069660
transform 1 0 132480 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1758069660
transform 1 0 137632 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1758069660
transform 1 0 142784 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1758069660
transform 1 0 147936 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1758069660
transform 1 0 153088 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1758069660
transform 1 0 158240 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1758069660
transform 1 0 163392 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1758069660
transform 1 0 168544 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1758069660
transform 1 0 173696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1758069660
transform 1 0 178848 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1758069660
transform 1 0 184000 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1758069660
transform 1 0 189152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1758069660
transform 1 0 194304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1758069660
transform 1 0 199456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1758069660
transform 1 0 204608 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1758069660
transform 1 0 209760 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1758069660
transform 1 0 214912 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1758069660
transform 1 0 220064 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1758069660
transform 1 0 225216 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1758069660
transform 1 0 230368 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1758069660
transform 1 0 235520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1758069660
transform 1 0 240672 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1758069660
transform 1 0 245824 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1758069660
transform 1 0 250976 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1758069660
transform 1 0 256128 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1758069660
transform 1 0 261280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1758069660
transform 1 0 266432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1758069660
transform 1 0 271584 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1758069660
transform 1 0 276736 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1758069660
transform 1 0 281888 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1758069660
transform 1 0 287040 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1758069660
transform 1 0 292192 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1758069660
transform 1 0 297344 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1758069660
transform 1 0 302496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1758069660
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1758069660
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1758069660
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1758069660
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1758069660
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1758069660
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1758069660
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1758069660
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1758069660
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1758069660
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1758069660
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1758069660
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1758069660
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1758069660
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1758069660
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1758069660
transform 1 0 83536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1758069660
transform 1 0 88688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1758069660
transform 1 0 93840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1758069660
transform 1 0 98992 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1758069660
transform 1 0 104144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1758069660
transform 1 0 109296 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1758069660
transform 1 0 114448 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1758069660
transform 1 0 119600 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1758069660
transform 1 0 124752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1758069660
transform 1 0 129904 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1758069660
transform 1 0 135056 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1758069660
transform 1 0 140208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1758069660
transform 1 0 145360 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1758069660
transform 1 0 150512 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1758069660
transform 1 0 155664 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1758069660
transform 1 0 160816 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1758069660
transform 1 0 165968 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1758069660
transform 1 0 171120 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1758069660
transform 1 0 176272 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1758069660
transform 1 0 181424 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1758069660
transform 1 0 186576 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1758069660
transform 1 0 191728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1758069660
transform 1 0 196880 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1758069660
transform 1 0 202032 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1758069660
transform 1 0 207184 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1758069660
transform 1 0 212336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1758069660
transform 1 0 217488 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1758069660
transform 1 0 222640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1758069660
transform 1 0 227792 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1758069660
transform 1 0 232944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1758069660
transform 1 0 238096 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1758069660
transform 1 0 243248 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1758069660
transform 1 0 248400 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1758069660
transform 1 0 253552 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1758069660
transform 1 0 258704 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1758069660
transform 1 0 263856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1758069660
transform 1 0 269008 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1758069660
transform 1 0 274160 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1758069660
transform 1 0 279312 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1758069660
transform 1 0 284464 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1758069660
transform 1 0 289616 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1758069660
transform 1 0 294768 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1758069660
transform 1 0 299920 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1758069660
transform 1 0 305072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1758069660
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1758069660
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1758069660
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1758069660
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1758069660
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1758069660
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1758069660
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1758069660
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1758069660
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1758069660
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1758069660
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1758069660
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1758069660
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1758069660
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1758069660
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1758069660
transform 1 0 80960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1758069660
transform 1 0 86112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1758069660
transform 1 0 91264 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1758069660
transform 1 0 96416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1758069660
transform 1 0 101568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1758069660
transform 1 0 106720 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1758069660
transform 1 0 111872 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1758069660
transform 1 0 117024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1758069660
transform 1 0 122176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1758069660
transform 1 0 127328 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1758069660
transform 1 0 132480 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1758069660
transform 1 0 137632 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1758069660
transform 1 0 142784 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1758069660
transform 1 0 147936 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1758069660
transform 1 0 153088 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1758069660
transform 1 0 158240 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1758069660
transform 1 0 163392 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1758069660
transform 1 0 168544 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1758069660
transform 1 0 173696 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1758069660
transform 1 0 178848 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1758069660
transform 1 0 184000 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1758069660
transform 1 0 189152 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1758069660
transform 1 0 194304 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1758069660
transform 1 0 199456 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1758069660
transform 1 0 204608 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1758069660
transform 1 0 209760 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1758069660
transform 1 0 214912 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1758069660
transform 1 0 220064 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1758069660
transform 1 0 225216 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1758069660
transform 1 0 230368 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1758069660
transform 1 0 235520 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1758069660
transform 1 0 240672 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1758069660
transform 1 0 245824 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1758069660
transform 1 0 250976 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1758069660
transform 1 0 256128 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1758069660
transform 1 0 261280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1758069660
transform 1 0 266432 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1758069660
transform 1 0 271584 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1758069660
transform 1 0 276736 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1758069660
transform 1 0 281888 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1758069660
transform 1 0 287040 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1758069660
transform 1 0 292192 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1758069660
transform 1 0 297344 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1758069660
transform 1 0 302496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1758069660
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1758069660
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1758069660
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1758069660
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1758069660
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1758069660
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1758069660
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1758069660
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1758069660
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1758069660
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1758069660
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1758069660
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1758069660
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1758069660
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1758069660
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1758069660
transform 1 0 83536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1758069660
transform 1 0 88688 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1758069660
transform 1 0 93840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1758069660
transform 1 0 98992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1758069660
transform 1 0 104144 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1758069660
transform 1 0 109296 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1758069660
transform 1 0 114448 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1758069660
transform 1 0 119600 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1758069660
transform 1 0 124752 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1758069660
transform 1 0 129904 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1758069660
transform 1 0 135056 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1758069660
transform 1 0 140208 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1758069660
transform 1 0 145360 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1758069660
transform 1 0 150512 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1758069660
transform 1 0 155664 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1758069660
transform 1 0 160816 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1758069660
transform 1 0 165968 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1758069660
transform 1 0 171120 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1758069660
transform 1 0 176272 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1758069660
transform 1 0 181424 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1758069660
transform 1 0 186576 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1758069660
transform 1 0 191728 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1758069660
transform 1 0 196880 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1758069660
transform 1 0 202032 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1758069660
transform 1 0 207184 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1758069660
transform 1 0 212336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1758069660
transform 1 0 217488 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1758069660
transform 1 0 222640 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1758069660
transform 1 0 227792 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1758069660
transform 1 0 232944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1758069660
transform 1 0 238096 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1758069660
transform 1 0 243248 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1758069660
transform 1 0 248400 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1758069660
transform 1 0 253552 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1758069660
transform 1 0 258704 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1758069660
transform 1 0 263856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1758069660
transform 1 0 269008 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1758069660
transform 1 0 274160 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1758069660
transform 1 0 279312 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1758069660
transform 1 0 284464 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1758069660
transform 1 0 289616 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1758069660
transform 1 0 294768 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1758069660
transform 1 0 299920 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1758069660
transform 1 0 305072 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1758069660
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1758069660
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1758069660
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1758069660
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1758069660
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1758069660
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1758069660
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1758069660
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1758069660
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1758069660
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1758069660
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1758069660
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1758069660
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1758069660
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1758069660
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1758069660
transform 1 0 80960 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1758069660
transform 1 0 86112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1758069660
transform 1 0 91264 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1758069660
transform 1 0 96416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1758069660
transform 1 0 101568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1758069660
transform 1 0 106720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1758069660
transform 1 0 111872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1758069660
transform 1 0 117024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1758069660
transform 1 0 122176 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1758069660
transform 1 0 127328 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1758069660
transform 1 0 132480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1758069660
transform 1 0 137632 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1758069660
transform 1 0 142784 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1758069660
transform 1 0 147936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1758069660
transform 1 0 153088 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1758069660
transform 1 0 158240 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1758069660
transform 1 0 163392 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1758069660
transform 1 0 168544 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1758069660
transform 1 0 173696 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1758069660
transform 1 0 178848 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1758069660
transform 1 0 184000 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1758069660
transform 1 0 189152 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1758069660
transform 1 0 194304 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1758069660
transform 1 0 199456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1758069660
transform 1 0 204608 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1758069660
transform 1 0 209760 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1758069660
transform 1 0 214912 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1758069660
transform 1 0 220064 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1758069660
transform 1 0 225216 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1758069660
transform 1 0 230368 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1758069660
transform 1 0 235520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1758069660
transform 1 0 240672 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1758069660
transform 1 0 245824 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1758069660
transform 1 0 250976 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1758069660
transform 1 0 256128 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1758069660
transform 1 0 261280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1758069660
transform 1 0 266432 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1758069660
transform 1 0 271584 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1758069660
transform 1 0 276736 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1758069660
transform 1 0 281888 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1758069660
transform 1 0 287040 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1758069660
transform 1 0 292192 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1758069660
transform 1 0 297344 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1758069660
transform 1 0 302496 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1758069660
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1758069660
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1758069660
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1758069660
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1758069660
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1758069660
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1758069660
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1758069660
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1758069660
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1758069660
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1758069660
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1758069660
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1758069660
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1758069660
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1758069660
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1758069660
transform 1 0 83536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1758069660
transform 1 0 88688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1758069660
transform 1 0 93840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1758069660
transform 1 0 98992 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1758069660
transform 1 0 104144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1758069660
transform 1 0 109296 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1758069660
transform 1 0 114448 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1758069660
transform 1 0 119600 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1758069660
transform 1 0 124752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1758069660
transform 1 0 129904 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1758069660
transform 1 0 135056 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1758069660
transform 1 0 140208 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1758069660
transform 1 0 145360 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1758069660
transform 1 0 150512 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1758069660
transform 1 0 155664 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1758069660
transform 1 0 160816 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1758069660
transform 1 0 165968 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1758069660
transform 1 0 171120 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1758069660
transform 1 0 176272 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1758069660
transform 1 0 181424 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1758069660
transform 1 0 186576 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1758069660
transform 1 0 191728 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1758069660
transform 1 0 196880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1758069660
transform 1 0 202032 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1758069660
transform 1 0 207184 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1758069660
transform 1 0 212336 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1758069660
transform 1 0 217488 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1758069660
transform 1 0 222640 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1758069660
transform 1 0 227792 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1758069660
transform 1 0 232944 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1758069660
transform 1 0 238096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1758069660
transform 1 0 243248 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1758069660
transform 1 0 248400 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1758069660
transform 1 0 253552 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1758069660
transform 1 0 258704 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1758069660
transform 1 0 263856 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1758069660
transform 1 0 269008 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1758069660
transform 1 0 274160 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1758069660
transform 1 0 279312 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1758069660
transform 1 0 284464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1758069660
transform 1 0 289616 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1758069660
transform 1 0 294768 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1758069660
transform 1 0 299920 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1758069660
transform 1 0 305072 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1758069660
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1758069660
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1758069660
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1758069660
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1758069660
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1758069660
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1758069660
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1758069660
transform 1 0 21712 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1758069660
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1758069660
transform 1 0 26864 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1758069660
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1758069660
transform 1 0 32016 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1758069660
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1758069660
transform 1 0 37168 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1758069660
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1758069660
transform 1 0 42320 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1758069660
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1758069660
transform 1 0 47472 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1758069660
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1758069660
transform 1 0 52624 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1758069660
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1758069660
transform 1 0 57776 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1758069660
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1758069660
transform 1 0 62928 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1758069660
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1758069660
transform 1 0 68080 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1758069660
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1758069660
transform 1 0 73232 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1758069660
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1758069660
transform 1 0 78384 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1758069660
transform 1 0 80960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1758069660
transform 1 0 83536 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1758069660
transform 1 0 86112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1758069660
transform 1 0 88688 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1758069660
transform 1 0 91264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1758069660
transform 1 0 93840 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1758069660
transform 1 0 96416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1758069660
transform 1 0 98992 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1758069660
transform 1 0 101568 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1758069660
transform 1 0 104144 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1758069660
transform 1 0 106720 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1758069660
transform 1 0 109296 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1758069660
transform 1 0 111872 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1758069660
transform 1 0 114448 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1758069660
transform 1 0 117024 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1758069660
transform 1 0 119600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1758069660
transform 1 0 122176 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1758069660
transform 1 0 124752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1758069660
transform 1 0 127328 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1758069660
transform 1 0 129904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1758069660
transform 1 0 132480 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1758069660
transform 1 0 135056 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1758069660
transform 1 0 137632 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1758069660
transform 1 0 140208 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1758069660
transform 1 0 142784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1758069660
transform 1 0 145360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1758069660
transform 1 0 147936 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1758069660
transform 1 0 150512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1758069660
transform 1 0 153088 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1758069660
transform 1 0 155664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1758069660
transform 1 0 158240 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1758069660
transform 1 0 160816 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1758069660
transform 1 0 163392 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1758069660
transform 1 0 165968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1758069660
transform 1 0 168544 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1758069660
transform 1 0 171120 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1758069660
transform 1 0 173696 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1758069660
transform 1 0 176272 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1758069660
transform 1 0 178848 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1758069660
transform 1 0 181424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1758069660
transform 1 0 184000 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1758069660
transform 1 0 186576 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1758069660
transform 1 0 189152 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1758069660
transform 1 0 191728 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1758069660
transform 1 0 194304 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1758069660
transform 1 0 196880 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1758069660
transform 1 0 199456 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1758069660
transform 1 0 202032 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1758069660
transform 1 0 204608 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1758069660
transform 1 0 207184 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1758069660
transform 1 0 209760 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1758069660
transform 1 0 212336 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1758069660
transform 1 0 214912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1758069660
transform 1 0 217488 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1758069660
transform 1 0 220064 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1758069660
transform 1 0 222640 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1758069660
transform 1 0 225216 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1758069660
transform 1 0 227792 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1758069660
transform 1 0 230368 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1758069660
transform 1 0 232944 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1758069660
transform 1 0 235520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1758069660
transform 1 0 238096 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1758069660
transform 1 0 240672 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1758069660
transform 1 0 243248 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1758069660
transform 1 0 245824 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1758069660
transform 1 0 248400 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1758069660
transform 1 0 250976 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1758069660
transform 1 0 253552 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1758069660
transform 1 0 256128 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1758069660
transform 1 0 258704 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1758069660
transform 1 0 261280 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1758069660
transform 1 0 263856 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1758069660
transform 1 0 266432 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1758069660
transform 1 0 269008 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1758069660
transform 1 0 271584 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1758069660
transform 1 0 274160 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1758069660
transform 1 0 276736 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1758069660
transform 1 0 279312 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1758069660
transform 1 0 281888 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1758069660
transform 1 0 284464 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1758069660
transform 1 0 287040 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1758069660
transform 1 0 289616 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1758069660
transform 1 0 292192 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1758069660
transform 1 0 294768 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1758069660
transform 1 0 297344 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1758069660
transform 1 0 299920 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1758069660
transform 1 0 302496 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1758069660
transform 1 0 305072 0 1 13056
box -38 -48 130 592
<< labels >>
rlabel metal4 s -1076 -4 -756 15780 4 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 -4 307988 316 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 15460 307988 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 307668 -4 307988 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 77142 -4 77462 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 153340 -4 153660 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 229538 -4 229858 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 4928 307988 5248 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 7840 307988 8160 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 10752 307988 11072 6 GND
port 0 nsew ground bidirectional
rlabel metal2 s 1490 15200 1546 16000 6 ROW_SEL[0]
port 1 nsew signal tristate
rlabel metal2 s 32126 15200 32182 16000 6 ROW_SEL[10]
port 2 nsew signal tristate
rlabel metal2 s 35254 15200 35310 16000 6 ROW_SEL[11]
port 3 nsew signal tristate
rlabel metal2 s 38290 15200 38346 16000 6 ROW_SEL[12]
port 4 nsew signal tristate
rlabel metal2 s 41326 15200 41382 16000 6 ROW_SEL[13]
port 5 nsew signal tristate
rlabel metal2 s 44454 15200 44510 16000 6 ROW_SEL[14]
port 6 nsew signal tristate
rlabel metal2 s 47490 15200 47546 16000 6 ROW_SEL[15]
port 7 nsew signal tristate
rlabel metal2 s 50526 15200 50582 16000 6 ROW_SEL[16]
port 8 nsew signal tristate
rlabel metal2 s 53654 15200 53710 16000 6 ROW_SEL[17]
port 9 nsew signal tristate
rlabel metal2 s 56690 15200 56746 16000 6 ROW_SEL[18]
port 10 nsew signal tristate
rlabel metal2 s 59818 15200 59874 16000 6 ROW_SEL[19]
port 11 nsew signal tristate
rlabel metal2 s 4526 15200 4582 16000 6 ROW_SEL[1]
port 12 nsew signal tristate
rlabel metal2 s 62854 15200 62910 16000 6 ROW_SEL[20]
port 13 nsew signal tristate
rlabel metal2 s 65890 15200 65946 16000 6 ROW_SEL[21]
port 14 nsew signal tristate
rlabel metal2 s 69018 15200 69074 16000 6 ROW_SEL[22]
port 15 nsew signal tristate
rlabel metal2 s 72054 15200 72110 16000 6 ROW_SEL[23]
port 16 nsew signal tristate
rlabel metal2 s 75090 15200 75146 16000 6 ROW_SEL[24]
port 17 nsew signal tristate
rlabel metal2 s 78218 15200 78274 16000 6 ROW_SEL[25]
port 18 nsew signal tristate
rlabel metal2 s 81254 15200 81310 16000 6 ROW_SEL[26]
port 19 nsew signal tristate
rlabel metal2 s 84290 15200 84346 16000 6 ROW_SEL[27]
port 20 nsew signal tristate
rlabel metal2 s 87418 15200 87474 16000 6 ROW_SEL[28]
port 21 nsew signal tristate
rlabel metal2 s 90454 15200 90510 16000 6 ROW_SEL[29]
port 22 nsew signal tristate
rlabel metal2 s 7562 15200 7618 16000 6 ROW_SEL[2]
port 23 nsew signal tristate
rlabel metal2 s 93582 15200 93638 16000 6 ROW_SEL[30]
port 24 nsew signal tristate
rlabel metal2 s 96618 15200 96674 16000 6 ROW_SEL[31]
port 25 nsew signal tristate
rlabel metal2 s 99654 15200 99710 16000 6 ROW_SEL[32]
port 26 nsew signal tristate
rlabel metal2 s 102782 15200 102838 16000 6 ROW_SEL[33]
port 27 nsew signal tristate
rlabel metal2 s 105818 15200 105874 16000 6 ROW_SEL[34]
port 28 nsew signal tristate
rlabel metal2 s 108854 15200 108910 16000 6 ROW_SEL[35]
port 29 nsew signal tristate
rlabel metal2 s 111982 15200 112038 16000 6 ROW_SEL[36]
port 30 nsew signal tristate
rlabel metal2 s 115018 15200 115074 16000 6 ROW_SEL[37]
port 31 nsew signal tristate
rlabel metal2 s 118146 15200 118202 16000 6 ROW_SEL[38]
port 32 nsew signal tristate
rlabel metal2 s 121182 15200 121238 16000 6 ROW_SEL[39]
port 33 nsew signal tristate
rlabel metal2 s 10690 15200 10746 16000 6 ROW_SEL[3]
port 34 nsew signal tristate
rlabel metal2 s 124218 15200 124274 16000 6 ROW_SEL[40]
port 35 nsew signal tristate
rlabel metal2 s 127346 15200 127402 16000 6 ROW_SEL[41]
port 36 nsew signal tristate
rlabel metal2 s 130382 15200 130438 16000 6 ROW_SEL[42]
port 37 nsew signal tristate
rlabel metal2 s 133418 15200 133474 16000 6 ROW_SEL[43]
port 38 nsew signal tristate
rlabel metal2 s 136546 15200 136602 16000 6 ROW_SEL[44]
port 39 nsew signal tristate
rlabel metal2 s 139582 15200 139638 16000 6 ROW_SEL[45]
port 40 nsew signal tristate
rlabel metal2 s 142710 15200 142766 16000 6 ROW_SEL[46]
port 41 nsew signal tristate
rlabel metal2 s 145746 15200 145802 16000 6 ROW_SEL[47]
port 42 nsew signal tristate
rlabel metal2 s 148782 15200 148838 16000 6 ROW_SEL[48]
port 43 nsew signal tristate
rlabel metal2 s 151910 15200 151966 16000 6 ROW_SEL[49]
port 44 nsew signal tristate
rlabel metal2 s 13726 15200 13782 16000 6 ROW_SEL[4]
port 45 nsew signal tristate
rlabel metal2 s 154946 15200 155002 16000 6 ROW_SEL[50]
port 46 nsew signal tristate
rlabel metal2 s 157982 15200 158038 16000 6 ROW_SEL[51]
port 47 nsew signal tristate
rlabel metal2 s 161110 15200 161166 16000 6 ROW_SEL[52]
port 48 nsew signal tristate
rlabel metal2 s 164146 15200 164202 16000 6 ROW_SEL[53]
port 49 nsew signal tristate
rlabel metal2 s 167182 15200 167238 16000 6 ROW_SEL[54]
port 50 nsew signal tristate
rlabel metal2 s 170310 15200 170366 16000 6 ROW_SEL[55]
port 51 nsew signal tristate
rlabel metal2 s 173346 15200 173402 16000 6 ROW_SEL[56]
port 52 nsew signal tristate
rlabel metal2 s 176474 15200 176530 16000 6 ROW_SEL[57]
port 53 nsew signal tristate
rlabel metal2 s 179510 15200 179566 16000 6 ROW_SEL[58]
port 54 nsew signal tristate
rlabel metal2 s 182546 15200 182602 16000 6 ROW_SEL[59]
port 55 nsew signal tristate
rlabel metal2 s 16762 15200 16818 16000 6 ROW_SEL[5]
port 56 nsew signal tristate
rlabel metal2 s 185674 15200 185730 16000 6 ROW_SEL[60]
port 57 nsew signal tristate
rlabel metal2 s 188710 15200 188766 16000 6 ROW_SEL[61]
port 58 nsew signal tristate
rlabel metal2 s 191746 15200 191802 16000 6 ROW_SEL[62]
port 59 nsew signal tristate
rlabel metal2 s 194874 15200 194930 16000 6 ROW_SEL[63]
port 60 nsew signal tristate
rlabel metal2 s 197910 15200 197966 16000 6 ROW_SEL[64]
port 61 nsew signal tristate
rlabel metal2 s 201038 15200 201094 16000 6 ROW_SEL[65]
port 62 nsew signal tristate
rlabel metal2 s 204074 15200 204130 16000 6 ROW_SEL[66]
port 63 nsew signal tristate
rlabel metal2 s 207110 15200 207166 16000 6 ROW_SEL[67]
port 64 nsew signal tristate
rlabel metal2 s 210238 15200 210294 16000 6 ROW_SEL[68]
port 65 nsew signal tristate
rlabel metal2 s 213274 15200 213330 16000 6 ROW_SEL[69]
port 66 nsew signal tristate
rlabel metal2 s 19890 15200 19946 16000 6 ROW_SEL[6]
port 67 nsew signal tristate
rlabel metal2 s 216310 15200 216366 16000 6 ROW_SEL[70]
port 68 nsew signal tristate
rlabel metal2 s 219438 15200 219494 16000 6 ROW_SEL[71]
port 69 nsew signal tristate
rlabel metal2 s 222474 15200 222530 16000 6 ROW_SEL[72]
port 70 nsew signal tristate
rlabel metal2 s 225602 15200 225658 16000 6 ROW_SEL[73]
port 71 nsew signal tristate
rlabel metal2 s 228638 15200 228694 16000 6 ROW_SEL[74]
port 72 nsew signal tristate
rlabel metal2 s 231674 15200 231730 16000 6 ROW_SEL[75]
port 73 nsew signal tristate
rlabel metal2 s 234802 15200 234858 16000 6 ROW_SEL[76]
port 74 nsew signal tristate
rlabel metal2 s 237838 15200 237894 16000 6 ROW_SEL[77]
port 75 nsew signal tristate
rlabel metal2 s 240874 15200 240930 16000 6 ROW_SEL[78]
port 76 nsew signal tristate
rlabel metal2 s 244002 15200 244058 16000 6 ROW_SEL[79]
port 77 nsew signal tristate
rlabel metal2 s 22926 15200 22982 16000 6 ROW_SEL[7]
port 78 nsew signal tristate
rlabel metal2 s 247038 15200 247094 16000 6 ROW_SEL[80]
port 79 nsew signal tristate
rlabel metal2 s 250074 15200 250130 16000 6 ROW_SEL[81]
port 80 nsew signal tristate
rlabel metal2 s 253202 15200 253258 16000 6 ROW_SEL[82]
port 81 nsew signal tristate
rlabel metal2 s 256238 15200 256294 16000 6 ROW_SEL[83]
port 82 nsew signal tristate
rlabel metal2 s 259366 15200 259422 16000 6 ROW_SEL[84]
port 83 nsew signal tristate
rlabel metal2 s 262402 15200 262458 16000 6 ROW_SEL[85]
port 84 nsew signal tristate
rlabel metal2 s 265438 15200 265494 16000 6 ROW_SEL[86]
port 85 nsew signal tristate
rlabel metal2 s 268566 15200 268622 16000 6 ROW_SEL[87]
port 86 nsew signal tristate
rlabel metal2 s 271602 15200 271658 16000 6 ROW_SEL[88]
port 87 nsew signal tristate
rlabel metal2 s 274638 15200 274694 16000 6 ROW_SEL[89]
port 88 nsew signal tristate
rlabel metal2 s 25962 15200 26018 16000 6 ROW_SEL[8]
port 89 nsew signal tristate
rlabel metal2 s 277766 15200 277822 16000 6 ROW_SEL[90]
port 90 nsew signal tristate
rlabel metal2 s 280802 15200 280858 16000 6 ROW_SEL[91]
port 91 nsew signal tristate
rlabel metal2 s 283930 15200 283986 16000 6 ROW_SEL[92]
port 92 nsew signal tristate
rlabel metal2 s 286966 15200 287022 16000 6 ROW_SEL[93]
port 93 nsew signal tristate
rlabel metal2 s 290002 15200 290058 16000 6 ROW_SEL[94]
port 94 nsew signal tristate
rlabel metal2 s 293130 15200 293186 16000 6 ROW_SEL[95]
port 95 nsew signal tristate
rlabel metal2 s 296166 15200 296222 16000 6 ROW_SEL[96]
port 96 nsew signal tristate
rlabel metal2 s 299202 15200 299258 16000 6 ROW_SEL[97]
port 97 nsew signal tristate
rlabel metal2 s 302330 15200 302386 16000 6 ROW_SEL[98]
port 98 nsew signal tristate
rlabel metal2 s 305366 15200 305422 16000 6 ROW_SEL[99]
port 99 nsew signal tristate
rlabel metal2 s 29090 15200 29146 16000 6 ROW_SEL[9]
port 100 nsew signal tristate
rlabel metal4 s -416 656 -96 15120 4 VDD
port 101 nsew power bidirectional
rlabel metal5 s -416 656 307328 976 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -416 14800 307328 15120 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 307008 656 307328 15120 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 39042 -4 39362 15780 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 115240 -4 115560 15780 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 191438 -4 191758 15780 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 267636 -4 267956 15780 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -1076 3472 307988 3792 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -1076 6384 307988 6704 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -1076 9296 307988 9616 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -1076 12208 307988 12528 6 VDD
port 101 nsew power bidirectional
rlabel metal3 s 306200 1912 307000 2032 6 clk
port 102 nsew signal input
rlabel metal3 s 306200 13880 307000 14000 6 data_in
port 103 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 data_out
port 104 nsew signal tristate
rlabel metal3 s 306200 5856 307000 5976 6 ena
port 105 nsew signal input
rlabel metal3 s 306200 9936 307000 10056 6 rst
port 106 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 307000 16000
<< end >>
