magic
tech sky130A
timestamp 1758222970
<< metal5 >>
rect 15800 54600 18800 55700
rect 35300 55400 35600 55700
rect 15800 52800 16300 54600
rect 15800 52300 16200 52800
rect 17200 48400 17500 54600
rect 18500 52300 18800 54600
rect 20600 53600 21500 53800
rect 23780 53600 24000 53620
rect 24600 53600 25400 53800
rect 27800 53600 28300 53800
rect 29000 53600 29600 53800
rect 31800 53600 32800 53800
rect 35200 53600 35600 55400
rect 42500 55100 43800 56200
rect 46700 55400 48000 55700
rect 48200 55400 48500 55700
rect 46400 55100 48600 55400
rect 39400 53600 40200 53800
rect 20400 53300 21800 53600
rect 23000 53460 24000 53600
rect 20200 53100 22100 53300
rect 23000 53100 23940 53460
rect 24200 53300 25700 53600
rect 26800 53300 27440 53600
rect 27600 53300 28600 53600
rect 28800 53300 29900 53600
rect 31600 53300 33000 53600
rect 24100 53100 25900 53300
rect 20000 52800 22200 53100
rect 23000 52800 26000 53100
rect 26600 52800 30000 53300
rect 31300 53100 33200 53300
rect 31200 52800 33400 53100
rect 34600 52800 37200 53600
rect 38900 53300 40400 53600
rect 38600 53100 40700 53300
rect 38600 52800 40800 53100
rect 19900 52500 20800 52800
rect 21400 52500 22300 52800
rect 23200 52500 24700 52800
rect 25300 52500 26200 52800
rect 26800 52500 28000 52800
rect 28200 52500 29200 52800
rect 29500 52500 30100 52800
rect 31100 52500 31900 52800
rect 32600 52500 33500 52800
rect 34700 52500 37100 52800
rect 38600 52500 39400 52800
rect 40100 52500 40800 52800
rect 19800 52300 20500 52500
rect 21600 52300 22400 52500
rect 19800 52000 20400 52300
rect 21800 52000 22400 52300
rect 23500 52300 24500 52500
rect 25600 52300 26300 52500
rect 23500 52000 24400 52300
rect 25700 52000 26300 52300
rect 27000 52300 27700 52500
rect 28300 52300 29000 52500
rect 19700 51800 20300 52000
rect 19700 51500 20200 51800
rect 22000 51500 22600 52000
rect 19600 51200 20200 51500
rect 19600 49900 20000 51200
rect 22100 51000 22600 51500
rect 23500 51800 24200 52000
rect 25800 51800 26400 52000
rect 23500 51500 24100 51800
rect 22100 50700 22700 51000
rect 22200 50200 22700 50700
rect 19600 49700 20200 49900
rect 19700 49400 20200 49700
rect 22100 49400 22600 50200
rect 19700 48900 20300 49400
rect 22000 49100 22600 49400
rect 23500 49900 24000 51500
rect 25900 51000 26400 51800
rect 26000 50700 26400 51000
rect 27000 51800 27600 52300
rect 28300 51800 28900 52300
rect 26000 50400 26500 50700
rect 23500 49700 24100 49900
rect 25900 49700 26400 50400
rect 23500 49100 24200 49700
rect 25800 49400 26400 49700
rect 25700 49100 26300 49400
rect 21800 48900 22400 49100
rect 19800 48600 20500 48900
rect 21700 48600 22400 48900
rect 23500 48900 24500 49100
rect 25600 48900 26300 49100
rect 23500 48600 24600 48900
rect 25300 48600 26200 48900
rect 19900 48400 20600 48600
rect 21500 48400 22300 48600
rect 23500 48400 26000 48600
rect 27000 48400 27500 51800
rect 28300 48400 28800 51800
rect 29600 48400 30100 52500
rect 31000 52300 31700 52500
rect 32900 52300 33600 52500
rect 30800 52000 31600 52300
rect 33000 52000 33600 52300
rect 30800 51800 31400 52000
rect 33100 51800 33700 52000
rect 30800 51500 31300 51800
rect 30700 51200 31300 51500
rect 33200 51200 33700 51800
rect 30700 50200 33800 51200
rect 30700 49700 31300 50200
rect 30800 49400 31300 49700
rect 30800 49100 31400 49400
rect 31000 48900 31600 49100
rect 33500 48900 33700 49100
rect 35200 48900 35600 52500
rect 38600 52300 38900 52500
rect 40300 52300 40900 52500
rect 39500 51200 40200 51500
rect 40400 51200 40900 52300
rect 38900 51000 40900 51200
rect 38600 50700 40900 51000
rect 38500 50400 40900 50700
rect 38400 50200 39400 50400
rect 40200 50200 40900 50400
rect 38400 49900 39100 50200
rect 38300 49700 38900 49900
rect 38300 48900 38800 49700
rect 40400 49100 40900 50200
rect 40200 48900 40900 49100
rect 31000 48600 31700 48900
rect 33200 48600 33800 48900
rect 35200 48600 35800 48900
rect 37200 48600 37600 48900
rect 38300 48600 38900 48900
rect 40100 48600 40900 48900
rect 31100 48400 31900 48600
rect 33000 48400 33800 48600
rect 35300 48400 35900 48600
rect 37000 48400 37600 48600
rect 16300 47600 18400 48400
rect 19900 48100 22200 48400
rect 20000 47800 22100 48100
rect 23500 47940 23940 48400
rect 24100 48100 25900 48400
rect 20300 47600 22000 47800
rect 20500 47300 21700 47600
rect 23500 45800 24000 47940
rect 24200 47800 25800 48100
rect 24500 47600 25400 47800
rect 26600 47600 27800 48400
rect 28300 47600 29200 48400
rect 29600 47600 30500 48400
rect 31200 48100 33700 48400
rect 35300 48100 37600 48400
rect 38400 48400 39000 48600
rect 39800 48400 40900 48600
rect 43300 48400 43800 55100
rect 46300 54900 48600 55100
rect 46200 54600 47200 54900
rect 47500 54600 48600 54900
rect 46200 54400 46800 54600
rect 47800 54400 48600 54600
rect 46100 54100 46700 54400
rect 46100 52800 46600 54100
rect 48000 53800 48600 54400
rect 48100 53100 48600 53800
rect 50500 53600 51500 53800
rect 50300 53300 51700 53600
rect 50000 53100 52000 53300
rect 49900 52800 52100 53100
rect 46100 52500 46700 52800
rect 49800 52500 50600 52800
rect 51400 52500 52200 52800
rect 46200 52300 46900 52500
rect 49700 52300 50400 52500
rect 51600 52300 52300 52500
rect 46200 52000 47400 52300
rect 49600 52000 50300 52300
rect 51700 52000 52300 52300
rect 46300 51800 48000 52000
rect 49600 51800 50200 52000
rect 51800 51800 52400 52000
rect 46600 51500 48200 51800
rect 49600 51500 50000 51800
rect 46900 51200 48500 51500
rect 49400 51200 50000 51500
rect 52000 51200 52400 51800
rect 47400 51000 48600 51200
rect 47900 50700 48600 51000
rect 48100 50400 48700 50700
rect 46000 49700 46300 50200
rect 46000 49100 46400 49700
rect 48200 49100 48700 50400
rect 49400 50200 52600 51200
rect 49400 49700 50000 50200
rect 49600 49400 50000 49700
rect 49600 49100 50200 49400
rect 46000 48900 46600 49100
rect 48100 48900 48700 49100
rect 49700 48900 50300 49100
rect 52200 48900 52400 49100
rect 46000 48600 46700 48900
rect 48000 48600 48600 48900
rect 49700 48600 50400 48900
rect 52000 48600 52600 48900
rect 46000 48400 46800 48600
rect 47800 48400 48600 48600
rect 49800 48400 50600 48600
rect 51700 48400 52600 48600
rect 38400 48100 41400 48400
rect 42200 48100 44900 48400
rect 46000 48100 47300 48400
rect 47460 48100 48500 48400
rect 49900 48100 52400 48400
rect 31300 47800 33600 48100
rect 35400 47800 37600 48100
rect 38500 47800 41400 48100
rect 42100 47800 45000 48100
rect 31400 47600 33500 47800
rect 35400 47600 37300 47800
rect 38600 47600 40240 47800
rect 40400 47600 41400 47800
rect 42200 47600 45000 47800
rect 46000 47800 48400 48100
rect 50000 47800 52300 48100
rect 46000 47600 46240 47800
rect 46400 47600 48200 47800
rect 50200 47600 52200 47800
rect 31700 47300 33100 47600
rect 35600 47300 37000 47600
rect 38800 47300 40000 47600
rect 46700 47300 48000 47600
rect 50400 47300 51800 47600
rect 23000 45000 24700 45800
rect 41400 42400 41900 42600
rect 14800 41600 16100 41800
rect 16300 41600 16700 41800
rect 14600 41300 16700 41600
rect 21800 41300 23200 42400
rect 41000 42100 42200 42400
rect 40900 41800 42400 42100
rect 40800 41600 42500 41800
rect 47300 41600 48200 42400
rect 51100 42100 52000 42400
rect 51000 41600 52000 42100
rect 40700 41300 41400 41600
rect 41800 41300 42600 41600
rect 47400 41300 48200 41600
rect 51100 41300 52000 41600
rect 14400 41100 16700 41300
rect 14300 40800 15200 41100
rect 15600 40800 16700 41100
rect 14300 40500 15000 40800
rect 16000 40500 16700 40800
rect 14200 40000 14800 40500
rect 16100 40300 16700 40500
rect 14200 39200 14600 40000
rect 16200 39500 16700 40300
rect 18700 39800 19600 40000
rect 18400 39500 19900 39800
rect 16300 39200 16700 39500
rect 18100 39200 20000 39500
rect 14200 39000 14800 39200
rect 18000 39000 20300 39200
rect 14200 38700 14900 39000
rect 17900 38700 18800 39000
rect 19400 38700 20400 39000
rect 14300 38400 15000 38700
rect 17900 38400 18600 38700
rect 19700 38400 20400 38700
rect 14400 38200 15500 38400
rect 14400 37900 16100 38200
rect 17800 37900 18400 38400
rect 19900 37900 20500 38400
rect 14600 37700 16400 37900
rect 17600 37700 18200 37900
rect 20000 37700 20600 37900
rect 15000 37400 16600 37700
rect 17600 37400 18100 37700
rect 20200 37400 20600 37700
rect 15600 37100 16700 37400
rect 16000 36900 16700 37100
rect 16200 36600 16800 36900
rect 14000 36100 14400 36400
rect 14000 35300 14500 36100
rect 16300 35300 16800 36600
rect 17600 36400 20600 37400
rect 17600 35800 18100 36400
rect 17600 35600 18200 35800
rect 14000 35100 14600 35300
rect 16200 35100 16800 35300
rect 17800 35100 18400 35600
rect 20300 35100 20500 35300
rect 14000 34800 14800 35100
rect 16100 34800 16800 35100
rect 17900 34800 18600 35100
rect 20200 34800 20600 35100
rect 14000 34500 15000 34800
rect 16000 34500 16700 34800
rect 17900 34500 18700 34800
rect 19800 34500 20600 34800
rect 22700 34500 23200 41300
rect 40600 41100 41300 41300
rect 42000 41100 42700 41300
rect 40600 40800 41200 41100
rect 42100 40800 42700 41100
rect 40600 40500 41000 40800
rect 40400 40000 41000 40500
rect 42200 40500 42700 40800
rect 42200 40300 42800 40500
rect 26200 39800 27000 40000
rect 30100 39800 31000 40000
rect 33700 39800 34400 40000
rect 25800 39500 27400 39800
rect 28900 39500 29600 39800
rect 29900 39500 31200 39800
rect 33200 39500 34800 39800
rect 25700 39200 27600 39500
rect 28800 39200 29600 39500
rect 29800 39200 31300 39500
rect 33000 39200 35000 39500
rect 25400 39000 27700 39200
rect 28800 39000 31400 39200
rect 32900 39000 35000 39200
rect 40400 39000 40900 40000
rect 42400 39800 42800 40300
rect 42400 39500 43000 39800
rect 43700 39500 45100 39800
rect 25400 38700 26300 39000
rect 27000 38700 27800 39000
rect 28900 38700 30200 39000
rect 30800 38700 31600 39000
rect 32900 38700 33700 39000
rect 34400 38700 35200 39000
rect 25300 38400 26000 38700
rect 27100 38400 28000 38700
rect 25200 38200 25900 38400
rect 27400 38200 28000 38400
rect 29300 38400 30100 38700
rect 31000 38400 31600 38700
rect 33000 38400 33200 38700
rect 34700 38400 35200 38700
rect 25200 37900 25800 38200
rect 25100 37400 25700 37900
rect 27500 37700 28100 38200
rect 27600 37400 28100 37700
rect 25100 36400 28100 37400
rect 29300 37900 29900 38400
rect 31100 38200 31600 38400
rect 31100 37900 31700 38200
rect 29300 37700 29800 37900
rect 25100 36100 25600 36400
rect 25100 35600 25700 36100
rect 25200 35300 25800 35600
rect 25200 35100 25900 35300
rect 27800 35100 28100 35300
rect 25300 34800 26000 35100
rect 27600 34800 28100 35100
rect 25400 34500 26300 34800
rect 27400 34500 28100 34800
rect 29300 34500 29600 37700
rect 31200 34500 31700 37900
rect 33800 37400 34400 37700
rect 34800 37400 35300 38400
rect 33200 37100 35300 37400
rect 33000 36900 35300 37100
rect 32900 36600 35300 36900
rect 32800 36400 33700 36600
rect 34600 36400 35300 36600
rect 32800 36100 33500 36400
rect 32600 35800 33200 36100
rect 32600 34800 33100 35800
rect 34800 35600 35300 36400
rect 40400 36600 40800 39000
rect 40400 35800 40900 36600
rect 42500 36400 43000 39500
rect 43600 39000 45100 39500
rect 45700 39000 47200 39800
rect 47800 39200 48200 41300
rect 48800 39800 49700 40000
rect 48600 39500 50000 39800
rect 48400 39200 50200 39500
rect 51600 39200 52000 41300
rect 52700 39800 53400 40000
rect 52300 39500 53800 39800
rect 52200 39200 53900 39500
rect 47800 39000 50300 39200
rect 51600 39000 54100 39200
rect 43700 38700 45000 39000
rect 45800 38700 47000 39000
rect 47800 38700 49000 39000
rect 49600 38700 50400 39000
rect 51600 38700 52800 39000
rect 53300 38700 54100 39000
rect 44000 38400 44600 38700
rect 46200 38400 46700 38700
rect 44200 38200 44600 38400
rect 46100 38200 46700 38400
rect 47800 38400 48800 38700
rect 49800 38400 50500 38700
rect 47800 38200 48600 38400
rect 49900 38200 50500 38400
rect 51600 38400 52600 38700
rect 53500 38400 54200 38700
rect 44200 37900 44800 38200
rect 46100 37900 46600 38200
rect 44300 37700 44800 37900
rect 44300 37400 44900 37700
rect 44400 37100 44900 37400
rect 46000 37400 46600 37900
rect 47800 37700 48500 38200
rect 50000 37900 50600 38200
rect 50200 37700 50600 37900
rect 51600 37900 52300 38400
rect 53600 38200 54400 38400
rect 53800 37900 54400 38200
rect 51600 37700 52200 37900
rect 53900 37700 54400 37900
rect 46000 37100 46400 37400
rect 44400 36900 45000 37100
rect 44500 36400 45000 36900
rect 45800 36900 46400 37100
rect 47800 37100 48400 37700
rect 50200 37100 50800 37700
rect 45800 36600 46300 36900
rect 45700 36400 46300 36600
rect 47800 36400 48200 37100
rect 40400 35600 41000 35800
rect 42400 35600 42800 36400
rect 44500 36100 45100 36400
rect 45700 36100 46200 36400
rect 44600 35800 45100 36100
rect 45600 35800 46200 36100
rect 44600 35600 45200 35800
rect 34700 35300 35300 35600
rect 34600 35100 35300 35300
rect 34400 34800 35300 35100
rect 40600 35300 41000 35600
rect 42200 35300 42800 35600
rect 44800 35300 45200 35600
rect 45600 35300 46100 35800
rect 40600 35100 41200 35300
rect 42200 35100 42700 35300
rect 44800 35100 45400 35300
rect 40600 34800 41300 35100
rect 42100 34800 42700 35100
rect 44900 34800 45400 35100
rect 45560 35100 46100 35300
rect 47800 35600 48400 36400
rect 50300 36100 50800 37100
rect 50200 35800 50800 36100
rect 51600 35800 52100 37700
rect 53900 37400 54500 37700
rect 54000 35800 54500 37400
rect 50200 35600 50600 35800
rect 47800 35300 48500 35600
rect 47800 35100 48600 35300
rect 50000 35100 50600 35600
rect 51600 35300 52200 35800
rect 53900 35600 54500 35800
rect 51600 35100 52300 35300
rect 53800 35100 54400 35600
rect 45560 34800 46000 35100
rect 32600 34500 33200 34800
rect 34200 34500 35300 34800
rect 40700 34500 41400 34800
rect 42000 34500 42600 34800
rect 44900 34500 46000 34800
rect 47800 34800 48700 35100
rect 49800 34800 50500 35100
rect 51600 34800 52400 35100
rect 53600 34800 54200 35100
rect 47800 34500 48800 34800
rect 49700 34500 50400 34800
rect 51600 34500 52600 34800
rect 53400 34500 54200 34800
rect 14000 34000 16600 34500
rect 18000 34300 20600 34500
rect 21600 34300 24200 34500
rect 25400 34300 28100 34500
rect 18100 34000 20500 34300
rect 21500 34000 24400 34300
rect 25700 34000 28000 34300
rect 14000 33800 14340 34000
rect 14500 33800 16300 34000
rect 18400 33800 20300 34000
rect 21600 33800 24400 34000
rect 25800 33800 27700 34000
rect 28800 33800 30100 34500
rect 30800 34300 31900 34500
rect 32800 34300 33600 34500
rect 33760 34300 35800 34500
rect 40700 34300 42600 34500
rect 30800 33800 32000 34300
rect 32800 34000 35800 34300
rect 40800 34000 42500 34300
rect 45000 34000 45800 34500
rect 47300 34300 50400 34500
rect 51100 34300 54100 34500
rect 32900 33800 34600 34000
rect 34800 33800 35800 34000
rect 40900 33800 42400 34000
rect 45000 33800 45700 34000
rect 47300 33800 48200 34300
rect 48400 34000 50300 34300
rect 48500 33800 50000 34000
rect 51000 33800 52000 34300
rect 52160 34000 54000 34300
rect 52200 33800 53900 34000
rect 14800 33500 16100 33800
rect 18600 33500 19900 33800
rect 26000 33500 27500 33800
rect 33100 33500 34300 33800
rect 41200 33500 42100 33800
rect 48700 33500 49800 33800
rect 52400 33500 53600 33800
rect 19600 27800 20800 28000
rect 21400 27800 22600 28000
rect 41800 27800 42700 28000
rect 19600 27200 20900 27800
rect 21400 27200 22700 27800
rect 41800 27500 42800 27800
rect 19700 27000 20800 27200
rect 21400 27000 22600 27200
rect 41800 27000 43000 27500
rect 43800 27200 45200 28000
rect 43900 27000 45200 27200
rect 46900 27000 47500 28800
rect 19900 24600 20300 27000
rect 21800 24600 22300 27000
rect 42200 26400 43100 27000
rect 24400 25900 25200 26200
rect 29300 25900 29600 26200
rect 33000 25900 33400 26200
rect 42200 25900 43200 26400
rect 23900 25700 25400 25900
rect 27400 25700 28300 25900
rect 28900 25700 30000 25900
rect 31100 25700 32000 25900
rect 32600 25700 33700 25900
rect 23600 25400 25700 25700
rect 23600 25100 25800 25400
rect 27200 25100 28300 25700
rect 28800 25400 30100 25700
rect 28600 25100 30200 25400
rect 31000 25100 32000 25700
rect 32500 25400 33800 25700
rect 32300 25100 34000 25400
rect 23600 24900 24400 25100
rect 25100 24900 25800 25100
rect 27400 24900 28300 25100
rect 28460 24900 29340 25100
rect 29500 24900 30200 25100
rect 31100 24900 32000 25100
rect 32200 24900 33100 25100
rect 33260 24900 34000 25100
rect 34600 25100 35800 25900
rect 36600 25100 37800 25900
rect 34600 24900 35600 25100
rect 36700 24900 37800 25100
rect 42200 25700 43300 25900
rect 42200 24940 42640 25700
rect 42800 25100 43400 25700
rect 23600 24600 23900 24900
rect 25300 24600 25900 24900
rect 19900 23600 22300 24600
rect 24500 23600 25200 23800
rect 25400 23600 25900 24600
rect 19900 20700 20300 23600
rect 21800 20700 22300 23600
rect 23900 23300 25900 23600
rect 23600 23100 25900 23300
rect 23500 22800 25900 23100
rect 23400 22500 24400 22800
rect 25200 22500 25900 22800
rect 23400 22300 24100 22500
rect 23300 22000 23900 22300
rect 23300 21200 23800 22000
rect 25400 21500 25900 22500
rect 25200 21200 25900 21500
rect 23300 21000 23900 21200
rect 25100 21000 25900 21200
rect 23400 20700 24000 21000
rect 24800 20700 25900 21000
rect 28000 24600 29200 24900
rect 29800 24600 30100 24900
rect 31700 24600 32900 24900
rect 33500 24600 33800 24900
rect 34800 24600 35400 24900
rect 28000 24400 28900 24600
rect 31700 24400 32600 24600
rect 34900 24400 35400 24600
rect 37000 24600 37600 24900
rect 37000 24400 37400 24600
rect 28000 24100 28800 24400
rect 31700 24100 32500 24400
rect 34900 24100 35500 24400
rect 28000 23800 28700 24100
rect 31700 23800 32400 24100
rect 35000 23800 35500 24100
rect 36800 24100 37400 24400
rect 36800 23800 37300 24100
rect 28000 23600 28600 23800
rect 31700 23600 32300 23800
rect 35000 23600 35600 23800
rect 28000 20700 28300 23600
rect 31700 20700 32000 23600
rect 35200 23300 35600 23600
rect 36700 23600 37300 23800
rect 36700 23300 37200 23600
rect 35200 23100 35800 23300
rect 35300 22800 35800 23100
rect 36600 23100 37200 23300
rect 36600 22800 37100 23100
rect 35300 22500 35900 22800
rect 35400 22300 35900 22500
rect 36500 22500 37100 22800
rect 36500 22300 37000 22500
rect 35400 22000 36000 22300
rect 35500 21800 36000 22000
rect 36400 22000 37000 22300
rect 36400 21800 36800 22000
rect 35500 21500 36100 21800
rect 35600 21200 36100 21500
rect 36260 21500 36800 21800
rect 36260 21200 36700 21500
rect 35600 21000 36700 21200
rect 19400 20400 20800 20700
rect 21400 20400 22700 20700
rect 23400 20400 26400 20700
rect 19400 19900 20900 20400
rect 21400 19900 22800 20400
rect 23500 20200 26400 20400
rect 23600 19900 25300 20200
rect 25460 19900 26400 20200
rect 27100 19900 29600 20700
rect 30800 19900 33400 20700
rect 35800 20400 36600 21000
rect 42200 20700 42700 24940
rect 43000 24900 43600 25100
rect 43100 24600 43600 24900
rect 43100 24400 43700 24600
rect 43200 23800 43800 24400
rect 43300 23600 43900 23800
rect 43400 23300 43900 23600
rect 43400 23100 44000 23300
rect 43600 22500 44200 23100
rect 43700 22300 44240 22500
rect 43800 22000 44240 22300
rect 44400 22000 44900 27000
rect 46200 24900 47500 25900
rect 43800 21800 44900 22000
rect 43900 21200 44900 21800
rect 44000 20700 44900 21200
rect 47000 20700 47500 24900
rect 35900 20200 36600 20400
rect 23800 19700 25000 19900
rect 35900 19700 36500 20200
rect 41900 19900 43300 20700
rect 44200 20400 44900 20700
rect 44300 19900 44900 20400
rect 46000 19900 48700 20700
rect 35800 19100 36400 19700
rect 35600 18600 36200 19100
rect 35600 18400 36100 18600
rect 35500 18100 36100 18400
rect 34600 17800 36500 18100
rect 34600 17600 36600 17800
rect 34600 17300 36500 17600
rect 10100 13900 12100 14200
rect 10000 13700 12500 13900
rect 10000 13400 12700 13700
rect 10100 13100 12800 13400
rect 26300 13100 26900 15000
rect 45100 14700 45600 15000
rect 52700 14700 53200 15000
rect 56400 14700 56900 15000
rect 44600 14400 46000 14700
rect 48100 14400 50200 14700
rect 52300 14400 53500 14700
rect 56000 14400 57200 14700
rect 42700 14200 42920 14220
rect 44500 14200 46200 14400
rect 37300 13900 38600 14200
rect 37100 13700 38840 13900
rect 39000 13700 39400 14200
rect 41000 13900 42400 14200
rect 42700 14060 43100 14200
rect 42760 13900 43100 14060
rect 44400 13900 46300 14200
rect 48100 13900 50300 14400
rect 52200 14200 53600 14400
rect 55900 14200 57500 14400
rect 52100 13900 53800 14200
rect 55800 13900 57600 14200
rect 40800 13700 42600 13900
rect 42760 13700 43200 13900
rect 44300 13700 45100 13900
rect 45600 13700 46400 13900
rect 37000 13400 39400 13700
rect 40700 13400 43200 13700
rect 36800 13100 37800 13400
rect 38200 13100 39400 13400
rect 40600 13100 41500 13400
rect 41900 13100 43200 13400
rect 44200 13400 44900 13700
rect 45800 13400 46400 13700
rect 48100 13700 50200 13900
rect 52000 13700 52700 13900
rect 53000 13700 53900 13900
rect 55800 13700 56500 13900
rect 56900 13700 57700 13900
rect 44200 13100 44800 13400
rect 46000 13100 46600 13400
rect 10600 10300 10900 13100
rect 12100 12900 12800 13100
rect 36700 12900 37400 13100
rect 38500 12900 39400 13100
rect 12200 12600 13000 12900
rect 12500 12400 13000 12600
rect 36600 12600 37300 12900
rect 38600 12600 39400 12900
rect 40400 12900 41300 13100
rect 42200 12900 43200 13100
rect 40400 12600 41000 12900
rect 42500 12600 43200 12900
rect 36600 12400 37200 12600
rect 38800 12400 39400 12600
rect 40300 12400 40900 12600
rect 12500 12100 13100 12400
rect 15000 12100 15800 12400
rect 18800 12100 19600 12400
rect 22700 12100 23500 12400
rect 30200 12100 31000 12400
rect 12600 11600 13100 12100
rect 14600 11800 16200 12100
rect 18500 11800 19900 12100
rect 20060 11800 20400 12100
rect 14400 11600 16300 11800
rect 18200 11600 20400 11800
rect 12500 11300 13100 11600
rect 14300 11300 16600 11600
rect 18100 11300 20400 11600
rect 21100 11600 22100 12100
rect 22300 11800 23800 12100
rect 22260 11600 24000 11800
rect 21100 11300 24100 11600
rect 25600 11300 26900 12100
rect 12500 11100 13000 11300
rect 12400 10800 13000 11100
rect 14200 11100 15100 11300
rect 15700 11100 16700 11300
rect 14200 10800 14900 11100
rect 16000 10800 16700 11100
rect 18000 11100 18800 11300
rect 19600 11100 20400 11300
rect 21200 11100 22800 11300
rect 23400 11100 24200 11300
rect 25700 11100 26900 11300
rect 28900 11800 29600 12100
rect 29900 11800 31200 12100
rect 36500 11800 37100 12400
rect 38900 11800 39400 12400
rect 28900 11300 31400 11800
rect 36400 11600 37000 11800
rect 39000 11600 39400 11800
rect 40200 11800 40800 12400
rect 42600 12100 43200 12600
rect 44000 12900 44600 13100
rect 44000 12400 44500 12900
rect 44200 12100 44400 12400
rect 28900 11100 30200 11300
rect 30800 11100 31600 11300
rect 18000 10800 18600 11100
rect 19800 10800 20400 11100
rect 12100 10500 13000 10800
rect 11500 10300 12800 10500
rect 14000 10300 14600 10800
rect 16200 10300 16800 10800
rect 18000 10300 18500 10800
rect 19900 10300 20400 10800
rect 10600 10000 12700 10300
rect 13900 10000 14500 10300
rect 16300 10000 16900 10300
rect 18000 10000 18600 10300
rect 20000 10000 20400 10300
rect 21600 10800 22600 11100
rect 23600 10800 24400 11100
rect 21600 10500 22400 10800
rect 23800 10500 24400 10800
rect 21600 10300 22300 10500
rect 23900 10300 24500 10500
rect 21600 10000 22200 10300
rect 10600 9800 12500 10000
rect 13900 9800 14400 10000
rect 16400 9800 16900 10000
rect 10600 9500 12400 9800
rect 10600 6900 10900 9500
rect 11600 9200 12500 9500
rect 11900 9000 12600 9200
rect 12000 8700 12700 9000
rect 13900 8700 16900 9800
rect 18100 9800 19000 10000
rect 18100 9500 19800 9800
rect 18200 9200 20000 9500
rect 18500 9000 20300 9200
rect 19100 8700 20400 9000
rect 12100 8400 12800 8700
rect 12200 8200 12800 8400
rect 13900 8200 14400 8700
rect 19700 8400 20500 8700
rect 19900 8200 20500 8400
rect 12400 7900 13000 8200
rect 13900 7900 14500 8200
rect 17900 7900 18200 8200
rect 12500 7400 13100 7900
rect 14000 7400 14600 7900
rect 16600 7400 16800 7700
rect 17900 7400 18400 7900
rect 20000 7400 20500 8200
rect 12600 6900 13200 7400
rect 14200 7100 14900 7400
rect 16400 7100 16900 7400
rect 14200 6900 15000 7100
rect 16100 6900 16900 7100
rect 10100 6600 11500 6900
rect 12700 6600 13600 6900
rect 14300 6600 16900 6900
rect 17900 7100 18500 7400
rect 19900 7100 20500 7400
rect 17900 6900 18600 7100
rect 19800 6900 20500 7100
rect 21600 8400 22100 10000
rect 24000 9500 24500 10300
rect 24100 9200 24500 9500
rect 24100 9000 24600 9200
rect 21600 8200 22200 8400
rect 24000 8200 24500 9000
rect 21600 7700 22300 8200
rect 23900 7900 24500 8200
rect 23800 7700 24400 7900
rect 21600 7400 22600 7700
rect 23600 7400 24400 7700
rect 21600 7100 22700 7400
rect 23400 7100 24200 7400
rect 21600 6900 24100 7100
rect 26500 6900 26900 11100
rect 29300 10800 30100 11100
rect 31000 10800 31600 11100
rect 29300 10500 30000 10800
rect 31100 10500 31700 10800
rect 29300 10300 29900 10500
rect 29300 6900 29800 10300
rect 31200 6900 31700 10500
rect 32800 9500 35600 10500
rect 36400 8700 36800 11600
rect 39100 11300 39260 11600
rect 40200 11300 40700 11800
rect 42700 11600 43200 12100
rect 46100 11600 46600 13100
rect 42800 11300 43100 11600
rect 46000 11300 46600 11600
rect 48100 11600 48600 13700
rect 51800 13400 52600 13700
rect 53300 13400 53900 13700
rect 55700 13400 56300 13700
rect 57100 13400 57700 13700
rect 51800 13100 52400 13400
rect 53400 13100 54000 13400
rect 55700 13100 56200 13400
rect 57200 13100 57800 13400
rect 51700 12600 52300 13100
rect 53500 12900 54000 13100
rect 55600 12900 56200 13100
rect 57400 12900 57800 13100
rect 51700 12100 52200 12600
rect 53500 12400 54100 12900
rect 51600 11800 52200 12100
rect 48800 11600 49700 11800
rect 48100 11300 49900 11600
rect 40100 8700 40600 11300
rect 45800 11100 46400 11300
rect 45700 10800 46400 11100
rect 48100 11100 50000 11300
rect 48100 10800 50200 11100
rect 45600 10500 46300 10800
rect 48100 10500 48800 10800
rect 49600 10500 50300 10800
rect 45500 10300 46200 10500
rect 48100 10300 48600 10500
rect 49700 10300 50400 10500
rect 45400 10000 46100 10300
rect 49800 10000 50400 10300
rect 45200 9800 46000 10000
rect 49900 9800 50400 10000
rect 45100 9500 45800 9800
rect 50000 9500 50400 9800
rect 45000 9200 45700 9500
rect 44900 9000 45600 9200
rect 44800 8700 45500 9000
rect 36400 8400 37000 8700
rect 36500 8200 37000 8400
rect 40200 8200 40700 8700
rect 44600 8400 45400 8700
rect 44500 8200 45200 8400
rect 50000 8200 50500 9500
rect 51600 8700 52100 11800
rect 53600 11600 54100 12400
rect 53800 9500 54100 11600
rect 55600 11100 56000 12900
rect 57400 12600 58000 12900
rect 57500 11800 58000 12600
rect 57500 11600 58100 11800
rect 57400 11100 58100 11600
rect 55600 10800 56200 11100
rect 57200 10800 58100 11100
rect 55700 10500 56300 10800
rect 57100 10500 58100 10800
rect 55700 10300 56400 10500
rect 57000 10300 58100 10500
rect 55800 10000 58100 10300
rect 55800 9800 57500 10000
rect 56000 9500 57400 9800
rect 57660 9640 58100 10000
rect 36500 7900 37100 8200
rect 39100 7900 39500 8200
rect 40200 7900 40800 8200
rect 43000 7900 43200 8200
rect 44400 7900 45100 8200
rect 36500 7700 37200 7900
rect 39000 7700 39500 7900
rect 36600 7400 37200 7700
rect 38900 7400 39500 7700
rect 40300 7700 40900 7900
rect 42700 7700 43200 7900
rect 44300 7700 45000 7900
rect 49900 7700 50400 8200
rect 51700 7900 52200 8700
rect 53600 8200 54100 9500
rect 56200 9200 57100 9500
rect 57600 9200 58100 9640
rect 57500 9000 58100 9200
rect 57500 8400 58000 9000
rect 57400 8200 58000 8400
rect 51700 7700 52300 7900
rect 53500 7700 54100 8200
rect 57200 7900 57800 8200
rect 57100 7700 57800 7900
rect 40300 7400 41000 7700
rect 42600 7400 43200 7700
rect 44200 7400 44900 7700
rect 47800 7400 48200 7700
rect 49800 7400 50400 7700
rect 51800 7400 52300 7700
rect 36700 7100 37400 7400
rect 38800 7100 39500 7400
rect 40400 7100 41200 7400
rect 42500 7100 43200 7400
rect 44000 7100 44800 7400
rect 46200 7100 46600 7400
rect 47800 7100 48500 7400
rect 49700 7100 50300 7400
rect 51800 7100 52400 7400
rect 53400 7100 54000 7700
rect 57000 7400 57700 7700
rect 56900 7100 57600 7400
rect 36800 6900 37600 7100
rect 38500 6900 39400 7100
rect 40600 6900 41400 7100
rect 42400 6900 43100 7100
rect 43900 6900 44600 7100
rect 46200 6900 46700 7100
rect 47800 6900 48600 7100
rect 49400 6900 50300 7100
rect 52000 6900 52600 7100
rect 53300 6900 53900 7100
rect 56600 6900 57600 7100
rect 17900 6600 19200 6900
rect 19360 6600 20400 6900
rect 10000 6400 11600 6600
rect 10100 6100 11600 6400
rect 12800 6100 13700 6600
rect 14400 6400 16800 6600
rect 17900 6400 20300 6600
rect 21600 6440 22040 6900
rect 22200 6600 24000 6900
rect 14600 6100 16600 6400
rect 17900 6100 20200 6400
rect 14900 5800 16200 6100
rect 18600 5800 19900 6100
rect 21600 4300 22100 6440
rect 22300 6400 23900 6600
rect 22600 6100 23500 6400
rect 25300 6100 28100 6900
rect 28800 6100 30100 6900
rect 30800 6100 32000 6900
rect 37000 6600 38000 6900
rect 38200 6600 39200 6900
rect 40700 6600 41800 6900
rect 41960 6600 43000 6900
rect 37100 6400 39100 6600
rect 40800 6400 42800 6600
rect 37200 6100 38900 6400
rect 40900 6100 42700 6400
rect 43900 6100 46700 6900
rect 47900 6600 50200 6900
rect 52000 6600 53800 6900
rect 48000 6400 50000 6600
rect 52100 6400 53800 6600
rect 55600 6600 57400 6900
rect 55600 6400 57200 6600
rect 48200 6100 49900 6400
rect 52200 6100 53500 6400
rect 55600 6100 57000 6400
rect 37400 5800 38600 6100
rect 41200 5800 42500 6100
rect 48500 5800 49700 6100
rect 52400 5800 53400 6100
rect 55700 5800 56800 6100
rect 21100 3500 22800 4300
<< properties >>
string GDS_END 2458154
string GDS_FILE /home/hni/TopmetalSe-Respin/mag/text.gds
string GDS_START 102
<< end >>
