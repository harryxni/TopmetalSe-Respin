magic
tech sky130A
timestamp 1758224170
<< metal5 >>
rect 18800 56200 21000 56400
rect 22700 56200 23000 56400
rect 51100 56200 51600 56400
rect 18400 55900 21500 56200
rect 22600 55900 23200 56200
rect 23900 55900 30700 56200
rect 18000 55700 21800 55900
rect 22400 55700 23200 55900
rect 23800 55700 30700 55900
rect 31700 55900 34100 56200
rect 31700 55700 34200 55900
rect 17800 55400 23200 55700
rect 23900 55400 30800 55700
rect 31700 55400 34300 55700
rect 37600 55400 40542 56200
rect 41491 55900 45600 56200
rect 41491 55700 46100 55900
rect 51100 55700 51700 56200
rect 41491 55400 46600 55700
rect 17500 55100 23200 55400
rect 24500 55100 30800 55400
rect 32300 55100 34400 55400
rect 38200 55100 40300 55400
rect 41500 55100 46800 55400
rect 51000 55100 51800 55700
rect 17400 54900 19300 55100
rect 20800 54900 23200 55100
rect 24700 54900 30800 55100
rect 32500 54900 34600 55100
rect 17200 54600 19100 54900
rect 21100 54600 23200 54900
rect 17000 54400 18700 54600
rect 21400 54400 23200 54600
rect 24800 54400 26400 54900
rect 29400 54600 30800 54900
rect 32600 54600 34600 54900
rect 38500 54900 40000 55100
rect 41900 54900 46900 55100
rect 38500 54600 39800 54900
rect 29900 54400 30800 54600
rect 32800 54400 34700 54600
rect 16900 54100 18600 54400
rect 21600 54100 23200 54400
rect 16800 53800 18400 54100
rect 21700 53800 23200 54100
rect 16700 53600 18200 53800
rect 21800 53600 23200 53800
rect 16600 53300 18100 53600
rect 22000 53300 23200 53600
rect 16400 53100 18000 53300
rect 22100 53100 23200 53300
rect 16300 52800 17900 53100
rect 16200 52500 17900 52800
rect 22200 52500 23200 53100
rect 16200 52300 17800 52500
rect 22300 52300 23200 52500
rect 16100 52000 17600 52300
rect 16000 51800 17600 52000
rect 22400 51800 23200 52300
rect 16000 51500 17500 51800
rect 15800 51000 17400 51500
rect 22600 51200 23200 51800
rect 15700 50700 17400 51000
rect 15700 50200 17300 50700
rect 22700 50400 23300 51200
rect 15600 49900 17300 50200
rect 22800 50200 23300 50400
rect 22800 49900 23200 50200
rect 15600 49400 17200 49900
rect 6400 48160 6600 49300
rect 6340 48000 6600 48160
rect 15500 48400 17200 49400
rect 6200 47200 6500 48000
rect 15500 47600 17000 48400
rect 6100 46560 6400 47200
rect 7800 46900 8400 47200
rect 7600 46857 8400 46900
rect 7600 46700 8500 46857
rect 6040 46400 6400 46560
rect 7400 46400 7800 46700
rect 6100 45400 6260 46400
rect 7200 46100 7700 46400
rect 7100 45900 7400 46100
rect 7000 45760 7300 45900
rect 8300 45760 8500 46700
rect 15400 46000 17000 47600
rect 6940 45600 7300 45760
rect 8240 45600 8500 45760
rect 6700 45400 7100 45600
rect 6100 45100 7000 45400
rect 6200 44800 6700 45100
rect 8200 44800 8400 45600
rect 8000 44600 8400 44800
rect 15500 45000 17000 46000
rect 25000 48100 26400 54400
rect 30000 54100 30800 54400
rect 30100 53300 30800 54100
rect 30200 52800 30800 53300
rect 30400 52000 30800 52800
rect 32900 54100 34800 54400
rect 38600 54100 39700 54600
rect 42000 54100 43600 54900
rect 44900 54600 47200 54900
rect 45400 54400 47400 54600
rect 50900 54400 52000 55100
rect 45600 54100 47400 54400
rect 32900 53800 34900 54100
rect 38800 53800 39700 54100
rect 32900 53600 35000 53800
rect 32900 53100 35200 53600
rect 32900 52800 35300 53100
rect 32900 52500 35400 52800
rect 32900 52300 35500 52500
rect 32900 52000 35600 52300
rect 32900 51640 33540 52000
rect 33700 51800 35600 52000
rect 29600 49900 30100 50700
rect 29500 49100 30100 49900
rect 32900 49400 33600 51640
rect 33800 51500 35800 51800
rect 34000 51200 35900 51500
rect 34100 51000 36000 51200
rect 34100 50700 36100 51000
rect 34200 50400 36100 50700
rect 34300 50200 36200 50400
rect 34400 49900 36400 50200
rect 34600 49700 36500 49900
rect 29400 48600 30100 49100
rect 29300 48400 30100 48600
rect 29200 48100 30100 48400
rect 25000 46800 30100 48100
rect 8000 44100 8300 44600
rect 9700 44300 10100 44600
rect 9500 44100 10300 44300
rect 15500 44200 17200 45000
rect 7900 43800 8300 44100
rect 9400 43800 10400 44100
rect 7900 42500 8200 43800
rect 9100 43500 9800 43800
rect 10000 43500 10400 43800
rect 9000 43300 9600 43500
rect 8900 43000 9400 43300
rect 10100 43000 10400 43500
rect 15600 43700 17200 44200
rect 15600 43400 17300 43700
rect 8600 42800 9200 43000
rect 8500 42500 9100 42800
rect 10000 42500 10400 43000
rect 15700 42900 17300 43400
rect 15700 42600 17400 42900
rect 7900 42200 8900 42500
rect 8000 42000 8600 42200
rect 10000 42000 10300 42500
rect 15800 42400 17400 42600
rect 15800 42100 17500 42400
rect 8200 41700 8400 42000
rect 9800 41400 10200 42000
rect 16000 41800 17500 42100
rect 11400 41400 12100 41700
rect 16000 41600 17600 41800
rect 9700 40700 10200 41400
rect 11300 41200 12200 41400
rect 16100 41300 17800 41600
rect 11000 40900 12200 41200
rect 16200 41100 17800 41300
rect 22900 41100 23300 41300
rect 10900 40700 12400 40900
rect 16200 40800 17900 41100
rect 22800 40800 23400 41100
rect 9700 39900 10100 40700
rect 10800 40400 11500 40700
rect 10600 40100 11400 40400
rect 11900 40100 12400 40700
rect 16300 40500 18000 40800
rect 22700 40500 23400 40800
rect 16400 40300 18100 40500
rect 22600 40300 23300 40500
rect 10400 39900 11200 40100
rect 11800 39900 12400 40100
rect 16600 40000 18200 40300
rect 22300 40000 23200 40300
rect 9700 39600 11000 39900
rect 9700 39400 10800 39600
rect 11800 39400 12200 39900
rect 16600 39800 18400 40000
rect 22200 39800 23000 40000
rect 16700 39500 18600 39800
rect 22000 39500 22900 39800
rect 9700 39100 10700 39400
rect 10000 38800 10400 39100
rect 11600 38800 12200 39400
rect 16800 39200 18700 39500
rect 21700 39200 22800 39500
rect 25000 39200 26400 46800
rect 28700 46500 30100 46800
rect 29200 46300 30100 46500
rect 29300 46000 30100 46300
rect 29400 45500 30100 46000
rect 29500 44700 30100 45500
rect 29600 44200 30100 44700
rect 29600 43900 30000 44200
rect 31100 42400 31400 42600
rect 31000 42100 31400 42400
rect 30800 41600 31400 42100
rect 30700 41300 31400 41600
rect 30700 41100 31300 41300
rect 33000 41100 33600 49400
rect 34700 49100 36600 49700
rect 34800 48900 36700 49100
rect 34900 48600 36800 48900
rect 35000 48400 37000 48600
rect 35200 48100 37000 48400
rect 35200 47800 37100 48100
rect 35300 47600 37200 47800
rect 35400 47300 37300 47600
rect 35500 47100 37400 47300
rect 35600 46500 37600 47100
rect 35800 46300 37700 46500
rect 35900 46000 37800 46300
rect 36000 45800 37900 46000
rect 36100 45200 38000 45800
rect 36200 45000 38200 45200
rect 36400 44700 38300 45000
rect 36500 44400 38300 44700
rect 36600 44200 38400 44400
rect 38800 44200 39600 53800
rect 42100 47800 43600 54100
rect 45700 53800 47500 54100
rect 50800 53800 52100 54400
rect 45800 53600 47600 53800
rect 46000 53300 47800 53600
rect 50600 53300 52200 53800
rect 46100 53100 47800 53300
rect 46200 52300 47900 53100
rect 50500 52500 52300 53300
rect 46300 49700 48000 52300
rect 50400 52000 52400 52500
rect 50300 51500 50940 52000
rect 51100 51500 52600 52000
rect 50300 51200 50900 51500
rect 50200 51000 50900 51200
rect 51200 51000 52700 51500
rect 50200 50700 50800 51000
rect 50000 50200 50800 50700
rect 51400 50700 52700 51000
rect 51400 50200 52800 50700
rect 49900 49700 50600 50200
rect 51500 49700 52900 50200
rect 46300 49400 47900 49700
rect 46200 48900 47900 49400
rect 49800 49400 50600 49700
rect 49800 48900 50500 49400
rect 51600 49100 53000 49700
rect 51600 48900 53200 49100
rect 46100 48400 47800 48900
rect 49700 48400 50400 48900
rect 51700 48400 53200 48900
rect 46000 48100 47600 48400
rect 49600 48100 50400 48400
rect 45800 47800 47500 48100
rect 42100 47100 43400 47800
rect 45700 47600 47400 47800
rect 49600 47600 50300 48100
rect 51800 47800 53300 48400
rect 45500 47300 47300 47600
rect 45100 47100 47200 47300
rect 49400 47100 50200 47600
rect 52000 47300 53400 47800
rect 52000 47100 53500 47300
rect 42100 46800 43900 47100
rect 44200 46800 46900 47100
rect 49300 46800 50200 47100
rect 52100 46800 53500 47100
rect 42100 46500 46700 46800
rect 49300 46500 50000 46800
rect 52100 46500 53600 46800
rect 42100 46300 46600 46500
rect 49200 46300 50000 46500
rect 42100 46000 46200 46300
rect 42100 45800 45700 46000
rect 49200 45800 49900 46300
rect 52200 46000 53600 46500
rect 42100 45500 43600 45800
rect 42100 45000 43400 45500
rect 49100 45200 49800 45800
rect 52300 45500 53800 46000
rect 52300 45200 53900 45500
rect 49000 45000 49800 45200
rect 52400 45000 53900 45200
rect 36600 43900 38500 44200
rect 36700 43700 38500 43900
rect 36800 43400 38600 43700
rect 38800 43400 39500 44200
rect 37000 43100 39500 43400
rect 37100 42900 39500 43100
rect 37200 42400 39500 42900
rect 37300 42100 39500 42400
rect 37400 41800 39500 42100
rect 37600 41300 39500 41800
rect 37700 41100 39500 41300
rect 30600 40800 31300 41100
rect 30500 40500 31300 40800
rect 30500 40300 31200 40500
rect 30400 40000 31200 40300
rect 30200 39800 31200 40000
rect 30000 39500 31200 39800
rect 32900 39500 33700 41100
rect 37800 40800 39500 41100
rect 37900 40500 39500 40800
rect 38000 40300 39500 40500
rect 38200 39800 39500 40300
rect 42100 39800 43600 45000
rect 49000 44700 54000 45000
rect 48800 44400 54000 44700
rect 48800 43900 54100 44400
rect 48700 43700 54100 43900
rect 48700 43400 49400 43700
rect 48600 42900 49400 43400
rect 52700 43100 54200 43700
rect 48500 42100 49300 42900
rect 52800 42600 54400 43100
rect 52900 42400 54400 42600
rect 48400 41600 49200 42100
rect 52900 41800 54500 42400
rect 48200 41300 49200 41600
rect 53000 41300 54600 41800
rect 48200 41100 49100 41300
rect 48100 40800 49100 41100
rect 53200 40800 54700 41300
rect 48100 40500 49000 40800
rect 48000 40300 49000 40500
rect 48000 40000 48800 40300
rect 53300 40000 54800 40800
rect 38300 39500 39500 39800
rect 29800 39200 31100 39500
rect 13400 38800 13900 39100
rect 17000 39000 19000 39200
rect 21500 39000 22700 39200
rect 24800 39000 26500 39200
rect 29300 39000 31100 39200
rect 32800 39000 33800 39500
rect 38400 39200 39500 39500
rect 38500 39000 39500 39200
rect 42000 39200 43600 39800
rect 47900 39500 48800 40000
rect 42000 39000 43700 39200
rect 47800 39000 48800 39500
rect 11600 38600 12100 38800
rect 13200 38600 14000 38800
rect 17200 38700 19400 39000
rect 21000 38700 22400 39000
rect 24700 38700 31100 39000
rect 32600 38700 34000 39000
rect 11500 38100 12100 38600
rect 13000 38300 14200 38600
rect 17300 38400 22300 38700
rect 24600 38400 31000 38700
rect 32400 38400 34200 38700
rect 38600 38400 39500 39000
rect 41900 38700 43700 39000
rect 47600 38700 48800 39000
rect 53400 39500 55000 40000
rect 53400 39200 55100 39500
rect 53400 38700 55200 39200
rect 41800 38400 43900 38700
rect 47400 38400 49000 38700
rect 53300 38400 55400 38700
rect 12800 38100 14200 38300
rect 17500 38200 22100 38400
rect 23900 38200 31000 38400
rect 31800 38200 34800 38400
rect 38800 38200 39500 38400
rect 11500 37500 12000 38100
rect 12700 37800 14300 38100
rect 17800 37900 21800 38200
rect 23800 37900 31000 38200
rect 12500 37500 13400 37800
rect 11400 37460 12000 37500
rect 11400 37000 11940 37460
rect 12400 37300 13300 37500
rect 13700 37300 14300 37800
rect 18000 37700 21600 37900
rect 23900 37700 31000 37900
rect 31700 37700 34800 38200
rect 38900 37900 39500 38200
rect 39000 37700 39500 37900
rect 41000 38200 44600 38400
rect 47000 38200 49600 38400
rect 52600 38200 55800 38400
rect 41000 37700 44800 38200
rect 46900 37700 49700 38200
rect 52600 37700 55900 38200
rect 18400 37400 21200 37700
rect 12100 37000 13100 37300
rect 13600 37000 14300 37300
rect 19000 37100 20800 37400
rect 39100 37100 39500 37700
rect 11400 36800 13000 37000
rect 11500 36500 12800 36800
rect 13600 36500 14200 37000
rect 11500 36200 12600 36500
rect 13400 36200 14200 36500
rect 11600 36000 12400 36200
rect 13400 35700 14000 36200
rect 13300 35200 14000 35700
rect 57500 36000 57700 36200
rect 57500 35700 58000 36000
rect 57500 35400 58300 35700
rect 57600 35200 58600 35400
rect 13300 34400 13900 35200
rect 57600 34900 58800 35200
rect 57700 34700 59200 34900
rect 57700 34400 59400 34700
rect 13300 34100 59600 34400
rect 13300 33900 59900 34100
rect 13200 33600 59800 33900
rect 13000 33400 59500 33600
rect 12800 33100 13700 33400
rect 57700 33100 59200 33400
rect 12700 32800 13600 33100
rect 57600 32800 58900 33100
rect 12600 32600 13400 32800
rect 57600 32600 58600 32800
rect 12400 32300 13200 32600
rect 57500 32300 58300 32600
rect 12200 32100 13100 32300
rect 57500 32100 58100 32300
rect 12100 31800 13000 32100
rect 57500 31800 57700 32100
rect 11900 31500 12800 31800
rect 11800 31300 12600 31500
rect 11600 31000 12500 31300
rect 11500 30800 12400 31000
rect 11300 30500 12100 30800
rect 11200 30200 12000 30500
rect 11000 30000 11900 30200
rect 10900 29700 11800 30000
rect 10700 29400 11500 29700
rect 10600 29200 11400 29400
rect 10400 28900 11300 29200
rect 10200 28700 11200 28900
rect 10100 28400 10900 28700
rect 10000 28100 10800 28400
rect 9800 27900 10700 28100
rect 9600 27600 10400 27900
rect 9500 27400 10300 27600
rect 9400 27100 10200 27400
rect 9200 26800 10100 27100
rect 9100 26600 10000 26800
rect 8900 26300 9700 26600
rect 8800 26100 9600 26300
rect 8600 25800 9500 26100
rect 8500 25500 9200 25800
rect 8300 25300 9100 25500
rect 8200 25000 9000 25300
rect 8000 24800 8900 25000
rect 7800 24500 8600 24800
rect 7700 24200 8500 24500
rect 7600 24000 8400 24200
rect 7400 23700 8200 24000
rect 7200 23400 8000 23700
rect 7100 23200 7900 23400
rect 7000 22900 7800 23200
rect 6700 22700 7600 22900
rect 6600 22400 7400 22700
rect 6500 22100 7300 22400
rect 6400 21900 7200 22100
rect 6100 21600 7000 21900
rect 6000 21400 6800 21600
rect 5900 21100 6700 21400
rect 5600 20800 6500 21100
rect 5500 20600 6400 20800
rect 4100 20100 4300 20600
rect 5400 20300 6200 20600
rect 5300 20100 6100 20300
rect 4000 19500 4300 20100
rect 5000 19800 5900 20100
rect 4900 19500 5800 19800
rect 3800 19000 4400 19500
rect 4800 19300 5600 19500
rect 4700 19000 5500 19300
rect 3700 18800 5300 19000
rect 3600 18500 5200 18800
rect 3600 18200 5000 18500
rect 3500 18000 4800 18200
rect 3500 17700 4900 18000
rect 3400 17400 5000 17700
rect 3400 17200 5300 17400
rect 3200 16900 5400 17200
rect 3200 16700 5300 16900
rect 3100 16400 4900 16700
rect 3000 16100 4400 16400
rect 3000 15900 4000 16100
rect 2900 15600 3600 15900
rect 2900 15400 3100 15600
<< end >>
