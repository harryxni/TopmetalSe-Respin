** sch_path: /home/hni/TopmetalSe-Respin/xschem/array100.sch
**.subckt array100 VDD GND SF_IB CSA_VREF VREF GRING ARRAY_OUT
*+ ROW_SEL[0],ROW_SEL[1],ROW_SEL[2],ROW_SEL[3],ROW_SEL[4],ROW_SEL[5],ROW_SEL[6],ROW_SEL[7],ROW_SEL[8],ROW_SEL[9],ROW_SEL[10],ROW_SEL[11],ROW_SEL[12],ROW_SEL[13],ROW_SEL[14],ROW_SEL[15],ROW_SEL[16],ROW_SEL[17],ROW_SEL[18],ROW_SEL[19],ROW_SEL[20],ROW_SEL[21],ROW_SEL[22],ROW_SEL[23],ROW_SEL[24],ROW_SEL[25],ROW_SEL[26],ROW_SEL[27],ROW_SEL[28],ROW_SEL[29],ROW_SEL[30],ROW_SEL[31],ROW_SEL[32],ROW_SEL[33],ROW_SEL[34],ROW_SEL[35],ROW_SEL[36],ROW_SEL[37],ROW_SEL[38],ROW_SEL[39],ROW_SEL[40],ROW_SEL[41],ROW_SEL[42],ROW_SEL[43],ROW_SEL[44],ROW_SEL[45],ROW_SEL[46],ROW_SEL[47],ROW_SEL[48],ROW_SEL[49],ROW_SEL[50],ROW_SEL[51],ROW_SEL[52],ROW_SEL[53],ROW_SEL[54],ROW_SEL[55],ROW_SEL[56],ROW_SEL[57],ROW_SEL[58],ROW_SEL[59],ROW_SEL[60],ROW_SEL[61],ROW_SEL[62],ROW_SEL[63],ROW_SEL[64],ROW_SEL[65],ROW_SEL[66],ROW_SEL[67],ROW_SEL[68],ROW_SEL[69],ROW_SEL[70],ROW_SEL[71],ROW_SEL[72],ROW_SEL[73],ROW_SEL[74],ROW_SEL[75],ROW_SEL[76],ROW_SEL[77],ROW_SEL[78],ROW_SEL[79],ROW_SEL[80],ROW_SEL[81],ROW_SEL[82],ROW_SEL[83],ROW_SEL[84],ROW_SEL[85],ROW_SEL[86],ROW_SEL[87],ROW_SEL[88],ROW_SEL[89],ROW_SEL[90],ROW_SEL[91],ROW_SEL[92],ROW_SEL[93],ROW_SEL[94],ROW_SEL[95],ROW_SEL[96],ROW_SEL[97],ROW_SEL[98],ROW_SEL[99] VBIAS IN NB1 NB2
*+ COL_SEL[0],COL_SEL[1],COL_SEL[2],COL_SEL[3],COL_SEL[4],COL_SEL[5],COL_SEL[6],COL_SEL[7],COL_SEL[8],COL_SEL[9],COL_SEL[10],COL_SEL[11],COL_SEL[12],COL_SEL[13],COL_SEL[14],COL_SEL[15],COL_SEL[16],COL_SEL[17],COL_SEL[18],COL_SEL[19],COL_SEL[20],COL_SEL[21],COL_SEL[22],COL_SEL[23],COL_SEL[24],COL_SEL[25],COL_SEL[26],COL_SEL[27],COL_SEL[28],COL_SEL[29],COL_SEL[30],COL_SEL[31],COL_SEL[32],COL_SEL[33],COL_SEL[34],COL_SEL[35],COL_SEL[36],COL_SEL[37],COL_SEL[38],COL_SEL[39],COL_SEL[40],COL_SEL[41],COL_SEL[42],COL_SEL[43],COL_SEL[44],COL_SEL[45],COL_SEL[46],COL_SEL[47],COL_SEL[48],COL_SEL[49],COL_SEL[50],COL_SEL[51],COL_SEL[52],COL_SEL[53],COL_SEL[54],COL_SEL[55],COL_SEL[56],COL_SEL[57],COL_SEL[58],COL_SEL[59],COL_SEL[60],COL_SEL[61],COL_SEL[62],COL_SEL[63],COL_SEL[64],COL_SEL[65],COL_SEL[66],COL_SEL[67],COL_SEL[68],COL_SEL[69],COL_SEL[70],COL_SEL[71],COL_SEL[72],COL_SEL[73],COL_SEL[74],COL_SEL[75],COL_SEL[76],COL_SEL[77],COL_SEL[78],COL_SEL[79],COL_SEL[80],COL_SEL[81],COL_SEL[82],COL_SEL[83],COL_SEL[84],COL_SEL[85],COL_SEL[86],COL_SEL[87],COL_SEL[88],COL_SEL[89],COL_SEL[90],COL_SEL[91],COL_SEL[92],COL_SEL[93],COL_SEL[94],COL_SEL[95],COL_SEL[96],COL_SEL[97],COL_SEL[98],COL_SEL[99]
*.ipin VDD
*.ipin GND
*.ipin SF_IB
*.ipin CSA_VREF
*.ipin VREF
*.ipin GRING
*.opin ARRAY_OUT
*.ipin
*+ ROW_SEL[0],ROW_SEL[1],ROW_SEL[2],ROW_SEL[3],ROW_SEL[4],ROW_SEL[5],ROW_SEL[6],ROW_SEL[7],ROW_SEL[8],ROW_SEL[9],ROW_SEL[10],ROW_SEL[11],ROW_SEL[12],ROW_SEL[13],ROW_SEL[14],ROW_SEL[15],ROW_SEL[16],ROW_SEL[17],ROW_SEL[18],ROW_SEL[19],ROW_SEL[20],ROW_SEL[21],ROW_SEL[22],ROW_SEL[23],ROW_SEL[24],ROW_SEL[25],ROW_SEL[26],ROW_SEL[27],ROW_SEL[28],ROW_SEL[29],ROW_SEL[30],ROW_SEL[31],ROW_SEL[32],ROW_SEL[33],ROW_SEL[34],ROW_SEL[35],ROW_SEL[36],ROW_SEL[37],ROW_SEL[38],ROW_SEL[39],ROW_SEL[40],ROW_SEL[41],ROW_SEL[42],ROW_SEL[43],ROW_SEL[44],ROW_SEL[45],ROW_SEL[46],ROW_SEL[47],ROW_SEL[48],ROW_SEL[49],ROW_SEL[50],ROW_SEL[51],ROW_SEL[52],ROW_SEL[53],ROW_SEL[54],ROW_SEL[55],ROW_SEL[56],ROW_SEL[57],ROW_SEL[58],ROW_SEL[59],ROW_SEL[60],ROW_SEL[61],ROW_SEL[62],ROW_SEL[63],ROW_SEL[64],ROW_SEL[65],ROW_SEL[66],ROW_SEL[67],ROW_SEL[68],ROW_SEL[69],ROW_SEL[70],ROW_SEL[71],ROW_SEL[72],ROW_SEL[73],ROW_SEL[74],ROW_SEL[75],ROW_SEL[76],ROW_SEL[77],ROW_SEL[78],ROW_SEL[79],ROW_SEL[80],ROW_SEL[81],ROW_SEL[82],ROW_SEL[83],ROW_SEL[84],ROW_SEL[85],ROW_SEL[86],ROW_SEL[87],ROW_SEL[88],ROW_SEL[89],ROW_SEL[90],ROW_SEL[91],ROW_SEL[92],ROW_SEL[93],ROW_SEL[94],ROW_SEL[95],ROW_SEL[96],ROW_SEL[97],ROW_SEL[98],ROW_SEL[99]
*.ipin VBIAS
*.ipin IN
*.ipin NB1
*.ipin NB2
*.ipin
*+ COL_SEL[0],COL_SEL[1],COL_SEL[2],COL_SEL[3],COL_SEL[4],COL_SEL[5],COL_SEL[6],COL_SEL[7],COL_SEL[8],COL_SEL[9],COL_SEL[10],COL_SEL[11],COL_SEL[12],COL_SEL[13],COL_SEL[14],COL_SEL[15],COL_SEL[16],COL_SEL[17],COL_SEL[18],COL_SEL[19],COL_SEL[20],COL_SEL[21],COL_SEL[22],COL_SEL[23],COL_SEL[24],COL_SEL[25],COL_SEL[26],COL_SEL[27],COL_SEL[28],COL_SEL[29],COL_SEL[30],COL_SEL[31],COL_SEL[32],COL_SEL[33],COL_SEL[34],COL_SEL[35],COL_SEL[36],COL_SEL[37],COL_SEL[38],COL_SEL[39],COL_SEL[40],COL_SEL[41],COL_SEL[42],COL_SEL[43],COL_SEL[44],COL_SEL[45],COL_SEL[46],COL_SEL[47],COL_SEL[48],COL_SEL[49],COL_SEL[50],COL_SEL[51],COL_SEL[52],COL_SEL[53],COL_SEL[54],COL_SEL[55],COL_SEL[56],COL_SEL[57],COL_SEL[58],COL_SEL[59],COL_SEL[60],COL_SEL[61],COL_SEL[62],COL_SEL[63],COL_SEL[64],COL_SEL[65],COL_SEL[66],COL_SEL[67],COL_SEL[68],COL_SEL[69],COL_SEL[70],COL_SEL[71],COL_SEL[72],COL_SEL[73],COL_SEL[74],COL_SEL[75],COL_SEL[76],COL_SEL[77],COL_SEL[78],COL_SEL[79],COL_SEL[80],COL_SEL[81],COL_SEL[82],COL_SEL[83],COL_SEL[84],COL_SEL[85],COL_SEL[86],COL_SEL[87],COL_SEL[88],COL_SEL[89],COL_SEL[90],COL_SEL[91],COL_SEL[92],COL_SEL[93],COL_SEL[94],COL_SEL[95],COL_SEL[96],COL_SEL[97],COL_SEL[98],COL_SEL[99]
xPix0 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix1 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix2 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix3 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix4 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix5 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix6 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix7 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix8 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix9 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix10 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix11 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix12 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix13 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix14 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix15 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix16 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix17 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix18 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix19 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix20 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix21 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix22 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix23 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix24 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix25 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix26 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix27 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix28 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix29 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix30 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix31 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix32 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix33 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix34 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix35 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix36 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix37 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix38 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix39 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix40 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix41 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix42 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix43 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix44 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix45 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix46 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix47 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix48 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix49 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix50 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix51 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix52 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix53 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix54 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix55 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix56 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix57 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix58 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix59 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix60 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix61 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix62 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix63 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix64 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix65 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix66 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix67 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix68 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix69 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix70 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix71 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix72 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix73 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix74 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix75 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix76 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix77 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix78 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix79 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix80 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix81 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix82 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix83 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix84 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix85 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix86 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix87 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix88 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix89 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix90 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix91 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix92 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix93 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix94 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix95 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix96 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix97 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix98 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix99 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[0] VBIAS IN NB1 NB2 pixel
xPix100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[1] VBIAS IN NB1 NB2 pixel
xPix200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[2] VBIAS IN NB1 NB2 pixel
xPix300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[3] VBIAS IN NB1 NB2 pixel
xPix400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[4] VBIAS IN NB1 NB2 pixel
xPix500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[5] VBIAS IN NB1 NB2 pixel
xPix600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[6] VBIAS IN NB1 NB2 pixel
xPix700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[7] VBIAS IN NB1 NB2 pixel
xPix800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[8] VBIAS IN NB1 NB2 pixel
xPix900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[9] VBIAS IN NB1 NB2 pixel
xPix1000 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1001 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1002 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1003 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1004 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1005 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1006 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1007 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1008 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1009 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1010 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1011 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1012 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1013 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1014 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1015 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1016 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1017 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1018 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1019 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1020 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1021 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1022 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1023 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1024 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1025 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1026 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1027 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1028 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1029 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1030 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1031 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1032 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1033 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1034 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1035 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1036 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1037 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1038 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1039 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1040 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1041 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1042 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1043 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1044 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1045 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1046 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1047 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1048 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1049 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1050 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1051 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1052 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1053 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1054 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1055 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1056 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1057 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1058 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1059 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1060 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1061 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1062 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1063 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1064 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1065 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1066 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1067 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1068 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1069 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1070 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1071 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1072 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1073 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1074 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1075 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1076 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1077 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1078 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1079 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1080 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1081 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1082 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1083 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1084 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1085 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1086 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1087 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1088 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1089 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1090 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1091 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1092 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1093 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1094 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1095 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1096 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1097 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1098 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1099 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[10] VBIAS IN NB1 NB2 pixel
xPix1100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[11] VBIAS IN NB1 NB2 pixel
xPix1200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[12] VBIAS IN NB1 NB2 pixel
xPix1300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[13] VBIAS IN NB1 NB2 pixel
xPix1400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[14] VBIAS IN NB1 NB2 pixel
xPix1500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[15] VBIAS IN NB1 NB2 pixel
xPix1600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[16] VBIAS IN NB1 NB2 pixel
xPix1700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[17] VBIAS IN NB1 NB2 pixel
xPix1800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[18] VBIAS IN NB1 NB2 pixel
xPix1900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix1999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[19] VBIAS IN NB1 NB2 pixel
xPix2000 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2001 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2002 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2003 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2004 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2005 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2006 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2007 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2008 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2009 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2010 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2011 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2012 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2013 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2014 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2015 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2016 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2017 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2018 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2019 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2020 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2021 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2022 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2023 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2024 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2025 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2026 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2027 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2028 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2029 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2030 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2031 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2032 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2033 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2034 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2035 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2036 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2037 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2038 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2039 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2040 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2041 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2042 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2043 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2044 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2045 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2046 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2047 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2048 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2049 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2050 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2051 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2052 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2053 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2054 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2055 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2056 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2057 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2058 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2059 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2060 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2061 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2062 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2063 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2064 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2065 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2066 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2067 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2068 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2069 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2070 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2071 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2072 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2073 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2074 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2075 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2076 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2077 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2078 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2079 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2080 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2081 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2082 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2083 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2084 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2085 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2086 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2087 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2088 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2089 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2090 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2091 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2092 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2093 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2094 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2095 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2096 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2097 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2098 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2099 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[20] VBIAS IN NB1 NB2 pixel
xPix2100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[21] VBIAS IN NB1 NB2 pixel
xPix2200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[22] VBIAS IN NB1 NB2 pixel
xPix2300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[23] VBIAS IN NB1 NB2 pixel
xPix2400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[24] VBIAS IN NB1 NB2 pixel
xPix2500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[25] VBIAS IN NB1 NB2 pixel
xPix2600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[26] VBIAS IN NB1 NB2 pixel
xPix2700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[27] VBIAS IN NB1 NB2 pixel
xPix2800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[28] VBIAS IN NB1 NB2 pixel
xPix2900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix2999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[29] VBIAS IN NB1 NB2 pixel
xPix3000 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3001 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3002 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3003 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3004 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3005 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3006 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3007 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3008 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3009 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3010 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3011 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3012 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3013 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3014 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3015 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3016 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3017 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3018 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3019 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3020 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3021 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3022 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3023 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3024 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3025 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3026 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3027 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3028 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3029 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3030 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3031 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3032 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3033 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3034 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3035 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3036 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3037 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3038 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3039 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3040 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3041 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3042 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3043 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3044 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3045 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3046 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3047 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3048 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3049 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3050 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3051 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3052 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3053 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3054 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3055 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3056 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3057 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3058 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3059 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3060 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3061 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3062 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3063 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3064 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3065 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3066 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3067 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3068 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3069 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3070 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3071 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3072 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3073 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3074 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3075 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3076 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3077 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3078 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3079 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3080 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3081 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3082 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3083 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3084 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3085 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3086 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3087 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3088 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3089 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3090 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3091 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3092 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3093 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3094 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3095 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3096 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3097 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3098 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3099 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[30] VBIAS IN NB1 NB2 pixel
xPix3100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[31] VBIAS IN NB1 NB2 pixel
xPix3200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[32] VBIAS IN NB1 NB2 pixel
xPix3300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[33] VBIAS IN NB1 NB2 pixel
xPix3400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[34] VBIAS IN NB1 NB2 pixel
xPix3500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[35] VBIAS IN NB1 NB2 pixel
xPix3600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[36] VBIAS IN NB1 NB2 pixel
xPix3700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[37] VBIAS IN NB1 NB2 pixel
xPix3800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[38] VBIAS IN NB1 NB2 pixel
xPix3900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix3999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[39] VBIAS IN NB1 NB2 pixel
xPix4000 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4001 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4002 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4003 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4004 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4005 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4006 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4007 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4008 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4009 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4010 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4011 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4012 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4013 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4014 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4015 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4016 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4017 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4018 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4019 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4020 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4021 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4022 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4023 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4024 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4025 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4026 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4027 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4028 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4029 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4030 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4031 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4032 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4033 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4034 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4035 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4036 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4037 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4038 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4039 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4040 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4041 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4042 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4043 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4044 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4045 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4046 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4047 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4048 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4049 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4050 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4051 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4052 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4053 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4054 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4055 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4056 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4057 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4058 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4059 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4060 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4061 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4062 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4063 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4064 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4065 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4066 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4067 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4068 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4069 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4070 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4071 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4072 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4073 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4074 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4075 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4076 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4077 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4078 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4079 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4080 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4081 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4082 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4083 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4084 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4085 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4086 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4087 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4088 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4089 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4090 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4091 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4092 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4093 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4094 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4095 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4096 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4097 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4098 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4099 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[40] VBIAS IN NB1 NB2 pixel
xPix4100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[41] VBIAS IN NB1 NB2 pixel
xPix4200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[42] VBIAS IN NB1 NB2 pixel
xPix4300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[43] VBIAS IN NB1 NB2 pixel
xPix4400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[44] VBIAS IN NB1 NB2 pixel
xPix4500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[45] VBIAS IN NB1 NB2 pixel
xPix4600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[46] VBIAS IN NB1 NB2 pixel
xPix4700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[47] VBIAS IN NB1 NB2 pixel
xPix4800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[48] VBIAS IN NB1 NB2 pixel
xPix4900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix4999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[49] VBIAS IN NB1 NB2 pixel
xPix5000 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5001 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5002 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5003 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5004 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5005 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5006 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5007 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5008 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5009 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5010 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5011 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5012 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5013 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5014 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5015 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5016 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5017 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5018 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5019 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5020 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5021 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5022 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5023 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5024 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5025 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5026 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5027 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5028 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5029 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5030 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5031 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5032 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5033 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5034 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5035 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5036 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5037 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5038 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5039 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5040 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5041 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5042 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5043 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5044 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5045 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5046 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5047 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5048 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5049 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5050 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5051 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5052 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5053 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5054 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5055 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5056 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5057 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5058 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5059 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5060 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5061 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5062 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5063 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5064 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5065 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5066 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5067 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5068 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5069 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5070 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5071 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5072 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5073 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5074 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5075 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5076 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5077 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5078 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5079 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5080 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5081 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5082 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5083 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5084 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5085 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5086 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5087 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5088 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5089 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5090 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5091 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5092 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5093 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5094 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5095 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5096 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5097 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5098 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5099 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[50] VBIAS IN NB1 NB2 pixel
xPix5100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[51] VBIAS IN NB1 NB2 pixel
xPix5200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[52] VBIAS IN NB1 NB2 pixel
xPix5300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[53] VBIAS IN NB1 NB2 pixel
xPix5400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[54] VBIAS IN NB1 NB2 pixel
xPix5500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[55] VBIAS IN NB1 NB2 pixel
xPix5600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[56] VBIAS IN NB1 NB2 pixel
xPix5700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[57] VBIAS IN NB1 NB2 pixel
xPix5800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[58] VBIAS IN NB1 NB2 pixel
xPix5900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix5999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[59] VBIAS IN NB1 NB2 pixel
xPix6000 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6001 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6002 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6003 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6004 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6005 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6006 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6007 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6008 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6009 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6010 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6011 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6012 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6013 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6014 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6015 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6016 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6017 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6018 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6019 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6020 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6021 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6022 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6023 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6024 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6025 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6026 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6027 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6028 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6029 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6030 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6031 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6032 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6033 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6034 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6035 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6036 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6037 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6038 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6039 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6040 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6041 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6042 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6043 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6044 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6045 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6046 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6047 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6048 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6049 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6050 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6051 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6052 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6053 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6054 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6055 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6056 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6057 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6058 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6059 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6060 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6061 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6062 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6063 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6064 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6065 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6066 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6067 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6068 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6069 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6070 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6071 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6072 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6073 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6074 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6075 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6076 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6077 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6078 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6079 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6080 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6081 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6082 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6083 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6084 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6085 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6086 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6087 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6088 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6089 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6090 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6091 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6092 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6093 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6094 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6095 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6096 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6097 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6098 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6099 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[60] VBIAS IN NB1 NB2 pixel
xPix6100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[61] VBIAS IN NB1 NB2 pixel
xPix6200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[62] VBIAS IN NB1 NB2 pixel
xPix6300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[63] VBIAS IN NB1 NB2 pixel
xPix6400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[64] VBIAS IN NB1 NB2 pixel
xPix6500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[65] VBIAS IN NB1 NB2 pixel
xPix6600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[66] VBIAS IN NB1 NB2 pixel
xPix6700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[67] VBIAS IN NB1 NB2 pixel
xPix6800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[68] VBIAS IN NB1 NB2 pixel
xPix6900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix6999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[69] VBIAS IN NB1 NB2 pixel
xPix7000 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7001 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7002 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7003 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7004 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7005 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7006 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7007 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7008 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7009 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7010 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7011 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7012 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7013 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7014 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7015 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7016 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7017 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7018 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7019 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7020 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7021 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7022 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7023 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7024 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7025 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7026 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7027 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7028 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7029 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7030 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7031 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7032 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7033 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7034 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7035 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7036 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7037 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7038 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7039 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7040 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7041 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7042 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7043 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7044 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7045 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7046 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7047 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7048 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7049 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7050 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7051 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7052 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7053 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7054 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7055 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7056 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7057 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7058 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7059 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7060 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7061 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7062 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7063 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7064 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7065 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7066 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7067 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7068 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7069 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7070 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7071 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7072 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7073 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7074 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7075 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7076 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7077 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7078 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7079 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7080 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7081 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7082 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7083 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7084 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7085 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7086 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7087 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7088 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7089 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7090 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7091 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7092 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7093 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7094 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7095 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7096 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7097 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7098 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7099 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[70] VBIAS IN NB1 NB2 pixel
xPix7100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[71] VBIAS IN NB1 NB2 pixel
xPix7200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[72] VBIAS IN NB1 NB2 pixel
xPix7300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[73] VBIAS IN NB1 NB2 pixel
xPix7400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[74] VBIAS IN NB1 NB2 pixel
xPix7500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[75] VBIAS IN NB1 NB2 pixel
xPix7600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[76] VBIAS IN NB1 NB2 pixel
xPix7700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[77] VBIAS IN NB1 NB2 pixel
xPix7800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[78] VBIAS IN NB1 NB2 pixel
xPix7900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix7999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[79] VBIAS IN NB1 NB2 pixel
xPix8000 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8001 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8002 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8003 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8004 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8005 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8006 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8007 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8008 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8009 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8010 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8011 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8012 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8013 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8014 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8015 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8016 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8017 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8018 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8019 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8020 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8021 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8022 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8023 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8024 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8025 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8026 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8027 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8028 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8029 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8030 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8031 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8032 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8033 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8034 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8035 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8036 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8037 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8038 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8039 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8040 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8041 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8042 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8043 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8044 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8045 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8046 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8047 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8048 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8049 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8050 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8051 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8052 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8053 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8054 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8055 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8056 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8057 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8058 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8059 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8060 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8061 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8062 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8063 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8064 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8065 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8066 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8067 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8068 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8069 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8070 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8071 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8072 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8073 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8074 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8075 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8076 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8077 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8078 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8079 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8080 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8081 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8082 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8083 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8084 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8085 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8086 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8087 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8088 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8089 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8090 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8091 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8092 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8093 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8094 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8095 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8096 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8097 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8098 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8099 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[80] VBIAS IN NB1 NB2 pixel
xPix8100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[81] VBIAS IN NB1 NB2 pixel
xPix8200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[82] VBIAS IN NB1 NB2 pixel
xPix8300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[83] VBIAS IN NB1 NB2 pixel
xPix8400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[84] VBIAS IN NB1 NB2 pixel
xPix8500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[85] VBIAS IN NB1 NB2 pixel
xPix8600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[86] VBIAS IN NB1 NB2 pixel
xPix8700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[87] VBIAS IN NB1 NB2 pixel
xPix8800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[88] VBIAS IN NB1 NB2 pixel
xPix8900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix8999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[89] VBIAS IN NB1 NB2 pixel
xPix9000 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9001 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9002 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9003 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9004 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9005 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9006 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9007 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9008 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9009 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9010 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9011 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9012 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9013 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9014 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9015 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9016 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9017 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9018 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9019 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9020 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9021 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9022 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9023 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9024 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9025 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9026 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9027 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9028 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9029 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9030 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9031 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9032 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9033 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9034 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9035 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9036 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9037 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9038 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9039 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9040 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9041 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9042 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9043 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9044 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9045 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9046 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9047 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9048 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9049 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9050 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9051 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9052 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9053 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9054 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9055 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9056 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9057 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9058 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9059 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9060 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9061 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9062 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9063 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9064 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9065 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9066 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9067 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9068 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9069 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9070 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9071 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9072 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9073 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9074 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9075 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9076 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9077 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9078 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9079 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9080 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9081 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9082 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9083 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9084 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9085 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9086 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9087 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9088 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9089 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9090 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9091 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9092 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9093 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9094 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9095 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9096 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9097 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9098 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9099 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[90] VBIAS IN NB1 NB2 pixel
xPix9100 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9101 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9102 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9103 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9104 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9105 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9106 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9107 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9108 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9109 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9110 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9111 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9112 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9113 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9114 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9115 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9116 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9117 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9118 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9119 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9120 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9121 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9122 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9123 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9124 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9125 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9126 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9127 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9128 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9129 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9130 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9131 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9132 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9133 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9134 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9135 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9136 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9137 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9138 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9139 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9140 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9141 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9142 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9143 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9144 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9145 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9146 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9147 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9148 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9149 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9150 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9151 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9152 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9153 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9154 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9155 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9156 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9157 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9158 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9159 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9160 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9161 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9162 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9163 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9164 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9165 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9166 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9167 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9168 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9169 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9170 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9171 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9172 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9173 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9174 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9175 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9176 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9177 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9178 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9179 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9180 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9181 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9182 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9183 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9184 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9185 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9186 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9187 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9188 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9189 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9190 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9191 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9192 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9193 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9194 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9195 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9196 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9197 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9198 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9199 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[91] VBIAS IN NB1 NB2 pixel
xPix9200 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9201 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9202 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9203 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9204 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9205 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9206 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9207 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9208 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9209 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9210 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9211 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9212 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9213 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9214 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9215 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9216 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9217 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9218 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9219 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9220 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9221 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9222 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9223 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9224 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9225 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9226 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9227 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9228 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9229 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9230 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9231 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9232 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9233 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9234 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9235 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9236 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9237 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9238 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9239 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9240 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9241 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9242 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9243 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9244 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9245 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9246 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9247 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9248 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9249 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9250 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9251 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9252 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9253 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9254 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9255 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9256 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9257 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9258 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9259 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9260 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9261 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9262 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9263 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9264 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9265 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9266 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9267 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9268 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9269 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9270 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9271 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9272 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9273 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9274 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9275 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9276 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9277 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9278 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9279 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9280 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9281 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9282 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9283 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9284 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9285 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9286 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9287 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9288 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9289 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9290 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9291 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9292 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9293 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9294 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9295 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9296 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9297 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9298 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9299 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[92] VBIAS IN NB1 NB2 pixel
xPix9300 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9301 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9302 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9303 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9304 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9305 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9306 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9307 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9308 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9309 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9310 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9311 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9312 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9313 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9314 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9315 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9316 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9317 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9318 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9319 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9320 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9321 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9322 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9323 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9324 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9325 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9326 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9327 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9328 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9329 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9330 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9331 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9332 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9333 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9334 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9335 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9336 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9337 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9338 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9339 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9340 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9341 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9342 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9343 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9344 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9345 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9346 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9347 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9348 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9349 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9350 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9351 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9352 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9353 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9354 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9355 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9356 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9357 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9358 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9359 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9360 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9361 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9362 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9363 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9364 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9365 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9366 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9367 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9368 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9369 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9370 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9371 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9372 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9373 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9374 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9375 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9376 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9377 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9378 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9379 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9380 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9381 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9382 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9383 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9384 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9385 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9386 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9387 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9388 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9389 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9390 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9391 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9392 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9393 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9394 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9395 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9396 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9397 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9398 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9399 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[93] VBIAS IN NB1 NB2 pixel
xPix9400 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9401 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9402 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9403 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9404 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9405 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9406 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9407 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9408 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9409 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9410 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9411 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9412 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9413 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9414 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9415 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9416 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9417 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9418 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9419 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9420 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9421 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9422 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9423 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9424 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9425 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9426 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9427 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9428 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9429 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9430 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9431 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9432 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9433 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9434 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9435 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9436 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9437 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9438 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9439 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9440 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9441 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9442 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9443 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9444 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9445 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9446 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9447 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9448 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9449 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9450 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9451 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9452 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9453 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9454 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9455 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9456 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9457 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9458 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9459 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9460 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9461 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9462 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9463 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9464 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9465 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9466 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9467 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9468 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9469 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9470 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9471 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9472 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9473 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9474 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9475 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9476 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9477 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9478 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9479 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9480 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9481 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9482 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9483 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9484 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9485 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9486 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9487 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9488 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9489 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9490 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9491 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9492 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9493 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9494 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9495 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9496 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9497 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9498 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9499 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[94] VBIAS IN NB1 NB2 pixel
xPix9500 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9501 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9502 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9503 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9504 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9505 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9506 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9507 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9508 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9509 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9510 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9511 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9512 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9513 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9514 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9515 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9516 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9517 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9518 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9519 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9520 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9521 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9522 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9523 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9524 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9525 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9526 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9527 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9528 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9529 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9530 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9531 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9532 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9533 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9534 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9535 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9536 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9537 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9538 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9539 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9540 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9541 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9542 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9543 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9544 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9545 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9546 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9547 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9548 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9549 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9550 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9551 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9552 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9553 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9554 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9555 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9556 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9557 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9558 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9559 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9560 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9561 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9562 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9563 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9564 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9565 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9566 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9567 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9568 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9569 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9570 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9571 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9572 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9573 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9574 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9575 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9576 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9577 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9578 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9579 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9580 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9581 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9582 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9583 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9584 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9585 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9586 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9587 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9588 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9589 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9590 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9591 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9592 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9593 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9594 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9595 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9596 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9597 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9598 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9599 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[95] VBIAS IN NB1 NB2 pixel
xPix9600 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9601 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9602 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9603 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9604 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9605 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9606 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9607 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9608 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9609 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9610 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9611 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9612 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9613 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9614 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9615 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9616 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9617 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9618 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9619 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9620 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9621 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9622 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9623 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9624 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9625 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9626 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9627 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9628 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9629 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9630 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9631 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9632 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9633 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9634 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9635 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9636 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9637 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9638 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9639 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9640 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9641 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9642 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9643 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9644 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9645 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9646 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9647 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9648 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9649 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9650 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9651 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9652 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9653 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9654 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9655 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9656 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9657 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9658 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9659 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9660 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9661 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9662 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9663 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9664 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9665 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9666 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9667 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9668 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9669 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9670 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9671 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9672 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9673 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9674 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9675 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9676 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9677 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9678 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9679 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9680 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9681 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9682 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9683 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9684 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9685 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9686 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9687 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9688 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9689 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9690 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9691 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9692 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9693 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9694 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9695 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9696 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9697 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9698 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9699 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[96] VBIAS IN NB1 NB2 pixel
xPix9700 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9701 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9702 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9703 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9704 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9705 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9706 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9707 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9708 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9709 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9710 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9711 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9712 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9713 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9714 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9715 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9716 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9717 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9718 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9719 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9720 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9721 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9722 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9723 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9724 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9725 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9726 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9727 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9728 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9729 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9730 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9731 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9732 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9733 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9734 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9735 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9736 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9737 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9738 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9739 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9740 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9741 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9742 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9743 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9744 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9745 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9746 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9747 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9748 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9749 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9750 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9751 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9752 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9753 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9754 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9755 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9756 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9757 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9758 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9759 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9760 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9761 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9762 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9763 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9764 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9765 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9766 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9767 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9768 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9769 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9770 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9771 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9772 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9773 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9774 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9775 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9776 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9777 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9778 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9779 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9780 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9781 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9782 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9783 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9784 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9785 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9786 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9787 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9788 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9789 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9790 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9791 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9792 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9793 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9794 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9795 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9796 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9797 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9798 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9799 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[97] VBIAS IN NB1 NB2 pixel
xPix9800 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9801 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9802 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9803 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9804 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9805 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9806 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9807 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9808 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9809 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9810 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9811 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9812 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9813 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9814 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9815 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9816 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9817 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9818 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9819 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9820 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9821 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9822 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9823 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9824 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9825 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9826 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9827 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9828 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9829 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9830 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9831 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9832 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9833 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9834 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9835 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9836 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9837 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9838 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9839 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9840 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9841 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9842 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9843 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9844 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9845 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9846 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9847 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9848 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9849 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9850 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9851 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9852 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9853 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9854 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9855 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9856 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9857 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9858 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9859 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9860 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9861 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9862 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9863 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9864 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9865 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9866 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9867 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9868 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9869 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9870 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9871 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9872 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9873 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9874 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9875 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9876 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9877 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9878 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9879 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9880 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9881 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9882 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9883 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9884 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9885 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9886 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9887 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9888 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9889 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9890 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9891 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9892 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9893 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9894 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9895 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9896 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9897 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9898 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9899 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[98] VBIAS IN NB1 NB2 pixel
xPix9900 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[0] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9901 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[1] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9902 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[2] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9903 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[3] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9904 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[4] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9905 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[5] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9906 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[6] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9907 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[7] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9908 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[8] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9909 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[9] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9910 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[10] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9911 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[11] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9912 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[12] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9913 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[13] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9914 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[14] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9915 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[15] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9916 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[16] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9917 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[17] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9918 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[18] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9919 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[19] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9920 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[20] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9921 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[21] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9922 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[22] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9923 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[23] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9924 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[24] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9925 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[25] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9926 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[26] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9927 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[27] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9928 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[28] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9929 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[29] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9930 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[30] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9931 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[31] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9932 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[32] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9933 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[33] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9934 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[34] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9935 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[35] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9936 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[36] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9937 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[37] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9938 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[38] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9939 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[39] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9940 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[40] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9941 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[41] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9942 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[42] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9943 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[43] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9944 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[44] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9945 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[45] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9946 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[46] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9947 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[47] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9948 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[48] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9949 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[49] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9950 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[50] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9951 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[51] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9952 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[52] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9953 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[53] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9954 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[54] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9955 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[55] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9956 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[56] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9957 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[57] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9958 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[58] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9959 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[59] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9960 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[60] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9961 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[61] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9962 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[62] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9963 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[63] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9964 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[64] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9965 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[65] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9966 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[66] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9967 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[67] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9968 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[68] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9969 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[69] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9970 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[70] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9971 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[71] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9972 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[72] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9973 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[73] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9974 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[74] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9975 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[75] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9976 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[76] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9977 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[77] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9978 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[78] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9979 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[79] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9980 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[80] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9981 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[81] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9982 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[82] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9983 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[83] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9984 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[84] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9985 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[85] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9986 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[86] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9987 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[87] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9988 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[88] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9989 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[89] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9990 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[90] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9991 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[91] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9992 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[92] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9993 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[93] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9994 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[94] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9995 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[95] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9996 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[96] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9997 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[97] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9998 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[98] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
xPix9999 VDD GND SF_IB CSA_VREF VREF GRING COL_OUT[99] ROW_SEL[99] VBIAS IN NB1 NB2 pixel
XM0 COL_OUT[0] COL_SEL[0] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 COL_OUT[1] COL_SEL[1] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 COL_OUT[2] COL_SEL[2] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 COL_OUT[3] COL_SEL[3] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 COL_OUT[4] COL_SEL[4] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 COL_OUT[5] COL_SEL[5] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 COL_OUT[6] COL_SEL[6] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 COL_OUT[7] COL_SEL[7] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 COL_OUT[8] COL_SEL[8] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 COL_OUT[9] COL_SEL[9] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 COL_OUT[10] COL_SEL[10] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 COL_OUT[11] COL_SEL[11] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 COL_OUT[12] COL_SEL[12] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 COL_OUT[13] COL_SEL[13] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 COL_OUT[14] COL_SEL[14] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 COL_OUT[15] COL_SEL[15] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 COL_OUT[16] COL_SEL[16] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 COL_OUT[17] COL_SEL[17] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 COL_OUT[18] COL_SEL[18] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM19 COL_OUT[19] COL_SEL[19] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20 COL_OUT[20] COL_SEL[20] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21 COL_OUT[21] COL_SEL[21] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM22 COL_OUT[22] COL_SEL[22] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23 COL_OUT[23] COL_SEL[23] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 COL_OUT[24] COL_SEL[24] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM25 COL_OUT[25] COL_SEL[25] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM26 COL_OUT[26] COL_SEL[26] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM27 COL_OUT[27] COL_SEL[27] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM28 COL_OUT[28] COL_SEL[28] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM29 COL_OUT[29] COL_SEL[29] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM30 COL_OUT[30] COL_SEL[30] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM31 COL_OUT[31] COL_SEL[31] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM32 COL_OUT[32] COL_SEL[32] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM33 COL_OUT[33] COL_SEL[33] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM34 COL_OUT[34] COL_SEL[34] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM35 COL_OUT[35] COL_SEL[35] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM36 COL_OUT[36] COL_SEL[36] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM37 COL_OUT[37] COL_SEL[37] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM38 COL_OUT[38] COL_SEL[38] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM39 COL_OUT[39] COL_SEL[39] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM40 COL_OUT[40] COL_SEL[40] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM41 COL_OUT[41] COL_SEL[41] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM42 COL_OUT[42] COL_SEL[42] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM43 COL_OUT[43] COL_SEL[43] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM44 COL_OUT[44] COL_SEL[44] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM45 COL_OUT[45] COL_SEL[45] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM46 COL_OUT[46] COL_SEL[46] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM47 COL_OUT[47] COL_SEL[47] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM48 COL_OUT[48] COL_SEL[48] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM49 COL_OUT[49] COL_SEL[49] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM50 COL_OUT[50] COL_SEL[50] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM51 COL_OUT[51] COL_SEL[51] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM52 COL_OUT[52] COL_SEL[52] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM53 COL_OUT[53] COL_SEL[53] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM54 COL_OUT[54] COL_SEL[54] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM55 COL_OUT[55] COL_SEL[55] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM56 COL_OUT[56] COL_SEL[56] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM57 COL_OUT[57] COL_SEL[57] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM58 COL_OUT[58] COL_SEL[58] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM59 COL_OUT[59] COL_SEL[59] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM60 COL_OUT[60] COL_SEL[60] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM61 COL_OUT[61] COL_SEL[61] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM62 COL_OUT[62] COL_SEL[62] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM63 COL_OUT[63] COL_SEL[63] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM64 COL_OUT[64] COL_SEL[64] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM65 COL_OUT[65] COL_SEL[65] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM66 COL_OUT[66] COL_SEL[66] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM67 COL_OUT[67] COL_SEL[67] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM68 COL_OUT[68] COL_SEL[68] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM69 COL_OUT[69] COL_SEL[69] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM70 COL_OUT[70] COL_SEL[70] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM71 COL_OUT[71] COL_SEL[71] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM72 COL_OUT[72] COL_SEL[72] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM73 COL_OUT[73] COL_SEL[73] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM74 COL_OUT[74] COL_SEL[74] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM75 COL_OUT[75] COL_SEL[75] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM76 COL_OUT[76] COL_SEL[76] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM77 COL_OUT[77] COL_SEL[77] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM78 COL_OUT[78] COL_SEL[78] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM79 COL_OUT[79] COL_SEL[79] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM80 COL_OUT[80] COL_SEL[80] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM81 COL_OUT[81] COL_SEL[81] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM82 COL_OUT[82] COL_SEL[82] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM83 COL_OUT[83] COL_SEL[83] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM84 COL_OUT[84] COL_SEL[84] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM85 COL_OUT[85] COL_SEL[85] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM86 COL_OUT[86] COL_SEL[86] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM87 COL_OUT[87] COL_SEL[87] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM88 COL_OUT[88] COL_SEL[88] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM89 COL_OUT[89] COL_SEL[89] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM90 COL_OUT[90] COL_SEL[90] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM91 COL_OUT[91] COL_SEL[91] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM92 COL_OUT[92] COL_SEL[92] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM93 COL_OUT[93] COL_SEL[93] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM94 COL_OUT[94] COL_SEL[94] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM95 COL_OUT[95] COL_SEL[95] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM96 COL_OUT[96] COL_SEL[96] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM97 COL_OUT[97] COL_SEL[97] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM98 COL_OUT[98] COL_SEL[98] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM99 COL_OUT[99] COL_SEL[99] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**.ends

* expanding   symbol:  pixel/pixel.sym # of pins=12
** sym_path: /home/hni/TopmetalSe-Respin/xschem/pixel/pixel.sym
** sch_path: /home/hni/TopmetalSe-Respin/xschem/pixel/pixel.sch
.subckt pixel VDD GND SF_IB CSA_VREF VREF GRING pix_out ROW_SEL VBIAS IN NB1 NB2
*.opin pix_out
*.ipin SF_IB
*.ipin ROW_SEL
*.ipin VREF
*.ipin AMP_IN
*.ipin NB1
*.ipin CSA_VREF
*.ipin VBIAS
*.ipin NB2
*.ipin VDD
*.ipin GND
XM2 net2 ROW_SEL pix_out GND sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 GND AMP_OUT net1 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 SF_IB VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 VDD net1 net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 VDD net6 AMP_OUT GND sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net5 net5 net7 VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net8 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net7 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 AMP_OUT NB2 GND GND sky130_fd_pr__nfet_01v8_lvt L=1.2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 net4 NB1 GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC3 AMP_IN AMP_OUT sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=1 m=1
XM4 net3 VREF net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 AMP_IN CSA_VREF AMP_OUT VDD sky130_fd_pr__pfet_01v8_lvt L=7.95 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net6 net5 net8 VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net5 VBIAS net3 GND sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net9 AMP_IN net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 net6 VBIAS net9 GND sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMD_4 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMD_1 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt L=1.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
