magic
tech sky130A
magscale 1 2
timestamp 1758045453
<< error_s >>
rect -12961 322586 -12952 322595
rect -12953 322531 -12952 322586
rect -12944 322577 -12943 322586
rect -13008 322530 -12952 322531
rect -12944 322530 -12943 322539
rect -12961 322521 -12952 322530
rect 299 319928 308 319931
rect -2006 319921 -1806 319922
rect 108 319921 308 319922
rect -2006 319722 -2005 319723
rect 307 319722 308 319921
rect 316 319913 317 319922
rect 316 319722 317 319731
rect 299 319713 308 319716
rect -15137 19998 -15128 20007
rect -15129 19943 -15128 19998
rect -15120 19989 -15119 19998
rect -15184 19942 -15181 19943
rect -15131 19942 -15128 19943
rect -15120 19942 -15119 19951
rect -15137 19933 -15128 19942
rect -14902 19735 -14867 19746
rect -14868 19701 -14867 19712
rect -11057 19538 -11048 19547
rect -11049 19483 -11048 19538
rect -11040 19536 -11039 19538
rect -11104 19482 -11101 19483
rect -11051 19482 -11048 19483
rect -11040 19482 -11039 19484
rect -11057 19473 -11048 19482
rect -5999 17942 -5998 17946
rect -6095 17941 -5994 17942
rect -5999 17755 -5998 17941
rect -6207 17746 -6198 17755
rect -5999 17746 -5989 17755
rect -6198 17737 -6189 17738
rect -6007 17737 -5998 17738
<< metal1 >>
rect 302508 324532 302708 324538
rect 302508 321358 302708 324332
rect 303926 321358 304246 321364
rect 302508 321038 303926 321358
rect 108 319922 308 320310
rect 302508 320098 302708 321038
rect 303926 321032 304246 321038
rect 102 319722 108 319922
rect 308 319722 314 319922
rect 102 319700 314 319722
rect 108 319450 308 319700
rect 303926 318358 304246 318364
rect 302536 318038 303926 318358
rect 303926 318032 304246 318038
rect 108 316922 308 317310
rect 102 316722 108 316922
rect 308 316722 314 316922
rect 102 316700 314 316722
rect 108 316450 308 316700
rect 303926 315358 304246 315364
rect 302536 315038 303926 315358
rect 303926 315032 304246 315038
rect 108 313922 308 314310
rect 102 313722 108 313922
rect 308 313722 314 313922
rect 102 313700 314 313722
rect 108 313450 308 313700
rect 303926 312358 304246 312364
rect 302536 312038 303926 312358
rect 303926 312032 304246 312038
rect 108 310922 308 311310
rect 102 310722 108 310922
rect 308 310722 314 310922
rect 102 310700 314 310722
rect 108 310450 308 310700
rect 303926 309358 304246 309364
rect 302536 309038 303926 309358
rect 303926 309032 304246 309038
rect 108 307922 308 308310
rect 102 307722 108 307922
rect 308 307722 314 307922
rect 102 307700 314 307722
rect 108 307450 308 307700
rect 303926 306358 304246 306364
rect 302536 306038 303926 306358
rect 303926 306032 304246 306038
rect 108 304922 308 305310
rect 102 304722 108 304922
rect 308 304722 314 304922
rect 102 304700 314 304722
rect 108 304450 308 304700
rect 303926 303358 304246 303364
rect 302536 303038 303926 303358
rect 303926 303032 304246 303038
rect 108 301922 308 302310
rect 102 301722 108 301922
rect 308 301722 314 301922
rect 102 301700 314 301722
rect 108 301450 308 301700
rect 303926 300358 304246 300364
rect 302536 300038 303926 300358
rect 303926 300032 304246 300038
rect 108 298922 308 299310
rect 102 298722 108 298922
rect 308 298722 314 298922
rect 102 298700 314 298722
rect 108 298450 308 298700
rect 303926 297358 304246 297364
rect 302536 297038 303926 297358
rect 303926 297032 304246 297038
rect 108 295922 308 296310
rect 102 295722 108 295922
rect 308 295722 314 295922
rect 102 295700 314 295722
rect 108 295450 308 295700
rect 303926 294358 304246 294364
rect 302536 294038 303926 294358
rect 303926 294032 304246 294038
rect 108 292922 308 293310
rect 102 292722 108 292922
rect 308 292722 314 292922
rect 102 292700 314 292722
rect 108 292450 308 292700
rect 303926 291358 304246 291364
rect 302536 291038 303926 291358
rect 303926 291032 304246 291038
rect 108 289922 308 290310
rect 102 289722 108 289922
rect 308 289722 314 289922
rect 102 289700 314 289722
rect 108 289450 308 289700
rect 303926 288358 304246 288364
rect 302536 288038 303926 288358
rect 303926 288032 304246 288038
rect 108 286922 308 287310
rect 102 286722 108 286922
rect 308 286722 314 286922
rect 102 286700 314 286722
rect 108 286450 308 286700
rect 303926 285358 304246 285364
rect 302536 285038 303926 285358
rect 303926 285032 304246 285038
rect 108 283922 308 284310
rect 102 283722 108 283922
rect 308 283722 314 283922
rect 102 283700 314 283722
rect 108 283450 308 283700
rect 303926 282358 304246 282364
rect 302536 282038 303926 282358
rect 303926 282032 304246 282038
rect 108 280922 308 281310
rect 102 280722 108 280922
rect 308 280722 314 280922
rect 102 280700 314 280722
rect 108 280450 308 280700
rect 303926 279358 304246 279364
rect 302536 279038 303926 279358
rect 303926 279032 304246 279038
rect 108 277922 308 278310
rect 102 277722 108 277922
rect 308 277722 314 277922
rect 102 277700 314 277722
rect 108 277450 308 277700
rect 303926 276358 304246 276364
rect 302536 276038 303926 276358
rect 303926 276032 304246 276038
rect 108 274922 308 275310
rect 102 274722 108 274922
rect 308 274722 314 274922
rect 102 274700 314 274722
rect 108 274450 308 274700
rect 303926 273358 304246 273364
rect 302536 273038 303926 273358
rect 303926 273032 304246 273038
rect 108 271922 308 272310
rect 102 271722 108 271922
rect 308 271722 314 271922
rect 102 271700 314 271722
rect 108 271450 308 271700
rect 303926 270358 304246 270364
rect 302536 270038 303926 270358
rect 303926 270032 304246 270038
rect 108 268922 308 269310
rect 102 268722 108 268922
rect 308 268722 314 268922
rect 102 268700 314 268722
rect 108 268450 308 268700
rect 303926 267358 304246 267364
rect 302536 267038 303926 267358
rect 303926 267032 304246 267038
rect 108 265922 308 266310
rect 102 265722 108 265922
rect 308 265722 314 265922
rect 102 265700 314 265722
rect 108 265450 308 265700
rect 303926 264358 304246 264364
rect 302536 264038 303926 264358
rect 303926 264032 304246 264038
rect 108 262922 308 263310
rect 102 262722 108 262922
rect 308 262722 314 262922
rect 102 262700 314 262722
rect 108 262450 308 262700
rect 303926 261358 304246 261364
rect 302536 261038 303926 261358
rect 303926 261032 304246 261038
rect 108 259922 308 260310
rect 102 259722 108 259922
rect 308 259722 314 259922
rect 102 259700 314 259722
rect 108 259450 308 259700
rect 303926 258358 304246 258364
rect 302536 258038 303926 258358
rect 303926 258032 304246 258038
rect 108 256922 308 257310
rect 102 256722 108 256922
rect 308 256722 314 256922
rect 102 256700 314 256722
rect 108 256450 308 256700
rect 303926 255358 304246 255364
rect 302536 255038 303926 255358
rect 303926 255032 304246 255038
rect 108 253922 308 254310
rect 102 253722 108 253922
rect 308 253722 314 253922
rect 102 253700 314 253722
rect 108 253450 308 253700
rect 303926 252358 304246 252364
rect 302536 252038 303926 252358
rect 303926 252032 304246 252038
rect 108 250922 308 251310
rect 102 250722 108 250922
rect 308 250722 314 250922
rect 102 250700 314 250722
rect 108 250450 308 250700
rect 303926 249358 304246 249364
rect 302536 249038 303926 249358
rect 303926 249032 304246 249038
rect 108 247922 308 248310
rect 102 247722 108 247922
rect 308 247722 314 247922
rect 102 247700 314 247722
rect 108 247450 308 247700
rect 303926 246358 304246 246364
rect 302536 246038 303926 246358
rect 303926 246032 304246 246038
rect 108 244922 308 245310
rect 102 244722 108 244922
rect 308 244722 314 244922
rect 102 244700 314 244722
rect 108 244450 308 244700
rect 303926 243358 304246 243364
rect 302536 243038 303926 243358
rect 303926 243032 304246 243038
rect 108 241922 308 242310
rect 102 241722 108 241922
rect 308 241722 314 241922
rect 102 241700 314 241722
rect 108 241450 308 241700
rect 303926 240358 304246 240364
rect 302536 240038 303926 240358
rect 303926 240032 304246 240038
rect 108 238922 308 239310
rect 102 238722 108 238922
rect 308 238722 314 238922
rect 102 238700 314 238722
rect 108 238450 308 238700
rect 303926 237358 304246 237364
rect 302536 237038 303926 237358
rect 303926 237032 304246 237038
rect 108 235922 308 236310
rect 102 235722 108 235922
rect 308 235722 314 235922
rect 102 235700 314 235722
rect 108 235450 308 235700
rect 303926 234358 304246 234364
rect 302536 234038 303926 234358
rect 303926 234032 304246 234038
rect 108 232922 308 233310
rect 102 232722 108 232922
rect 308 232722 314 232922
rect 102 232700 314 232722
rect 108 232450 308 232700
rect 303926 231358 304246 231364
rect 302536 231038 303926 231358
rect 303926 231032 304246 231038
rect 108 229922 308 230310
rect 102 229722 108 229922
rect 308 229722 314 229922
rect 102 229700 314 229722
rect 108 229450 308 229700
rect 303926 228358 304246 228364
rect 302536 228038 303926 228358
rect 303926 228032 304246 228038
rect 108 226922 308 227310
rect 102 226722 108 226922
rect 308 226722 314 226922
rect 102 226700 314 226722
rect 108 226450 308 226700
rect 303926 225358 304246 225364
rect 302536 225038 303926 225358
rect 303926 225032 304246 225038
rect 108 223922 308 224310
rect 102 223722 108 223922
rect 308 223722 314 223922
rect 102 223700 314 223722
rect 108 223450 308 223700
rect 303926 222358 304246 222364
rect 302536 222038 303926 222358
rect 303926 222032 304246 222038
rect 108 220922 308 221310
rect 102 220722 108 220922
rect 308 220722 314 220922
rect 102 220700 314 220722
rect 108 220450 308 220700
rect 303926 219358 304246 219364
rect 302536 219038 303926 219358
rect 303926 219032 304246 219038
rect 108 217922 308 218310
rect 102 217722 108 217922
rect 308 217722 314 217922
rect 102 217700 314 217722
rect 108 217450 308 217700
rect 303926 216358 304246 216364
rect 302536 216038 303926 216358
rect 303926 216032 304246 216038
rect 108 214922 308 215310
rect 102 214722 108 214922
rect 308 214722 314 214922
rect 102 214700 314 214722
rect 108 214450 308 214700
rect 303926 213358 304246 213364
rect 302536 213038 303926 213358
rect 303926 213032 304246 213038
rect 108 211922 308 212310
rect 102 211722 108 211922
rect 308 211722 314 211922
rect 102 211700 314 211722
rect 108 211450 308 211700
rect 303926 210358 304246 210364
rect 302536 210038 303926 210358
rect 303926 210032 304246 210038
rect 108 208922 308 209310
rect 102 208722 108 208922
rect 308 208722 314 208922
rect 102 208700 314 208722
rect 108 208450 308 208700
rect 303926 207358 304246 207364
rect 302536 207038 303926 207358
rect 303926 207032 304246 207038
rect 108 205922 308 206310
rect 102 205722 108 205922
rect 308 205722 314 205922
rect 102 205700 314 205722
rect 108 205450 308 205700
rect 303926 204358 304246 204364
rect 302536 204038 303926 204358
rect 303926 204032 304246 204038
rect 108 202922 308 203310
rect 102 202722 108 202922
rect 308 202722 314 202922
rect 102 202700 314 202722
rect 108 202450 308 202700
rect 303926 201358 304246 201364
rect 302536 201038 303926 201358
rect 303926 201032 304246 201038
rect 108 199922 308 200310
rect 102 199722 108 199922
rect 308 199722 314 199922
rect 102 199700 314 199722
rect 108 199450 308 199700
rect 303926 198358 304246 198364
rect 302536 198038 303926 198358
rect 303926 198032 304246 198038
rect 108 196922 308 197310
rect 102 196722 108 196922
rect 308 196722 314 196922
rect 102 196700 314 196722
rect 108 196450 308 196700
rect 303926 195358 304246 195364
rect 302536 195038 303926 195358
rect 303926 195032 304246 195038
rect 108 193922 308 194310
rect 102 193722 108 193922
rect 308 193722 314 193922
rect 102 193700 314 193722
rect 108 193450 308 193700
rect 303926 192358 304246 192364
rect 302536 192038 303926 192358
rect 303926 192032 304246 192038
rect 108 190922 308 191310
rect 102 190722 108 190922
rect 308 190722 314 190922
rect 102 190700 314 190722
rect 108 190450 308 190700
rect 303926 189358 304246 189364
rect 302536 189038 303926 189358
rect 303926 189032 304246 189038
rect 108 187922 308 188310
rect 102 187722 108 187922
rect 308 187722 314 187922
rect 102 187700 314 187722
rect 108 187450 308 187700
rect 303926 186358 304246 186364
rect 302536 186038 303926 186358
rect 303926 186032 304246 186038
rect 108 184922 308 185310
rect 102 184722 108 184922
rect 308 184722 314 184922
rect 102 184700 314 184722
rect 108 184450 308 184700
rect 303926 183358 304246 183364
rect 302536 183038 303926 183358
rect 303926 183032 304246 183038
rect 108 181922 308 182310
rect 102 181722 108 181922
rect 308 181722 314 181922
rect 102 181700 314 181722
rect 108 181450 308 181700
rect 303926 180358 304246 180364
rect 302536 180038 303926 180358
rect 303926 180032 304246 180038
rect 108 178922 308 179310
rect 102 178722 108 178922
rect 308 178722 314 178922
rect 102 178700 314 178722
rect 108 178450 308 178700
rect 303926 177358 304246 177364
rect 302536 177038 303926 177358
rect 303926 177032 304246 177038
rect 108 175922 308 176310
rect 102 175722 108 175922
rect 308 175722 314 175922
rect 102 175700 314 175722
rect 108 175450 308 175700
rect 303926 174358 304246 174364
rect 302536 174038 303926 174358
rect 303926 174032 304246 174038
rect 108 172922 308 173310
rect 102 172722 108 172922
rect 308 172722 314 172922
rect 102 172700 314 172722
rect 108 172450 308 172700
rect 303926 171358 304246 171364
rect 302536 171038 303926 171358
rect 303926 171032 304246 171038
rect 108 169922 308 170310
rect 102 169722 108 169922
rect 308 169722 314 169922
rect 102 169700 314 169722
rect 108 169450 308 169700
rect 303926 168358 304246 168364
rect 302536 168038 303926 168358
rect 303926 168032 304246 168038
rect 108 166922 308 167310
rect 102 166722 108 166922
rect 308 166722 314 166922
rect 102 166700 314 166722
rect 108 166450 308 166700
rect 303926 165358 304246 165364
rect 302536 165038 303926 165358
rect 303926 165032 304246 165038
rect 108 163922 308 164310
rect 102 163722 108 163922
rect 308 163722 314 163922
rect 102 163700 314 163722
rect 108 163450 308 163700
rect 303926 162358 304246 162364
rect 302536 162038 303926 162358
rect 303926 162032 304246 162038
rect 108 160922 308 161310
rect 102 160722 108 160922
rect 308 160722 314 160922
rect 102 160700 314 160722
rect 108 160450 308 160700
rect 303926 159358 304246 159364
rect 302536 159038 303926 159358
rect 303926 159032 304246 159038
rect 108 157922 308 158310
rect 102 157722 108 157922
rect 308 157722 314 157922
rect 102 157700 314 157722
rect 108 157450 308 157700
rect 303926 156358 304246 156364
rect 302536 156038 303926 156358
rect 303926 156032 304246 156038
rect 108 154922 308 155310
rect 102 154722 108 154922
rect 308 154722 314 154922
rect 102 154700 314 154722
rect 108 154450 308 154700
rect 303926 153358 304246 153364
rect 302536 153038 303926 153358
rect 303926 153032 304246 153038
rect 108 151922 308 152310
rect 102 151722 108 151922
rect 308 151722 314 151922
rect 102 151700 314 151722
rect 108 151450 308 151700
rect 303926 150358 304246 150364
rect 302536 150038 303926 150358
rect 303926 150032 304246 150038
rect 108 148922 308 149310
rect 102 148722 108 148922
rect 308 148722 314 148922
rect 102 148700 314 148722
rect 108 148450 308 148700
rect 303926 147358 304246 147364
rect 302536 147038 303926 147358
rect 303926 147032 304246 147038
rect 108 145922 308 146310
rect 102 145722 108 145922
rect 308 145722 314 145922
rect 102 145700 314 145722
rect 108 145450 308 145700
rect 303926 144358 304246 144364
rect 302536 144038 303926 144358
rect 303926 144032 304246 144038
rect 108 142922 308 143310
rect 102 142722 108 142922
rect 308 142722 314 142922
rect 102 142700 314 142722
rect 108 142450 308 142700
rect 303926 141358 304246 141364
rect 302536 141038 303926 141358
rect 303926 141032 304246 141038
rect 108 139922 308 140310
rect 102 139722 108 139922
rect 308 139722 314 139922
rect 102 139700 314 139722
rect 108 139450 308 139700
rect 303926 138358 304246 138364
rect 302536 138038 303926 138358
rect 303926 138032 304246 138038
rect 108 136922 308 137310
rect 102 136722 108 136922
rect 308 136722 314 136922
rect 102 136700 314 136722
rect 108 136450 308 136700
rect 303926 135358 304246 135364
rect 302536 135038 303926 135358
rect 303926 135032 304246 135038
rect 108 133922 308 134310
rect 102 133722 108 133922
rect 308 133722 314 133922
rect 102 133700 314 133722
rect 108 133450 308 133700
rect 303926 132358 304246 132364
rect 302536 132038 303926 132358
rect 303926 132032 304246 132038
rect 108 130922 308 131310
rect 102 130722 108 130922
rect 308 130722 314 130922
rect 102 130700 314 130722
rect 108 130450 308 130700
rect 303926 129358 304246 129364
rect 302536 129038 303926 129358
rect 303926 129032 304246 129038
rect 108 127922 308 128310
rect 102 127722 108 127922
rect 308 127722 314 127922
rect 102 127700 314 127722
rect 108 127450 308 127700
rect 303926 126358 304246 126364
rect 302536 126038 303926 126358
rect 303926 126032 304246 126038
rect 108 124922 308 125310
rect 102 124722 108 124922
rect 308 124722 314 124922
rect 102 124700 314 124722
rect 108 124450 308 124700
rect 303926 123358 304246 123364
rect 302536 123038 303926 123358
rect 303926 123032 304246 123038
rect 108 121922 308 122310
rect 102 121722 108 121922
rect 308 121722 314 121922
rect 102 121700 314 121722
rect 108 121450 308 121700
rect 303926 120358 304246 120364
rect 302536 120038 303926 120358
rect 303926 120032 304246 120038
rect 108 118922 308 119310
rect 102 118722 108 118922
rect 308 118722 314 118922
rect 102 118700 314 118722
rect 108 118450 308 118700
rect 303926 117358 304246 117364
rect 302536 117038 303926 117358
rect 303926 117032 304246 117038
rect 108 115922 308 116310
rect 102 115722 108 115922
rect 308 115722 314 115922
rect 102 115700 314 115722
rect 108 115450 308 115700
rect 303926 114358 304246 114364
rect 302536 114038 303926 114358
rect 303926 114032 304246 114038
rect 108 112922 308 113310
rect 102 112722 108 112922
rect 308 112722 314 112922
rect 102 112700 314 112722
rect 108 112450 308 112700
rect 303926 111358 304246 111364
rect 302536 111038 303926 111358
rect 303926 111032 304246 111038
rect 108 109922 308 110310
rect 102 109722 108 109922
rect 308 109722 314 109922
rect 102 109700 314 109722
rect 108 109450 308 109700
rect 303926 108358 304246 108364
rect 302536 108038 303926 108358
rect 303926 108032 304246 108038
rect 108 106922 308 107310
rect 102 106722 108 106922
rect 308 106722 314 106922
rect 102 106700 314 106722
rect 108 106450 308 106700
rect 303926 105358 304246 105364
rect 302536 105038 303926 105358
rect 303926 105032 304246 105038
rect 108 103922 308 104310
rect 102 103722 108 103922
rect 308 103722 314 103922
rect 102 103700 314 103722
rect 108 103450 308 103700
rect 303926 102358 304246 102364
rect 302536 102038 303926 102358
rect 303926 102032 304246 102038
rect 108 100922 308 101310
rect 102 100722 108 100922
rect 308 100722 314 100922
rect 102 100700 314 100722
rect 108 100450 308 100700
rect 303926 99358 304246 99364
rect 302536 99038 303926 99358
rect 303926 99032 304246 99038
rect 108 97922 308 98310
rect 102 97722 108 97922
rect 308 97722 314 97922
rect 102 97700 314 97722
rect 108 97450 308 97700
rect 303926 96358 304246 96364
rect 302536 96038 303926 96358
rect 303926 96032 304246 96038
rect 108 94922 308 95310
rect 102 94722 108 94922
rect 308 94722 314 94922
rect 102 94700 314 94722
rect 108 94450 308 94700
rect 303926 93358 304246 93364
rect 302536 93038 303926 93358
rect 303926 93032 304246 93038
rect 108 91922 308 92310
rect 102 91722 108 91922
rect 308 91722 314 91922
rect 102 91700 314 91722
rect 108 91450 308 91700
rect 303926 90358 304246 90364
rect 302536 90038 303926 90358
rect 303926 90032 304246 90038
rect 108 88922 308 89310
rect 102 88722 108 88922
rect 308 88722 314 88922
rect 102 88700 314 88722
rect 108 88450 308 88700
rect 303926 87358 304246 87364
rect 302536 87038 303926 87358
rect 303926 87032 304246 87038
rect 108 85922 308 86310
rect 102 85722 108 85922
rect 308 85722 314 85922
rect 102 85700 314 85722
rect 108 85450 308 85700
rect 303926 84358 304246 84364
rect 302536 84038 303926 84358
rect 303926 84032 304246 84038
rect 108 82922 308 83310
rect 102 82722 108 82922
rect 308 82722 314 82922
rect 102 82700 314 82722
rect 108 82450 308 82700
rect 303926 81358 304246 81364
rect 302536 81038 303926 81358
rect 303926 81032 304246 81038
rect 108 79922 308 80310
rect 102 79722 108 79922
rect 308 79722 314 79922
rect 102 79700 314 79722
rect 108 79450 308 79700
rect 303926 78358 304246 78364
rect 302536 78038 303926 78358
rect 303926 78032 304246 78038
rect 108 76922 308 77310
rect 102 76722 108 76922
rect 308 76722 314 76922
rect 102 76700 314 76722
rect 108 76450 308 76700
rect 303926 75358 304246 75364
rect 302536 75038 303926 75358
rect 303926 75032 304246 75038
rect 108 73922 308 74310
rect 102 73722 108 73922
rect 308 73722 314 73922
rect 102 73700 314 73722
rect 108 73450 308 73700
rect 303926 72358 304246 72364
rect 302536 72038 303926 72358
rect 303926 72032 304246 72038
rect 108 70922 308 71310
rect 102 70722 108 70922
rect 308 70722 314 70922
rect 102 70700 314 70722
rect 108 70450 308 70700
rect 303926 69358 304246 69364
rect 302536 69038 303926 69358
rect 303926 69032 304246 69038
rect 108 67922 308 68310
rect 102 67722 108 67922
rect 308 67722 314 67922
rect 102 67700 314 67722
rect 108 67450 308 67700
rect 303926 66358 304246 66364
rect 302536 66038 303926 66358
rect 303926 66032 304246 66038
rect 108 64922 308 65310
rect 102 64722 108 64922
rect 308 64722 314 64922
rect 102 64700 314 64722
rect 108 64450 308 64700
rect 303926 63358 304246 63364
rect 302536 63038 303926 63358
rect 303926 63032 304246 63038
rect 108 61922 308 62310
rect 102 61722 108 61922
rect 308 61722 314 61922
rect 102 61700 314 61722
rect 108 61450 308 61700
rect 303926 60358 304246 60364
rect 302536 60038 303926 60358
rect 303926 60032 304246 60038
rect 108 58922 308 59310
rect 102 58722 108 58922
rect 308 58722 314 58922
rect 102 58700 314 58722
rect 108 58450 308 58700
rect 303926 57358 304246 57364
rect 302536 57038 303926 57358
rect 303926 57032 304246 57038
rect 108 55922 308 56310
rect 102 55722 108 55922
rect 308 55722 314 55922
rect 102 55700 314 55722
rect 108 55450 308 55700
rect 303926 54358 304246 54364
rect 302536 54038 303926 54358
rect 303926 54032 304246 54038
rect 108 52922 308 53310
rect 102 52722 108 52922
rect 308 52722 314 52922
rect 102 52700 314 52722
rect 108 52450 308 52700
rect 303926 51358 304246 51364
rect 302536 51038 303926 51358
rect 303926 51032 304246 51038
rect 108 49922 308 50310
rect 102 49722 108 49922
rect 308 49722 314 49922
rect 102 49700 314 49722
rect 108 49450 308 49700
rect 303926 48358 304246 48364
rect 302536 48038 303926 48358
rect 303926 48032 304246 48038
rect 108 46922 308 47310
rect 102 46722 108 46922
rect 308 46722 314 46922
rect 102 46700 314 46722
rect 108 46450 308 46700
rect 303926 45358 304246 45364
rect 302536 45038 303926 45358
rect 303926 45032 304246 45038
rect 108 43922 308 44310
rect 102 43722 108 43922
rect 308 43722 314 43922
rect 102 43700 314 43722
rect 108 43450 308 43700
rect 303926 42358 304246 42364
rect 302536 42038 303926 42358
rect 303926 42032 304246 42038
rect 108 40922 308 41310
rect 102 40722 108 40922
rect 308 40722 314 40922
rect 102 40700 314 40722
rect 108 40450 308 40700
rect 303926 39358 304246 39364
rect 302536 39038 303926 39358
rect 303926 39032 304246 39038
rect 108 37922 308 38310
rect 102 37722 108 37922
rect 308 37722 314 37922
rect 102 37700 314 37722
rect 108 37450 308 37700
rect 303926 36358 304246 36364
rect 302536 36038 303926 36358
rect 303926 36032 304246 36038
rect 108 34922 308 35310
rect 102 34722 108 34922
rect 308 34722 314 34922
rect 102 34700 314 34722
rect 108 34450 308 34700
rect 303926 33358 304246 33364
rect 302536 33038 303926 33358
rect 303926 33032 304246 33038
rect 108 31922 308 32310
rect 102 31722 108 31922
rect 308 31722 314 31922
rect 102 31700 314 31722
rect 108 31450 308 31700
rect 303926 30358 304246 30364
rect 302536 30038 303926 30358
rect 303926 30032 304246 30038
rect 108 28922 308 29310
rect 102 28722 108 28922
rect 308 28722 314 28922
rect 102 28700 314 28722
rect 108 28450 308 28700
rect 303926 27358 304246 27364
rect 302536 27038 303926 27358
rect 303926 27032 304246 27038
rect 108 25922 308 26310
rect 102 25722 108 25922
rect 308 25722 314 25922
rect 102 25700 314 25722
rect 108 25450 308 25700
rect 303926 24358 304246 24364
rect 302536 24038 303926 24358
rect 303926 24032 304246 24038
rect 108 22922 308 23310
rect 102 22722 108 22922
rect 308 22722 314 22922
rect 102 22700 314 22722
rect 108 22450 308 22700
rect 303926 21358 304246 21364
rect 302536 21038 303926 21358
rect 303926 21032 304246 21038
rect 108 19900 308 20808
rect 302508 20408 302828 20608
rect 102 19700 314 19900
rect 108 17946 308 19700
rect 3658 18440 3664 18760
rect 3984 18440 3990 18760
rect 18082 18440 18088 18760
rect 18408 18440 18414 18760
rect 32908 18440 32914 18760
rect 33234 18440 33240 18760
rect 64250 18440 64256 18760
rect 64576 18440 64582 18760
rect 121672 18440 121678 18760
rect 121998 18440 122004 18760
rect 167542 18440 167548 18760
rect 167868 18440 167874 18760
rect 180542 18440 180548 18760
rect 180868 18440 180874 18760
rect 189542 18440 189548 18760
rect 189868 18440 189874 18760
rect 198542 18440 198548 18760
rect 198868 18440 198874 18760
rect 204542 18440 204548 18760
rect 204868 18440 204874 18760
rect 211542 18440 211548 18760
rect 211868 18440 211874 18760
rect 223542 18440 223548 18760
rect 223868 18440 223874 18760
rect 232542 18440 232548 18760
rect 232868 18440 232874 18760
rect 238542 18440 238548 18760
rect 238868 18440 238874 18760
rect 250542 18440 250548 18760
rect 250868 18440 250874 18760
rect 263942 18440 263948 18760
rect 264268 18440 264274 18760
rect 269942 18440 269948 18760
rect 270268 18440 270274 18760
rect 272942 18440 272948 18760
rect 273268 18440 273274 18760
rect 275942 18440 275948 18760
rect 276268 18440 276274 18760
rect 281942 18440 281948 18760
rect 282268 18440 282274 18760
rect 285942 18440 285948 18760
rect 286268 18440 286274 18760
rect 293942 18440 293948 18760
rect 294268 18440 294274 18760
rect 296942 18440 296948 18760
rect 297268 18440 297274 18760
rect 299942 18440 299948 18760
rect 300268 18440 300274 18760
rect 302942 18440 302948 18760
rect 303268 18440 303274 18760
rect -6204 17746 -6198 17946
rect -5998 17746 308 17946
rect 3664 17938 3984 18440
rect 18088 17938 18408 18440
rect 32914 17938 33234 18440
rect 64256 17938 64576 18440
rect 121678 17938 121998 18440
rect 167548 17938 167868 18440
rect 180548 17938 180868 18440
rect 189548 17938 189868 18440
rect 198548 17938 198868 18440
rect 204548 17938 204868 18440
rect 211548 17938 211868 18440
rect 223548 17938 223868 18440
rect 232548 17938 232868 18440
rect 238548 17938 238868 18440
rect 250548 17938 250868 18440
rect 263948 17938 264268 18440
rect 269948 17938 270268 18440
rect 272948 17938 273268 18440
rect 275948 17938 276268 18440
rect 281948 17938 282268 18440
rect 285948 17938 286268 18440
rect 293948 17938 294268 18440
rect 296948 17938 297268 18440
rect 299948 17938 300268 18440
rect 302948 18258 303268 18440
rect 108 15588 308 17746
rect 302946 16416 303268 18258
rect 302946 16088 303268 16094
rect 108 15382 308 15388
<< via1 >>
rect 302508 324332 302708 324532
rect 303926 321038 304246 321358
rect 108 319722 308 319922
rect 303926 318038 304246 318358
rect 108 316722 308 316922
rect 303926 315038 304246 315358
rect 108 313722 308 313922
rect 303926 312038 304246 312358
rect 108 310722 308 310922
rect 303926 309038 304246 309358
rect 108 307722 308 307922
rect 303926 306038 304246 306358
rect 108 304722 308 304922
rect 303926 303038 304246 303358
rect 108 301722 308 301922
rect 303926 300038 304246 300358
rect 108 298722 308 298922
rect 303926 297038 304246 297358
rect 108 295722 308 295922
rect 303926 294038 304246 294358
rect 108 292722 308 292922
rect 303926 291038 304246 291358
rect 108 289722 308 289922
rect 303926 288038 304246 288358
rect 108 286722 308 286922
rect 303926 285038 304246 285358
rect 108 283722 308 283922
rect 303926 282038 304246 282358
rect 108 280722 308 280922
rect 303926 279038 304246 279358
rect 108 277722 308 277922
rect 303926 276038 304246 276358
rect 108 274722 308 274922
rect 303926 273038 304246 273358
rect 108 271722 308 271922
rect 303926 270038 304246 270358
rect 108 268722 308 268922
rect 303926 267038 304246 267358
rect 108 265722 308 265922
rect 303926 264038 304246 264358
rect 108 262722 308 262922
rect 303926 261038 304246 261358
rect 108 259722 308 259922
rect 303926 258038 304246 258358
rect 108 256722 308 256922
rect 303926 255038 304246 255358
rect 108 253722 308 253922
rect 303926 252038 304246 252358
rect 108 250722 308 250922
rect 303926 249038 304246 249358
rect 108 247722 308 247922
rect 303926 246038 304246 246358
rect 108 244722 308 244922
rect 303926 243038 304246 243358
rect 108 241722 308 241922
rect 303926 240038 304246 240358
rect 108 238722 308 238922
rect 303926 237038 304246 237358
rect 108 235722 308 235922
rect 303926 234038 304246 234358
rect 108 232722 308 232922
rect 303926 231038 304246 231358
rect 108 229722 308 229922
rect 303926 228038 304246 228358
rect 108 226722 308 226922
rect 303926 225038 304246 225358
rect 108 223722 308 223922
rect 303926 222038 304246 222358
rect 108 220722 308 220922
rect 303926 219038 304246 219358
rect 108 217722 308 217922
rect 303926 216038 304246 216358
rect 108 214722 308 214922
rect 303926 213038 304246 213358
rect 108 211722 308 211922
rect 303926 210038 304246 210358
rect 108 208722 308 208922
rect 303926 207038 304246 207358
rect 108 205722 308 205922
rect 303926 204038 304246 204358
rect 108 202722 308 202922
rect 303926 201038 304246 201358
rect 108 199722 308 199922
rect 303926 198038 304246 198358
rect 108 196722 308 196922
rect 303926 195038 304246 195358
rect 108 193722 308 193922
rect 303926 192038 304246 192358
rect 108 190722 308 190922
rect 303926 189038 304246 189358
rect 108 187722 308 187922
rect 303926 186038 304246 186358
rect 108 184722 308 184922
rect 303926 183038 304246 183358
rect 108 181722 308 181922
rect 303926 180038 304246 180358
rect 108 178722 308 178922
rect 303926 177038 304246 177358
rect 108 175722 308 175922
rect 303926 174038 304246 174358
rect 108 172722 308 172922
rect 303926 171038 304246 171358
rect 108 169722 308 169922
rect 303926 168038 304246 168358
rect 108 166722 308 166922
rect 303926 165038 304246 165358
rect 108 163722 308 163922
rect 303926 162038 304246 162358
rect 108 160722 308 160922
rect 303926 159038 304246 159358
rect 108 157722 308 157922
rect 303926 156038 304246 156358
rect 108 154722 308 154922
rect 303926 153038 304246 153358
rect 108 151722 308 151922
rect 303926 150038 304246 150358
rect 108 148722 308 148922
rect 303926 147038 304246 147358
rect 108 145722 308 145922
rect 303926 144038 304246 144358
rect 108 142722 308 142922
rect 303926 141038 304246 141358
rect 108 139722 308 139922
rect 303926 138038 304246 138358
rect 108 136722 308 136922
rect 303926 135038 304246 135358
rect 108 133722 308 133922
rect 303926 132038 304246 132358
rect 108 130722 308 130922
rect 303926 129038 304246 129358
rect 108 127722 308 127922
rect 303926 126038 304246 126358
rect 108 124722 308 124922
rect 303926 123038 304246 123358
rect 108 121722 308 121922
rect 303926 120038 304246 120358
rect 108 118722 308 118922
rect 303926 117038 304246 117358
rect 108 115722 308 115922
rect 303926 114038 304246 114358
rect 108 112722 308 112922
rect 303926 111038 304246 111358
rect 108 109722 308 109922
rect 303926 108038 304246 108358
rect 108 106722 308 106922
rect 303926 105038 304246 105358
rect 108 103722 308 103922
rect 303926 102038 304246 102358
rect 108 100722 308 100922
rect 303926 99038 304246 99358
rect 108 97722 308 97922
rect 303926 96038 304246 96358
rect 108 94722 308 94922
rect 303926 93038 304246 93358
rect 108 91722 308 91922
rect 303926 90038 304246 90358
rect 108 88722 308 88922
rect 303926 87038 304246 87358
rect 108 85722 308 85922
rect 303926 84038 304246 84358
rect 108 82722 308 82922
rect 303926 81038 304246 81358
rect 108 79722 308 79922
rect 303926 78038 304246 78358
rect 108 76722 308 76922
rect 303926 75038 304246 75358
rect 108 73722 308 73922
rect 303926 72038 304246 72358
rect 108 70722 308 70922
rect 303926 69038 304246 69358
rect 108 67722 308 67922
rect 303926 66038 304246 66358
rect 108 64722 308 64922
rect 303926 63038 304246 63358
rect 108 61722 308 61922
rect 303926 60038 304246 60358
rect 108 58722 308 58922
rect 303926 57038 304246 57358
rect 108 55722 308 55922
rect 303926 54038 304246 54358
rect 108 52722 308 52922
rect 303926 51038 304246 51358
rect 108 49722 308 49922
rect 303926 48038 304246 48358
rect 108 46722 308 46922
rect 303926 45038 304246 45358
rect 108 43722 308 43922
rect 303926 42038 304246 42358
rect 108 40722 308 40922
rect 303926 39038 304246 39358
rect 108 37722 308 37922
rect 303926 36038 304246 36358
rect 108 34722 308 34922
rect 303926 33038 304246 33358
rect 108 31722 308 31922
rect 303926 30038 304246 30358
rect 108 28722 308 28922
rect 303926 27038 304246 27358
rect 108 25722 308 25922
rect 303926 24038 304246 24358
rect 108 22722 308 22922
rect 303926 21038 304246 21358
rect 3664 18440 3984 18760
rect 18088 18440 18408 18760
rect 32914 18440 33234 18760
rect 64256 18440 64576 18760
rect 121678 18440 121998 18760
rect 167548 18440 167868 18760
rect 180548 18440 180868 18760
rect 189548 18440 189868 18760
rect 198548 18440 198868 18760
rect 204548 18440 204868 18760
rect 211548 18440 211868 18760
rect 223548 18440 223868 18760
rect 232548 18440 232868 18760
rect 238548 18440 238868 18760
rect 250548 18440 250868 18760
rect 263948 18440 264268 18760
rect 269948 18440 270268 18760
rect 272948 18440 273268 18760
rect 275948 18440 276268 18760
rect 281948 18440 282268 18760
rect 285948 18440 286268 18760
rect 293948 18440 294268 18760
rect 296948 18440 297268 18760
rect 299948 18440 300268 18760
rect 302948 18440 303268 18760
rect -6198 17746 -5998 17946
rect 302946 16094 303268 16416
rect 108 15388 308 15588
<< metal2 >>
rect -8166 325380 -1626 325490
rect -5180 322442 -2032 322532
rect -5132 319402 -2402 319458
rect -5168 316366 -2742 316422
rect -5148 313238 -3102 313294
rect -3534 310258 -3444 310274
rect -5148 310202 -3444 310258
rect -5138 307166 -3932 307222
rect -5158 304038 -4342 304094
rect -4398 302338 -4342 304038
rect -3988 303948 -3932 307166
rect -3534 306948 -3444 310202
rect -3158 309948 -3102 313238
rect -2798 312948 -2742 316366
rect -2458 315930 -2402 319402
rect -2122 318948 -2032 322442
rect -1736 320838 -1626 325380
rect 1358 321238 1468 327120
rect 2118 321418 2228 326996
rect 302508 324532 302708 324542
rect 302502 324332 302508 324532
rect 302708 324332 302714 324532
rect 302508 324324 302708 324332
rect 303930 321358 304240 321362
rect 303920 321038 303926 321358
rect 304246 321038 304252 321358
rect 303930 321034 304240 321038
rect -1736 320728 -782 320838
rect 108 319922 308 319928
rect 98 319722 108 319922
rect 308 319722 316 319922
rect 108 319716 308 319722
rect -2122 318858 -802 318948
rect 303930 318358 304240 318362
rect 303920 318038 303926 318358
rect 304246 318038 304252 318358
rect 303930 318034 304240 318038
rect 108 316922 308 316928
rect 98 316722 108 316922
rect 308 316722 316 316922
rect 108 316716 308 316722
rect -2458 315874 -578 315930
rect 303930 315358 304240 315362
rect 303920 315038 303926 315358
rect 304246 315038 304252 315358
rect 303930 315034 304240 315038
rect 108 313922 308 313928
rect 98 313722 108 313922
rect 308 313722 316 313922
rect 108 313716 308 313722
rect -2798 312892 -622 312948
rect 303930 312358 304240 312362
rect 303920 312038 303926 312358
rect 304246 312038 304252 312358
rect 303930 312034 304240 312038
rect 108 310922 308 310928
rect 98 310722 108 310922
rect 308 310722 316 310922
rect 108 310716 308 310722
rect -3164 309858 -754 309948
rect 303930 309358 304240 309362
rect 303920 309038 303926 309358
rect 304246 309038 304252 309358
rect 303930 309034 304240 309038
rect 108 307922 308 307928
rect 98 307722 108 307922
rect 308 307722 316 307922
rect 108 307716 308 307722
rect -3534 306858 -802 306948
rect 303930 306358 304240 306362
rect 303920 306038 303926 306358
rect 304246 306038 304252 306358
rect 303930 306034 304240 306038
rect 108 304922 308 304928
rect 98 304722 108 304922
rect 308 304722 316 304922
rect 108 304716 308 304722
rect -4004 303858 -774 303948
rect 303930 303358 304240 303362
rect 303920 303038 303926 303358
rect 304246 303038 304252 303358
rect 303930 303034 304240 303038
rect -4398 302282 -692 302338
rect -1484 301058 -1004 301064
rect -5128 301002 -1004 301058
rect -1484 300974 -1004 301002
rect -5148 297966 -1542 298022
rect -1634 294948 -1544 297966
rect -1094 297948 -1004 300974
rect -834 300858 -744 302282
rect 108 301922 308 301928
rect 98 301722 108 301922
rect 308 301722 316 301922
rect 108 301716 308 301722
rect 303930 300358 304240 300362
rect 303920 300038 303926 300358
rect 304246 300038 304252 300358
rect 303930 300034 304240 300038
rect 108 298922 308 298928
rect 98 298722 108 298922
rect 308 298722 316 298922
rect 108 298716 308 298722
rect -1094 297858 -744 297948
rect 303930 297358 304240 297362
rect 303920 297038 303926 297358
rect 304246 297038 304252 297358
rect 303930 297034 304240 297038
rect 108 295922 308 295928
rect 98 295722 108 295922
rect 308 295722 316 295922
rect 108 295716 308 295722
rect -5148 294838 -2152 294894
rect -1634 294858 -724 294948
rect -3094 291858 -3004 292054
rect -2208 291918 -2152 294838
rect 303930 294358 304240 294362
rect 303920 294038 303926 294358
rect 304246 294038 304252 294358
rect 303930 294034 304240 294038
rect 108 292922 308 292928
rect 98 292722 108 292922
rect 308 292722 316 292922
rect 108 292716 308 292722
rect -2208 291862 -452 291918
rect -5148 291802 -3004 291858
rect -3094 288948 -3004 291802
rect 303930 291358 304240 291362
rect 303920 291038 303926 291358
rect 304246 291038 304252 291358
rect 303930 291034 304240 291038
rect 108 289922 308 289928
rect 98 289722 108 289922
rect 308 289722 316 289922
rect 108 289716 308 289722
rect -3094 288858 -784 288948
rect -3914 288730 -3824 288814
rect -5148 288674 -3824 288730
rect -3914 285948 -3824 288674
rect 303930 288358 304240 288362
rect 303920 288038 303926 288358
rect 304246 288038 304252 288358
rect 303930 288034 304240 288038
rect 108 286922 308 286928
rect 98 286722 108 286922
rect 308 286722 316 286922
rect 108 286716 308 286722
rect -3914 285858 -764 285948
rect -5138 285638 -4232 285694
rect -4288 284088 -4232 285638
rect 303930 285358 304240 285362
rect 303920 285038 303926 285358
rect 304246 285038 304252 285358
rect 303930 285034 304240 285038
rect -1104 284088 -1014 284104
rect -4288 284032 -962 284088
rect -1104 282948 -1014 284032
rect 108 283922 308 283928
rect 98 283722 108 283922
rect 308 283722 316 283922
rect 108 283716 308 283722
rect -1104 282858 -802 282948
rect -2204 282658 -2114 282764
rect -5158 282602 -2114 282658
rect -2204 279948 -2114 282602
rect 303930 282358 304240 282362
rect 303920 282038 303926 282358
rect 304246 282038 304252 282358
rect 303930 282034 304240 282038
rect 108 280922 308 280928
rect 98 280722 108 280922
rect 308 280722 316 280922
rect 108 280716 308 280722
rect -2204 279858 -802 279948
rect -5218 279474 -1962 279530
rect -2054 276948 -1964 279474
rect 303930 279358 304240 279362
rect 303920 279038 303926 279358
rect 304246 279038 304252 279358
rect 303930 279034 304240 279038
rect 108 277922 308 277928
rect 98 277722 108 277922
rect 308 277722 316 277922
rect 108 277716 308 277722
rect -2054 276858 -784 276948
rect -892 276494 -802 276524
rect -5188 276438 -802 276494
rect -892 273858 -802 276438
rect 303930 276358 304240 276362
rect 303920 276038 303926 276358
rect 304246 276038 304252 276358
rect 303930 276034 304240 276038
rect 108 274922 308 274928
rect 98 274722 108 274922
rect 308 274722 316 274922
rect 108 274716 308 274722
rect -3964 273458 -3874 273584
rect -5228 273402 -3874 273458
rect -3964 270948 -3874 273402
rect 303930 273358 304240 273362
rect 303920 273038 303926 273358
rect 304246 273038 304252 273358
rect 303930 273034 304240 273038
rect 108 271922 308 271928
rect 98 271722 108 271922
rect 308 271722 316 271922
rect 108 271716 308 271722
rect -3964 270858 -802 270948
rect 303930 270358 304240 270362
rect -5168 270274 -4582 270330
rect -4638 267948 -4582 270274
rect 303920 270038 303926 270358
rect 304246 270038 304252 270358
rect 303930 270034 304240 270038
rect 108 268922 308 268928
rect 98 268722 108 268922
rect 308 268722 316 268922
rect 108 268716 308 268722
rect -4638 267882 -802 267948
rect -4614 267858 -802 267882
rect -4284 267294 -4194 267424
rect 303930 267358 304240 267362
rect -5148 267238 -4194 267294
rect -4284 264948 -4194 267238
rect 303920 267038 303926 267358
rect 304246 267038 304252 267358
rect 303930 267034 304240 267038
rect 108 265922 308 265928
rect 98 265722 108 265922
rect 308 265722 316 265922
rect 108 265716 308 265722
rect -4284 264858 -802 264948
rect 303930 264358 304240 264362
rect -5148 264110 -1932 264166
rect -1988 261948 -1932 264110
rect 303920 264038 303926 264358
rect 304246 264038 304252 264358
rect 303930 264034 304240 264038
rect 108 262922 308 262928
rect 98 262722 108 262922
rect 308 262722 316 262922
rect 108 262716 308 262722
rect -1988 261858 -802 261948
rect -1988 261812 -1932 261858
rect 303930 261358 304240 261362
rect -5178 261074 -1092 261130
rect -1148 258948 -1092 261074
rect 303920 261038 303926 261358
rect 304246 261038 304252 261358
rect 303930 261034 304240 261038
rect 108 259922 308 259928
rect 98 259722 108 259922
rect 308 259722 316 259922
rect 108 259716 308 259722
rect -1148 258858 -774 258948
rect -1148 258822 -1092 258858
rect 303930 258358 304240 258362
rect -5218 258038 -1112 258094
rect 303920 258038 303926 258358
rect 304246 258038 304252 258358
rect -1168 255948 -1112 258038
rect 303930 258034 304240 258038
rect 108 256922 308 256928
rect 98 256722 108 256922
rect 308 256722 316 256922
rect 108 256716 308 256722
rect -1168 255858 -802 255948
rect -1168 255842 -1112 255858
rect 303930 255358 304240 255362
rect 303920 255038 303926 255358
rect 304246 255038 304252 255358
rect 303930 255034 304240 255038
rect -5168 254910 -1172 254966
rect -1228 252948 -1172 254910
rect 108 253922 308 253928
rect 98 253722 108 253922
rect 308 253722 316 253922
rect 108 253716 308 253722
rect -1228 252858 -802 252948
rect -1228 252852 -1172 252858
rect 303930 252358 304240 252362
rect 303920 252038 303926 252358
rect 304246 252038 304252 252358
rect 303930 252034 304240 252038
rect -5208 251874 -1402 251930
rect -1458 249948 -1402 251874
rect 108 250922 308 250928
rect 98 250722 108 250922
rect 308 250722 316 250922
rect 108 250716 308 250722
rect -1458 249892 -794 249948
rect -1434 249858 -794 249892
rect 303930 249358 304240 249362
rect -884 248894 -794 249084
rect 303920 249038 303926 249358
rect 304246 249038 304252 249358
rect 303930 249034 304240 249038
rect -5128 248838 -792 248894
rect -884 246858 -794 248838
rect 108 247922 308 247928
rect 98 247722 108 247922
rect 308 247722 316 247922
rect 108 247716 308 247722
rect 303930 246358 304240 246362
rect 303920 246038 303926 246358
rect 304246 246038 304252 246358
rect 303930 246034 304240 246038
rect -892 245766 -802 245884
rect -5268 245710 -802 245766
rect -892 243858 -802 245710
rect 108 244922 308 244928
rect 98 244722 108 244922
rect 308 244722 316 244922
rect 108 244716 308 244722
rect 303930 243358 304240 243362
rect 303920 243038 303926 243358
rect 304246 243038 304252 243358
rect 303930 243034 304240 243038
rect -5228 242674 -832 242730
rect -888 240852 -832 242674
rect 108 241922 308 241928
rect 98 241722 108 241922
rect 308 241722 316 241922
rect 108 241716 308 241722
rect 303930 240358 304240 240362
rect 303920 240038 303926 240358
rect 304246 240038 304252 240358
rect 303930 240034 304240 240038
rect -5158 239638 -812 239694
rect -868 237892 -812 239638
rect 108 238922 308 238928
rect 98 238722 108 238922
rect 308 238722 316 238922
rect 108 238716 308 238722
rect 303930 237358 304240 237362
rect 303920 237038 303926 237358
rect 304246 237038 304252 237358
rect 303930 237034 304240 237038
rect -892 236566 -802 236724
rect -5188 236510 -802 236566
rect -892 234858 -802 236510
rect 108 235922 308 235928
rect 98 235722 108 235922
rect 308 235722 316 235922
rect 108 235716 308 235722
rect 303930 234358 304240 234362
rect 303920 234038 303926 234358
rect 304246 234038 304252 234358
rect 303930 234034 304240 234038
rect -5168 233474 -892 233530
rect -948 231852 -892 233474
rect 108 232922 308 232928
rect 98 232722 108 232922
rect 308 232722 316 232922
rect 108 232716 308 232722
rect 303930 231358 304240 231362
rect 303920 231038 303926 231358
rect 304246 231038 304252 231358
rect 303930 231034 304240 231038
rect -5168 228948 -5112 230402
rect 108 229922 308 229928
rect 98 229722 108 229922
rect 308 229722 316 229922
rect 108 229716 308 229722
rect -5168 228892 -784 228948
rect -5154 228858 -784 228892
rect 303930 228358 304240 228362
rect 303920 228038 303926 228358
rect 304246 228038 304252 228358
rect 303930 228034 304240 228038
rect -5138 227310 -612 227366
rect -834 225858 -744 227310
rect 108 226922 308 226928
rect 98 226722 108 226922
rect 308 226722 316 226922
rect 108 226716 308 226722
rect 303930 225358 304240 225362
rect 303920 225038 303926 225358
rect 304246 225038 304252 225358
rect 303930 225034 304240 225038
rect -5194 224264 -802 224354
rect -892 222858 -802 224264
rect 108 223922 308 223928
rect 98 223722 108 223922
rect 308 223722 316 223922
rect 108 223716 308 223722
rect 303930 222358 304240 222362
rect 303920 222038 303926 222358
rect 304246 222038 304252 222358
rect 303930 222034 304240 222038
rect -5148 221146 -808 221202
rect -864 219882 -808 221146
rect 108 220922 308 220928
rect 98 220722 108 220922
rect 308 220722 316 220922
rect 108 220716 308 220722
rect 303930 219358 304240 219362
rect 303920 219038 303926 219358
rect 304246 219038 304252 219358
rect 303930 219034 304240 219038
rect -808 218178 -752 218202
rect -5128 218122 -752 218178
rect -808 216872 -752 218122
rect 108 217922 308 217928
rect 98 217722 108 217922
rect 308 217722 316 217922
rect 108 217716 308 217722
rect 303930 216358 304240 216362
rect 303920 216038 303926 216358
rect 304246 216038 304252 216358
rect 303930 216034 304240 216038
rect -5128 215082 -752 215138
rect -808 213858 -752 215082
rect 108 214922 308 214928
rect 98 214722 108 214922
rect 308 214722 316 214922
rect 108 214716 308 214722
rect 303930 213358 304240 213362
rect 303920 213038 303926 213358
rect 304246 213038 304252 213358
rect 303930 213034 304240 213038
rect -5134 211914 -802 212004
rect 108 211922 308 211928
rect -892 210858 -802 211914
rect 98 211722 108 211922
rect 308 211722 316 211922
rect 108 211716 308 211722
rect 303930 210358 304240 210362
rect 303920 210038 303926 210358
rect 304246 210038 304252 210358
rect 303930 210034 304240 210038
rect -5128 208910 -732 208966
rect 108 208922 308 208928
rect -892 207872 -732 208910
rect 98 208722 108 208922
rect 308 208722 316 208922
rect 108 208716 308 208722
rect -892 207858 -764 207872
rect 303930 207358 304240 207362
rect 303920 207038 303926 207358
rect 304246 207038 304252 207358
rect 303930 207034 304240 207038
rect 108 205922 308 205928
rect -5168 205782 -802 205838
rect -858 204842 -802 205782
rect 98 205722 108 205922
rect 308 205722 316 205922
rect 108 205716 308 205722
rect 303930 204358 304240 204362
rect 303920 204038 303926 204358
rect 304246 204038 304252 204358
rect 303930 204034 304240 204038
rect 108 202922 308 202928
rect -5158 202746 -762 202802
rect -884 201858 -794 202746
rect 98 202722 108 202922
rect 308 202722 316 202922
rect 108 202716 308 202722
rect 303930 201358 304240 201362
rect 303920 201038 303926 201358
rect 304246 201038 304252 201358
rect 303930 201034 304240 201038
rect 108 199922 308 199928
rect -5208 199710 -722 199766
rect 98 199722 108 199922
rect 308 199722 316 199922
rect 108 199716 308 199722
rect -778 198852 -722 199710
rect 303930 198358 304240 198362
rect 303920 198038 303926 198358
rect 304246 198038 304252 198358
rect 303930 198034 304240 198038
rect 108 196922 308 196928
rect 98 196722 108 196922
rect 308 196722 316 196922
rect 108 196716 308 196722
rect -5144 196582 -1202 196638
rect -1258 195948 -1202 196582
rect -1258 195858 -792 195948
rect -1258 195804 -1202 195858
rect 303930 195358 304240 195362
rect 303920 195038 303926 195358
rect 304246 195038 304252 195358
rect 303930 195034 304240 195038
rect 108 193922 308 193928
rect 98 193722 108 193922
rect 308 193722 316 193922
rect 108 193716 308 193722
rect -5144 193552 -4890 193642
rect -4980 192948 -4890 193552
rect -4980 192858 -782 192948
rect 303930 192358 304240 192362
rect 303920 192038 303926 192358
rect 304246 192038 304252 192358
rect 303930 192034 304240 192038
rect 108 190922 308 190928
rect 98 190722 108 190922
rect 308 190722 316 190922
rect 108 190716 308 190722
rect -5134 190510 -736 190566
rect -792 189806 -736 190510
rect 303930 189358 304240 189362
rect 303920 189038 303926 189358
rect 304246 189038 304252 189358
rect 303930 189034 304240 189038
rect 108 187922 308 187928
rect 98 187722 108 187922
rect 308 187722 316 187922
rect 108 187716 308 187722
rect -5140 186948 -5050 187460
rect -5140 186858 -792 186948
rect 303930 186358 304240 186362
rect 303920 186038 303926 186358
rect 304246 186038 304252 186358
rect 303930 186034 304240 186038
rect 108 184922 308 184928
rect 98 184722 108 184922
rect 308 184722 316 184922
rect 108 184716 308 184722
rect -5140 183948 -5050 184424
rect -5140 183858 -578 183948
rect 303930 183358 304240 183362
rect 303920 183038 303926 183358
rect 304246 183038 304252 183358
rect 303930 183034 304240 183038
rect 108 181922 308 181928
rect 98 181722 108 181922
rect 308 181722 316 181922
rect 108 181716 308 181722
rect -5184 180948 -5094 181338
rect -5184 180858 -802 180948
rect 303930 180358 304240 180362
rect 303920 180038 303926 180358
rect 304246 180038 304252 180358
rect 303930 180034 304240 180038
rect 108 178922 308 178928
rect 98 178722 108 178922
rect 308 178722 316 178922
rect 108 178716 308 178722
rect -5168 177948 -5078 178234
rect -5168 177858 -572 177948
rect 303930 177358 304240 177362
rect 303920 177038 303926 177358
rect 304246 177038 304252 177358
rect 303930 177034 304240 177038
rect 108 175922 308 175928
rect 98 175722 108 175922
rect 308 175722 316 175922
rect 108 175716 308 175722
rect -5128 174948 -5072 175202
rect -5128 174858 -690 174948
rect -5128 174790 -5072 174858
rect 303930 174358 304240 174362
rect 303920 174038 303926 174358
rect 304246 174038 304252 174358
rect 303930 174034 304240 174038
rect 108 172922 308 172928
rect 98 172722 108 172922
rect 308 172722 316 172922
rect 108 172716 308 172722
rect -5208 171948 -5118 172064
rect -5208 171858 -782 171948
rect 303930 171358 304240 171362
rect 303920 171038 303926 171358
rect 304246 171038 304252 171358
rect 303930 171034 304240 171038
rect 108 169922 308 169928
rect 98 169722 108 169922
rect 308 169722 316 169922
rect 108 169716 308 169722
rect -5156 168948 -5066 169080
rect -5156 168858 -802 168948
rect 303930 168358 304240 168362
rect 303920 168038 303926 168358
rect 304246 168038 304252 168358
rect 303930 168034 304240 168038
rect 108 166922 308 166928
rect 98 166722 108 166922
rect 308 166722 316 166922
rect 108 166716 308 166722
rect -5144 165948 -5054 166032
rect -5144 165858 -730 165948
rect 303930 165358 304240 165362
rect 303920 165038 303926 165358
rect 304246 165038 304252 165358
rect 303930 165034 304240 165038
rect 108 163922 308 163928
rect 98 163722 108 163922
rect 308 163722 316 163922
rect 108 163716 308 163722
rect -5144 162858 -770 162948
rect 303930 162358 304240 162362
rect 303920 162038 303926 162358
rect 304246 162038 304252 162358
rect 303930 162034 304240 162038
rect 108 160922 308 160928
rect 98 160722 108 160922
rect 308 160722 316 160922
rect 108 160716 308 160722
rect -5922 159858 -798 159948
rect -5922 159778 -816 159858
rect 303930 159358 304240 159362
rect 303920 159038 303926 159358
rect 304246 159038 304252 159358
rect 303930 159034 304240 159038
rect 108 157922 308 157928
rect 98 157722 108 157922
rect 308 157722 316 157922
rect 108 157716 308 157722
rect -826 156900 -736 156948
rect -5162 156856 -736 156900
rect -5168 156742 -736 156856
rect 303930 156358 304240 156362
rect 303920 156038 303926 156358
rect 304246 156038 304252 156358
rect 303930 156034 304240 156038
rect 108 154922 308 154928
rect 98 154722 108 154922
rect 308 154722 316 154922
rect 108 154716 308 154722
rect -882 153678 -792 153948
rect -5134 153588 -792 153678
rect 303930 153358 304240 153362
rect 303920 153038 303926 153358
rect 304246 153038 304252 153358
rect 303930 153034 304240 153038
rect 108 151922 308 151928
rect 98 151722 108 151922
rect 308 151722 316 151922
rect 108 151716 308 151722
rect -5242 150584 -5010 150658
rect -892 150584 -802 150948
rect -5242 150568 -802 150584
rect -5100 150494 -802 150568
rect 303930 150358 304240 150362
rect 303920 150038 303926 150358
rect 304246 150038 304252 150358
rect 303930 150034 304240 150038
rect 108 148922 308 148928
rect 98 148722 108 148922
rect 308 148722 316 148922
rect 108 148716 308 148722
rect -5122 147428 -5032 147554
rect -882 147428 -792 147948
rect -5122 147338 -792 147428
rect 303930 147358 304240 147362
rect 303920 147038 303926 147358
rect 304246 147038 304252 147358
rect 303930 147034 304240 147038
rect 108 145922 308 145928
rect 98 145722 108 145922
rect 308 145722 316 145922
rect 108 145716 308 145722
rect -882 144568 -792 144948
rect -5178 144478 -792 144568
rect -5178 144416 -838 144478
rect 303930 144358 304240 144362
rect 303920 144038 303926 144358
rect 304246 144038 304252 144358
rect 303930 144034 304240 144038
rect 108 142922 308 142928
rect 98 142722 108 142922
rect 308 142722 316 142922
rect 108 142716 308 142722
rect -866 141504 -776 141948
rect -5140 141414 -776 141504
rect -5140 141352 -816 141414
rect 303930 141358 304240 141362
rect 303920 141038 303926 141358
rect 304246 141038 304252 141358
rect 303930 141034 304240 141038
rect 108 139922 308 139928
rect 98 139722 108 139922
rect 308 139722 316 139922
rect 108 139716 308 139722
rect -860 138338 -770 138948
rect 303930 138358 304240 138362
rect -5178 138248 -770 138338
rect 303920 138038 303926 138358
rect 304246 138038 304252 138358
rect 303930 138034 304240 138038
rect 108 136922 308 136928
rect 98 136722 108 136922
rect 308 136722 316 136922
rect 108 136716 308 136722
rect -892 135340 -802 135948
rect 303930 135358 304240 135362
rect -5190 135250 -802 135340
rect -5134 135182 -804 135250
rect 303920 135038 303926 135358
rect 304246 135038 304252 135358
rect 303930 135034 304240 135038
rect 108 133922 308 133928
rect 98 133722 108 133922
rect 308 133722 316 133922
rect 108 133716 308 133722
rect -848 132368 -758 132948
rect -5174 132278 -758 132368
rect 303930 132358 304240 132362
rect -5174 132186 -5084 132278
rect 303920 132038 303926 132358
rect 304246 132038 304252 132358
rect 303930 132034 304240 132038
rect 108 130922 308 130928
rect 98 130722 108 130922
rect 308 130722 316 130922
rect 108 130716 308 130722
rect -880 129084 -790 129948
rect 303930 129358 304240 129362
rect -5186 128936 -790 129084
rect 303920 129038 303926 129358
rect 304246 129038 304252 129358
rect 303930 129034 304240 129038
rect 108 127922 308 127928
rect 98 127722 108 127922
rect 308 127722 316 127922
rect 108 127716 308 127722
rect -852 126084 -762 126948
rect 303930 126358 304240 126362
rect -5198 125938 -762 126084
rect 303920 126038 303926 126358
rect 304246 126038 304252 126358
rect 303930 126034 304240 126038
rect 108 124922 308 124928
rect 98 124722 108 124922
rect 308 124722 316 124922
rect 108 124716 308 124722
rect -892 122976 -802 123948
rect 303930 123358 304240 123362
rect 303920 123038 303926 123358
rect 304246 123038 304252 123358
rect 303930 123034 304240 123038
rect -5140 122790 -802 122976
rect 108 121922 308 121928
rect 98 121722 108 121922
rect 308 121722 316 121922
rect 108 121716 308 121722
rect -5128 120948 -5072 121158
rect -5140 120858 -762 120948
rect -5128 119854 -5072 120858
rect 303930 120358 304240 120362
rect 303920 120038 303926 120358
rect 304246 120038 304252 120358
rect 303930 120034 304240 120038
rect 108 118922 308 118928
rect 98 118722 108 118922
rect 308 118722 316 118922
rect 108 118716 308 118722
rect -5186 117858 -802 117948
rect -5186 116774 -5096 117858
rect 303930 117358 304240 117362
rect 303920 117038 303926 117358
rect 304246 117038 304252 117358
rect 303930 117034 304240 117038
rect 108 115922 308 115928
rect 98 115722 108 115922
rect 308 115722 316 115922
rect 108 115716 308 115722
rect -5158 114858 -614 114948
rect -5158 113650 -5068 114858
rect 303930 114358 304240 114362
rect 303920 114038 303926 114358
rect 304246 114038 304252 114358
rect 303930 114034 304240 114038
rect 108 112922 308 112928
rect 98 112722 108 112922
rect 308 112722 316 112922
rect 108 112716 308 112722
rect -5192 111858 -768 111948
rect -5192 110632 -5102 111858
rect 303930 111358 304240 111362
rect 303920 111038 303926 111358
rect 304246 111038 304252 111358
rect 303930 111034 304240 111038
rect 108 109922 308 109928
rect 98 109722 108 109922
rect 308 109722 316 109922
rect 108 109716 308 109722
rect -5124 108858 -802 108948
rect -5124 107622 -5034 108858
rect 303930 108358 304240 108362
rect 303920 108038 303926 108358
rect 304246 108038 304252 108358
rect 303930 108034 304240 108038
rect 108 106922 308 106928
rect 98 106722 108 106922
rect 308 106722 316 106922
rect 108 106716 308 106722
rect -836 104588 -746 105948
rect 303930 105358 304240 105362
rect 303920 105038 303926 105358
rect 304246 105038 304252 105358
rect 303930 105034 304240 105038
rect -5164 104498 -746 104588
rect -5164 104490 -768 104498
rect 108 103922 308 103928
rect 98 103722 108 103922
rect 308 103722 316 103922
rect 108 103716 308 103722
rect -892 101548 -802 102948
rect 303930 102358 304240 102362
rect 303920 102038 303926 102358
rect 304246 102038 304252 102358
rect 303930 102034 304240 102038
rect -5174 101458 -802 101548
rect -892 101258 -802 101458
rect 108 100922 308 100928
rect 98 100722 108 100922
rect 308 100722 316 100922
rect 108 100716 308 100722
rect -892 98428 -802 99948
rect 303930 99358 304240 99362
rect 303920 99038 303926 99358
rect 304246 99038 304252 99358
rect 303930 99034 304240 99038
rect -5208 98338 -802 98428
rect -892 98076 -802 98338
rect 108 97922 308 97928
rect 98 97722 108 97922
rect 308 97722 316 97922
rect 108 97716 308 97722
rect -880 95396 -790 96948
rect 303930 96358 304240 96362
rect 303920 96038 303926 96358
rect 304246 96038 304252 96358
rect 303930 96034 304240 96038
rect -5180 95306 -790 95396
rect -880 95008 -790 95306
rect 108 94922 308 94928
rect 98 94722 108 94922
rect 308 94722 316 94922
rect 108 94716 308 94722
rect -870 92316 -780 93948
rect 303930 93358 304240 93362
rect 303920 93038 303926 93358
rect 304246 93038 304252 93358
rect 303930 93034 304240 93038
rect -5232 92226 -780 92316
rect -870 91912 -780 92226
rect 108 91922 308 91928
rect 98 91722 108 91922
rect 308 91722 316 91922
rect 108 91716 308 91722
rect -852 89208 -762 90948
rect 303930 90358 304240 90362
rect 303920 90038 303926 90358
rect 304246 90038 304252 90358
rect 303930 90034 304240 90038
rect -5192 89118 -762 89208
rect -852 89016 -762 89118
rect 108 88922 308 88928
rect 98 88722 108 88922
rect 308 88722 316 88922
rect 108 88716 308 88722
rect -836 86198 -746 87948
rect 303930 87358 304240 87362
rect 303920 87038 303926 87358
rect 304246 87038 304252 87358
rect 303930 87034 304240 87038
rect -5128 86108 -746 86198
rect -836 85976 -746 86108
rect 108 85922 308 85928
rect 98 85722 108 85922
rect 308 85722 316 85922
rect 108 85716 308 85722
rect -796 83152 -706 84948
rect 303930 84358 304240 84362
rect 303920 84038 303926 84358
rect 304246 84038 304252 84358
rect 303930 84034 304240 84038
rect -5220 83062 -706 83152
rect -796 82720 -706 83062
rect 108 82922 308 82928
rect 98 82722 108 82922
rect 308 82722 316 82922
rect 108 82716 308 82722
rect -880 80022 -790 81948
rect 303930 81358 304240 81362
rect 303920 81038 303926 81358
rect 304246 81038 304252 81358
rect 303930 81034 304240 81038
rect -5202 79932 -790 80022
rect -880 79526 -790 79932
rect 108 79922 308 79928
rect 98 79722 108 79922
rect 308 79722 316 79922
rect 108 79716 308 79722
rect -858 76948 -768 78948
rect 303930 78358 304240 78362
rect 303920 78038 303926 78358
rect 304246 78038 304252 78358
rect 303930 78034 304240 78038
rect -5208 76858 -768 76948
rect 108 76922 308 76928
rect -858 76390 -768 76858
rect 98 76722 108 76922
rect 308 76722 316 76922
rect 108 76716 308 76722
rect -5164 73772 -5074 74058
rect -790 73772 -700 75948
rect 303930 75358 304240 75362
rect 303920 75038 303926 75358
rect 304246 75038 304252 75358
rect 303930 75034 304240 75038
rect 108 73922 308 73928
rect -5164 73682 -700 73772
rect 98 73722 108 73922
rect 308 73722 316 73922
rect 108 73716 308 73722
rect -790 73476 -700 73682
rect -830 70796 -740 72948
rect 303930 72358 304240 72362
rect 303920 72038 303926 72358
rect 304246 72038 304252 72358
rect 303930 72034 304240 72038
rect 108 70922 308 70928
rect -5152 70706 -740 70796
rect 98 70722 108 70922
rect 308 70722 316 70922
rect 108 70716 308 70722
rect -830 70580 -740 70706
rect -5168 67654 -5078 67774
rect -892 67654 -802 69948
rect 303930 69358 304240 69362
rect 303920 69038 303926 69358
rect 304246 69038 304252 69358
rect 303930 69034 304240 69038
rect 108 67922 308 67928
rect 98 67722 108 67922
rect 308 67722 316 67922
rect 108 67716 308 67722
rect -5168 67564 -802 67654
rect -892 67370 -802 67564
rect -608 64618 -552 66924
rect 303930 66358 304240 66362
rect 303920 66038 303926 66358
rect 304246 66038 304252 66358
rect 303930 66034 304240 66038
rect 108 64922 308 64928
rect 98 64722 108 64922
rect 308 64722 316 64922
rect 108 64716 308 64722
rect -5226 64562 -552 64618
rect -5208 63858 -642 63948
rect -5208 61354 -5118 63858
rect 303930 63358 304240 63362
rect 303920 63038 303926 63358
rect 304246 63038 304252 63358
rect 303930 63034 304240 63038
rect 108 61922 308 61928
rect 98 61722 108 61922
rect 308 61722 316 61922
rect 108 61716 308 61722
rect -5242 60858 -700 60948
rect -5242 58378 -5152 60858
rect 303930 60358 304240 60362
rect 303920 60038 303926 60358
rect 304246 60038 304252 60358
rect 303930 60034 304240 60038
rect 108 58922 308 58928
rect 98 58722 108 58922
rect 308 58722 316 58922
rect 108 58716 308 58722
rect -5214 57858 -774 57948
rect -5214 55224 -5124 57858
rect 303930 57358 304240 57362
rect 303920 57038 303926 57358
rect 304246 57038 304252 57358
rect 303930 57034 304240 57038
rect 108 55922 308 55928
rect 98 55722 108 55922
rect 308 55722 316 55922
rect 108 55716 308 55722
rect -5242 54858 -774 54948
rect -5242 52316 -5152 54858
rect 303930 54358 304240 54362
rect 303920 54038 303926 54358
rect 304246 54038 304252 54358
rect 303930 54034 304240 54038
rect 108 52922 308 52928
rect 98 52722 108 52922
rect 308 52722 316 52922
rect 108 52716 308 52722
rect -322 49346 -266 52178
rect 303930 51358 304240 51362
rect 303920 51038 303926 51358
rect 304246 51038 304252 51358
rect 303930 51034 304240 51038
rect 108 49922 308 49928
rect 98 49722 108 49922
rect 308 49722 316 49922
rect 108 49716 308 49722
rect -5146 49290 -266 49346
rect -5226 48858 -488 48948
rect -5226 45970 -5136 48858
rect 303930 48358 304240 48362
rect 303920 48038 303926 48358
rect 304246 48038 304252 48358
rect 303930 48034 304240 48038
rect 108 46922 308 46928
rect 98 46722 108 46922
rect 308 46722 316 46922
rect 108 46716 308 46722
rect -3540 45858 -802 45948
rect -3540 43182 -3450 45858
rect 303930 45358 304240 45362
rect 303920 45038 303926 45358
rect 304246 45038 304252 45358
rect 303930 45034 304240 45038
rect 108 43922 308 43928
rect 98 43722 108 43922
rect 308 43722 316 43922
rect 108 43716 308 43722
rect -5188 43126 -3342 43182
rect -3540 42490 -3450 43126
rect -2360 42948 -2304 43190
rect -2458 42858 -802 42948
rect -2360 40054 -2304 42858
rect 303930 42358 304240 42362
rect 303920 42038 303926 42358
rect 304246 42038 304252 42358
rect 303930 42034 304240 42038
rect 108 40922 308 40928
rect 98 40722 108 40922
rect 308 40722 316 40922
rect 108 40716 308 40722
rect -5256 39998 -2304 40054
rect -750 38442 -660 39948
rect 303930 39358 304240 39362
rect 303920 39038 303926 39358
rect 304246 39038 304252 39358
rect 303930 39034 304240 39038
rect -1990 38386 -496 38442
rect -1990 37018 -1934 38386
rect -750 38280 -660 38386
rect 108 37922 308 37928
rect 98 37722 108 37922
rect 308 37722 316 37922
rect 108 37716 308 37722
rect -5130 36962 -1934 37018
rect -462 35564 -372 36948
rect 303930 36358 304240 36362
rect 303920 36038 303926 36358
rect 304246 36038 304252 36358
rect 303930 36034 304240 36038
rect -2434 35508 -372 35564
rect -2434 33982 -2378 35508
rect -462 35254 -372 35508
rect 108 34922 308 34928
rect 98 34722 108 34922
rect 308 34722 316 34922
rect 108 34716 308 34722
rect -5144 33926 -2378 33982
rect -772 32850 -716 34558
rect 303930 33358 304240 33362
rect 303920 33038 303926 33358
rect 304246 33038 304252 33358
rect 303930 33034 304240 33038
rect -3298 32794 -716 32850
rect -3298 30854 -3242 32794
rect 108 31922 308 31928
rect 98 31722 108 31922
rect 308 31722 316 31922
rect 108 31716 308 31722
rect -5174 30798 -3242 30854
rect -720 29740 -630 30948
rect 303930 30358 304240 30362
rect 303920 30038 303926 30358
rect 304246 30038 304252 30358
rect 303930 30034 304240 30038
rect -2904 29684 -584 29740
rect -2904 27818 -2848 29684
rect -720 29384 -584 29684
rect -720 29260 -630 29384
rect 108 28922 308 28928
rect 98 28722 108 28922
rect 308 28722 316 28922
rect 108 28716 308 28722
rect -5174 27762 -2848 27818
rect -756 26900 -666 27948
rect 303930 27358 304240 27362
rect 303920 27038 303926 27358
rect 304246 27038 304252 27358
rect 303930 27034 304240 27038
rect -2592 26844 -628 26900
rect -2592 24782 -2536 26844
rect -756 26590 -666 26844
rect 108 25922 308 25928
rect 98 25722 108 25922
rect 308 25722 316 25922
rect 108 25716 308 25722
rect -5188 24726 -2536 24782
rect -764 23910 -674 24948
rect 303930 24358 304240 24362
rect 303920 24038 303926 24358
rect 304246 24038 304252 24358
rect 303930 24034 304240 24038
rect -5244 23854 -458 23910
rect -5244 21598 -5188 23854
rect -764 23518 -674 23854
rect 108 22922 308 22928
rect 98 22722 108 22922
rect 308 22722 316 22922
rect 108 22716 308 22722
rect -4016 21858 -736 21948
rect -4016 18618 -3926 21858
rect 303930 21358 304240 21362
rect 303920 21038 303926 21358
rect 304246 21038 304252 21358
rect 303930 21034 304240 21038
rect 302848 19472 303028 19478
rect 302848 19292 307364 19472
rect 302848 19278 303028 19292
rect 38312 19214 38562 19226
rect 19850 19188 20100 19202
rect 19850 18978 19874 19188
rect 20084 18978 20100 19188
rect 29084 19062 29304 19070
rect 13790 18930 14040 18950
rect 19850 18944 20100 18978
rect 25908 19006 26226 19028
rect 13650 18924 14040 18930
rect 7470 18886 7720 18910
rect 5316 18784 5566 18810
rect 4518 18780 5566 18784
rect 3664 18760 3984 18766
rect -5180 18510 -3804 18618
rect -5180 18496 -3926 18510
rect 2316 18440 2566 18466
rect 3660 18444 3664 18754
rect 3984 18444 3988 18754
rect 4518 18570 5332 18780
rect 5542 18570 5566 18780
rect 7470 18676 7486 18886
rect 7696 18676 7720 18886
rect 7470 18652 7720 18676
rect 10692 18830 10942 18858
rect 4518 18564 5566 18570
rect 1498 18434 2566 18440
rect 3664 18434 3984 18440
rect 1498 18224 2332 18434
rect 2542 18224 2566 18434
rect 1498 18220 2566 18224
rect -6198 17946 -5998 17956
rect -6198 17738 -5998 17746
rect 1498 16556 1718 18220
rect 2316 18208 2566 18220
rect 4518 16430 4738 18564
rect 5316 18552 5566 18564
rect 7482 16456 7702 18652
rect 10692 18620 10716 18830
rect 10926 18620 10942 18830
rect 10692 18600 10942 18620
rect 13650 18714 13806 18924
rect 14016 18714 14040 18924
rect 13650 18692 14040 18714
rect 16900 18812 17150 18824
rect 10710 16526 10930 18600
rect 13650 16450 13870 18692
rect 16900 18602 16916 18812
rect 17126 18602 17150 18812
rect 18088 18760 18408 18766
rect 16900 18566 17150 18602
rect 16910 16694 17130 18566
rect 18084 18444 18088 18754
rect 18408 18444 18412 18754
rect 18088 18434 18408 18440
rect 16746 16474 17130 16694
rect 19868 16482 20088 18944
rect 25908 18796 25948 19006
rect 26158 18796 26226 19006
rect 29074 18842 29084 19052
rect 29304 18842 29312 19052
rect 35298 19050 35584 19066
rect 32332 18986 32542 18990
rect 32124 18982 32548 18986
rect 25908 18762 26226 18796
rect 22872 18654 23188 18672
rect 22872 18444 22902 18654
rect 23112 18444 23188 18654
rect 22872 18406 23188 18444
rect 22896 16456 23116 18406
rect 25942 16450 26162 18762
rect 29084 16482 29304 18842
rect 32124 18772 32332 18982
rect 32542 18772 32548 18982
rect 35298 18840 35332 19050
rect 35542 18840 35584 19050
rect 38312 19004 38332 19214
rect 38542 19004 38562 19214
rect 56594 19158 56844 19178
rect 38312 18968 38562 19004
rect 47318 19126 47568 19144
rect 35298 18828 35584 18840
rect 32124 18766 32548 18772
rect 32124 18762 32542 18766
rect 32124 16526 32344 18762
rect 32914 18760 33234 18766
rect 32910 18444 32914 18754
rect 33234 18444 33238 18754
rect 32914 18434 33234 18440
rect 35328 17248 35548 18828
rect 35196 17028 35548 17248
rect 35196 16482 35416 17028
rect 38328 16512 38548 18968
rect 44320 18918 44570 18936
rect 41318 18868 41568 18892
rect 41318 18658 41332 18868
rect 41542 18658 41568 18868
rect 44320 18708 44332 18918
rect 44542 18708 44570 18918
rect 47318 18916 47332 19126
rect 47542 18916 47568 19126
rect 53520 19038 53770 19064
rect 47318 18886 47568 18916
rect 50500 19006 50750 19022
rect 44320 18678 44570 18708
rect 41318 18634 41568 18658
rect 41328 16456 41548 18634
rect 44328 16424 44548 18678
rect 47328 17632 47548 18886
rect 50500 18796 50520 19006
rect 50730 18796 50750 19006
rect 53520 18828 53542 19038
rect 53752 18828 53770 19038
rect 56594 18948 56620 19158
rect 56830 18948 56844 19158
rect 174366 19130 174586 19136
rect 75052 19026 75346 19044
rect 108900 19028 109120 19032
rect 68554 18952 68764 18956
rect 56594 18920 56844 18948
rect 68550 18948 69258 18952
rect 53520 18806 53770 18828
rect 50500 18764 50750 18796
rect 47328 17412 47734 17632
rect 47514 16506 47734 17412
rect 50516 16474 50736 18764
rect 53536 17810 53756 18806
rect 53536 17590 53888 17810
rect 53668 16506 53888 17590
rect 56614 16444 56834 18920
rect 59608 18866 59858 18886
rect 65736 18876 66010 18892
rect 59608 18862 60000 18866
rect 59608 18652 59634 18862
rect 59844 18652 60000 18862
rect 59608 18628 60000 18652
rect 59780 16494 60000 18628
rect 62620 18790 62870 18802
rect 62620 18786 62996 18790
rect 62620 18576 62636 18786
rect 62846 18576 62996 18786
rect 64256 18760 64576 18766
rect 62620 18544 62996 18576
rect 62776 16468 62996 18544
rect 64252 18444 64256 18754
rect 64576 18444 64580 18754
rect 65736 18666 65746 18876
rect 65956 18666 66010 18876
rect 68550 18738 68554 18948
rect 68764 18738 69258 18948
rect 75052 18816 75082 19026
rect 75292 18816 75346 19026
rect 96452 18870 96672 18876
rect 90412 18832 90632 18838
rect 75052 18782 75346 18816
rect 68550 18732 69258 18738
rect 68554 18728 68764 18732
rect 65736 18610 66010 18666
rect 64256 18434 64576 18440
rect 65946 16498 66002 18610
rect 69038 16506 69258 18732
rect 71928 18520 72148 18524
rect 71924 18310 71932 18520
rect 72142 18310 72152 18520
rect 71928 17006 72148 18310
rect 71928 16786 72278 17006
rect 72058 16506 72278 16786
rect 75078 16416 75298 18782
rect 81190 18706 81410 18710
rect 81186 18496 81194 18706
rect 81404 18496 81414 18706
rect 90408 18622 90416 18832
rect 90626 18622 90636 18832
rect 93556 18788 93776 18794
rect 78102 18082 78312 18086
rect 78098 18076 78318 18082
rect 78098 17866 78102 18076
rect 78312 17866 78318 18076
rect 78098 17154 78318 17866
rect 78098 16934 78452 17154
rect 78232 16492 78452 16934
rect 81190 16478 81410 18496
rect 87334 18310 87554 18314
rect 87330 18100 87340 18310
rect 87550 18100 87558 18310
rect 84274 17980 84494 17984
rect 84270 17770 84278 17980
rect 84488 17770 84498 17980
rect 84274 16492 84494 17770
rect 87334 16380 87554 18100
rect 90412 16440 90632 18622
rect 93552 18578 93560 18788
rect 93770 18578 93780 18788
rect 96448 18660 96458 18870
rect 96668 18660 96676 18870
rect 108896 18818 108906 19028
rect 109116 18818 109124 19028
rect 157842 18992 158062 18998
rect 114952 18980 115172 18984
rect 111948 18930 112168 18936
rect 105674 18750 105894 18756
rect 102710 18736 102930 18740
rect 93556 16448 93776 18578
rect 96452 17026 96672 18660
rect 102706 18526 102716 18736
rect 102926 18526 102934 18736
rect 105670 18540 105680 18750
rect 105890 18540 105898 18750
rect 99602 18502 99812 18506
rect 99596 18496 99816 18502
rect 99596 18286 99602 18496
rect 99812 18286 99816 18496
rect 96452 16806 96814 17026
rect 96594 16478 96814 16806
rect 99596 16514 99816 18286
rect 102710 16410 102930 18526
rect 105674 16996 105894 18540
rect 105674 16776 106014 16996
rect 105794 16462 106014 16776
rect 108900 16454 109120 18818
rect 111944 18720 111952 18930
rect 112162 18720 112172 18930
rect 114948 18770 114958 18980
rect 115168 18770 115176 18980
rect 117960 18972 118202 18992
rect 111948 16514 112168 18720
rect 114952 16452 115172 18770
rect 117960 18762 117972 18972
rect 118182 18762 118202 18972
rect 127240 18938 127460 18942
rect 117960 18746 118202 18762
rect 121128 18860 121382 18878
rect 117968 17904 118188 18746
rect 121128 18650 121154 18860
rect 121364 18650 121382 18860
rect 124118 18852 124338 18860
rect 124114 18842 124118 18846
rect 121678 18760 121998 18766
rect 121128 18614 121382 18650
rect 117968 17684 118368 17904
rect 118148 16482 118368 17684
rect 121150 16460 121370 18614
rect 121674 18444 121678 18754
rect 121998 18444 122002 18754
rect 124108 18632 124118 18842
rect 124338 18842 124342 18846
rect 124338 18632 124346 18842
rect 127236 18728 127246 18938
rect 127456 18728 127464 18938
rect 133412 18866 133632 18876
rect 133408 18856 133412 18862
rect 130250 18808 130470 18814
rect 121678 18434 121998 18440
rect 124118 16552 124338 18632
rect 127240 16460 127460 18728
rect 130246 18598 130254 18808
rect 130464 18598 130474 18808
rect 133402 18646 133412 18856
rect 133632 18856 133636 18862
rect 133632 18646 133640 18856
rect 154792 18854 155012 18858
rect 145578 18838 145798 18844
rect 148754 18838 148974 18844
rect 142598 18664 142818 18668
rect 130250 16476 130470 18598
rect 133412 16460 133632 18646
rect 139552 18596 139772 18600
rect 139548 18386 139556 18596
rect 139766 18386 139776 18596
rect 142594 18454 142604 18664
rect 142814 18454 142822 18664
rect 145574 18628 145582 18838
rect 145792 18628 145802 18838
rect 148750 18628 148758 18838
rect 148968 18628 148978 18838
rect 151772 18770 151992 18774
rect 136466 18236 136686 18242
rect 136462 18026 136472 18236
rect 136682 18026 136690 18236
rect 136466 16400 136686 18026
rect 139552 16484 139772 18386
rect 142598 16468 142818 18454
rect 145578 16946 145798 18628
rect 145578 16726 145918 16946
rect 145698 16452 145918 16726
rect 148754 16406 148974 18628
rect 151768 18560 151776 18770
rect 151986 18560 151996 18770
rect 154788 18644 154796 18854
rect 155006 18644 155016 18854
rect 157838 18782 157848 18992
rect 158058 18782 158066 18992
rect 174362 18920 174370 19130
rect 174580 18920 174590 19130
rect 305384 19094 305604 19100
rect 290332 18956 290542 18960
rect 290328 18950 293618 18956
rect 229658 18934 229878 18940
rect 151772 16372 151992 18560
rect 154792 17614 155012 18644
rect 154792 17394 155166 17614
rect 154946 16464 155166 17394
rect 157842 17038 158062 18782
rect 167548 18760 167868 18766
rect 160886 18754 161106 18758
rect 160882 18544 160890 18754
rect 161100 18544 161110 18754
rect 160886 17192 161106 18544
rect 163242 18460 163452 18464
rect 163238 18454 164318 18460
rect 163238 18244 163242 18454
rect 163452 18244 164318 18454
rect 167544 18444 167548 18754
rect 167868 18444 167872 18754
rect 173066 18484 173336 18534
rect 167548 18434 167868 18440
rect 163238 18240 164318 18244
rect 163242 18236 163452 18240
rect 164098 17688 164318 18240
rect 173066 18274 173086 18484
rect 173296 18274 173336 18484
rect 173066 18238 173336 18274
rect 165932 18174 166142 18178
rect 165928 18170 167322 18174
rect 165928 17960 165932 18170
rect 166142 17960 167322 18170
rect 165928 17954 167322 17960
rect 165932 17950 166142 17954
rect 164052 17332 164318 17688
rect 157842 16818 158224 17038
rect 160886 16972 161244 17192
rect 158004 16494 158224 16818
rect 161024 16540 161244 16972
rect 164052 16440 164272 17332
rect 167102 16440 167322 17954
rect 173082 17606 173302 18238
rect 168868 17422 169078 17426
rect 168862 17416 170482 17422
rect 168862 17206 168868 17416
rect 169078 17206 170482 17416
rect 173082 17386 173510 17606
rect 168862 17202 170482 17206
rect 168868 17198 169078 17202
rect 170262 16502 170482 17202
rect 173290 16464 173510 17386
rect 174366 17560 174586 18920
rect 176310 18812 176564 18822
rect 176310 18808 179212 18812
rect 176310 18598 176332 18808
rect 176542 18598 179212 18808
rect 180548 18760 180868 18766
rect 189548 18760 189868 18766
rect 198548 18760 198868 18766
rect 204548 18760 204868 18766
rect 211548 18760 211868 18766
rect 223548 18760 223868 18766
rect 176310 18592 179212 18598
rect 176310 18578 176564 18592
rect 174366 17340 176668 17560
rect 176448 16456 176668 17340
rect 178992 17290 179212 18592
rect 180544 18444 180548 18754
rect 180868 18444 180872 18754
rect 189544 18444 189548 18754
rect 189868 18444 189872 18754
rect 198544 18444 198548 18754
rect 198868 18444 198872 18754
rect 204544 18444 204548 18754
rect 204868 18444 204872 18754
rect 206332 18456 206542 18460
rect 206328 18450 208700 18456
rect 180548 18434 180868 18440
rect 189548 18434 189868 18440
rect 198548 18434 198868 18440
rect 204548 18434 204868 18440
rect 206328 18240 206332 18450
rect 206542 18240 208700 18450
rect 211544 18444 211548 18754
rect 211868 18444 211872 18754
rect 215332 18564 215542 18568
rect 215328 18558 219616 18564
rect 211548 18434 211868 18440
rect 215328 18348 215332 18558
rect 215542 18348 219616 18558
rect 223544 18444 223548 18754
rect 223868 18444 223872 18754
rect 229654 18724 229662 18934
rect 229872 18724 229882 18934
rect 232548 18760 232868 18766
rect 238548 18760 238868 18766
rect 250548 18760 250868 18766
rect 263948 18760 264268 18766
rect 269948 18760 270268 18766
rect 272948 18760 273268 18766
rect 275948 18760 276268 18766
rect 281948 18760 282268 18766
rect 285948 18760 286268 18766
rect 223548 18434 223868 18440
rect 227194 18424 227414 18428
rect 215328 18344 219616 18348
rect 215332 18340 215542 18344
rect 206328 18236 208700 18240
rect 206332 18232 206542 18236
rect 185332 18036 185542 18040
rect 185328 18032 188126 18036
rect 182472 17854 182692 17860
rect 182468 17644 182478 17854
rect 182688 17644 182696 17854
rect 185328 17822 185332 18032
rect 185542 17822 188126 18032
rect 200914 17952 201134 17956
rect 196792 17924 197012 17930
rect 185328 17816 188126 17822
rect 185332 17812 185542 17816
rect 178992 17070 179704 17290
rect 179484 16494 179704 17070
rect 182472 16480 182692 17644
rect 184014 17152 184224 17156
rect 184010 17148 185874 17152
rect 184010 16938 184014 17148
rect 184224 16938 185874 17148
rect 184010 16932 185874 16938
rect 184014 16928 184224 16932
rect 185654 16456 185874 16932
rect 187906 16884 188126 17816
rect 196788 17714 196798 17924
rect 197008 17714 197016 17924
rect 200910 17742 200920 17952
rect 201130 17742 201138 17952
rect 206998 17746 207218 17752
rect 188332 17660 188542 17664
rect 188328 17654 191876 17660
rect 188328 17444 188332 17654
rect 188542 17444 191876 17654
rect 188328 17440 191876 17444
rect 188332 17436 188542 17440
rect 187906 16664 188840 16884
rect 188620 16448 188840 16664
rect 191656 16486 191876 17440
rect 193470 17020 193680 17024
rect 196792 17020 197012 17714
rect 193464 17014 195050 17020
rect 193464 16804 193470 17014
rect 193680 16804 195050 17014
rect 193464 16800 195050 16804
rect 196792 16800 198136 17020
rect 193470 16796 193680 16800
rect 194830 16452 195050 16800
rect 197916 16380 198136 16800
rect 200914 16470 201134 17742
rect 206994 17536 207004 17746
rect 207214 17536 207222 17746
rect 202008 16894 202218 16898
rect 202002 16890 204256 16894
rect 202002 16680 202008 16890
rect 202218 16680 204256 16890
rect 202002 16674 204256 16680
rect 202008 16670 202218 16674
rect 204036 16514 204256 16674
rect 206998 16522 207218 17536
rect 208480 17090 208700 18236
rect 213154 18094 213374 18098
rect 213150 17884 213160 18094
rect 213370 17884 213378 18094
rect 208480 16870 210430 17090
rect 210210 16506 210430 16870
rect 213154 16434 213374 17884
rect 213908 17270 214118 17274
rect 213904 17264 216496 17270
rect 213904 17054 213908 17264
rect 214118 17054 216496 17264
rect 213904 17050 216496 17054
rect 213908 17046 214118 17050
rect 216276 16372 216496 17050
rect 219396 16434 219616 18344
rect 227190 18214 227198 18424
rect 227408 18214 227418 18424
rect 221332 17712 221542 17716
rect 221328 17706 225720 17712
rect 221328 17496 221332 17706
rect 221542 17496 225720 17706
rect 221328 17492 225720 17496
rect 221332 17488 221542 17492
rect 220692 17228 220902 17232
rect 220688 17224 222682 17228
rect 220688 17014 220692 17224
rect 220902 17014 222682 17224
rect 220688 17008 222682 17014
rect 220692 17004 220902 17008
rect 222462 16426 222682 17008
rect 225500 16498 225720 17492
rect 227194 17524 227414 18214
rect 227194 17304 228838 17524
rect 228618 16480 228838 17304
rect 229658 17434 229878 18724
rect 232544 18444 232548 18754
rect 232868 18444 232872 18754
rect 233332 18690 233542 18694
rect 233328 18684 237602 18690
rect 233328 18474 233332 18684
rect 233542 18680 237602 18684
rect 233542 18474 237948 18680
rect 233328 18470 237948 18474
rect 233332 18466 233542 18470
rect 237356 18460 237948 18470
rect 232548 18434 232868 18440
rect 234650 18298 235040 18304
rect 234646 18088 234654 18298
rect 234864 18088 235040 18298
rect 234650 18084 235040 18088
rect 229658 17214 231876 17434
rect 231656 16542 231876 17214
rect 234820 16506 235040 18084
rect 237728 17960 237948 18460
rect 238544 18444 238548 18754
rect 238868 18444 238872 18754
rect 242332 18570 242542 18574
rect 242328 18566 245088 18570
rect 241672 18530 241892 18534
rect 238548 18434 238868 18440
rect 241668 18320 241676 18530
rect 241886 18320 241896 18530
rect 242328 18356 242332 18566
rect 242542 18356 245088 18566
rect 250544 18444 250548 18754
rect 250868 18444 250872 18754
rect 254332 18700 254542 18704
rect 254328 18696 257536 18700
rect 253924 18504 254144 18510
rect 250548 18434 250868 18440
rect 242328 18350 245088 18356
rect 242332 18346 242542 18350
rect 240916 18010 241136 18016
rect 237706 17778 237948 17960
rect 240912 17800 240920 18010
rect 241130 17800 241140 18010
rect 237706 16426 237926 17778
rect 240916 16484 241136 17800
rect 241672 17214 241892 18320
rect 241672 16994 244150 17214
rect 243930 16320 244150 16994
rect 244868 16986 245088 18350
rect 253920 18294 253930 18504
rect 254140 18294 254148 18504
rect 254328 18486 254332 18696
rect 254542 18486 257536 18696
rect 254328 18480 257536 18486
rect 254332 18476 254542 18480
rect 249644 17860 249924 17882
rect 249644 17856 253346 17860
rect 249644 17646 249672 17856
rect 249882 17646 253346 17856
rect 249644 17640 253346 17646
rect 249644 17622 249924 17640
rect 248716 17078 248926 17082
rect 248710 17072 250268 17078
rect 244868 16766 247272 16986
rect 248710 16862 248716 17072
rect 248926 16862 250268 17072
rect 248710 16858 250268 16862
rect 248716 16854 248926 16858
rect 247052 16520 247272 16766
rect 250048 16420 250268 16858
rect 253126 16520 253346 17640
rect 253924 17354 254144 18294
rect 257316 17358 257536 18480
rect 263944 18444 263948 18754
rect 264268 18444 264272 18754
rect 269032 18556 269252 18560
rect 263948 18434 264268 18440
rect 269028 18346 269036 18556
rect 269246 18346 269256 18556
rect 269944 18444 269948 18754
rect 270268 18444 270272 18754
rect 272944 18444 272948 18754
rect 273268 18444 273272 18754
rect 275944 18444 275948 18754
rect 276268 18444 276272 18754
rect 279676 18694 279896 18698
rect 279672 18484 279680 18694
rect 279890 18484 279900 18694
rect 269948 18434 270268 18440
rect 272948 18434 273268 18440
rect 275948 18434 276268 18440
rect 261048 18126 261258 18130
rect 261044 18120 265648 18126
rect 261044 17910 261048 18120
rect 261258 17910 265648 18120
rect 265874 17964 266084 17968
rect 261044 17906 265648 17910
rect 261048 17902 261258 17906
rect 259366 17358 259586 17386
rect 253924 17134 256416 17354
rect 257316 17138 259608 17358
rect 260058 17246 260268 17250
rect 260052 17242 262606 17246
rect 256196 16438 256416 17134
rect 259366 16506 259586 17138
rect 260052 17032 260058 17242
rect 260268 17032 262606 17242
rect 260052 17026 262606 17032
rect 260058 17022 260268 17026
rect 262386 16480 262606 17026
rect 265428 16438 265648 17906
rect 265870 17958 267378 17964
rect 265870 17748 265874 17958
rect 266084 17748 267378 17958
rect 265870 17744 267378 17748
rect 265874 17740 266084 17744
rect 267158 17370 267378 17744
rect 267158 17150 268752 17370
rect 267158 17148 267378 17150
rect 268532 16388 268752 17150
rect 269032 17090 269252 18346
rect 269332 18268 269542 18272
rect 269328 18264 274812 18268
rect 269328 18054 269332 18264
rect 269542 18054 274812 18264
rect 278878 18202 279098 18206
rect 269328 18048 274812 18054
rect 269332 18044 269542 18048
rect 269032 16870 271810 17090
rect 271590 16406 271810 16870
rect 274592 16502 274812 18048
rect 278874 17992 278882 18202
rect 279092 17992 279102 18202
rect 277692 17578 277912 17582
rect 277688 17368 277698 17578
rect 277908 17368 277916 17578
rect 277692 16482 277912 17368
rect 278878 17146 279098 17992
rect 279676 17916 279896 18484
rect 281944 18444 281948 18754
rect 282268 18444 282272 18754
rect 285944 18444 285948 18754
rect 286268 18444 286272 18754
rect 290328 18740 290332 18950
rect 290542 18740 293618 18950
rect 305380 18884 305390 19094
rect 305600 18884 305608 19094
rect 293948 18760 294268 18766
rect 296948 18760 297268 18766
rect 299948 18760 300268 18766
rect 302948 18760 303268 18766
rect 290328 18736 293618 18740
rect 290332 18732 290542 18736
rect 281948 18434 282268 18440
rect 285948 18434 286268 18440
rect 292406 18222 292626 18228
rect 284332 18138 284542 18142
rect 284328 18132 287822 18138
rect 284328 17922 284332 18132
rect 284542 17922 287822 18132
rect 292402 18012 292412 18222
rect 292622 18012 292630 18222
rect 284328 17918 287822 17922
rect 279676 17696 284112 17916
rect 284332 17914 284542 17918
rect 278878 16926 280970 17146
rect 280750 16364 280970 16926
rect 283892 16454 284112 17696
rect 286928 17508 287148 17512
rect 286924 17298 286934 17508
rect 287144 17298 287152 17508
rect 286928 16446 287148 17298
rect 287602 16980 287822 17918
rect 287602 16760 290186 16980
rect 289966 16488 290186 16760
rect 292406 16924 292626 18012
rect 293398 17354 293618 18736
rect 293944 18444 293948 18754
rect 294268 18444 294272 18754
rect 296944 18444 296948 18754
rect 297268 18444 297272 18754
rect 299944 18444 299948 18754
rect 300268 18444 300272 18754
rect 302944 18444 302948 18754
rect 303268 18444 303272 18754
rect 293948 18434 294268 18440
rect 296948 18434 297268 18440
rect 299948 18434 300268 18440
rect 302948 18434 303268 18440
rect 299258 17718 299478 17724
rect 299254 17508 299262 17718
rect 299472 17508 299482 17718
rect 293398 17134 296406 17354
rect 292406 16704 293306 16924
rect 293086 16446 293306 16704
rect 296186 16460 296406 17134
rect 299258 16890 299478 17508
rect 300256 17106 300466 17110
rect 299146 16670 299478 16890
rect 300250 17100 302500 17106
rect 300250 16890 300256 17100
rect 300466 16890 302500 17100
rect 300250 16886 302500 16890
rect 300256 16882 300466 16886
rect 299146 16398 299366 16670
rect 302280 16510 302500 16886
rect 305384 16504 305604 18884
rect 302946 16416 303268 16424
rect 302940 16094 302946 16416
rect 303268 16094 303274 16416
rect 302946 16084 303268 16094
rect 18088 15712 18408 15720
rect 3664 15694 3984 15702
rect 108 15588 308 15596
rect 102 15388 108 15588
rect 308 15388 314 15588
rect 108 15378 308 15388
rect 3658 15374 3664 15694
rect 3984 15374 3990 15694
rect 18082 15392 18088 15712
rect 18408 15392 18414 15712
rect 121678 15710 121998 15718
rect 167548 15712 167868 15720
rect 180548 15712 180868 15720
rect 189548 15712 189868 15720
rect 198548 15712 198868 15720
rect 204548 15712 204868 15720
rect 211548 15712 211868 15720
rect 223548 15712 223868 15720
rect 232548 15712 232868 15720
rect 238548 15712 238868 15720
rect 250548 15712 250868 15720
rect 263948 15712 264268 15720
rect 269948 15712 270268 15720
rect 272948 15712 273268 15720
rect 275948 15712 276268 15720
rect 281948 15712 282268 15720
rect 285948 15712 286268 15720
rect 293948 15712 294268 15720
rect 296948 15712 297268 15720
rect 299948 15712 300268 15720
rect 302948 15712 303268 15720
rect 64256 15696 64576 15704
rect 32914 15688 33234 15696
rect 18088 15382 18408 15392
rect 3664 15364 3984 15374
rect 32908 15368 32914 15688
rect 33234 15368 33240 15688
rect 64250 15376 64256 15696
rect 64576 15376 64582 15696
rect 121672 15390 121678 15710
rect 121998 15390 122004 15710
rect 167542 15392 167548 15712
rect 167868 15392 167874 15712
rect 180542 15392 180548 15712
rect 180868 15392 180874 15712
rect 189542 15392 189548 15712
rect 189868 15392 189874 15712
rect 198542 15392 198548 15712
rect 198868 15392 198874 15712
rect 204542 15392 204548 15712
rect 204868 15392 204874 15712
rect 211542 15392 211548 15712
rect 211868 15392 211874 15712
rect 223542 15392 223548 15712
rect 223868 15392 223874 15712
rect 232542 15392 232548 15712
rect 232868 15392 232874 15712
rect 238542 15392 238548 15712
rect 238868 15392 238874 15712
rect 250542 15392 250548 15712
rect 250868 15392 250874 15712
rect 263942 15392 263948 15712
rect 264268 15392 264274 15712
rect 269942 15392 269948 15712
rect 270268 15392 270274 15712
rect 272942 15392 272948 15712
rect 273268 15392 273274 15712
rect 275942 15392 275948 15712
rect 276268 15392 276274 15712
rect 281942 15392 281948 15712
rect 282268 15392 282274 15712
rect 285942 15392 285948 15712
rect 286268 15392 286274 15712
rect 293942 15392 293948 15712
rect 294268 15392 294274 15712
rect 296942 15392 296948 15712
rect 297268 15392 297274 15712
rect 299942 15392 299948 15712
rect 300268 15392 300274 15712
rect 302942 15392 302948 15712
rect 303268 15392 303274 15712
rect 121678 15380 121998 15390
rect 167548 15382 167868 15392
rect 180548 15382 180868 15392
rect 189548 15382 189868 15392
rect 198548 15382 198868 15392
rect 204548 15382 204868 15392
rect 211548 15382 211868 15392
rect 223548 15382 223868 15392
rect 232548 15382 232868 15392
rect 238548 15382 238868 15392
rect 250548 15382 250868 15392
rect 263948 15382 264268 15392
rect 269948 15382 270268 15392
rect 272948 15382 273268 15392
rect 275948 15382 276268 15392
rect 281948 15382 282268 15392
rect 285948 15382 286268 15392
rect 293948 15382 294268 15392
rect 296948 15382 297268 15392
rect 299948 15382 300268 15392
rect 302948 15382 303268 15392
rect 32914 15358 33234 15368
rect 64256 15366 64576 15376
<< via2 >>
rect 302508 324332 302708 324532
rect 303930 321042 304240 321352
rect 108 319722 308 319922
rect 303930 318042 304240 318352
rect 108 316722 308 316922
rect 303930 315042 304240 315352
rect 108 313722 308 313922
rect 303930 312042 304240 312352
rect 108 310722 308 310922
rect 303930 309042 304240 309352
rect 108 307722 308 307922
rect 303930 306042 304240 306352
rect 108 304722 308 304922
rect 303930 303042 304240 303352
rect 108 301722 308 301922
rect 303930 300042 304240 300352
rect 108 298722 308 298922
rect 303930 297042 304240 297352
rect 108 295722 308 295922
rect 303930 294042 304240 294352
rect 108 292722 308 292922
rect 303930 291042 304240 291352
rect 108 289722 308 289922
rect 303930 288042 304240 288352
rect 108 286722 308 286922
rect 303930 285042 304240 285352
rect 108 283722 308 283922
rect 303930 282042 304240 282352
rect 108 280722 308 280922
rect 303930 279042 304240 279352
rect 108 277722 308 277922
rect 303930 276042 304240 276352
rect 108 274722 308 274922
rect 303930 273042 304240 273352
rect 108 271722 308 271922
rect 303930 270042 304240 270352
rect 108 268722 308 268922
rect 303930 267042 304240 267352
rect 108 265722 308 265922
rect 303930 264042 304240 264352
rect 108 262722 308 262922
rect 303930 261042 304240 261352
rect 108 259722 308 259922
rect 303930 258042 304240 258352
rect 108 256722 308 256922
rect 303930 255042 304240 255352
rect 108 253722 308 253922
rect 303930 252042 304240 252352
rect 108 250722 308 250922
rect 303930 249042 304240 249352
rect 108 247722 308 247922
rect 303930 246042 304240 246352
rect 108 244722 308 244922
rect 303930 243042 304240 243352
rect 108 241722 308 241922
rect 303930 240042 304240 240352
rect 108 238722 308 238922
rect 303930 237042 304240 237352
rect 108 235722 308 235922
rect 303930 234042 304240 234352
rect 108 232722 308 232922
rect 303930 231042 304240 231352
rect 108 229722 308 229922
rect 303930 228042 304240 228352
rect 108 226722 308 226922
rect 303930 225042 304240 225352
rect 108 223722 308 223922
rect 303930 222042 304240 222352
rect 108 220722 308 220922
rect 303930 219042 304240 219352
rect 108 217722 308 217922
rect 303930 216042 304240 216352
rect 108 214722 308 214922
rect 303930 213042 304240 213352
rect 108 211722 308 211922
rect 303930 210042 304240 210352
rect 108 208722 308 208922
rect 303930 207042 304240 207352
rect 108 205722 308 205922
rect 303930 204042 304240 204352
rect 108 202722 308 202922
rect 303930 201042 304240 201352
rect 108 199722 308 199922
rect 303930 198042 304240 198352
rect 108 196722 308 196922
rect 303930 195042 304240 195352
rect 108 193722 308 193922
rect 303930 192042 304240 192352
rect 108 190722 308 190922
rect 303930 189042 304240 189352
rect 108 187722 308 187922
rect 303930 186042 304240 186352
rect 108 184722 308 184922
rect 303930 183042 304240 183352
rect 108 181722 308 181922
rect 303930 180042 304240 180352
rect 108 178722 308 178922
rect 303930 177042 304240 177352
rect 108 175722 308 175922
rect 303930 174042 304240 174352
rect 108 172722 308 172922
rect 303930 171042 304240 171352
rect 108 169722 308 169922
rect 303930 168042 304240 168352
rect 108 166722 308 166922
rect 303930 165042 304240 165352
rect 108 163722 308 163922
rect 303930 162042 304240 162352
rect 108 160722 308 160922
rect 303930 159042 304240 159352
rect 108 157722 308 157922
rect 303930 156042 304240 156352
rect 108 154722 308 154922
rect 303930 153042 304240 153352
rect 108 151722 308 151922
rect 303930 150042 304240 150352
rect 108 148722 308 148922
rect 303930 147042 304240 147352
rect 108 145722 308 145922
rect 303930 144042 304240 144352
rect 108 142722 308 142922
rect 303930 141042 304240 141352
rect 108 139722 308 139922
rect 303930 138042 304240 138352
rect 108 136722 308 136922
rect 303930 135042 304240 135352
rect 108 133722 308 133922
rect 303930 132042 304240 132352
rect 108 130722 308 130922
rect 303930 129042 304240 129352
rect 108 127722 308 127922
rect 303930 126042 304240 126352
rect 108 124722 308 124922
rect 303930 123042 304240 123352
rect 108 121722 308 121922
rect 303930 120042 304240 120352
rect 108 118722 308 118922
rect 303930 117042 304240 117352
rect 108 115722 308 115922
rect 303930 114042 304240 114352
rect 108 112722 308 112922
rect 303930 111042 304240 111352
rect 108 109722 308 109922
rect 303930 108042 304240 108352
rect 108 106722 308 106922
rect 303930 105042 304240 105352
rect 108 103722 308 103922
rect 303930 102042 304240 102352
rect 108 100722 308 100922
rect 303930 99042 304240 99352
rect 108 97722 308 97922
rect 303930 96042 304240 96352
rect 108 94722 308 94922
rect 303930 93042 304240 93352
rect 108 91722 308 91922
rect 303930 90042 304240 90352
rect 108 88722 308 88922
rect 303930 87042 304240 87352
rect 108 85722 308 85922
rect 303930 84042 304240 84352
rect 108 82722 308 82922
rect 303930 81042 304240 81352
rect 108 79722 308 79922
rect 303930 78042 304240 78352
rect 108 76722 308 76922
rect 303930 75042 304240 75352
rect 108 73722 308 73922
rect 303930 72042 304240 72352
rect 108 70722 308 70922
rect 303930 69042 304240 69352
rect 108 67722 308 67922
rect 303930 66042 304240 66352
rect 108 64722 308 64922
rect 303930 63042 304240 63352
rect 108 61722 308 61922
rect 303930 60042 304240 60352
rect 108 58722 308 58922
rect 303930 57042 304240 57352
rect 108 55722 308 55922
rect 303930 54042 304240 54352
rect 108 52722 308 52922
rect 303930 51042 304240 51352
rect 108 49722 308 49922
rect 303930 48042 304240 48352
rect 108 46722 308 46922
rect 303930 45042 304240 45352
rect 108 43722 308 43922
rect 303930 42042 304240 42352
rect 108 40722 308 40922
rect 303930 39042 304240 39352
rect 108 37722 308 37922
rect 303930 36042 304240 36352
rect 108 34722 308 34922
rect 303930 33042 304240 33352
rect 108 31722 308 31922
rect 303930 30042 304240 30352
rect 108 28722 308 28922
rect 303930 27042 304240 27352
rect 108 25722 308 25922
rect 303930 24042 304240 24352
rect 108 22722 308 22922
rect 303930 21042 304240 21352
rect 19874 18978 20084 19188
rect 3668 18444 3978 18754
rect 5332 18570 5542 18780
rect 7486 18676 7696 18886
rect 2332 18224 2542 18434
rect -6198 17746 -5998 17946
rect 10716 18620 10926 18830
rect 13806 18714 14016 18924
rect 16916 18602 17126 18812
rect 18092 18444 18402 18754
rect 25948 18796 26158 19006
rect 29084 18842 29304 19062
rect 22902 18444 23112 18654
rect 32332 18772 32542 18982
rect 35332 18840 35542 19050
rect 38332 19004 38542 19214
rect 32918 18444 33228 18754
rect 41332 18658 41542 18868
rect 44332 18708 44542 18918
rect 47332 18916 47542 19126
rect 50520 18796 50730 19006
rect 53542 18828 53752 19038
rect 56620 18948 56830 19158
rect 59634 18652 59844 18862
rect 62636 18576 62846 18786
rect 64260 18444 64570 18754
rect 65746 18666 65956 18876
rect 68554 18738 68764 18948
rect 75082 18816 75292 19026
rect 71932 18310 72142 18520
rect 81194 18496 81404 18706
rect 90416 18622 90626 18832
rect 78102 17866 78312 18076
rect 87340 18100 87550 18310
rect 84278 17770 84488 17980
rect 93560 18578 93770 18788
rect 96458 18660 96668 18870
rect 108906 18818 109116 19028
rect 102716 18526 102926 18736
rect 105680 18540 105890 18750
rect 99602 18286 99812 18496
rect 111952 18720 112162 18930
rect 114958 18770 115168 18980
rect 117972 18762 118182 18972
rect 121154 18650 121364 18860
rect 121682 18444 121992 18754
rect 124118 18632 124338 18852
rect 127246 18728 127456 18938
rect 130254 18598 130464 18808
rect 133412 18646 133632 18866
rect 139556 18386 139766 18596
rect 142604 18454 142814 18664
rect 145582 18628 145792 18838
rect 148758 18628 148968 18838
rect 136472 18026 136682 18236
rect 151776 18560 151986 18770
rect 154796 18644 155006 18854
rect 157848 18782 158058 18992
rect 174370 18920 174580 19130
rect 160890 18544 161100 18754
rect 163242 18244 163452 18454
rect 167552 18444 167862 18754
rect 173086 18274 173296 18484
rect 165932 17960 166142 18170
rect 168868 17206 169078 17416
rect 176332 18598 176542 18808
rect 180552 18444 180862 18754
rect 189552 18444 189862 18754
rect 198552 18444 198862 18754
rect 204552 18444 204862 18754
rect 206332 18240 206542 18450
rect 211552 18444 211862 18754
rect 215332 18348 215542 18558
rect 223552 18444 223862 18754
rect 229662 18724 229872 18934
rect 182478 17644 182688 17854
rect 185332 17822 185542 18032
rect 184014 16938 184224 17148
rect 196798 17714 197008 17924
rect 200920 17742 201130 17952
rect 188332 17444 188542 17654
rect 193470 16804 193680 17014
rect 207004 17536 207214 17746
rect 202008 16680 202218 16890
rect 213160 17884 213370 18094
rect 213908 17054 214118 17264
rect 227198 18214 227408 18424
rect 221332 17496 221542 17706
rect 220692 17014 220902 17224
rect 232552 18444 232862 18754
rect 233332 18474 233542 18684
rect 234654 18088 234864 18298
rect 238552 18444 238862 18754
rect 241676 18320 241886 18530
rect 242332 18356 242542 18566
rect 250552 18444 250862 18754
rect 240920 17800 241130 18010
rect 253930 18294 254140 18504
rect 254332 18486 254542 18696
rect 249672 17646 249882 17856
rect 248716 16862 248926 17072
rect 263952 18444 264262 18754
rect 269036 18346 269246 18556
rect 269952 18444 270262 18754
rect 272952 18444 273262 18754
rect 275952 18444 276262 18754
rect 279680 18484 279890 18694
rect 261048 17910 261258 18120
rect 260058 17032 260268 17242
rect 265874 17748 266084 17958
rect 269332 18054 269542 18264
rect 278882 17992 279092 18202
rect 277698 17368 277908 17578
rect 281952 18444 282262 18754
rect 285952 18444 286262 18754
rect 290332 18740 290542 18950
rect 305390 18884 305600 19094
rect 284332 17922 284542 18132
rect 292412 18012 292622 18222
rect 286934 17298 287144 17508
rect 293952 18444 294262 18754
rect 296952 18444 297262 18754
rect 299952 18444 300262 18754
rect 302952 18444 303262 18754
rect 299262 17508 299472 17718
rect 300256 16890 300466 17100
rect 302946 16094 303268 16416
rect 108 15388 308 15588
rect 3664 15374 3984 15694
rect 18088 15392 18408 15712
rect 32914 15368 33234 15688
rect 64256 15376 64576 15696
rect 121678 15390 121998 15710
rect 167548 15392 167868 15712
rect 180548 15392 180868 15712
rect 189548 15392 189868 15712
rect 198548 15392 198868 15712
rect 204548 15392 204868 15712
rect 211548 15392 211868 15712
rect 223548 15392 223868 15712
rect 232548 15392 232868 15712
rect 238548 15392 238868 15712
rect 250548 15392 250868 15712
rect 263948 15392 264268 15712
rect 269948 15392 270268 15712
rect 272948 15392 273268 15712
rect 275948 15392 276268 15712
rect 281948 15392 282268 15712
rect 285948 15392 286268 15712
rect 293948 15392 294268 15712
rect 296948 15392 297268 15712
rect 299948 15392 300268 15712
rect 302948 15392 303268 15712
<< metal3 >>
rect -13040 323508 -12920 323868
rect 908 322280 998 327366
rect 302502 324538 302712 324544
rect 302502 324332 302508 324338
rect 302708 324332 302712 324338
rect 302502 324328 302712 324332
rect 303926 321358 304244 321362
rect 303926 321356 304246 321358
rect 304244 321038 304246 321356
rect 303926 321032 304244 321038
rect 102 319922 312 319926
rect -2012 319722 -2006 319922
rect -1806 319722 108 319922
rect 308 319722 312 319922
rect 102 319716 312 319722
rect 303926 318358 304244 318362
rect 303926 318356 304246 318358
rect 304244 318038 304246 318356
rect 303926 318032 304244 318038
rect 102 316922 312 316926
rect -2012 316722 -2006 316922
rect -1806 316722 108 316922
rect 308 316722 312 316922
rect 102 316716 312 316722
rect 303926 315358 304244 315362
rect 303926 315356 304246 315358
rect 304244 315038 304246 315356
rect 303926 315032 304244 315038
rect 102 313922 312 313926
rect -2012 313722 -2006 313922
rect -1806 313722 108 313922
rect 308 313722 312 313922
rect 102 313716 312 313722
rect 303926 312358 304244 312362
rect 303926 312356 304246 312358
rect 304244 312038 304246 312356
rect 303926 312032 304244 312038
rect 102 310922 312 310926
rect -2012 310722 -2006 310922
rect -1806 310722 108 310922
rect 308 310722 312 310922
rect 102 310716 312 310722
rect 303926 309358 304244 309362
rect 303926 309356 304246 309358
rect 304244 309038 304246 309356
rect 303926 309032 304244 309038
rect 102 307922 312 307926
rect -2012 307722 -2006 307922
rect -1806 307722 108 307922
rect 308 307722 312 307922
rect 102 307716 312 307722
rect 303926 306358 304244 306362
rect 303926 306356 304246 306358
rect 304244 306038 304246 306356
rect 303926 306032 304244 306038
rect 102 304922 312 304926
rect -2012 304722 -2006 304922
rect -1806 304722 108 304922
rect 308 304722 312 304922
rect 102 304716 312 304722
rect 303926 303358 304244 303362
rect 303926 303356 304246 303358
rect 304244 303038 304246 303356
rect 303926 303032 304244 303038
rect 102 301922 312 301926
rect -2012 301722 -2006 301922
rect -1806 301722 108 301922
rect 308 301722 312 301922
rect 102 301716 312 301722
rect 303926 300358 304244 300362
rect 303926 300356 304246 300358
rect 304244 300038 304246 300356
rect 303926 300032 304244 300038
rect 102 298922 312 298926
rect -2012 298722 -2006 298922
rect -1806 298722 108 298922
rect 308 298722 312 298922
rect 102 298716 312 298722
rect 303926 297358 304244 297362
rect 303926 297356 304246 297358
rect 304244 297038 304246 297356
rect 303926 297032 304244 297038
rect 102 295922 312 295926
rect -2012 295722 -2006 295922
rect -1806 295722 108 295922
rect 308 295722 312 295922
rect 102 295716 312 295722
rect 303926 294358 304244 294362
rect 303926 294356 304246 294358
rect 304244 294038 304246 294356
rect 303926 294032 304244 294038
rect 102 292922 312 292926
rect -2012 292722 -2006 292922
rect -1806 292722 108 292922
rect 308 292722 312 292922
rect 102 292716 312 292722
rect 303926 291358 304244 291362
rect 303926 291356 304246 291358
rect 304244 291038 304246 291356
rect 303926 291032 304244 291038
rect 102 289922 312 289926
rect -2012 289722 -2006 289922
rect -1806 289722 108 289922
rect 308 289722 312 289922
rect 102 289716 312 289722
rect 303926 288358 304244 288362
rect 303926 288356 304246 288358
rect 304244 288038 304246 288356
rect 303926 288032 304244 288038
rect 102 286922 312 286926
rect -2012 286722 -2006 286922
rect -1806 286722 108 286922
rect 308 286722 312 286922
rect 102 286716 312 286722
rect 303926 285358 304244 285362
rect 303926 285356 304246 285358
rect 304244 285038 304246 285356
rect 303926 285032 304244 285038
rect 102 283922 312 283926
rect -2012 283722 -2006 283922
rect -1806 283722 108 283922
rect 308 283722 312 283922
rect 102 283716 312 283722
rect 303926 282358 304244 282362
rect 303926 282356 304246 282358
rect 304244 282038 304246 282356
rect 303926 282032 304244 282038
rect 102 280922 312 280926
rect -2012 280722 -2006 280922
rect -1806 280722 108 280922
rect 308 280722 312 280922
rect 102 280716 312 280722
rect 303926 279358 304244 279362
rect 303926 279356 304246 279358
rect 304244 279038 304246 279356
rect 303926 279032 304244 279038
rect 102 277922 312 277926
rect -2012 277722 -2006 277922
rect -1806 277722 108 277922
rect 308 277722 312 277922
rect 102 277716 312 277722
rect 303926 276358 304244 276362
rect 303926 276356 304246 276358
rect 304244 276038 304246 276356
rect 303926 276032 304244 276038
rect 102 274922 312 274926
rect -2012 274722 -2006 274922
rect -1806 274722 108 274922
rect 308 274722 312 274922
rect 102 274716 312 274722
rect 303926 273358 304244 273362
rect 303926 273356 304246 273358
rect 304244 273038 304246 273356
rect 303926 273032 304244 273038
rect 102 271922 312 271926
rect -2012 271722 -2006 271922
rect -1806 271722 108 271922
rect 308 271722 312 271922
rect 102 271716 312 271722
rect 303926 270358 304244 270362
rect 303926 270356 304246 270358
rect 304244 270038 304246 270356
rect 303926 270032 304244 270038
rect 102 268922 312 268926
rect -2012 268722 -2006 268922
rect -1806 268722 108 268922
rect 308 268722 312 268922
rect 102 268716 312 268722
rect 303926 267358 304244 267362
rect 303926 267356 304246 267358
rect 304244 267038 304246 267356
rect 303926 267032 304244 267038
rect 102 265922 312 265926
rect -2012 265722 -2006 265922
rect -1806 265722 108 265922
rect 308 265722 312 265922
rect 102 265716 312 265722
rect 303926 264358 304244 264362
rect 303926 264356 304246 264358
rect 304244 264038 304246 264356
rect 303926 264032 304244 264038
rect 102 262922 312 262926
rect -2012 262722 -2006 262922
rect -1806 262722 108 262922
rect 308 262722 312 262922
rect 102 262716 312 262722
rect 303926 261358 304244 261362
rect 303926 261356 304246 261358
rect 304244 261038 304246 261356
rect 303926 261032 304244 261038
rect 102 259922 312 259926
rect -2012 259722 -2006 259922
rect -1806 259722 108 259922
rect 308 259722 312 259922
rect 102 259716 312 259722
rect 303926 258358 304244 258362
rect 303926 258356 304246 258358
rect 304244 258038 304246 258356
rect 303926 258032 304244 258038
rect 102 256922 312 256926
rect -2012 256722 -2006 256922
rect -1806 256722 108 256922
rect 308 256722 312 256922
rect 102 256716 312 256722
rect 303926 255358 304244 255362
rect 303926 255356 304246 255358
rect 304244 255038 304246 255356
rect 303926 255032 304244 255038
rect 102 253922 312 253926
rect -2012 253722 -2006 253922
rect -1806 253722 108 253922
rect 308 253722 312 253922
rect 102 253716 312 253722
rect 303926 252358 304244 252362
rect 303926 252356 304246 252358
rect 304244 252038 304246 252356
rect 303926 252032 304244 252038
rect 102 250922 312 250926
rect -2012 250722 -2006 250922
rect -1806 250722 108 250922
rect 308 250722 312 250922
rect 102 250716 312 250722
rect 303926 249358 304244 249362
rect 303926 249356 304246 249358
rect 304244 249038 304246 249356
rect 303926 249032 304244 249038
rect 102 247922 312 247926
rect -2012 247722 -2006 247922
rect -1806 247722 108 247922
rect 308 247722 312 247922
rect 102 247716 312 247722
rect 303926 246358 304244 246362
rect 303926 246356 304246 246358
rect 304244 246038 304246 246356
rect 303926 246032 304244 246038
rect 102 244922 312 244926
rect -2012 244722 -2006 244922
rect -1806 244722 108 244922
rect 308 244722 312 244922
rect 102 244716 312 244722
rect 303926 243358 304244 243362
rect 303926 243356 304246 243358
rect 304244 243038 304246 243356
rect 303926 243032 304244 243038
rect 102 241922 312 241926
rect -2012 241722 -2006 241922
rect -1806 241722 108 241922
rect 308 241722 312 241922
rect 102 241716 312 241722
rect 303926 240358 304244 240362
rect 303926 240356 304246 240358
rect 304244 240038 304246 240356
rect 303926 240032 304244 240038
rect 102 238922 312 238926
rect -2012 238722 -2006 238922
rect -1806 238722 108 238922
rect 308 238722 312 238922
rect 102 238716 312 238722
rect 303926 237358 304244 237362
rect 303926 237356 304246 237358
rect 304244 237038 304246 237356
rect 303926 237032 304244 237038
rect 102 235922 312 235926
rect -2012 235722 -2006 235922
rect -1806 235722 108 235922
rect 308 235722 312 235922
rect 102 235716 312 235722
rect 303926 234358 304244 234362
rect 303926 234356 304246 234358
rect 304244 234038 304246 234356
rect 303926 234032 304244 234038
rect 102 232922 312 232926
rect -2012 232722 -2006 232922
rect -1806 232722 108 232922
rect 308 232722 312 232922
rect 102 232716 312 232722
rect 303926 231358 304244 231362
rect 303926 231356 304246 231358
rect 304244 231038 304246 231356
rect 303926 231032 304244 231038
rect 102 229922 312 229926
rect -2012 229722 -2006 229922
rect -1806 229722 108 229922
rect 308 229722 312 229922
rect 102 229716 312 229722
rect 303926 228358 304244 228362
rect 303926 228356 304246 228358
rect 304244 228038 304246 228356
rect 303926 228032 304244 228038
rect 102 226922 312 226926
rect -2012 226722 -2006 226922
rect -1806 226722 108 226922
rect 308 226722 312 226922
rect 102 226716 312 226722
rect 303926 225358 304244 225362
rect 303926 225356 304246 225358
rect 304244 225038 304246 225356
rect 303926 225032 304244 225038
rect 102 223922 312 223926
rect -2012 223722 -2006 223922
rect -1806 223722 108 223922
rect 308 223722 312 223922
rect 102 223716 312 223722
rect 303926 222358 304244 222362
rect 303926 222356 304246 222358
rect 304244 222038 304246 222356
rect 303926 222032 304244 222038
rect 102 220922 312 220926
rect -2012 220722 -2006 220922
rect -1806 220722 108 220922
rect 308 220722 312 220922
rect 102 220716 312 220722
rect 303926 219358 304244 219362
rect 303926 219356 304246 219358
rect 304244 219038 304246 219356
rect 303926 219032 304244 219038
rect 102 217922 312 217926
rect -2012 217722 -2006 217922
rect -1806 217722 108 217922
rect 308 217722 312 217922
rect 102 217716 312 217722
rect 303926 216358 304244 216362
rect 303926 216356 304246 216358
rect 304244 216038 304246 216356
rect 303926 216032 304244 216038
rect 102 214922 312 214926
rect -2012 214722 -2006 214922
rect -1806 214722 108 214922
rect 308 214722 312 214922
rect 102 214716 312 214722
rect 303926 213358 304244 213362
rect 303926 213356 304246 213358
rect 304244 213038 304246 213356
rect 303926 213032 304244 213038
rect 102 211922 312 211926
rect -2012 211722 -2006 211922
rect -1806 211722 108 211922
rect 308 211722 312 211922
rect 102 211716 312 211722
rect 303926 210358 304244 210362
rect 303926 210356 304246 210358
rect 304244 210038 304246 210356
rect 303926 210032 304244 210038
rect 102 208922 312 208926
rect -2012 208722 -2006 208922
rect -1806 208722 108 208922
rect 308 208722 312 208922
rect 102 208716 312 208722
rect 303926 207358 304244 207362
rect 303926 207356 304246 207358
rect 304244 207038 304246 207356
rect 303926 207032 304244 207038
rect 102 205922 312 205926
rect -2012 205722 -2006 205922
rect -1806 205722 108 205922
rect 308 205722 312 205922
rect 102 205716 312 205722
rect 303926 204358 304244 204362
rect 303926 204356 304246 204358
rect 304244 204038 304246 204356
rect 303926 204032 304244 204038
rect 102 202922 312 202926
rect -2012 202722 -2006 202922
rect -1806 202722 108 202922
rect 308 202722 312 202922
rect 102 202716 312 202722
rect 303926 201358 304244 201362
rect 303926 201356 304246 201358
rect 304244 201038 304246 201356
rect 303926 201032 304244 201038
rect 102 199922 312 199926
rect -2012 199722 -2006 199922
rect -1806 199722 108 199922
rect 308 199722 312 199922
rect 102 199716 312 199722
rect 303926 198358 304244 198362
rect 303926 198356 304246 198358
rect 304244 198038 304246 198356
rect 303926 198032 304244 198038
rect 102 196922 312 196926
rect -2012 196722 -2006 196922
rect -1806 196722 108 196922
rect 308 196722 312 196922
rect 102 196716 312 196722
rect 303926 195358 304244 195362
rect 303926 195356 304246 195358
rect 304244 195038 304246 195356
rect 303926 195032 304244 195038
rect 102 193922 312 193926
rect -2012 193722 -2006 193922
rect -1806 193722 108 193922
rect 308 193722 312 193922
rect 102 193716 312 193722
rect 303926 192358 304244 192362
rect 303926 192356 304246 192358
rect 304244 192038 304246 192356
rect 303926 192032 304244 192038
rect 102 190922 312 190926
rect -2012 190722 -2006 190922
rect -1806 190722 108 190922
rect 308 190722 312 190922
rect 102 190716 312 190722
rect 303926 189358 304244 189362
rect 303926 189356 304246 189358
rect 304244 189038 304246 189356
rect 303926 189032 304244 189038
rect 102 187922 312 187926
rect -2012 187722 -2006 187922
rect -1806 187722 108 187922
rect 308 187722 312 187922
rect 102 187716 312 187722
rect 303926 186358 304244 186362
rect 303926 186356 304246 186358
rect 304244 186038 304246 186356
rect 303926 186032 304244 186038
rect 102 184922 312 184926
rect -2012 184722 -2006 184922
rect -1806 184722 108 184922
rect 308 184722 312 184922
rect 102 184716 312 184722
rect 303926 183358 304244 183362
rect 303926 183356 304246 183358
rect 304244 183038 304246 183356
rect 303926 183032 304244 183038
rect 102 181922 312 181926
rect -2012 181722 -2006 181922
rect -1806 181722 108 181922
rect 308 181722 312 181922
rect 102 181716 312 181722
rect 303926 180358 304244 180362
rect 303926 180356 304246 180358
rect 304244 180038 304246 180356
rect 303926 180032 304244 180038
rect 102 178922 312 178926
rect -2012 178722 -2006 178922
rect -1806 178722 108 178922
rect 308 178722 312 178922
rect 102 178716 312 178722
rect 303926 177358 304244 177362
rect 303926 177356 304246 177358
rect 304244 177038 304246 177356
rect 303926 177032 304244 177038
rect 102 175922 312 175926
rect -2012 175722 -2006 175922
rect -1806 175722 108 175922
rect 308 175722 312 175922
rect 102 175716 312 175722
rect 303926 174358 304244 174362
rect 303926 174356 304246 174358
rect 304244 174038 304246 174356
rect 303926 174032 304244 174038
rect 102 172922 312 172926
rect -2012 172722 -2006 172922
rect -1806 172722 108 172922
rect 308 172722 312 172922
rect 102 172716 312 172722
rect 303926 171358 304244 171362
rect 303926 171356 304246 171358
rect 304244 171038 304246 171356
rect 303926 171032 304244 171038
rect 102 169922 312 169926
rect -2012 169722 -2006 169922
rect -1806 169722 108 169922
rect 308 169722 312 169922
rect 102 169716 312 169722
rect 303926 168358 304244 168362
rect 303926 168356 304246 168358
rect 304244 168038 304246 168356
rect 303926 168032 304244 168038
rect 102 166922 312 166926
rect -2012 166722 -2006 166922
rect -1806 166722 108 166922
rect 308 166722 312 166922
rect 102 166716 312 166722
rect 303926 165358 304244 165362
rect 303926 165356 304246 165358
rect 304244 165038 304246 165356
rect 303926 165032 304244 165038
rect 102 163922 312 163926
rect -2012 163722 -2006 163922
rect -1806 163722 108 163922
rect 308 163722 312 163922
rect 102 163716 312 163722
rect 303926 162358 304244 162362
rect 303926 162356 304246 162358
rect 304244 162038 304246 162356
rect 303926 162032 304244 162038
rect 102 160922 312 160926
rect -2012 160722 -2006 160922
rect -1806 160722 108 160922
rect 308 160722 312 160922
rect 102 160716 312 160722
rect 303926 159358 304244 159362
rect 303926 159356 304246 159358
rect 304244 159038 304246 159356
rect 303926 159032 304244 159038
rect 102 157922 312 157926
rect -2012 157722 -2006 157922
rect -1806 157722 108 157922
rect 308 157722 312 157922
rect 102 157716 312 157722
rect 303926 156358 304244 156362
rect 303926 156356 304246 156358
rect 304244 156038 304246 156356
rect 303926 156032 304244 156038
rect 102 154922 312 154926
rect -2012 154722 -2006 154922
rect -1806 154722 108 154922
rect 308 154722 312 154922
rect 102 154716 312 154722
rect 303926 153358 304244 153362
rect 303926 153356 304246 153358
rect 304244 153038 304246 153356
rect 303926 153032 304244 153038
rect 102 151922 312 151926
rect -2012 151722 -2006 151922
rect -1806 151722 108 151922
rect 308 151722 312 151922
rect 102 151716 312 151722
rect 303926 150358 304244 150362
rect 303926 150356 304246 150358
rect 304244 150038 304246 150356
rect 303926 150032 304244 150038
rect 102 148922 312 148926
rect -2012 148722 -2006 148922
rect -1806 148722 108 148922
rect 308 148722 312 148922
rect 102 148716 312 148722
rect 303926 147358 304244 147362
rect 303926 147356 304246 147358
rect 304244 147038 304246 147356
rect 303926 147032 304244 147038
rect 102 145922 312 145926
rect -2012 145722 -2006 145922
rect -1806 145722 108 145922
rect 308 145722 312 145922
rect 102 145716 312 145722
rect 303926 144358 304244 144362
rect 303926 144356 304246 144358
rect 304244 144038 304246 144356
rect 303926 144032 304244 144038
rect 102 142922 312 142926
rect -2012 142722 -2006 142922
rect -1806 142722 108 142922
rect 308 142722 312 142922
rect 102 142716 312 142722
rect 303926 141358 304244 141362
rect 303926 141356 304246 141358
rect 304244 141038 304246 141356
rect 303926 141032 304244 141038
rect 102 139922 312 139926
rect -2012 139722 -2006 139922
rect -1806 139722 108 139922
rect 308 139722 312 139922
rect 102 139716 312 139722
rect 303926 138358 304244 138362
rect 303926 138356 304246 138358
rect 304244 138038 304246 138356
rect 303926 138032 304244 138038
rect 102 136922 312 136926
rect -2012 136722 -2006 136922
rect -1806 136722 108 136922
rect 308 136722 312 136922
rect 102 136716 312 136722
rect 303926 135358 304244 135362
rect 303926 135356 304246 135358
rect 304244 135038 304246 135356
rect 303926 135032 304244 135038
rect 102 133922 312 133926
rect -2012 133722 -2006 133922
rect -1806 133722 108 133922
rect 308 133722 312 133922
rect 102 133716 312 133722
rect 303926 132358 304244 132362
rect 303926 132356 304246 132358
rect 304244 132038 304246 132356
rect 303926 132032 304244 132038
rect 102 130922 312 130926
rect -2012 130722 -2006 130922
rect -1806 130722 108 130922
rect 308 130722 312 130922
rect 102 130716 312 130722
rect 303926 129358 304244 129362
rect 303926 129356 304246 129358
rect 304244 129038 304246 129356
rect 303926 129032 304244 129038
rect 102 127922 312 127926
rect -2012 127722 -2006 127922
rect -1806 127722 108 127922
rect 308 127722 312 127922
rect 102 127716 312 127722
rect 303926 126358 304244 126362
rect 303926 126356 304246 126358
rect 304244 126038 304246 126356
rect 303926 126032 304244 126038
rect 102 124922 312 124926
rect -2012 124722 -2006 124922
rect -1806 124722 108 124922
rect 308 124722 312 124922
rect 102 124716 312 124722
rect 303926 123358 304244 123362
rect 303926 123356 304246 123358
rect 304244 123038 304246 123356
rect 303926 123032 304244 123038
rect 102 121922 312 121926
rect -2012 121722 -2006 121922
rect -1806 121722 108 121922
rect 308 121722 312 121922
rect 102 121716 312 121722
rect 303926 120358 304244 120362
rect 303926 120356 304246 120358
rect 304244 120038 304246 120356
rect 303926 120032 304244 120038
rect 102 118922 312 118926
rect -2012 118722 -2006 118922
rect -1806 118722 108 118922
rect 308 118722 312 118922
rect 102 118716 312 118722
rect 303926 117358 304244 117362
rect 303926 117356 304246 117358
rect 304244 117038 304246 117356
rect 303926 117032 304244 117038
rect 102 115922 312 115926
rect -2012 115722 -2006 115922
rect -1806 115722 108 115922
rect 308 115722 312 115922
rect 102 115716 312 115722
rect 303926 114358 304244 114362
rect 303926 114356 304246 114358
rect 304244 114038 304246 114356
rect 303926 114032 304244 114038
rect 102 112922 312 112926
rect -2012 112722 -2006 112922
rect -1806 112722 108 112922
rect 308 112722 312 112922
rect 102 112716 312 112722
rect 303926 111358 304244 111362
rect 303926 111356 304246 111358
rect 304244 111038 304246 111356
rect 303926 111032 304244 111038
rect 102 109922 312 109926
rect -2012 109722 -2006 109922
rect -1806 109722 108 109922
rect 308 109722 312 109922
rect 102 109716 312 109722
rect 303926 108358 304244 108362
rect 303926 108356 304246 108358
rect 304244 108038 304246 108356
rect 303926 108032 304244 108038
rect 102 106922 312 106926
rect -2012 106722 -2006 106922
rect -1806 106722 108 106922
rect 308 106722 312 106922
rect 102 106716 312 106722
rect 303926 105358 304244 105362
rect 303926 105356 304246 105358
rect 304244 105038 304246 105356
rect 303926 105032 304244 105038
rect 102 103922 312 103926
rect -2012 103722 -2006 103922
rect -1806 103722 108 103922
rect 308 103722 312 103922
rect 102 103716 312 103722
rect 303926 102358 304244 102362
rect 303926 102356 304246 102358
rect 304244 102038 304246 102356
rect 303926 102032 304244 102038
rect 102 100922 312 100926
rect -2012 100722 -2006 100922
rect -1806 100722 108 100922
rect 308 100722 312 100922
rect 102 100716 312 100722
rect 303926 99358 304244 99362
rect 303926 99356 304246 99358
rect 304244 99038 304246 99356
rect 303926 99032 304244 99038
rect 102 97922 312 97926
rect -2012 97722 -2006 97922
rect -1806 97722 108 97922
rect 308 97722 312 97922
rect 102 97716 312 97722
rect 303926 96358 304244 96362
rect 303926 96356 304246 96358
rect 304244 96038 304246 96356
rect 303926 96032 304244 96038
rect 102 94922 312 94926
rect -2012 94722 -2006 94922
rect -1806 94722 108 94922
rect 308 94722 312 94922
rect 102 94716 312 94722
rect 303926 93358 304244 93362
rect 303926 93356 304246 93358
rect 304244 93038 304246 93356
rect 303926 93032 304244 93038
rect 102 91922 312 91926
rect -2012 91722 -2006 91922
rect -1806 91722 108 91922
rect 308 91722 312 91922
rect 102 91716 312 91722
rect 303926 90358 304244 90362
rect 303926 90356 304246 90358
rect 304244 90038 304246 90356
rect 303926 90032 304244 90038
rect 102 88922 312 88926
rect -2012 88722 -2006 88922
rect -1806 88722 108 88922
rect 308 88722 312 88922
rect 102 88716 312 88722
rect 303926 87358 304244 87362
rect 303926 87356 304246 87358
rect 304244 87038 304246 87356
rect 303926 87032 304244 87038
rect 102 85922 312 85926
rect -2012 85722 -2006 85922
rect -1806 85722 108 85922
rect 308 85722 312 85922
rect 102 85716 312 85722
rect 303926 84358 304244 84362
rect 303926 84356 304246 84358
rect 304244 84038 304246 84356
rect 303926 84032 304244 84038
rect 102 82922 312 82926
rect -2012 82722 -2006 82922
rect -1806 82722 108 82922
rect 308 82722 312 82922
rect 102 82716 312 82722
rect 303926 81358 304244 81362
rect 303926 81356 304246 81358
rect 304244 81038 304246 81356
rect 303926 81032 304244 81038
rect 102 79922 312 79926
rect -2012 79722 -2006 79922
rect -1806 79722 108 79922
rect 308 79722 312 79922
rect 102 79716 312 79722
rect 303926 78358 304244 78362
rect 303926 78356 304246 78358
rect 304244 78038 304246 78356
rect 303926 78032 304244 78038
rect 102 76922 312 76926
rect -2012 76722 -2006 76922
rect -1806 76722 108 76922
rect 308 76722 312 76922
rect 102 76716 312 76722
rect 303926 75358 304244 75362
rect 303926 75356 304246 75358
rect 304244 75038 304246 75356
rect 303926 75032 304244 75038
rect 102 73922 312 73926
rect -2012 73722 -2006 73922
rect -1806 73722 108 73922
rect 308 73722 312 73922
rect 102 73716 312 73722
rect 303926 72358 304244 72362
rect 303926 72356 304246 72358
rect 304244 72038 304246 72356
rect 303926 72032 304244 72038
rect 102 70922 312 70926
rect -2012 70722 -2006 70922
rect -1806 70722 108 70922
rect 308 70722 312 70922
rect 102 70716 312 70722
rect 303926 69358 304244 69362
rect 303926 69356 304246 69358
rect 304244 69038 304246 69356
rect 303926 69032 304244 69038
rect 102 67922 312 67926
rect -2012 67722 -2006 67922
rect -1806 67722 108 67922
rect 308 67722 312 67922
rect 102 67716 312 67722
rect 303926 66358 304244 66362
rect 303926 66356 304246 66358
rect 304244 66038 304246 66356
rect 303926 66032 304244 66038
rect 102 64922 312 64926
rect -2012 64722 -2006 64922
rect -1806 64722 108 64922
rect 308 64722 312 64922
rect 102 64716 312 64722
rect 303926 63358 304244 63362
rect 303926 63356 304246 63358
rect 304244 63038 304246 63356
rect 303926 63032 304244 63038
rect 102 61922 312 61926
rect -2012 61722 -2006 61922
rect -1806 61722 108 61922
rect 308 61722 312 61922
rect 102 61716 312 61722
rect 303926 60358 304244 60362
rect 303926 60356 304246 60358
rect 304244 60038 304246 60356
rect 303926 60032 304244 60038
rect 102 58922 312 58926
rect -2012 58722 -2006 58922
rect -1806 58722 108 58922
rect 308 58722 312 58922
rect 102 58716 312 58722
rect 303926 57358 304244 57362
rect 303926 57356 304246 57358
rect 304244 57038 304246 57356
rect 303926 57032 304244 57038
rect 102 55922 312 55926
rect -2012 55722 -2006 55922
rect -1806 55722 108 55922
rect 308 55722 312 55922
rect 102 55716 312 55722
rect 303926 54358 304244 54362
rect 303926 54356 304246 54358
rect 304244 54038 304246 54356
rect 303926 54032 304244 54038
rect 102 52922 312 52926
rect -2012 52722 -2006 52922
rect -1806 52722 108 52922
rect 308 52722 312 52922
rect 102 52716 312 52722
rect 303926 51358 304244 51362
rect 303926 51356 304246 51358
rect 304244 51038 304246 51356
rect 303926 51032 304244 51038
rect 102 49922 312 49926
rect -2012 49722 -2006 49922
rect -1806 49722 108 49922
rect 308 49722 312 49922
rect 102 49716 312 49722
rect 303926 48358 304244 48362
rect 303926 48356 304246 48358
rect 304244 48038 304246 48356
rect 303926 48032 304244 48038
rect 102 46922 312 46926
rect -2012 46722 -2006 46922
rect -1806 46722 108 46922
rect 308 46722 312 46922
rect 102 46716 312 46722
rect 303926 45358 304244 45362
rect 303926 45356 304246 45358
rect 304244 45038 304246 45356
rect 303926 45032 304244 45038
rect 102 43922 312 43926
rect -2012 43722 -2006 43922
rect -1806 43722 108 43922
rect 308 43722 312 43922
rect 102 43716 312 43722
rect 303926 42358 304244 42362
rect 303926 42356 304246 42358
rect 304244 42038 304246 42356
rect 303926 42032 304244 42038
rect 102 40922 312 40926
rect -2012 40722 -2006 40922
rect -1806 40722 108 40922
rect 308 40722 312 40922
rect 102 40716 312 40722
rect 303926 39358 304244 39362
rect 303926 39356 304246 39358
rect 304244 39038 304246 39356
rect 303926 39032 304244 39038
rect 102 37922 312 37926
rect -2012 37722 -2006 37922
rect -1806 37722 108 37922
rect 308 37722 312 37922
rect 102 37716 312 37722
rect 303926 36358 304244 36362
rect 303926 36356 304246 36358
rect 304244 36038 304246 36356
rect 303926 36032 304244 36038
rect 102 34922 312 34926
rect -2012 34722 -2006 34922
rect -1806 34722 108 34922
rect 308 34722 312 34922
rect 102 34716 312 34722
rect 303926 33358 304244 33362
rect 303926 33356 304246 33358
rect 304244 33038 304246 33356
rect 303926 33032 304244 33038
rect 102 31922 312 31926
rect -2012 31722 -2006 31922
rect -1806 31722 108 31922
rect 308 31722 312 31922
rect 102 31716 312 31722
rect 303926 30358 304244 30362
rect 303926 30356 304246 30358
rect 304244 30038 304246 30356
rect 303926 30032 304244 30038
rect 102 28922 312 28926
rect -2012 28722 -2006 28922
rect -1806 28722 108 28922
rect 308 28722 312 28922
rect 102 28716 312 28722
rect 303926 27358 304244 27362
rect 303926 27356 304246 27358
rect 304244 27038 304246 27356
rect 303926 27032 304244 27038
rect 102 25922 312 25926
rect -2012 25722 -2006 25922
rect -1806 25722 108 25922
rect 308 25722 312 25922
rect 102 25716 312 25722
rect 303926 24358 304244 24362
rect 303926 24356 304246 24358
rect 304244 24038 304246 24356
rect 303926 24032 304244 24038
rect 102 22922 312 22926
rect -2012 22722 -2006 22922
rect -1806 22722 108 22922
rect 308 22722 312 22922
rect 102 22716 312 22722
rect 303926 21358 304244 21362
rect 303926 21356 304246 21358
rect 304244 21038 304246 21356
rect 303926 21032 304244 21038
rect 19870 19194 20088 19198
rect 19868 19192 20088 19194
rect 19868 18974 19870 19192
rect 29078 19062 29308 19066
rect 25944 19012 26162 19016
rect 19870 18968 20088 18974
rect 25942 19010 26162 19012
rect 13802 18930 14020 18934
rect 13800 18928 14020 18930
rect 7482 18890 7702 18892
rect 5328 18784 5546 18790
rect 3664 18758 3984 18760
rect 3658 18440 3664 18758
rect 3982 18440 3988 18758
rect 5546 18566 5548 18784
rect 7476 18672 7482 18890
rect 7700 18672 7706 18890
rect 10712 18836 10930 18840
rect 10710 18834 10930 18836
rect 10710 18616 10712 18834
rect 13800 18710 13802 18928
rect 16912 18816 17130 18822
rect 13802 18704 14020 18710
rect 10712 18610 10930 18616
rect 16910 18598 16912 18816
rect 25942 18792 25944 19010
rect 29078 18842 29084 19062
rect 29304 18842 29308 19062
rect 35328 19054 35548 19056
rect 29078 18836 29308 18842
rect 32328 18986 32546 18992
rect 25944 18786 26162 18792
rect 32546 18768 32548 18986
rect 35322 18836 35328 19054
rect 35546 18836 35552 19054
rect 38322 19000 38328 19218
rect 38546 19000 38552 19218
rect 56616 19162 56834 19168
rect 38328 18998 38548 19000
rect 44328 18922 44548 18924
rect 32328 18766 32548 18768
rect 32328 18762 32546 18766
rect 18088 18758 18408 18760
rect 32914 18758 33234 18760
rect 16910 18596 17130 18598
rect 16912 18592 17130 18596
rect 5328 18564 5548 18566
rect 5328 18560 5546 18564
rect 18082 18440 18088 18758
rect 18406 18440 18412 18758
rect 22898 18658 23116 18664
rect 22896 18440 22898 18658
rect 32908 18440 32914 18758
rect 33232 18440 33238 18758
rect 41322 18654 41328 18872
rect 41546 18654 41552 18872
rect 44322 18704 44328 18922
rect 44546 18704 44552 18922
rect 47322 18912 47328 19130
rect 47546 18912 47552 19130
rect 53538 19042 53756 19048
rect 50516 19012 50734 19016
rect 50516 19010 50736 19012
rect 47328 18910 47548 18912
rect 50734 18792 50736 19010
rect 53536 18824 53538 19042
rect 56614 18944 56616 19162
rect 174366 19134 174586 19136
rect 71928 19060 72146 19066
rect 56614 18942 56834 18944
rect 56616 18938 56834 18942
rect 65742 18882 65960 18886
rect 65742 18880 65962 18882
rect 53536 18822 53756 18824
rect 53538 18818 53756 18822
rect 59630 18866 59848 18872
rect 50516 18786 50734 18792
rect 41328 18652 41548 18654
rect 59848 18648 59850 18866
rect 59630 18646 59850 18648
rect 62632 18790 62850 18796
rect 59630 18642 59848 18646
rect 62850 18572 62852 18790
rect 64256 18758 64576 18760
rect 62632 18570 62852 18572
rect 62632 18566 62850 18570
rect 64250 18440 64256 18758
rect 64574 18440 64580 18758
rect 65960 18662 65962 18880
rect 68322 18734 68328 18952
rect 68546 18948 68770 18952
rect 68546 18738 68554 18948
rect 68764 18738 68770 18948
rect 68546 18734 68770 18738
rect 68328 18732 68770 18734
rect 72146 18842 72148 19060
rect 65742 18656 65960 18662
rect 71928 18520 72148 18842
rect 75078 19030 75296 19036
rect 108902 19032 109120 19038
rect 75296 18812 75298 19030
rect 81190 18904 81410 18906
rect 75078 18810 75298 18812
rect 75078 18806 75296 18810
rect 81184 18686 81190 18904
rect 81408 18686 81414 18904
rect 96452 18874 96672 18876
rect 90412 18836 90632 18838
rect 2328 18438 2548 18440
rect 22896 18438 23116 18440
rect 2322 18220 2328 18438
rect 2546 18220 2552 18438
rect 22898 18434 23116 18438
rect 71928 18310 71932 18520
rect 72142 18310 72148 18520
rect 81190 18496 81194 18686
rect 81404 18496 81410 18686
rect 90406 18618 90412 18836
rect 90630 18618 90636 18836
rect 93556 18792 93776 18794
rect 93550 18574 93556 18792
rect 93774 18574 93780 18792
rect 96448 18656 96454 18874
rect 96672 18656 96678 18874
rect 108900 18814 108902 19032
rect 157844 18998 158062 19002
rect 157842 18996 158062 18998
rect 114954 18984 115172 18990
rect 108900 18812 109120 18814
rect 108902 18808 109120 18812
rect 111948 18936 112166 18940
rect 111948 18934 112168 18936
rect 105674 18754 105894 18756
rect 102712 18740 102930 18746
rect 102710 18522 102712 18740
rect 105670 18536 105676 18754
rect 105894 18536 105900 18754
rect 112166 18716 112168 18934
rect 114952 18766 114954 18984
rect 114952 18764 115172 18766
rect 114954 18760 115172 18764
rect 117968 18978 118186 18982
rect 117968 18976 118188 18978
rect 118186 18758 118188 18976
rect 127242 18942 127460 18948
rect 121150 18864 121368 18870
rect 117968 18752 118186 18758
rect 111948 18710 112166 18716
rect 121368 18646 121370 18864
rect 124112 18852 124342 18856
rect 121678 18758 121998 18760
rect 121150 18644 121370 18646
rect 121150 18640 121368 18644
rect 102710 18520 102930 18522
rect 102712 18516 102930 18520
rect 99598 18502 99816 18506
rect 81190 18490 81410 18496
rect 99596 18500 99816 18502
rect 84274 18404 84492 18408
rect 84274 18402 84494 18404
rect 71928 18304 72148 18310
rect 78098 18306 78316 18312
rect 78316 18088 78318 18306
rect 78098 18076 78318 18088
rect -6204 17946 -5994 17952
rect -6204 17942 -6198 17946
rect -5998 17942 -5994 17946
rect 78098 17866 78102 18076
rect 78312 17866 78318 18076
rect 78098 17862 78318 17866
rect 84492 18184 84494 18402
rect 87336 18314 87554 18320
rect 84274 17980 84494 18184
rect 87334 18096 87336 18314
rect 99596 18282 99598 18500
rect 121672 18440 121678 18758
rect 121996 18440 122002 18758
rect 124112 18632 124118 18852
rect 124338 18632 124342 18852
rect 127240 18724 127242 18942
rect 133406 18866 133636 18872
rect 127240 18722 127460 18724
rect 127242 18718 127460 18722
rect 130250 18814 130468 18818
rect 130250 18812 130470 18814
rect 124112 18626 124342 18632
rect 130468 18594 130470 18812
rect 133406 18646 133412 18866
rect 133632 18646 133636 18866
rect 154792 18858 155010 18864
rect 145578 18844 145796 18848
rect 148754 18844 148972 18848
rect 145578 18842 145798 18844
rect 142600 18668 142818 18674
rect 133406 18642 133636 18646
rect 139552 18600 139770 18606
rect 130250 18588 130468 18594
rect 139770 18382 139772 18600
rect 142598 18450 142600 18668
rect 145796 18624 145798 18842
rect 148754 18842 148974 18844
rect 148972 18624 148974 18842
rect 151772 18774 151990 18780
rect 145578 18618 145796 18624
rect 148754 18618 148972 18624
rect 151990 18556 151992 18774
rect 155010 18640 155012 18858
rect 157842 18778 157844 18996
rect 174360 18916 174366 19134
rect 174584 18916 174590 19134
rect 305386 19100 305604 19104
rect 305384 19098 305604 19100
rect 290328 18956 290546 18960
rect 290328 18954 290548 18956
rect 229658 18938 229878 18940
rect 157844 18772 158062 18778
rect 167548 18758 167868 18760
rect 154792 18638 155012 18640
rect 154792 18634 155010 18638
rect 151772 18554 151992 18556
rect 151772 18550 151990 18554
rect 160880 18540 160886 18758
rect 161104 18540 161110 18758
rect 160886 18538 161106 18540
rect 163238 18458 163458 18460
rect 142598 18448 142818 18450
rect 142600 18444 142818 18448
rect 139552 18380 139772 18382
rect 139552 18376 139770 18380
rect 99598 18276 99816 18282
rect 136466 18240 136686 18242
rect 163232 18240 163238 18458
rect 163456 18240 163462 18458
rect 167542 18440 167548 18758
rect 167866 18440 167872 18758
rect 176322 18594 176328 18812
rect 176546 18594 176552 18812
rect 180548 18758 180868 18760
rect 189548 18758 189868 18760
rect 198548 18758 198868 18760
rect 204548 18758 204868 18760
rect 211548 18758 211868 18760
rect 223548 18758 223868 18760
rect 176328 18592 176548 18594
rect 173082 18490 173300 18494
rect 173082 18488 173302 18490
rect 173300 18270 173302 18488
rect 180542 18440 180548 18758
rect 180866 18440 180872 18758
rect 189542 18440 189548 18758
rect 189866 18440 189872 18758
rect 198542 18440 198548 18758
rect 198866 18440 198872 18758
rect 204542 18440 204548 18758
rect 204866 18440 204872 18758
rect 206328 18456 206546 18460
rect 206328 18454 206548 18456
rect 173082 18264 173300 18270
rect 87334 18094 87554 18096
rect 87336 18090 87554 18094
rect 136462 18022 136468 18240
rect 136686 18022 136692 18240
rect 206546 18236 206548 18454
rect 211542 18440 211548 18758
rect 211866 18440 211872 18758
rect 215328 18564 215546 18568
rect 215328 18562 215548 18564
rect 215546 18344 215548 18562
rect 223542 18440 223548 18758
rect 223866 18440 223872 18758
rect 229652 18720 229658 18938
rect 229876 18720 229882 18938
rect 232548 18758 232868 18760
rect 238548 18758 238868 18760
rect 250548 18758 250868 18760
rect 263948 18758 264268 18760
rect 269948 18758 270268 18760
rect 272948 18758 273268 18760
rect 275948 18758 276268 18760
rect 281948 18758 282268 18760
rect 285948 18758 286268 18760
rect 232542 18440 232548 18758
rect 232866 18440 232872 18758
rect 233328 18690 233546 18694
rect 233328 18688 233548 18690
rect 233546 18470 233548 18688
rect 233328 18464 233546 18470
rect 238542 18440 238548 18758
rect 238866 18440 238872 18758
rect 242328 18570 242546 18576
rect 241672 18534 241890 18540
rect 215328 18338 215546 18344
rect 206328 18230 206546 18236
rect 227188 18210 227194 18428
rect 227412 18210 227418 18428
rect 241890 18316 241892 18534
rect 242546 18352 242548 18570
rect 250542 18440 250548 18758
rect 250866 18440 250872 18758
rect 254328 18700 254546 18706
rect 253924 18508 254144 18510
rect 242328 18350 242548 18352
rect 242328 18346 242546 18350
rect 241672 18314 241892 18316
rect 241672 18310 241890 18314
rect 234650 18302 234870 18304
rect 227194 18208 227414 18210
rect 165928 18174 166146 18180
rect 84274 17770 84278 17980
rect 84488 17770 84494 17980
rect 166146 17956 166148 18174
rect 213156 18098 213374 18104
rect 165928 17954 166148 17956
rect 185328 18036 185546 18042
rect 165928 17950 166146 17954
rect 182472 17858 182692 17860
rect 84274 17764 84494 17770
rect -6204 17736 -5994 17742
rect -19160 17346 -19040 17596
rect -15216 17346 -15096 17624
rect -11136 17394 -11016 17688
rect -7192 17338 -7072 17696
rect 182468 17640 182474 17858
rect 182692 17640 182698 17858
rect 185546 17818 185548 18036
rect 200916 17956 201134 17962
rect 196792 17928 197012 17930
rect 185328 17816 185548 17818
rect 185328 17812 185546 17816
rect 196788 17710 196794 17928
rect 197012 17710 197018 17928
rect 200914 17738 200916 17956
rect 213154 17880 213156 18098
rect 234644 18084 234650 18302
rect 234868 18084 234874 18302
rect 253920 18290 253926 18508
rect 254144 18290 254150 18508
rect 254546 18482 254548 18700
rect 254328 18480 254548 18482
rect 254328 18476 254546 18480
rect 263942 18440 263948 18758
rect 264266 18440 264272 18758
rect 269026 18342 269032 18560
rect 269250 18342 269256 18560
rect 269942 18440 269948 18758
rect 270266 18440 270272 18758
rect 272942 18440 272948 18758
rect 273266 18440 273272 18758
rect 275942 18440 275948 18758
rect 276266 18440 276272 18758
rect 279670 18480 279676 18698
rect 279894 18480 279900 18698
rect 279676 18478 279896 18480
rect 281942 18440 281948 18758
rect 282266 18440 282272 18758
rect 285942 18440 285948 18758
rect 286266 18440 286272 18758
rect 290546 18736 290548 18954
rect 305384 18880 305386 19098
rect 305386 18874 305604 18880
rect 293948 18758 294268 18760
rect 296948 18758 297268 18760
rect 299948 18758 300268 18760
rect 302948 18758 303268 18760
rect 290328 18730 290546 18736
rect 293942 18440 293948 18758
rect 294266 18440 294272 18758
rect 296942 18440 296948 18758
rect 297266 18440 297272 18758
rect 299942 18440 299948 18758
rect 300266 18440 300272 18758
rect 302942 18440 302948 18758
rect 303266 18440 303272 18758
rect 269032 18340 269252 18342
rect 269328 18268 269546 18274
rect 261044 18126 261262 18130
rect 261044 18124 261264 18126
rect 213154 17878 213374 17880
rect 213156 17874 213374 17878
rect 240916 18016 241134 18020
rect 240916 18014 241136 18016
rect 241134 17796 241136 18014
rect 261262 17906 261264 18124
rect 269546 18050 269548 18268
rect 292406 18226 292626 18228
rect 269328 18048 269548 18050
rect 269328 18044 269546 18048
rect 278872 17988 278878 18206
rect 279096 17988 279102 18206
rect 284328 18138 284546 18142
rect 284328 18136 284548 18138
rect 278878 17986 279098 17988
rect 265870 17964 266088 17968
rect 265870 17962 266090 17964
rect 261044 17900 261262 17906
rect 240916 17790 241134 17796
rect 207000 17752 207218 17756
rect 200914 17736 201134 17738
rect 200916 17732 201134 17736
rect 206998 17750 207218 17752
rect 188328 17660 188546 17664
rect 188328 17658 188548 17660
rect 188546 17440 188548 17658
rect 206998 17532 207000 17750
rect 207000 17526 207218 17532
rect 221328 17712 221546 17716
rect 221328 17710 221548 17712
rect 221546 17492 221548 17710
rect 249662 17642 249668 17860
rect 249886 17642 249892 17860
rect 266088 17744 266090 17962
rect 284546 17918 284548 18136
rect 292402 18008 292408 18226
rect 292626 18008 292632 18226
rect 284328 17912 284546 17918
rect 265870 17738 266088 17744
rect 299258 17724 299476 17728
rect 299258 17722 299478 17724
rect 249666 17640 249886 17642
rect 221328 17486 221546 17492
rect 188328 17434 188546 17440
rect 168864 17422 169082 17426
rect 168862 17420 169082 17422
rect 168862 17202 168864 17420
rect 277688 17364 277694 17582
rect 277912 17364 277918 17582
rect 286930 17512 287148 17518
rect 277692 17362 277912 17364
rect 286928 17294 286930 17512
rect 299476 17504 299478 17722
rect 299258 17498 299476 17504
rect 286928 17292 287148 17294
rect 286930 17288 287148 17292
rect 168864 17196 169082 17202
rect 213904 17270 214122 17274
rect 213904 17268 214124 17270
rect 184010 17152 184228 17158
rect 184228 16934 184230 17152
rect 214122 17050 214124 17268
rect 260054 17246 260272 17252
rect 220688 17228 220906 17234
rect 213904 17044 214122 17050
rect 193466 17020 193684 17024
rect 184010 16932 184230 16934
rect 193464 17018 193684 17020
rect 184010 16928 184228 16932
rect 193464 16800 193466 17018
rect 220906 17010 220908 17228
rect 248712 17078 248930 17082
rect 220688 17008 220908 17010
rect 248710 17076 248930 17078
rect 220688 17004 220906 17008
rect 202004 16894 202222 16900
rect 193466 16794 193684 16800
rect 202002 16676 202004 16894
rect 248710 16858 248712 17076
rect 260052 17028 260054 17246
rect 300252 17106 300470 17110
rect 260052 17026 260272 17028
rect 260054 17022 260272 17026
rect 300250 17104 300470 17106
rect 300250 16886 300252 17104
rect 300252 16880 300470 16886
rect 248712 16852 248930 16858
rect 202002 16674 202222 16676
rect 202004 16670 202222 16674
rect 302942 16416 303274 16420
rect 302942 16410 302946 16416
rect 303268 16410 303274 16416
rect 302942 16082 303274 16088
rect 18082 15712 18412 15716
rect 18082 15706 18088 15712
rect 18408 15706 18412 15712
rect 3658 15694 3988 15698
rect 3658 15688 3664 15694
rect 3984 15688 3988 15694
rect 102 15588 312 15592
rect 102 15582 108 15588
rect 308 15582 312 15588
rect 102 15376 312 15382
rect 121672 15710 122002 15714
rect 121672 15704 121678 15710
rect 121998 15704 122002 15710
rect 64250 15696 64580 15700
rect 18082 15380 18412 15386
rect 32908 15688 33238 15692
rect 32908 15682 32914 15688
rect 33234 15682 33238 15688
rect 3658 15362 3988 15368
rect 64250 15690 64256 15696
rect 64576 15690 64580 15696
rect 121672 15378 122002 15384
rect 167542 15712 167872 15716
rect 167542 15706 167548 15712
rect 167868 15706 167872 15712
rect 167542 15380 167872 15386
rect 180542 15712 180872 15716
rect 180542 15706 180548 15712
rect 180868 15706 180872 15712
rect 180542 15380 180872 15386
rect 189542 15712 189872 15716
rect 189542 15706 189548 15712
rect 189868 15706 189872 15712
rect 189542 15380 189872 15386
rect 198542 15712 198872 15716
rect 198542 15706 198548 15712
rect 198868 15706 198872 15712
rect 198542 15380 198872 15386
rect 204542 15712 204872 15716
rect 204542 15706 204548 15712
rect 204868 15706 204872 15712
rect 204542 15380 204872 15386
rect 211542 15712 211872 15716
rect 211542 15706 211548 15712
rect 211868 15706 211872 15712
rect 211542 15380 211872 15386
rect 223542 15712 223872 15716
rect 223542 15706 223548 15712
rect 223868 15706 223872 15712
rect 223542 15380 223872 15386
rect 232542 15712 232872 15716
rect 232542 15706 232548 15712
rect 232868 15706 232872 15712
rect 232542 15380 232872 15386
rect 238542 15712 238872 15716
rect 238542 15706 238548 15712
rect 238868 15706 238872 15712
rect 238542 15380 238872 15386
rect 250542 15712 250872 15716
rect 250542 15706 250548 15712
rect 250868 15706 250872 15712
rect 250542 15380 250872 15386
rect 263942 15712 264272 15716
rect 263942 15706 263948 15712
rect 264268 15706 264272 15712
rect 263942 15380 264272 15386
rect 269942 15712 270272 15716
rect 269942 15706 269948 15712
rect 270268 15706 270272 15712
rect 269942 15380 270272 15386
rect 272942 15712 273272 15716
rect 272942 15706 272948 15712
rect 273268 15706 273272 15712
rect 272942 15380 273272 15386
rect 275942 15712 276272 15716
rect 275942 15706 275948 15712
rect 276268 15706 276272 15712
rect 275942 15380 276272 15386
rect 281942 15712 282272 15716
rect 281942 15706 281948 15712
rect 282268 15706 282272 15712
rect 281942 15380 282272 15386
rect 285942 15712 286272 15716
rect 285942 15706 285948 15712
rect 286268 15706 286272 15712
rect 285942 15380 286272 15386
rect 293942 15712 294272 15716
rect 293942 15706 293948 15712
rect 294268 15706 294272 15712
rect 293942 15380 294272 15386
rect 296942 15712 297272 15716
rect 296942 15706 296948 15712
rect 297268 15706 297272 15712
rect 296942 15380 297272 15386
rect 299942 15712 300272 15716
rect 299942 15706 299948 15712
rect 300268 15706 300272 15712
rect 299942 15380 300272 15386
rect 302942 15712 303272 15716
rect 302942 15706 302948 15712
rect 303268 15706 303272 15712
rect 302942 15380 303272 15386
rect 64250 15364 64580 15370
rect 32908 15356 33238 15362
rect 306608 14470 306790 14590
rect 306628 10526 306844 10646
rect 114 8622 316 8742
rect 306712 6446 306920 6566
rect 306596 2502 306806 2622
<< via3 >>
rect 302502 324532 302712 324538
rect 302502 324338 302508 324532
rect 302508 324338 302708 324532
rect 302708 324338 302712 324532
rect 303926 321352 304244 321356
rect 303926 321042 303930 321352
rect 303930 321042 304240 321352
rect 304240 321042 304244 321352
rect 303926 321038 304244 321042
rect -2006 319722 -1806 319922
rect 303926 318352 304244 318356
rect 303926 318042 303930 318352
rect 303930 318042 304240 318352
rect 304240 318042 304244 318352
rect 303926 318038 304244 318042
rect -2006 316722 -1806 316922
rect 303926 315352 304244 315356
rect 303926 315042 303930 315352
rect 303930 315042 304240 315352
rect 304240 315042 304244 315352
rect 303926 315038 304244 315042
rect -2006 313722 -1806 313922
rect 303926 312352 304244 312356
rect 303926 312042 303930 312352
rect 303930 312042 304240 312352
rect 304240 312042 304244 312352
rect 303926 312038 304244 312042
rect -2006 310722 -1806 310922
rect 303926 309352 304244 309356
rect 303926 309042 303930 309352
rect 303930 309042 304240 309352
rect 304240 309042 304244 309352
rect 303926 309038 304244 309042
rect -2006 307722 -1806 307922
rect 303926 306352 304244 306356
rect 303926 306042 303930 306352
rect 303930 306042 304240 306352
rect 304240 306042 304244 306352
rect 303926 306038 304244 306042
rect -2006 304722 -1806 304922
rect 303926 303352 304244 303356
rect 303926 303042 303930 303352
rect 303930 303042 304240 303352
rect 304240 303042 304244 303352
rect 303926 303038 304244 303042
rect -2006 301722 -1806 301922
rect 303926 300352 304244 300356
rect 303926 300042 303930 300352
rect 303930 300042 304240 300352
rect 304240 300042 304244 300352
rect 303926 300038 304244 300042
rect -2006 298722 -1806 298922
rect 303926 297352 304244 297356
rect 303926 297042 303930 297352
rect 303930 297042 304240 297352
rect 304240 297042 304244 297352
rect 303926 297038 304244 297042
rect -2006 295722 -1806 295922
rect 303926 294352 304244 294356
rect 303926 294042 303930 294352
rect 303930 294042 304240 294352
rect 304240 294042 304244 294352
rect 303926 294038 304244 294042
rect -2006 292722 -1806 292922
rect 303926 291352 304244 291356
rect 303926 291042 303930 291352
rect 303930 291042 304240 291352
rect 304240 291042 304244 291352
rect 303926 291038 304244 291042
rect -2006 289722 -1806 289922
rect 303926 288352 304244 288356
rect 303926 288042 303930 288352
rect 303930 288042 304240 288352
rect 304240 288042 304244 288352
rect 303926 288038 304244 288042
rect -2006 286722 -1806 286922
rect 303926 285352 304244 285356
rect 303926 285042 303930 285352
rect 303930 285042 304240 285352
rect 304240 285042 304244 285352
rect 303926 285038 304244 285042
rect -2006 283722 -1806 283922
rect 303926 282352 304244 282356
rect 303926 282042 303930 282352
rect 303930 282042 304240 282352
rect 304240 282042 304244 282352
rect 303926 282038 304244 282042
rect -2006 280722 -1806 280922
rect 303926 279352 304244 279356
rect 303926 279042 303930 279352
rect 303930 279042 304240 279352
rect 304240 279042 304244 279352
rect 303926 279038 304244 279042
rect -2006 277722 -1806 277922
rect 303926 276352 304244 276356
rect 303926 276042 303930 276352
rect 303930 276042 304240 276352
rect 304240 276042 304244 276352
rect 303926 276038 304244 276042
rect -2006 274722 -1806 274922
rect 303926 273352 304244 273356
rect 303926 273042 303930 273352
rect 303930 273042 304240 273352
rect 304240 273042 304244 273352
rect 303926 273038 304244 273042
rect -2006 271722 -1806 271922
rect 303926 270352 304244 270356
rect 303926 270042 303930 270352
rect 303930 270042 304240 270352
rect 304240 270042 304244 270352
rect 303926 270038 304244 270042
rect -2006 268722 -1806 268922
rect 303926 267352 304244 267356
rect 303926 267042 303930 267352
rect 303930 267042 304240 267352
rect 304240 267042 304244 267352
rect 303926 267038 304244 267042
rect -2006 265722 -1806 265922
rect 303926 264352 304244 264356
rect 303926 264042 303930 264352
rect 303930 264042 304240 264352
rect 304240 264042 304244 264352
rect 303926 264038 304244 264042
rect -2006 262722 -1806 262922
rect 303926 261352 304244 261356
rect 303926 261042 303930 261352
rect 303930 261042 304240 261352
rect 304240 261042 304244 261352
rect 303926 261038 304244 261042
rect -2006 259722 -1806 259922
rect 303926 258352 304244 258356
rect 303926 258042 303930 258352
rect 303930 258042 304240 258352
rect 304240 258042 304244 258352
rect 303926 258038 304244 258042
rect -2006 256722 -1806 256922
rect 303926 255352 304244 255356
rect 303926 255042 303930 255352
rect 303930 255042 304240 255352
rect 304240 255042 304244 255352
rect 303926 255038 304244 255042
rect -2006 253722 -1806 253922
rect 303926 252352 304244 252356
rect 303926 252042 303930 252352
rect 303930 252042 304240 252352
rect 304240 252042 304244 252352
rect 303926 252038 304244 252042
rect -2006 250722 -1806 250922
rect 303926 249352 304244 249356
rect 303926 249042 303930 249352
rect 303930 249042 304240 249352
rect 304240 249042 304244 249352
rect 303926 249038 304244 249042
rect -2006 247722 -1806 247922
rect 303926 246352 304244 246356
rect 303926 246042 303930 246352
rect 303930 246042 304240 246352
rect 304240 246042 304244 246352
rect 303926 246038 304244 246042
rect -2006 244722 -1806 244922
rect 303926 243352 304244 243356
rect 303926 243042 303930 243352
rect 303930 243042 304240 243352
rect 304240 243042 304244 243352
rect 303926 243038 304244 243042
rect -2006 241722 -1806 241922
rect 303926 240352 304244 240356
rect 303926 240042 303930 240352
rect 303930 240042 304240 240352
rect 304240 240042 304244 240352
rect 303926 240038 304244 240042
rect -2006 238722 -1806 238922
rect 303926 237352 304244 237356
rect 303926 237042 303930 237352
rect 303930 237042 304240 237352
rect 304240 237042 304244 237352
rect 303926 237038 304244 237042
rect -2006 235722 -1806 235922
rect 303926 234352 304244 234356
rect 303926 234042 303930 234352
rect 303930 234042 304240 234352
rect 304240 234042 304244 234352
rect 303926 234038 304244 234042
rect -2006 232722 -1806 232922
rect 303926 231352 304244 231356
rect 303926 231042 303930 231352
rect 303930 231042 304240 231352
rect 304240 231042 304244 231352
rect 303926 231038 304244 231042
rect -2006 229722 -1806 229922
rect 303926 228352 304244 228356
rect 303926 228042 303930 228352
rect 303930 228042 304240 228352
rect 304240 228042 304244 228352
rect 303926 228038 304244 228042
rect -2006 226722 -1806 226922
rect 303926 225352 304244 225356
rect 303926 225042 303930 225352
rect 303930 225042 304240 225352
rect 304240 225042 304244 225352
rect 303926 225038 304244 225042
rect -2006 223722 -1806 223922
rect 303926 222352 304244 222356
rect 303926 222042 303930 222352
rect 303930 222042 304240 222352
rect 304240 222042 304244 222352
rect 303926 222038 304244 222042
rect -2006 220722 -1806 220922
rect 303926 219352 304244 219356
rect 303926 219042 303930 219352
rect 303930 219042 304240 219352
rect 304240 219042 304244 219352
rect 303926 219038 304244 219042
rect -2006 217722 -1806 217922
rect 303926 216352 304244 216356
rect 303926 216042 303930 216352
rect 303930 216042 304240 216352
rect 304240 216042 304244 216352
rect 303926 216038 304244 216042
rect -2006 214722 -1806 214922
rect 303926 213352 304244 213356
rect 303926 213042 303930 213352
rect 303930 213042 304240 213352
rect 304240 213042 304244 213352
rect 303926 213038 304244 213042
rect -2006 211722 -1806 211922
rect 303926 210352 304244 210356
rect 303926 210042 303930 210352
rect 303930 210042 304240 210352
rect 304240 210042 304244 210352
rect 303926 210038 304244 210042
rect -2006 208722 -1806 208922
rect 303926 207352 304244 207356
rect 303926 207042 303930 207352
rect 303930 207042 304240 207352
rect 304240 207042 304244 207352
rect 303926 207038 304244 207042
rect -2006 205722 -1806 205922
rect 303926 204352 304244 204356
rect 303926 204042 303930 204352
rect 303930 204042 304240 204352
rect 304240 204042 304244 204352
rect 303926 204038 304244 204042
rect -2006 202722 -1806 202922
rect 303926 201352 304244 201356
rect 303926 201042 303930 201352
rect 303930 201042 304240 201352
rect 304240 201042 304244 201352
rect 303926 201038 304244 201042
rect -2006 199722 -1806 199922
rect 303926 198352 304244 198356
rect 303926 198042 303930 198352
rect 303930 198042 304240 198352
rect 304240 198042 304244 198352
rect 303926 198038 304244 198042
rect -2006 196722 -1806 196922
rect 303926 195352 304244 195356
rect 303926 195042 303930 195352
rect 303930 195042 304240 195352
rect 304240 195042 304244 195352
rect 303926 195038 304244 195042
rect -2006 193722 -1806 193922
rect 303926 192352 304244 192356
rect 303926 192042 303930 192352
rect 303930 192042 304240 192352
rect 304240 192042 304244 192352
rect 303926 192038 304244 192042
rect -2006 190722 -1806 190922
rect 303926 189352 304244 189356
rect 303926 189042 303930 189352
rect 303930 189042 304240 189352
rect 304240 189042 304244 189352
rect 303926 189038 304244 189042
rect -2006 187722 -1806 187922
rect 303926 186352 304244 186356
rect 303926 186042 303930 186352
rect 303930 186042 304240 186352
rect 304240 186042 304244 186352
rect 303926 186038 304244 186042
rect -2006 184722 -1806 184922
rect 303926 183352 304244 183356
rect 303926 183042 303930 183352
rect 303930 183042 304240 183352
rect 304240 183042 304244 183352
rect 303926 183038 304244 183042
rect -2006 181722 -1806 181922
rect 303926 180352 304244 180356
rect 303926 180042 303930 180352
rect 303930 180042 304240 180352
rect 304240 180042 304244 180352
rect 303926 180038 304244 180042
rect -2006 178722 -1806 178922
rect 303926 177352 304244 177356
rect 303926 177042 303930 177352
rect 303930 177042 304240 177352
rect 304240 177042 304244 177352
rect 303926 177038 304244 177042
rect -2006 175722 -1806 175922
rect 303926 174352 304244 174356
rect 303926 174042 303930 174352
rect 303930 174042 304240 174352
rect 304240 174042 304244 174352
rect 303926 174038 304244 174042
rect -2006 172722 -1806 172922
rect 303926 171352 304244 171356
rect 303926 171042 303930 171352
rect 303930 171042 304240 171352
rect 304240 171042 304244 171352
rect 303926 171038 304244 171042
rect -2006 169722 -1806 169922
rect 303926 168352 304244 168356
rect 303926 168042 303930 168352
rect 303930 168042 304240 168352
rect 304240 168042 304244 168352
rect 303926 168038 304244 168042
rect -2006 166722 -1806 166922
rect 303926 165352 304244 165356
rect 303926 165042 303930 165352
rect 303930 165042 304240 165352
rect 304240 165042 304244 165352
rect 303926 165038 304244 165042
rect -2006 163722 -1806 163922
rect 303926 162352 304244 162356
rect 303926 162042 303930 162352
rect 303930 162042 304240 162352
rect 304240 162042 304244 162352
rect 303926 162038 304244 162042
rect -2006 160722 -1806 160922
rect 303926 159352 304244 159356
rect 303926 159042 303930 159352
rect 303930 159042 304240 159352
rect 304240 159042 304244 159352
rect 303926 159038 304244 159042
rect -2006 157722 -1806 157922
rect 303926 156352 304244 156356
rect 303926 156042 303930 156352
rect 303930 156042 304240 156352
rect 304240 156042 304244 156352
rect 303926 156038 304244 156042
rect -2006 154722 -1806 154922
rect 303926 153352 304244 153356
rect 303926 153042 303930 153352
rect 303930 153042 304240 153352
rect 304240 153042 304244 153352
rect 303926 153038 304244 153042
rect -2006 151722 -1806 151922
rect 303926 150352 304244 150356
rect 303926 150042 303930 150352
rect 303930 150042 304240 150352
rect 304240 150042 304244 150352
rect 303926 150038 304244 150042
rect -2006 148722 -1806 148922
rect 303926 147352 304244 147356
rect 303926 147042 303930 147352
rect 303930 147042 304240 147352
rect 304240 147042 304244 147352
rect 303926 147038 304244 147042
rect -2006 145722 -1806 145922
rect 303926 144352 304244 144356
rect 303926 144042 303930 144352
rect 303930 144042 304240 144352
rect 304240 144042 304244 144352
rect 303926 144038 304244 144042
rect -2006 142722 -1806 142922
rect 303926 141352 304244 141356
rect 303926 141042 303930 141352
rect 303930 141042 304240 141352
rect 304240 141042 304244 141352
rect 303926 141038 304244 141042
rect -2006 139722 -1806 139922
rect 303926 138352 304244 138356
rect 303926 138042 303930 138352
rect 303930 138042 304240 138352
rect 304240 138042 304244 138352
rect 303926 138038 304244 138042
rect -2006 136722 -1806 136922
rect 303926 135352 304244 135356
rect 303926 135042 303930 135352
rect 303930 135042 304240 135352
rect 304240 135042 304244 135352
rect 303926 135038 304244 135042
rect -2006 133722 -1806 133922
rect 303926 132352 304244 132356
rect 303926 132042 303930 132352
rect 303930 132042 304240 132352
rect 304240 132042 304244 132352
rect 303926 132038 304244 132042
rect -2006 130722 -1806 130922
rect 303926 129352 304244 129356
rect 303926 129042 303930 129352
rect 303930 129042 304240 129352
rect 304240 129042 304244 129352
rect 303926 129038 304244 129042
rect -2006 127722 -1806 127922
rect 303926 126352 304244 126356
rect 303926 126042 303930 126352
rect 303930 126042 304240 126352
rect 304240 126042 304244 126352
rect 303926 126038 304244 126042
rect -2006 124722 -1806 124922
rect 303926 123352 304244 123356
rect 303926 123042 303930 123352
rect 303930 123042 304240 123352
rect 304240 123042 304244 123352
rect 303926 123038 304244 123042
rect -2006 121722 -1806 121922
rect 303926 120352 304244 120356
rect 303926 120042 303930 120352
rect 303930 120042 304240 120352
rect 304240 120042 304244 120352
rect 303926 120038 304244 120042
rect -2006 118722 -1806 118922
rect 303926 117352 304244 117356
rect 303926 117042 303930 117352
rect 303930 117042 304240 117352
rect 304240 117042 304244 117352
rect 303926 117038 304244 117042
rect -2006 115722 -1806 115922
rect 303926 114352 304244 114356
rect 303926 114042 303930 114352
rect 303930 114042 304240 114352
rect 304240 114042 304244 114352
rect 303926 114038 304244 114042
rect -2006 112722 -1806 112922
rect 303926 111352 304244 111356
rect 303926 111042 303930 111352
rect 303930 111042 304240 111352
rect 304240 111042 304244 111352
rect 303926 111038 304244 111042
rect -2006 109722 -1806 109922
rect 303926 108352 304244 108356
rect 303926 108042 303930 108352
rect 303930 108042 304240 108352
rect 304240 108042 304244 108352
rect 303926 108038 304244 108042
rect -2006 106722 -1806 106922
rect 303926 105352 304244 105356
rect 303926 105042 303930 105352
rect 303930 105042 304240 105352
rect 304240 105042 304244 105352
rect 303926 105038 304244 105042
rect -2006 103722 -1806 103922
rect 303926 102352 304244 102356
rect 303926 102042 303930 102352
rect 303930 102042 304240 102352
rect 304240 102042 304244 102352
rect 303926 102038 304244 102042
rect -2006 100722 -1806 100922
rect 303926 99352 304244 99356
rect 303926 99042 303930 99352
rect 303930 99042 304240 99352
rect 304240 99042 304244 99352
rect 303926 99038 304244 99042
rect -2006 97722 -1806 97922
rect 303926 96352 304244 96356
rect 303926 96042 303930 96352
rect 303930 96042 304240 96352
rect 304240 96042 304244 96352
rect 303926 96038 304244 96042
rect -2006 94722 -1806 94922
rect 303926 93352 304244 93356
rect 303926 93042 303930 93352
rect 303930 93042 304240 93352
rect 304240 93042 304244 93352
rect 303926 93038 304244 93042
rect -2006 91722 -1806 91922
rect 303926 90352 304244 90356
rect 303926 90042 303930 90352
rect 303930 90042 304240 90352
rect 304240 90042 304244 90352
rect 303926 90038 304244 90042
rect -2006 88722 -1806 88922
rect 303926 87352 304244 87356
rect 303926 87042 303930 87352
rect 303930 87042 304240 87352
rect 304240 87042 304244 87352
rect 303926 87038 304244 87042
rect -2006 85722 -1806 85922
rect 303926 84352 304244 84356
rect 303926 84042 303930 84352
rect 303930 84042 304240 84352
rect 304240 84042 304244 84352
rect 303926 84038 304244 84042
rect -2006 82722 -1806 82922
rect 303926 81352 304244 81356
rect 303926 81042 303930 81352
rect 303930 81042 304240 81352
rect 304240 81042 304244 81352
rect 303926 81038 304244 81042
rect -2006 79722 -1806 79922
rect 303926 78352 304244 78356
rect 303926 78042 303930 78352
rect 303930 78042 304240 78352
rect 304240 78042 304244 78352
rect 303926 78038 304244 78042
rect -2006 76722 -1806 76922
rect 303926 75352 304244 75356
rect 303926 75042 303930 75352
rect 303930 75042 304240 75352
rect 304240 75042 304244 75352
rect 303926 75038 304244 75042
rect -2006 73722 -1806 73922
rect 303926 72352 304244 72356
rect 303926 72042 303930 72352
rect 303930 72042 304240 72352
rect 304240 72042 304244 72352
rect 303926 72038 304244 72042
rect -2006 70722 -1806 70922
rect 303926 69352 304244 69356
rect 303926 69042 303930 69352
rect 303930 69042 304240 69352
rect 304240 69042 304244 69352
rect 303926 69038 304244 69042
rect -2006 67722 -1806 67922
rect 303926 66352 304244 66356
rect 303926 66042 303930 66352
rect 303930 66042 304240 66352
rect 304240 66042 304244 66352
rect 303926 66038 304244 66042
rect -2006 64722 -1806 64922
rect 303926 63352 304244 63356
rect 303926 63042 303930 63352
rect 303930 63042 304240 63352
rect 304240 63042 304244 63352
rect 303926 63038 304244 63042
rect -2006 61722 -1806 61922
rect 303926 60352 304244 60356
rect 303926 60042 303930 60352
rect 303930 60042 304240 60352
rect 304240 60042 304244 60352
rect 303926 60038 304244 60042
rect -2006 58722 -1806 58922
rect 303926 57352 304244 57356
rect 303926 57042 303930 57352
rect 303930 57042 304240 57352
rect 304240 57042 304244 57352
rect 303926 57038 304244 57042
rect -2006 55722 -1806 55922
rect 303926 54352 304244 54356
rect 303926 54042 303930 54352
rect 303930 54042 304240 54352
rect 304240 54042 304244 54352
rect 303926 54038 304244 54042
rect -2006 52722 -1806 52922
rect 303926 51352 304244 51356
rect 303926 51042 303930 51352
rect 303930 51042 304240 51352
rect 304240 51042 304244 51352
rect 303926 51038 304244 51042
rect -2006 49722 -1806 49922
rect 303926 48352 304244 48356
rect 303926 48042 303930 48352
rect 303930 48042 304240 48352
rect 304240 48042 304244 48352
rect 303926 48038 304244 48042
rect -2006 46722 -1806 46922
rect 303926 45352 304244 45356
rect 303926 45042 303930 45352
rect 303930 45042 304240 45352
rect 304240 45042 304244 45352
rect 303926 45038 304244 45042
rect -2006 43722 -1806 43922
rect 303926 42352 304244 42356
rect 303926 42042 303930 42352
rect 303930 42042 304240 42352
rect 304240 42042 304244 42352
rect 303926 42038 304244 42042
rect -2006 40722 -1806 40922
rect 303926 39352 304244 39356
rect 303926 39042 303930 39352
rect 303930 39042 304240 39352
rect 304240 39042 304244 39352
rect 303926 39038 304244 39042
rect -2006 37722 -1806 37922
rect 303926 36352 304244 36356
rect 303926 36042 303930 36352
rect 303930 36042 304240 36352
rect 304240 36042 304244 36352
rect 303926 36038 304244 36042
rect -2006 34722 -1806 34922
rect 303926 33352 304244 33356
rect 303926 33042 303930 33352
rect 303930 33042 304240 33352
rect 304240 33042 304244 33352
rect 303926 33038 304244 33042
rect -2006 31722 -1806 31922
rect 303926 30352 304244 30356
rect 303926 30042 303930 30352
rect 303930 30042 304240 30352
rect 304240 30042 304244 30352
rect 303926 30038 304244 30042
rect -2006 28722 -1806 28922
rect 303926 27352 304244 27356
rect 303926 27042 303930 27352
rect 303930 27042 304240 27352
rect 304240 27042 304244 27352
rect 303926 27038 304244 27042
rect -2006 25722 -1806 25922
rect 303926 24352 304244 24356
rect 303926 24042 303930 24352
rect 303930 24042 304240 24352
rect 304240 24042 304244 24352
rect 303926 24038 304244 24042
rect -2006 22722 -1806 22922
rect 303926 21352 304244 21356
rect 303926 21042 303930 21352
rect 303930 21042 304240 21352
rect 304240 21042 304244 21352
rect 303926 21038 304244 21042
rect 19870 19188 20088 19192
rect 19870 18978 19874 19188
rect 19874 18978 20084 19188
rect 20084 18978 20088 19188
rect 19870 18974 20088 18978
rect 5328 18780 5546 18784
rect 3664 18754 3982 18758
rect 3664 18444 3668 18754
rect 3668 18444 3978 18754
rect 3978 18444 3982 18754
rect 3664 18440 3982 18444
rect 5328 18570 5332 18780
rect 5332 18570 5542 18780
rect 5542 18570 5546 18780
rect 5328 18566 5546 18570
rect 7482 18886 7700 18890
rect 7482 18676 7486 18886
rect 7486 18676 7696 18886
rect 7696 18676 7700 18886
rect 7482 18672 7700 18676
rect 10712 18830 10930 18834
rect 10712 18620 10716 18830
rect 10716 18620 10926 18830
rect 10926 18620 10930 18830
rect 13802 18924 14020 18928
rect 13802 18714 13806 18924
rect 13806 18714 14016 18924
rect 14016 18714 14020 18924
rect 13802 18710 14020 18714
rect 10712 18616 10930 18620
rect 16912 18812 17130 18816
rect 16912 18602 16916 18812
rect 16916 18602 17126 18812
rect 17126 18602 17130 18812
rect 25944 19006 26162 19010
rect 25944 18796 25948 19006
rect 25948 18796 26158 19006
rect 26158 18796 26162 19006
rect 29084 18842 29302 19060
rect 32328 18982 32546 18986
rect 25944 18792 26162 18796
rect 32328 18772 32332 18982
rect 32332 18772 32542 18982
rect 32542 18772 32546 18982
rect 32328 18768 32546 18772
rect 35328 19050 35546 19054
rect 35328 18840 35332 19050
rect 35332 18840 35542 19050
rect 35542 18840 35546 19050
rect 35328 18836 35546 18840
rect 38328 19214 38546 19218
rect 38328 19004 38332 19214
rect 38332 19004 38542 19214
rect 38542 19004 38546 19214
rect 38328 19000 38546 19004
rect 16912 18598 17130 18602
rect 18088 18754 18406 18758
rect 18088 18444 18092 18754
rect 18092 18444 18402 18754
rect 18402 18444 18406 18754
rect 18088 18440 18406 18444
rect 22898 18654 23116 18658
rect 22898 18444 22902 18654
rect 22902 18444 23112 18654
rect 23112 18444 23116 18654
rect 22898 18440 23116 18444
rect 32914 18754 33232 18758
rect 32914 18444 32918 18754
rect 32918 18444 33228 18754
rect 33228 18444 33232 18754
rect 32914 18440 33232 18444
rect 41328 18868 41546 18872
rect 41328 18658 41332 18868
rect 41332 18658 41542 18868
rect 41542 18658 41546 18868
rect 41328 18654 41546 18658
rect 44328 18918 44546 18922
rect 44328 18708 44332 18918
rect 44332 18708 44542 18918
rect 44542 18708 44546 18918
rect 44328 18704 44546 18708
rect 47328 19126 47546 19130
rect 47328 18916 47332 19126
rect 47332 18916 47542 19126
rect 47542 18916 47546 19126
rect 47328 18912 47546 18916
rect 50516 19006 50734 19010
rect 50516 18796 50520 19006
rect 50520 18796 50730 19006
rect 50730 18796 50734 19006
rect 50516 18792 50734 18796
rect 53538 19038 53756 19042
rect 53538 18828 53542 19038
rect 53542 18828 53752 19038
rect 53752 18828 53756 19038
rect 56616 19158 56834 19162
rect 56616 18948 56620 19158
rect 56620 18948 56830 19158
rect 56830 18948 56834 19158
rect 56616 18944 56834 18948
rect 65742 18876 65960 18880
rect 53538 18824 53756 18828
rect 59630 18862 59848 18866
rect 59630 18652 59634 18862
rect 59634 18652 59844 18862
rect 59844 18652 59848 18862
rect 59630 18648 59848 18652
rect 62632 18786 62850 18790
rect 62632 18576 62636 18786
rect 62636 18576 62846 18786
rect 62846 18576 62850 18786
rect 62632 18572 62850 18576
rect 64256 18754 64574 18758
rect 64256 18444 64260 18754
rect 64260 18444 64570 18754
rect 64570 18444 64574 18754
rect 64256 18440 64574 18444
rect 65742 18666 65746 18876
rect 65746 18666 65956 18876
rect 65956 18666 65960 18876
rect 65742 18662 65960 18666
rect 68328 18734 68546 18952
rect 71928 18842 72146 19060
rect 75078 19026 75296 19030
rect 75078 18816 75082 19026
rect 75082 18816 75292 19026
rect 75292 18816 75296 19026
rect 75078 18812 75296 18816
rect 81190 18706 81408 18904
rect 81190 18686 81194 18706
rect 81194 18686 81404 18706
rect 81404 18686 81408 18706
rect 2328 18434 2546 18438
rect 2328 18224 2332 18434
rect 2332 18224 2542 18434
rect 2542 18224 2546 18434
rect 2328 18220 2546 18224
rect 90412 18832 90630 18836
rect 90412 18622 90416 18832
rect 90416 18622 90626 18832
rect 90626 18622 90630 18832
rect 90412 18618 90630 18622
rect 93556 18788 93774 18792
rect 93556 18578 93560 18788
rect 93560 18578 93770 18788
rect 93770 18578 93774 18788
rect 93556 18574 93774 18578
rect 96454 18870 96672 18874
rect 96454 18660 96458 18870
rect 96458 18660 96668 18870
rect 96668 18660 96672 18870
rect 96454 18656 96672 18660
rect 108902 19028 109120 19032
rect 108902 18818 108906 19028
rect 108906 18818 109116 19028
rect 109116 18818 109120 19028
rect 108902 18814 109120 18818
rect 111948 18930 112166 18934
rect 102712 18736 102930 18740
rect 102712 18526 102716 18736
rect 102716 18526 102926 18736
rect 102926 18526 102930 18736
rect 105676 18750 105894 18754
rect 105676 18540 105680 18750
rect 105680 18540 105890 18750
rect 105890 18540 105894 18750
rect 105676 18536 105894 18540
rect 111948 18720 111952 18930
rect 111952 18720 112162 18930
rect 112162 18720 112166 18930
rect 111948 18716 112166 18720
rect 114954 18980 115172 18984
rect 114954 18770 114958 18980
rect 114958 18770 115168 18980
rect 115168 18770 115172 18980
rect 114954 18766 115172 18770
rect 117968 18972 118186 18976
rect 117968 18762 117972 18972
rect 117972 18762 118182 18972
rect 118182 18762 118186 18972
rect 117968 18758 118186 18762
rect 121150 18860 121368 18864
rect 121150 18650 121154 18860
rect 121154 18650 121364 18860
rect 121364 18650 121368 18860
rect 121150 18646 121368 18650
rect 102712 18522 102930 18526
rect 78098 18088 78316 18306
rect -6204 17746 -6198 17942
rect -6198 17746 -5998 17942
rect -5998 17746 -5994 17942
rect 84274 18184 84492 18402
rect 87336 18310 87554 18314
rect 87336 18100 87340 18310
rect 87340 18100 87550 18310
rect 87550 18100 87554 18310
rect 99598 18496 99816 18500
rect 99598 18286 99602 18496
rect 99602 18286 99812 18496
rect 99812 18286 99816 18496
rect 121678 18754 121996 18758
rect 121678 18444 121682 18754
rect 121682 18444 121992 18754
rect 121992 18444 121996 18754
rect 121678 18440 121996 18444
rect 124118 18632 124336 18850
rect 127242 18938 127460 18942
rect 127242 18728 127246 18938
rect 127246 18728 127456 18938
rect 127456 18728 127460 18938
rect 127242 18724 127460 18728
rect 130250 18808 130468 18812
rect 130250 18598 130254 18808
rect 130254 18598 130464 18808
rect 130464 18598 130468 18808
rect 130250 18594 130468 18598
rect 133412 18648 133630 18866
rect 154792 18854 155010 18858
rect 145578 18838 145796 18842
rect 139552 18596 139770 18600
rect 139552 18386 139556 18596
rect 139556 18386 139766 18596
rect 139766 18386 139770 18596
rect 139552 18382 139770 18386
rect 142600 18664 142818 18668
rect 142600 18454 142604 18664
rect 142604 18454 142814 18664
rect 142814 18454 142818 18664
rect 145578 18628 145582 18838
rect 145582 18628 145792 18838
rect 145792 18628 145796 18838
rect 145578 18624 145796 18628
rect 148754 18838 148972 18842
rect 148754 18628 148758 18838
rect 148758 18628 148968 18838
rect 148968 18628 148972 18838
rect 148754 18624 148972 18628
rect 151772 18770 151990 18774
rect 151772 18560 151776 18770
rect 151776 18560 151986 18770
rect 151986 18560 151990 18770
rect 151772 18556 151990 18560
rect 154792 18644 154796 18854
rect 154796 18644 155006 18854
rect 155006 18644 155010 18854
rect 154792 18640 155010 18644
rect 157844 18992 158062 18996
rect 157844 18782 157848 18992
rect 157848 18782 158058 18992
rect 158058 18782 158062 18992
rect 174366 19130 174584 19134
rect 174366 18920 174370 19130
rect 174370 18920 174580 19130
rect 174580 18920 174584 19130
rect 174366 18916 174584 18920
rect 290328 18950 290546 18954
rect 157844 18778 158062 18782
rect 160886 18754 161104 18758
rect 160886 18544 160890 18754
rect 160890 18544 161100 18754
rect 161100 18544 161104 18754
rect 160886 18540 161104 18544
rect 142600 18450 142818 18454
rect 99598 18282 99816 18286
rect 163238 18454 163456 18458
rect 163238 18244 163242 18454
rect 163242 18244 163452 18454
rect 163452 18244 163456 18454
rect 163238 18240 163456 18244
rect 167548 18754 167866 18758
rect 167548 18444 167552 18754
rect 167552 18444 167862 18754
rect 167862 18444 167866 18754
rect 167548 18440 167866 18444
rect 176328 18808 176546 18812
rect 176328 18598 176332 18808
rect 176332 18598 176542 18808
rect 176542 18598 176546 18808
rect 176328 18594 176546 18598
rect 173082 18484 173300 18488
rect 173082 18274 173086 18484
rect 173086 18274 173296 18484
rect 173296 18274 173300 18484
rect 173082 18270 173300 18274
rect 180548 18754 180866 18758
rect 180548 18444 180552 18754
rect 180552 18444 180862 18754
rect 180862 18444 180866 18754
rect 180548 18440 180866 18444
rect 189548 18754 189866 18758
rect 189548 18444 189552 18754
rect 189552 18444 189862 18754
rect 189862 18444 189866 18754
rect 189548 18440 189866 18444
rect 198548 18754 198866 18758
rect 198548 18444 198552 18754
rect 198552 18444 198862 18754
rect 198862 18444 198866 18754
rect 198548 18440 198866 18444
rect 204548 18754 204866 18758
rect 204548 18444 204552 18754
rect 204552 18444 204862 18754
rect 204862 18444 204866 18754
rect 204548 18440 204866 18444
rect 206328 18450 206546 18454
rect 206328 18240 206332 18450
rect 206332 18240 206542 18450
rect 206542 18240 206546 18450
rect 87336 18096 87554 18100
rect 136468 18236 136686 18240
rect 136468 18026 136472 18236
rect 136472 18026 136682 18236
rect 136682 18026 136686 18236
rect 136468 18022 136686 18026
rect 206328 18236 206546 18240
rect 211548 18754 211866 18758
rect 211548 18444 211552 18754
rect 211552 18444 211862 18754
rect 211862 18444 211866 18754
rect 211548 18440 211866 18444
rect 215328 18558 215546 18562
rect 215328 18348 215332 18558
rect 215332 18348 215542 18558
rect 215542 18348 215546 18558
rect 215328 18344 215546 18348
rect 223548 18754 223866 18758
rect 223548 18444 223552 18754
rect 223552 18444 223862 18754
rect 223862 18444 223866 18754
rect 223548 18440 223866 18444
rect 229658 18934 229876 18938
rect 229658 18724 229662 18934
rect 229662 18724 229872 18934
rect 229872 18724 229876 18934
rect 229658 18720 229876 18724
rect 232548 18754 232866 18758
rect 232548 18444 232552 18754
rect 232552 18444 232862 18754
rect 232862 18444 232866 18754
rect 232548 18440 232866 18444
rect 233328 18684 233546 18688
rect 233328 18474 233332 18684
rect 233332 18474 233542 18684
rect 233542 18474 233546 18684
rect 233328 18470 233546 18474
rect 238548 18754 238866 18758
rect 238548 18444 238552 18754
rect 238552 18444 238862 18754
rect 238862 18444 238866 18754
rect 238548 18440 238866 18444
rect 242328 18566 242546 18570
rect 241672 18530 241890 18534
rect 227194 18424 227412 18428
rect 227194 18214 227198 18424
rect 227198 18214 227408 18424
rect 227408 18214 227412 18424
rect 227194 18210 227412 18214
rect 241672 18320 241676 18530
rect 241676 18320 241886 18530
rect 241886 18320 241890 18530
rect 241672 18316 241890 18320
rect 242328 18356 242332 18566
rect 242332 18356 242542 18566
rect 242542 18356 242546 18566
rect 242328 18352 242546 18356
rect 250548 18754 250866 18758
rect 250548 18444 250552 18754
rect 250552 18444 250862 18754
rect 250862 18444 250866 18754
rect 250548 18440 250866 18444
rect 254328 18696 254546 18700
rect 165928 18170 166146 18174
rect 165928 17960 165932 18170
rect 165932 17960 166142 18170
rect 166142 17960 166146 18170
rect 165928 17956 166146 17960
rect 185328 18032 185546 18036
rect -6204 17742 -5994 17746
rect 182474 17854 182692 17858
rect 182474 17644 182478 17854
rect 182478 17644 182688 17854
rect 182688 17644 182692 17854
rect 182474 17640 182692 17644
rect 185328 17822 185332 18032
rect 185332 17822 185542 18032
rect 185542 17822 185546 18032
rect 185328 17818 185546 17822
rect 196794 17924 197012 17928
rect 196794 17714 196798 17924
rect 196798 17714 197008 17924
rect 197008 17714 197012 17924
rect 196794 17710 197012 17714
rect 200916 17952 201134 17956
rect 200916 17742 200920 17952
rect 200920 17742 201130 17952
rect 201130 17742 201134 17952
rect 213156 18094 213374 18098
rect 213156 17884 213160 18094
rect 213160 17884 213370 18094
rect 213370 17884 213374 18094
rect 234650 18298 234868 18302
rect 234650 18088 234654 18298
rect 234654 18088 234864 18298
rect 234864 18088 234868 18298
rect 234650 18084 234868 18088
rect 253926 18504 254144 18508
rect 253926 18294 253930 18504
rect 253930 18294 254140 18504
rect 254140 18294 254144 18504
rect 253926 18290 254144 18294
rect 254328 18486 254332 18696
rect 254332 18486 254542 18696
rect 254542 18486 254546 18696
rect 254328 18482 254546 18486
rect 263948 18754 264266 18758
rect 263948 18444 263952 18754
rect 263952 18444 264262 18754
rect 264262 18444 264266 18754
rect 263948 18440 264266 18444
rect 269032 18556 269250 18560
rect 269032 18346 269036 18556
rect 269036 18346 269246 18556
rect 269246 18346 269250 18556
rect 269032 18342 269250 18346
rect 269948 18754 270266 18758
rect 269948 18444 269952 18754
rect 269952 18444 270262 18754
rect 270262 18444 270266 18754
rect 269948 18440 270266 18444
rect 272948 18754 273266 18758
rect 272948 18444 272952 18754
rect 272952 18444 273262 18754
rect 273262 18444 273266 18754
rect 272948 18440 273266 18444
rect 275948 18754 276266 18758
rect 275948 18444 275952 18754
rect 275952 18444 276262 18754
rect 276262 18444 276266 18754
rect 275948 18440 276266 18444
rect 279676 18694 279894 18698
rect 279676 18484 279680 18694
rect 279680 18484 279890 18694
rect 279890 18484 279894 18694
rect 279676 18480 279894 18484
rect 281948 18754 282266 18758
rect 281948 18444 281952 18754
rect 281952 18444 282262 18754
rect 282262 18444 282266 18754
rect 281948 18440 282266 18444
rect 285948 18754 286266 18758
rect 285948 18444 285952 18754
rect 285952 18444 286262 18754
rect 286262 18444 286266 18754
rect 285948 18440 286266 18444
rect 290328 18740 290332 18950
rect 290332 18740 290542 18950
rect 290542 18740 290546 18950
rect 290328 18736 290546 18740
rect 305386 19094 305604 19098
rect 305386 18884 305390 19094
rect 305390 18884 305600 19094
rect 305600 18884 305604 19094
rect 305386 18880 305604 18884
rect 293948 18754 294266 18758
rect 293948 18444 293952 18754
rect 293952 18444 294262 18754
rect 294262 18444 294266 18754
rect 293948 18440 294266 18444
rect 296948 18754 297266 18758
rect 296948 18444 296952 18754
rect 296952 18444 297262 18754
rect 297262 18444 297266 18754
rect 296948 18440 297266 18444
rect 299948 18754 300266 18758
rect 299948 18444 299952 18754
rect 299952 18444 300262 18754
rect 300262 18444 300266 18754
rect 299948 18440 300266 18444
rect 302948 18754 303266 18758
rect 302948 18444 302952 18754
rect 302952 18444 303262 18754
rect 303262 18444 303266 18754
rect 302948 18440 303266 18444
rect 269328 18264 269546 18268
rect 261044 18120 261262 18124
rect 213156 17880 213374 17884
rect 240916 18010 241134 18014
rect 240916 17800 240920 18010
rect 240920 17800 241130 18010
rect 241130 17800 241134 18010
rect 240916 17796 241134 17800
rect 261044 17910 261048 18120
rect 261048 17910 261258 18120
rect 261258 17910 261262 18120
rect 261044 17906 261262 17910
rect 269328 18054 269332 18264
rect 269332 18054 269542 18264
rect 269542 18054 269546 18264
rect 269328 18050 269546 18054
rect 278878 18202 279096 18206
rect 278878 17992 278882 18202
rect 278882 17992 279092 18202
rect 279092 17992 279096 18202
rect 278878 17988 279096 17992
rect 284328 18132 284546 18136
rect 265870 17958 266088 17962
rect 200916 17738 201134 17742
rect 188328 17654 188546 17658
rect 188328 17444 188332 17654
rect 188332 17444 188542 17654
rect 188542 17444 188546 17654
rect 188328 17440 188546 17444
rect 207000 17746 207218 17750
rect 207000 17536 207004 17746
rect 207004 17536 207214 17746
rect 207214 17536 207218 17746
rect 207000 17532 207218 17536
rect 221328 17706 221546 17710
rect 221328 17496 221332 17706
rect 221332 17496 221542 17706
rect 221542 17496 221546 17706
rect 221328 17492 221546 17496
rect 249668 17856 249886 17860
rect 249668 17646 249672 17856
rect 249672 17646 249882 17856
rect 249882 17646 249886 17856
rect 249668 17642 249886 17646
rect 265870 17748 265874 17958
rect 265874 17748 266084 17958
rect 266084 17748 266088 17958
rect 265870 17744 266088 17748
rect 284328 17922 284332 18132
rect 284332 17922 284542 18132
rect 284542 17922 284546 18132
rect 284328 17918 284546 17922
rect 292408 18222 292626 18226
rect 292408 18012 292412 18222
rect 292412 18012 292622 18222
rect 292622 18012 292626 18222
rect 292408 18008 292626 18012
rect 299258 17718 299476 17722
rect 168864 17416 169082 17420
rect 168864 17206 168868 17416
rect 168868 17206 169078 17416
rect 169078 17206 169082 17416
rect 277694 17578 277912 17582
rect 277694 17368 277698 17578
rect 277698 17368 277908 17578
rect 277908 17368 277912 17578
rect 277694 17364 277912 17368
rect 286930 17508 287148 17512
rect 286930 17298 286934 17508
rect 286934 17298 287144 17508
rect 287144 17298 287148 17508
rect 299258 17508 299262 17718
rect 299262 17508 299472 17718
rect 299472 17508 299476 17718
rect 299258 17504 299476 17508
rect 286930 17294 287148 17298
rect 168864 17202 169082 17206
rect 213904 17264 214122 17268
rect 184010 17148 184228 17152
rect 184010 16938 184014 17148
rect 184014 16938 184224 17148
rect 184224 16938 184228 17148
rect 184010 16934 184228 16938
rect 213904 17054 213908 17264
rect 213908 17054 214118 17264
rect 214118 17054 214122 17264
rect 213904 17050 214122 17054
rect 220688 17224 220906 17228
rect 193466 17014 193684 17018
rect 193466 16804 193470 17014
rect 193470 16804 193680 17014
rect 193680 16804 193684 17014
rect 220688 17014 220692 17224
rect 220692 17014 220902 17224
rect 220902 17014 220906 17224
rect 220688 17010 220906 17014
rect 193466 16800 193684 16804
rect 202004 16890 202222 16894
rect 202004 16680 202008 16890
rect 202008 16680 202218 16890
rect 202218 16680 202222 16890
rect 248712 17072 248930 17076
rect 248712 16862 248716 17072
rect 248716 16862 248926 17072
rect 248926 16862 248930 17072
rect 260054 17242 260272 17246
rect 260054 17032 260058 17242
rect 260058 17032 260268 17242
rect 260268 17032 260272 17242
rect 260054 17028 260272 17032
rect 300252 17100 300470 17104
rect 300252 16890 300256 17100
rect 300256 16890 300466 17100
rect 300466 16890 300470 17100
rect 300252 16886 300470 16890
rect 248712 16858 248930 16862
rect 202004 16676 202222 16680
rect 302942 16094 302946 16410
rect 302946 16094 303268 16410
rect 303268 16094 303274 16410
rect 302942 16088 303274 16094
rect 102 15388 108 15582
rect 108 15388 308 15582
rect 308 15388 312 15582
rect 102 15382 312 15388
rect 3658 15374 3664 15688
rect 3664 15374 3984 15688
rect 3984 15374 3988 15688
rect 18082 15392 18088 15706
rect 18088 15392 18408 15706
rect 18408 15392 18412 15706
rect 18082 15386 18412 15392
rect 3658 15368 3988 15374
rect 32908 15368 32914 15682
rect 32914 15368 33234 15682
rect 33234 15368 33238 15682
rect 32908 15362 33238 15368
rect 64250 15376 64256 15690
rect 64256 15376 64576 15690
rect 64576 15376 64580 15690
rect 121672 15390 121678 15704
rect 121678 15390 121998 15704
rect 121998 15390 122002 15704
rect 121672 15384 122002 15390
rect 167542 15392 167548 15706
rect 167548 15392 167868 15706
rect 167868 15392 167872 15706
rect 167542 15386 167872 15392
rect 180542 15392 180548 15706
rect 180548 15392 180868 15706
rect 180868 15392 180872 15706
rect 180542 15386 180872 15392
rect 189542 15392 189548 15706
rect 189548 15392 189868 15706
rect 189868 15392 189872 15706
rect 189542 15386 189872 15392
rect 198542 15392 198548 15706
rect 198548 15392 198868 15706
rect 198868 15392 198872 15706
rect 198542 15386 198872 15392
rect 204542 15392 204548 15706
rect 204548 15392 204868 15706
rect 204868 15392 204872 15706
rect 204542 15386 204872 15392
rect 211542 15392 211548 15706
rect 211548 15392 211868 15706
rect 211868 15392 211872 15706
rect 211542 15386 211872 15392
rect 223542 15392 223548 15706
rect 223548 15392 223868 15706
rect 223868 15392 223872 15706
rect 223542 15386 223872 15392
rect 232542 15392 232548 15706
rect 232548 15392 232868 15706
rect 232868 15392 232872 15706
rect 232542 15386 232872 15392
rect 238542 15392 238548 15706
rect 238548 15392 238868 15706
rect 238868 15392 238872 15706
rect 238542 15386 238872 15392
rect 250542 15392 250548 15706
rect 250548 15392 250868 15706
rect 250868 15392 250872 15706
rect 250542 15386 250872 15392
rect 263942 15392 263948 15706
rect 263948 15392 264268 15706
rect 264268 15392 264272 15706
rect 263942 15386 264272 15392
rect 269942 15392 269948 15706
rect 269948 15392 270268 15706
rect 270268 15392 270272 15706
rect 269942 15386 270272 15392
rect 272942 15392 272948 15706
rect 272948 15392 273268 15706
rect 273268 15392 273272 15706
rect 272942 15386 273272 15392
rect 275942 15392 275948 15706
rect 275948 15392 276268 15706
rect 276268 15392 276272 15706
rect 275942 15386 276272 15392
rect 281942 15392 281948 15706
rect 281948 15392 282268 15706
rect 282268 15392 282272 15706
rect 281942 15386 282272 15392
rect 285942 15392 285948 15706
rect 285948 15392 286268 15706
rect 286268 15392 286272 15706
rect 285942 15386 286272 15392
rect 293942 15392 293948 15706
rect 293948 15392 294268 15706
rect 294268 15392 294272 15706
rect 293942 15386 294272 15392
rect 296942 15392 296948 15706
rect 296948 15392 297268 15706
rect 297268 15392 297272 15706
rect 296942 15386 297272 15392
rect 299942 15392 299948 15706
rect 299948 15392 300268 15706
rect 300268 15392 300272 15706
rect 299942 15386 300272 15392
rect 302942 15392 302948 15706
rect 302948 15392 303268 15706
rect 303268 15392 303272 15706
rect 302942 15386 303272 15392
rect 64250 15370 64580 15376
<< metal4 >>
rect -7596 325866 -762 325976
rect -5202 322052 -1206 322076
rect -5202 321780 -1502 322052
rect -1230 321780 -1206 322052
rect -5202 321760 -1206 321780
rect -5202 321756 -1526 321760
rect -872 320928 -762 325866
rect 303926 321356 304246 321358
rect 304244 321038 304246 321356
rect -5974 319800 -3762 320120
rect -2674 319722 -2006 319922
rect -1806 319722 -1804 319922
rect -2006 319720 -1804 319722
rect -5202 319052 -1206 319076
rect -5202 318780 -1502 319052
rect -1230 318780 -1206 319052
rect -5202 318760 -1206 318780
rect -5202 318756 -1526 318760
rect 303926 318356 304246 318358
rect 304244 318038 304246 318356
rect -5974 316800 -3762 317120
rect -2674 316722 -2006 316922
rect -1806 316722 -1804 316922
rect -2006 316720 -1804 316722
rect -5202 316052 -1206 316076
rect -5202 315780 -1502 316052
rect -1230 315780 -1206 316052
rect -5202 315760 -1206 315780
rect -5202 315756 -1526 315760
rect 303926 315356 304246 315358
rect 304244 315038 304246 315356
rect -5974 313800 -3762 314120
rect -2674 313722 -2006 313922
rect -1806 313722 -1804 313922
rect -2006 313720 -1804 313722
rect -5202 313052 -1206 313076
rect -5202 312780 -1502 313052
rect -1230 312780 -1206 313052
rect -5202 312760 -1206 312780
rect -5202 312756 -1526 312760
rect 303926 312356 304246 312358
rect 304244 312038 304246 312356
rect -5974 310800 -3762 311120
rect -2674 310722 -2006 310922
rect -1806 310722 -1804 310922
rect -2006 310720 -1804 310722
rect -5202 310052 -1206 310076
rect -5202 309780 -1502 310052
rect -1230 309780 -1206 310052
rect -5202 309760 -1206 309780
rect -5202 309756 -1526 309760
rect 303926 309356 304246 309358
rect 304244 309038 304246 309356
rect -5974 307800 -3762 308120
rect -2674 307722 -2006 307922
rect -1806 307722 -1804 307922
rect -2006 307720 -1804 307722
rect -5202 307052 -1206 307076
rect -5202 306780 -1502 307052
rect -1230 306780 -1206 307052
rect -5202 306760 -1206 306780
rect -5202 306756 -1526 306760
rect 303926 306356 304246 306358
rect 304244 306038 304246 306356
rect -5974 304800 -3762 305120
rect -2674 304722 -2006 304922
rect -1806 304722 -1804 304922
rect -2006 304720 -1804 304722
rect -5202 304052 -1206 304076
rect -5202 303780 -1502 304052
rect -1230 303780 -1206 304052
rect -5202 303760 -1206 303780
rect -5202 303756 -1526 303760
rect 303926 303356 304246 303358
rect 304244 303038 304246 303356
rect -5974 301800 -3762 302120
rect -2674 301722 -2006 301922
rect -1806 301722 -1804 301922
rect -2006 301720 -1804 301722
rect -5202 301052 -1206 301076
rect -5202 300780 -1502 301052
rect -1230 300780 -1206 301052
rect -5202 300760 -1206 300780
rect -5202 300756 -1526 300760
rect 303926 300356 304246 300358
rect 304244 300038 304246 300356
rect -5974 298800 -3762 299120
rect -2674 298722 -2006 298922
rect -1806 298722 -1804 298922
rect -2006 298720 -1804 298722
rect -5202 298052 -1206 298076
rect -5202 297780 -1502 298052
rect -1230 297780 -1206 298052
rect -5202 297760 -1206 297780
rect -5202 297756 -1526 297760
rect 303926 297356 304246 297358
rect 304244 297038 304246 297356
rect -5974 295800 -3762 296120
rect -2674 295722 -2006 295922
rect -1806 295722 -1804 295922
rect -2006 295720 -1804 295722
rect -5202 295052 -1206 295076
rect -5202 294780 -1502 295052
rect -1230 294780 -1206 295052
rect -5202 294760 -1206 294780
rect -5202 294756 -1526 294760
rect 303926 294356 304246 294358
rect 304244 294038 304246 294356
rect -5974 292800 -3762 293120
rect -2674 292722 -2006 292922
rect -1806 292722 -1804 292922
rect -2006 292720 -1804 292722
rect -5202 292052 -1206 292076
rect -5202 291780 -1502 292052
rect -1230 291780 -1206 292052
rect -5202 291760 -1206 291780
rect -5202 291756 -1526 291760
rect 303926 291356 304246 291358
rect 304244 291038 304246 291356
rect -5974 289800 -3762 290120
rect -2674 289722 -2006 289922
rect -1806 289722 -1804 289922
rect -2006 289720 -1804 289722
rect -5202 289052 -1206 289076
rect -5202 288780 -1502 289052
rect -1230 288780 -1206 289052
rect -5202 288760 -1206 288780
rect -5202 288756 -1526 288760
rect 303926 288356 304246 288358
rect 304244 288038 304246 288356
rect -5974 286800 -3762 287120
rect -2674 286722 -2006 286922
rect -1806 286722 -1804 286922
rect -2006 286720 -1804 286722
rect -5202 286052 -1206 286076
rect -5202 285780 -1502 286052
rect -1230 285780 -1206 286052
rect -5202 285760 -1206 285780
rect -5202 285756 -1526 285760
rect 303926 285356 304246 285358
rect 304244 285038 304246 285356
rect -5974 283800 -3762 284120
rect -2674 283722 -2006 283922
rect -1806 283722 -1804 283922
rect -2006 283720 -1804 283722
rect -5202 283052 -1206 283076
rect -5202 282780 -1502 283052
rect -1230 282780 -1206 283052
rect -5202 282760 -1206 282780
rect -5202 282756 -1526 282760
rect 303926 282356 304246 282358
rect 304244 282038 304246 282356
rect -5974 280800 -3762 281120
rect -2674 280722 -2006 280922
rect -1806 280722 -1804 280922
rect -2006 280720 -1804 280722
rect -5202 280052 -1206 280076
rect -5202 279780 -1502 280052
rect -1230 279780 -1206 280052
rect -5202 279760 -1206 279780
rect -5202 279756 -1526 279760
rect 303926 279356 304246 279358
rect 304244 279038 304246 279356
rect -5974 277800 -3762 278120
rect -2674 277722 -2006 277922
rect -1806 277722 -1804 277922
rect -2006 277720 -1804 277722
rect -5202 277052 -1206 277076
rect -5202 276780 -1502 277052
rect -1230 276780 -1206 277052
rect -5202 276760 -1206 276780
rect -5202 276756 -1526 276760
rect 303926 276356 304246 276358
rect 304244 276038 304246 276356
rect -5974 274800 -3762 275120
rect -2674 274722 -2006 274922
rect -1806 274722 -1804 274922
rect -2006 274720 -1804 274722
rect -5202 274052 -1206 274076
rect -5202 273780 -1502 274052
rect -1230 273780 -1206 274052
rect -5202 273760 -1206 273780
rect -5202 273756 -1526 273760
rect 303926 273356 304246 273358
rect 304244 273038 304246 273356
rect -5974 271800 -3762 272120
rect -2674 271722 -2006 271922
rect -1806 271722 -1804 271922
rect -2006 271720 -1804 271722
rect -5202 271052 -1206 271076
rect -5202 270780 -1502 271052
rect -1230 270780 -1206 271052
rect -5202 270760 -1206 270780
rect -5202 270756 -1526 270760
rect 303926 270356 304246 270358
rect 304244 270038 304246 270356
rect -5974 268800 -3762 269120
rect -2674 268722 -2006 268922
rect -1806 268722 -1804 268922
rect -2006 268720 -1804 268722
rect -5202 268052 -1206 268076
rect -5202 267780 -1502 268052
rect -1230 267780 -1206 268052
rect -5202 267760 -1206 267780
rect -5202 267756 -1526 267760
rect 303926 267356 304246 267358
rect 304244 267038 304246 267356
rect -5974 265800 -3762 266120
rect -2674 265722 -2006 265922
rect -1806 265722 -1804 265922
rect -2006 265720 -1804 265722
rect -5202 265052 -1206 265076
rect -5202 264780 -1502 265052
rect -1230 264780 -1206 265052
rect -5202 264760 -1206 264780
rect -5202 264756 -1526 264760
rect 303926 264356 304246 264358
rect 304244 264038 304246 264356
rect -5974 262800 -3762 263120
rect -2674 262722 -2006 262922
rect -1806 262722 -1804 262922
rect -2006 262720 -1804 262722
rect -5202 262052 -1206 262076
rect -5202 261780 -1502 262052
rect -1230 261780 -1206 262052
rect -5202 261760 -1206 261780
rect -5202 261756 -1526 261760
rect 303926 261356 304246 261358
rect 304244 261038 304246 261356
rect -5974 259800 -3762 260120
rect -2674 259722 -2006 259922
rect -1806 259722 -1804 259922
rect -2006 259720 -1804 259722
rect -5202 259052 -1206 259076
rect -5202 258780 -1502 259052
rect -1230 258780 -1206 259052
rect -5202 258760 -1206 258780
rect -5202 258756 -1526 258760
rect 303926 258356 304246 258358
rect 304244 258038 304246 258356
rect -5974 256800 -3762 257120
rect -2674 256722 -2006 256922
rect -1806 256722 -1804 256922
rect -2006 256720 -1804 256722
rect -5202 256052 -1206 256076
rect -5202 255780 -1502 256052
rect -1230 255780 -1206 256052
rect -5202 255760 -1206 255780
rect -5202 255756 -1526 255760
rect 303926 255356 304246 255358
rect 304244 255038 304246 255356
rect -5974 253800 -3762 254120
rect -2674 253722 -2006 253922
rect -1806 253722 -1804 253922
rect -2006 253720 -1804 253722
rect -5202 253052 -1206 253076
rect -5202 252780 -1502 253052
rect -1230 252780 -1206 253052
rect -5202 252760 -1206 252780
rect -5202 252756 -1526 252760
rect 303926 252356 304246 252358
rect 304244 252038 304246 252356
rect -5974 250800 -3762 251120
rect -2674 250722 -2006 250922
rect -1806 250722 -1804 250922
rect -2006 250720 -1804 250722
rect -5202 250052 -1206 250076
rect -5202 249780 -1502 250052
rect -1230 249780 -1206 250052
rect -5202 249760 -1206 249780
rect -5202 249756 -1526 249760
rect 303926 249356 304246 249358
rect 304244 249038 304246 249356
rect -5974 247800 -3762 248120
rect -2674 247722 -2006 247922
rect -1806 247722 -1804 247922
rect -2006 247720 -1804 247722
rect 303926 246356 304246 246358
rect 304244 246038 304246 246356
rect -5974 244800 -3762 245120
rect -2674 244722 -2006 244922
rect -1806 244722 -1804 244922
rect -2006 244720 -1804 244722
rect -5202 244052 -1206 244076
rect -5202 243780 -1502 244052
rect -1230 243780 -1206 244052
rect -5202 243760 -1206 243780
rect -5202 243756 -1526 243760
rect 303926 243356 304246 243358
rect 304244 243038 304246 243356
rect -5974 241800 -3762 242120
rect -2674 241722 -2006 241922
rect -1806 241722 -1804 241922
rect -2006 241720 -1804 241722
rect -5202 241052 -1206 241076
rect -5202 240780 -1502 241052
rect -1230 240780 -1206 241052
rect -5202 240760 -1206 240780
rect -5202 240756 -1526 240760
rect 303926 240356 304246 240358
rect 304244 240038 304246 240356
rect -5974 238800 -3762 239120
rect -2674 238722 -2006 238922
rect -1806 238722 -1804 238922
rect -2006 238720 -1804 238722
rect -5202 238052 -1206 238076
rect -5202 237780 -1502 238052
rect -1230 237780 -1206 238052
rect -5202 237760 -1206 237780
rect -5202 237756 -1526 237760
rect 303926 237356 304246 237358
rect 304244 237038 304246 237356
rect -5974 235800 -3762 236120
rect -2674 235722 -2006 235922
rect -1806 235722 -1804 235922
rect -2006 235720 -1804 235722
rect -5202 235052 -1206 235076
rect -5202 234780 -1502 235052
rect -1230 234780 -1206 235052
rect -5202 234760 -1206 234780
rect -5202 234756 -1526 234760
rect 303926 234356 304246 234358
rect 304244 234038 304246 234356
rect -5974 232800 -3762 233120
rect -2674 232722 -2006 232922
rect -1806 232722 -1804 232922
rect -2006 232720 -1804 232722
rect -5202 232052 -1206 232076
rect -5202 231780 -1502 232052
rect -1230 231780 -1206 232052
rect -5202 231760 -1206 231780
rect -5202 231756 -1526 231760
rect 303926 231356 304246 231358
rect 304244 231038 304246 231356
rect -5974 229800 -3762 230120
rect -2674 229722 -2006 229922
rect -1806 229722 -1804 229922
rect -2006 229720 -1804 229722
rect -5202 229052 -1206 229076
rect -5202 228780 -1502 229052
rect -1230 228780 -1206 229052
rect -5202 228760 -1206 228780
rect -5202 228756 -1526 228760
rect 303926 228356 304246 228358
rect 304244 228038 304246 228356
rect -5974 226800 -3762 227120
rect -2674 226722 -2006 226922
rect -1806 226722 -1804 226922
rect -2006 226720 -1804 226722
rect -5202 226052 -1206 226076
rect -5202 225780 -1502 226052
rect -1230 225780 -1206 226052
rect -5202 225760 -1206 225780
rect -5202 225756 -1526 225760
rect 303926 225356 304246 225358
rect 304244 225038 304246 225356
rect -5974 223800 -3762 224120
rect -2674 223722 -2006 223922
rect -1806 223722 -1804 223922
rect -2006 223720 -1804 223722
rect -5202 223052 -1206 223076
rect -5202 222780 -1502 223052
rect -1230 222780 -1206 223052
rect -5202 222760 -1206 222780
rect -5202 222756 -1526 222760
rect 303926 222356 304246 222358
rect 304244 222038 304246 222356
rect -5974 220800 -3762 221120
rect -2674 220722 -2006 220922
rect -1806 220722 -1804 220922
rect -2006 220720 -1804 220722
rect -5202 220052 -1206 220076
rect -5202 219780 -1502 220052
rect -1230 219780 -1206 220052
rect -5202 219760 -1206 219780
rect -5202 219756 -1526 219760
rect 303926 219356 304246 219358
rect 304244 219038 304246 219356
rect -5974 217800 -3762 218120
rect -2674 217722 -2006 217922
rect -1806 217722 -1804 217922
rect -2006 217720 -1804 217722
rect -5202 217052 -1206 217076
rect -5202 216780 -1502 217052
rect -1230 216780 -1206 217052
rect -5202 216760 -1206 216780
rect -5202 216756 -1526 216760
rect 303926 216356 304246 216358
rect 304244 216038 304246 216356
rect -5974 214800 -3762 215120
rect -2674 214722 -2006 214922
rect -1806 214722 -1804 214922
rect -2006 214720 -1804 214722
rect -5202 214052 -1206 214076
rect -5202 213780 -1502 214052
rect -1230 213780 -1206 214052
rect -5202 213760 -1206 213780
rect -5202 213756 -1526 213760
rect 303926 213356 304246 213358
rect 304244 213038 304246 213356
rect -5974 211800 -3762 212120
rect -2674 211722 -2006 211922
rect -1806 211722 -1804 211922
rect -2006 211720 -1804 211722
rect -5202 211052 -1206 211076
rect -5202 210780 -1502 211052
rect -1230 210780 -1206 211052
rect -5202 210760 -1206 210780
rect -5202 210756 -1526 210760
rect 303926 210356 304246 210358
rect 304244 210038 304246 210356
rect -2674 208722 -2006 208922
rect -1806 208722 -1804 208922
rect -2006 208720 -1804 208722
rect -5202 208052 -1206 208076
rect -5202 207780 -1502 208052
rect -1230 207780 -1206 208052
rect -5202 207760 -1206 207780
rect -5202 207756 -1526 207760
rect 303926 207356 304246 207358
rect 304244 207038 304246 207356
rect -5974 205800 -3762 206120
rect -2674 205722 -2006 205922
rect -1806 205722 -1804 205922
rect -2006 205720 -1804 205722
rect -5202 205052 -1206 205076
rect -5202 204780 -1502 205052
rect -1230 204780 -1206 205052
rect -5202 204760 -1206 204780
rect -5202 204756 -1526 204760
rect 303926 204356 304246 204358
rect 304244 204038 304246 204356
rect -5974 202800 -3762 203120
rect -2674 202722 -2006 202922
rect -1806 202722 -1804 202922
rect -2006 202720 -1804 202722
rect -5202 202052 -1206 202076
rect -5202 201780 -1502 202052
rect -1230 201780 -1206 202052
rect -5202 201760 -1206 201780
rect -5202 201756 -1526 201760
rect 303926 201356 304246 201358
rect 304244 201038 304246 201356
rect -5974 199800 -3762 200120
rect -2674 199722 -2006 199922
rect -1806 199722 -1804 199922
rect -2006 199720 -1804 199722
rect -5202 199052 -1206 199076
rect -5202 198780 -1502 199052
rect -1230 198780 -1206 199052
rect -5202 198760 -1206 198780
rect -5202 198756 -1526 198760
rect 303926 198356 304246 198358
rect 304244 198038 304246 198356
rect -5974 196800 -3762 197120
rect -2674 196722 -2006 196922
rect -1806 196722 -1804 196922
rect -2006 196720 -1804 196722
rect -5202 196052 -1206 196076
rect -5202 195780 -1502 196052
rect -1230 195780 -1206 196052
rect -5202 195760 -1206 195780
rect -5202 195756 -1526 195760
rect 303926 195356 304246 195358
rect 304244 195038 304246 195356
rect -5974 193800 -3762 194120
rect -2674 193722 -2006 193922
rect -1806 193722 -1804 193922
rect -2006 193720 -1804 193722
rect -5202 193052 -1206 193076
rect -5202 192780 -1502 193052
rect -1230 192780 -1206 193052
rect -5202 192760 -1206 192780
rect -5202 192756 -1526 192760
rect 303926 192356 304246 192358
rect 304244 192038 304246 192356
rect -5974 190800 -3762 191120
rect -2674 190722 -2006 190922
rect -1806 190722 -1804 190922
rect -2006 190720 -1804 190722
rect -5202 190052 -1206 190076
rect -5202 189780 -1502 190052
rect -1230 189780 -1206 190052
rect -5202 189760 -1206 189780
rect -5202 189756 -1526 189760
rect 303926 189356 304246 189358
rect 304244 189038 304246 189356
rect -5974 187800 -3762 188120
rect -2674 187722 -2006 187922
rect -1806 187722 -1804 187922
rect -2006 187720 -1804 187722
rect -5202 187052 -1206 187076
rect -5202 186780 -1502 187052
rect -1230 186780 -1206 187052
rect -5202 186760 -1206 186780
rect -5202 186756 -1526 186760
rect 303926 186356 304246 186358
rect 304244 186038 304246 186356
rect -5974 184800 -3762 185120
rect -2674 184722 -2006 184922
rect -1806 184722 -1804 184922
rect -2006 184720 -1804 184722
rect -5202 184052 -1206 184076
rect -5202 183780 -1502 184052
rect -1230 183780 -1206 184052
rect -5202 183760 -1206 183780
rect -5202 183756 -1526 183760
rect 303926 183356 304246 183358
rect 304244 183038 304246 183356
rect -5974 181800 -3762 182120
rect -2674 181722 -2006 181922
rect -1806 181722 -1804 181922
rect -2006 181720 -1804 181722
rect -5202 181052 -1206 181076
rect -5202 180780 -1502 181052
rect -1230 180780 -1206 181052
rect -5202 180760 -1206 180780
rect -5202 180756 -1526 180760
rect 303926 180356 304246 180358
rect 304244 180038 304246 180356
rect -5974 178800 -3762 179120
rect -2674 178722 -2006 178922
rect -1806 178722 -1804 178922
rect -2006 178720 -1804 178722
rect -5202 178052 -1206 178076
rect -5202 177780 -1502 178052
rect -1230 177780 -1206 178052
rect -5202 177760 -1206 177780
rect -5202 177756 -1526 177760
rect 303926 177356 304246 177358
rect 304244 177038 304246 177356
rect -5974 175800 -3762 176120
rect -2674 175722 -2006 175922
rect -1806 175722 -1804 175922
rect -2006 175720 -1804 175722
rect -5202 175052 -1206 175076
rect -5202 174780 -1502 175052
rect -1230 174780 -1206 175052
rect -5202 174760 -1206 174780
rect -5202 174756 -1526 174760
rect 303926 174356 304246 174358
rect 304244 174038 304246 174356
rect -5974 172800 -3762 173120
rect -2674 172722 -2006 172922
rect -1806 172722 -1804 172922
rect -2006 172720 -1804 172722
rect -5202 172052 -1206 172076
rect -5202 171780 -1502 172052
rect -1230 171780 -1206 172052
rect -5202 171760 -1206 171780
rect -5202 171756 -1526 171760
rect 303926 171356 304246 171358
rect 304244 171038 304246 171356
rect -5974 169800 -3762 170120
rect -2674 169722 -2006 169922
rect -1806 169722 -1804 169922
rect -2006 169720 -1804 169722
rect -5202 169052 -1206 169076
rect -5202 168780 -1502 169052
rect -1230 168780 -1206 169052
rect -5202 168760 -1206 168780
rect -5202 168756 -1526 168760
rect 303926 168356 304246 168358
rect 304244 168038 304246 168356
rect -5974 166800 -3762 167120
rect -2674 166722 -2006 166922
rect -1806 166722 -1804 166922
rect -2006 166720 -1804 166722
rect -5202 166052 -1206 166076
rect -5202 165780 -1502 166052
rect -1230 165780 -1206 166052
rect -5202 165760 -1206 165780
rect -5202 165756 -1526 165760
rect 303926 165356 304246 165358
rect 304244 165038 304246 165356
rect -5974 163800 -3762 164120
rect -2674 163722 -2006 163922
rect -1806 163722 -1804 163922
rect -2006 163720 -1804 163722
rect -5202 163052 -1206 163076
rect -5202 162780 -1502 163052
rect -1230 162780 -1206 163052
rect -5202 162760 -1206 162780
rect -5202 162756 -1526 162760
rect 303926 162356 304246 162358
rect 304244 162038 304246 162356
rect -5974 160800 -3762 161120
rect -2674 160722 -2006 160922
rect -1806 160722 -1804 160922
rect -2006 160720 -1804 160722
rect -5202 160052 -1206 160076
rect -5202 159780 -1502 160052
rect -1230 159780 -1206 160052
rect -5202 159760 -1206 159780
rect -5202 159756 -1526 159760
rect 303926 159356 304246 159358
rect 304244 159038 304246 159356
rect -5974 157800 -3762 158120
rect -2674 157722 -2006 157922
rect -1806 157722 -1804 157922
rect -2006 157720 -1804 157722
rect -5202 157052 -1206 157076
rect -5202 156780 -1502 157052
rect -1230 156780 -1206 157052
rect -5202 156760 -1206 156780
rect -5202 156756 -1526 156760
rect 303926 156356 304246 156358
rect 304244 156038 304246 156356
rect -5974 154800 -3762 155120
rect -2674 154722 -2006 154922
rect -1806 154722 -1804 154922
rect -2006 154720 -1804 154722
rect -5202 154052 -1206 154076
rect -5202 153780 -1502 154052
rect -1230 153780 -1206 154052
rect -5202 153760 -1206 153780
rect -5202 153756 -1526 153760
rect 303926 153356 304246 153358
rect 304244 153038 304246 153356
rect -5974 151800 -3762 152120
rect -2674 151722 -2006 151922
rect -1806 151722 -1804 151922
rect -2006 151720 -1804 151722
rect -5202 151052 -1206 151076
rect -5202 150780 -1502 151052
rect -1230 150780 -1206 151052
rect -5202 150760 -1206 150780
rect -5202 150756 -1526 150760
rect 303926 150356 304246 150358
rect 304244 150038 304246 150356
rect -5974 148800 -3762 149120
rect -2674 148722 -2006 148922
rect -1806 148722 -1804 148922
rect -2006 148720 -1804 148722
rect -5202 148052 -1206 148076
rect -5202 147780 -1502 148052
rect -1230 147780 -1206 148052
rect -5202 147760 -1206 147780
rect -5202 147756 -1526 147760
rect 303926 147356 304246 147358
rect 304244 147038 304246 147356
rect -5974 145800 -3762 146120
rect -2674 145722 -2006 145922
rect -1806 145722 -1804 145922
rect -2006 145720 -1804 145722
rect -5202 145052 -1206 145076
rect -5202 144780 -1502 145052
rect -1230 144780 -1206 145052
rect -5202 144760 -1206 144780
rect -5202 144756 -1526 144760
rect 303926 144356 304246 144358
rect 304244 144038 304246 144356
rect -5974 142800 -3762 143120
rect -2674 142722 -2006 142922
rect -1806 142722 -1804 142922
rect -2006 142720 -1804 142722
rect -5202 142052 -1206 142076
rect -5202 141780 -1502 142052
rect -1230 141780 -1206 142052
rect -5202 141760 -1206 141780
rect -5202 141756 -1526 141760
rect 303926 141356 304246 141358
rect 304244 141038 304246 141356
rect -5974 139800 -3762 140120
rect -2674 139722 -2006 139922
rect -1806 139722 -1804 139922
rect -2006 139720 -1804 139722
rect -5202 139052 -1206 139076
rect -5202 138780 -1502 139052
rect -1230 138780 -1206 139052
rect -5202 138760 -1206 138780
rect -5202 138756 -1526 138760
rect 303926 138356 304246 138358
rect 304244 138038 304246 138356
rect -5974 136800 -3762 137120
rect -2674 136722 -2006 136922
rect -1806 136722 -1804 136922
rect -2006 136720 -1804 136722
rect -5202 136052 -1206 136076
rect -5202 135780 -1502 136052
rect -1230 135780 -1206 136052
rect -5202 135760 -1206 135780
rect -5202 135756 -1526 135760
rect 303926 135356 304246 135358
rect 304244 135038 304246 135356
rect -5974 133800 -3762 134120
rect -2674 133722 -2006 133922
rect -1806 133722 -1804 133922
rect -2006 133720 -1804 133722
rect -5202 133052 -1206 133076
rect -5202 132780 -1502 133052
rect -1230 132780 -1206 133052
rect -5202 132760 -1206 132780
rect -5202 132756 -1526 132760
rect 303926 132356 304246 132358
rect 304244 132038 304246 132356
rect -5974 130800 -3762 131120
rect -2674 130722 -2006 130922
rect -1806 130722 -1804 130922
rect -2006 130720 -1804 130722
rect -5202 130052 -1206 130076
rect -5202 129780 -1502 130052
rect -1230 129780 -1206 130052
rect -5202 129760 -1206 129780
rect -5202 129756 -1526 129760
rect 303926 129356 304246 129358
rect 304244 129038 304246 129356
rect -5974 127800 -3762 128120
rect -2674 127722 -2006 127922
rect -1806 127722 -1804 127922
rect -2006 127720 -1804 127722
rect -5202 127052 -1206 127076
rect -5202 126780 -1502 127052
rect -1230 126780 -1206 127052
rect -5202 126760 -1206 126780
rect -5202 126756 -1526 126760
rect 303926 126356 304246 126358
rect 304244 126038 304246 126356
rect -5974 124800 -3762 125120
rect -2674 124722 -2006 124922
rect -1806 124722 -1804 124922
rect -2006 124720 -1804 124722
rect -5202 124052 -1206 124076
rect -5202 123780 -1502 124052
rect -1230 123780 -1206 124052
rect -5202 123760 -1206 123780
rect -5202 123756 -1526 123760
rect 303926 123356 304246 123358
rect 304244 123038 304246 123356
rect -5974 121800 -3762 122120
rect -2674 121722 -2006 121922
rect -1806 121722 -1804 121922
rect -2006 121720 -1804 121722
rect -5202 121052 -1206 121076
rect -5202 120780 -1502 121052
rect -1230 120780 -1206 121052
rect -5202 120760 -1206 120780
rect -5202 120756 -1526 120760
rect 303926 120356 304246 120358
rect 304244 120038 304246 120356
rect -5974 118800 -3762 119120
rect -2674 118722 -2006 118922
rect -1806 118722 -1804 118922
rect -2006 118720 -1804 118722
rect -5202 118052 -1206 118076
rect -5202 117780 -1502 118052
rect -1230 117780 -1206 118052
rect -5202 117760 -1206 117780
rect -5202 117756 -1526 117760
rect 303926 117356 304246 117358
rect 304244 117038 304246 117356
rect -5974 115800 -3762 116120
rect -2674 115722 -2006 115922
rect -1806 115722 -1804 115922
rect -2006 115720 -1804 115722
rect -5202 115052 -1206 115076
rect -5202 114780 -1502 115052
rect -1230 114780 -1206 115052
rect -5202 114760 -1206 114780
rect -5202 114756 -1526 114760
rect 303926 114356 304246 114358
rect 304244 114038 304246 114356
rect -5974 112800 -3762 113120
rect -2674 112722 -2006 112922
rect -1806 112722 -1804 112922
rect -2006 112720 -1804 112722
rect -5202 112052 -1206 112076
rect -5202 111780 -1502 112052
rect -1230 111780 -1206 112052
rect -5202 111760 -1206 111780
rect -5202 111756 -1526 111760
rect 303926 111356 304246 111358
rect 304244 111038 304246 111356
rect -5974 109800 -3762 110120
rect -2674 109722 -2006 109922
rect -1806 109722 -1804 109922
rect -2006 109720 -1804 109722
rect -5202 109052 -1206 109076
rect -5202 108780 -1502 109052
rect -1230 108780 -1206 109052
rect -5202 108760 -1206 108780
rect -5202 108756 -1526 108760
rect 303926 108356 304246 108358
rect 304244 108038 304246 108356
rect -5974 106800 -3762 107120
rect -2674 106722 -2006 106922
rect -1806 106722 -1804 106922
rect -2006 106720 -1804 106722
rect -5202 106052 -1206 106076
rect -5202 105780 -1502 106052
rect -1230 105780 -1206 106052
rect -5202 105760 -1206 105780
rect -5202 105756 -1526 105760
rect 303926 105356 304246 105358
rect 304244 105038 304246 105356
rect -5974 103800 -3762 104120
rect -2674 103722 -2006 103922
rect -1806 103722 -1804 103922
rect -2006 103720 -1804 103722
rect -5202 103052 -1206 103076
rect -5202 102780 -1502 103052
rect -1230 102780 -1206 103052
rect -5202 102760 -1206 102780
rect -5202 102756 -1526 102760
rect 303926 102356 304246 102358
rect 304244 102038 304246 102356
rect -5974 100800 -3762 101120
rect -2674 100722 -2006 100922
rect -1806 100722 -1804 100922
rect -2006 100720 -1804 100722
rect -5202 100052 -1206 100076
rect -5202 99780 -1502 100052
rect -1230 99780 -1206 100052
rect -5202 99760 -1206 99780
rect -5202 99756 -1526 99760
rect 303926 99356 304246 99358
rect 304244 99038 304246 99356
rect -5974 97800 -3762 98120
rect -2674 97722 -2006 97922
rect -1806 97722 -1804 97922
rect -2006 97720 -1804 97722
rect -5202 97052 -1206 97076
rect -5202 96780 -1502 97052
rect -1230 96780 -1206 97052
rect -5202 96760 -1206 96780
rect -5202 96756 -1526 96760
rect 303926 96356 304246 96358
rect 304244 96038 304246 96356
rect -5974 94800 -3762 95120
rect -2674 94722 -2006 94922
rect -1806 94722 -1804 94922
rect -2006 94720 -1804 94722
rect 303926 93356 304246 93358
rect 304244 93038 304246 93356
rect -5974 91800 -3762 92120
rect -2674 91722 -2006 91922
rect -1806 91722 -1804 91922
rect -2006 91720 -1804 91722
rect -5202 91052 -1206 91076
rect -5202 90780 -1502 91052
rect -1230 90780 -1206 91052
rect -5202 90760 -1206 90780
rect -5202 90756 -1526 90760
rect 303926 90356 304246 90358
rect 304244 90038 304246 90356
rect -5974 88800 -3762 89120
rect -2674 88722 -2006 88922
rect -1806 88722 -1804 88922
rect -2006 88720 -1804 88722
rect -5202 88052 -1206 88076
rect -5202 87780 -1502 88052
rect -1230 87780 -1206 88052
rect -5202 87760 -1206 87780
rect -5202 87756 -1526 87760
rect 303926 87356 304246 87358
rect 304244 87038 304246 87356
rect -5974 85800 -3762 86120
rect -2674 85722 -2006 85922
rect -1806 85722 -1804 85922
rect -2006 85720 -1804 85722
rect -5202 85052 -1206 85076
rect -5202 84780 -1502 85052
rect -1230 84780 -1206 85052
rect -5202 84760 -1206 84780
rect -5202 84756 -1526 84760
rect 303926 84356 304246 84358
rect 304244 84038 304246 84356
rect -5974 82800 -3762 83120
rect -2674 82722 -2006 82922
rect -1806 82722 -1804 82922
rect -2006 82720 -1804 82722
rect -5202 82052 -1206 82076
rect -5202 81780 -1502 82052
rect -1230 81780 -1206 82052
rect -5202 81760 -1206 81780
rect -5202 81756 -1526 81760
rect 303926 81356 304246 81358
rect 304244 81038 304246 81356
rect -5974 79800 -3762 80120
rect -2674 79722 -2006 79922
rect -1806 79722 -1804 79922
rect -2006 79720 -1804 79722
rect -5202 79052 -1206 79076
rect -5202 78780 -1502 79052
rect -1230 78780 -1206 79052
rect -5202 78760 -1206 78780
rect -5202 78756 -1526 78760
rect 303926 78356 304246 78358
rect 304244 78038 304246 78356
rect -5974 76800 -3762 77120
rect -2674 76722 -2006 76922
rect -1806 76722 -1804 76922
rect -2006 76720 -1804 76722
rect -5202 76052 -1206 76076
rect -5202 75780 -1502 76052
rect -1230 75780 -1206 76052
rect -5202 75760 -1206 75780
rect -5202 75756 -1526 75760
rect 303926 75356 304246 75358
rect 304244 75038 304246 75356
rect -5974 73800 -3762 74120
rect -2674 73722 -2006 73922
rect -1806 73722 -1804 73922
rect -2006 73720 -1804 73722
rect -5202 73052 -1206 73076
rect -5202 72780 -1502 73052
rect -1230 72780 -1206 73052
rect -5202 72760 -1206 72780
rect -5202 72756 -1526 72760
rect 303926 72356 304246 72358
rect 304244 72038 304246 72356
rect -5974 70800 -3762 71120
rect -2674 70722 -2006 70922
rect -1806 70722 -1804 70922
rect -2006 70720 -1804 70722
rect -5202 70052 -1206 70076
rect -5202 69780 -1502 70052
rect -1230 69780 -1206 70052
rect -5202 69760 -1206 69780
rect -5202 69756 -1526 69760
rect 303926 69356 304246 69358
rect 304244 69038 304246 69356
rect -5974 67800 -3762 68120
rect -2674 67722 -2006 67922
rect -1806 67722 -1804 67922
rect -2006 67720 -1804 67722
rect -5202 67052 -1206 67076
rect -5202 66780 -1502 67052
rect -1230 66780 -1206 67052
rect -5202 66760 -1206 66780
rect -5202 66756 -1526 66760
rect 303926 66356 304246 66358
rect 304244 66038 304246 66356
rect -5974 64800 -3762 65120
rect -2674 64722 -2006 64922
rect -1806 64722 -1804 64922
rect -2006 64720 -1804 64722
rect -5202 64052 -1206 64076
rect -5202 63780 -1502 64052
rect -1230 63780 -1206 64052
rect -5202 63760 -1206 63780
rect -5202 63756 -1526 63760
rect 303926 63356 304246 63358
rect 304244 63038 304246 63356
rect -5974 61800 -3762 62120
rect -2674 61722 -2006 61922
rect -1806 61722 -1804 61922
rect -2006 61720 -1804 61722
rect -5202 61052 -1206 61076
rect -5202 60780 -1502 61052
rect -1230 60780 -1206 61052
rect -5202 60760 -1206 60780
rect -5202 60756 -1526 60760
rect 303926 60356 304246 60358
rect 304244 60038 304246 60356
rect -5974 58800 -3762 59120
rect -2674 58722 -2006 58922
rect -1806 58722 -1804 58922
rect -2006 58720 -1804 58722
rect -5202 58052 -1206 58076
rect -5202 57780 -1502 58052
rect -1230 57780 -1206 58052
rect -5202 57760 -1206 57780
rect -5202 57756 -1526 57760
rect 303926 57356 304246 57358
rect 304244 57038 304246 57356
rect -2674 55722 -2006 55922
rect -1806 55722 -1804 55922
rect -2006 55720 -1804 55722
rect -5202 55052 -1206 55076
rect -5202 54780 -1502 55052
rect -1230 54780 -1206 55052
rect -5202 54760 -1206 54780
rect -5202 54756 -1526 54760
rect 303926 54356 304246 54358
rect 304244 54038 304246 54356
rect -5974 52800 -3762 53120
rect -2674 52722 -2006 52922
rect -1806 52722 -1804 52922
rect -2006 52720 -1804 52722
rect -5202 52052 -1206 52076
rect -5202 51780 -1502 52052
rect -1230 51780 -1206 52052
rect -5202 51760 -1206 51780
rect -5202 51756 -1526 51760
rect 303926 51356 304246 51358
rect 304244 51038 304246 51356
rect -5974 49800 -3762 50120
rect -2674 49722 -2006 49922
rect -1806 49722 -1804 49922
rect -2006 49720 -1804 49722
rect -5202 49052 -1206 49076
rect -5202 48780 -1502 49052
rect -1230 48780 -1206 49052
rect -5202 48760 -1206 48780
rect -5202 48756 -1526 48760
rect 303926 48356 304246 48358
rect 304244 48038 304246 48356
rect -5974 46800 -3762 47120
rect -2674 46722 -2006 46922
rect -1806 46722 -1804 46922
rect -2006 46720 -1804 46722
rect -5202 46052 -1206 46076
rect -5202 45780 -1502 46052
rect -1230 45780 -1206 46052
rect -5202 45760 -1206 45780
rect -5202 45756 -1526 45760
rect 303926 45356 304246 45358
rect 304244 45038 304246 45356
rect -5974 43800 -3762 44120
rect -2674 43722 -2006 43922
rect -1806 43722 -1804 43922
rect -2006 43720 -1804 43722
rect -5202 43052 -1206 43076
rect -5202 42780 -1502 43052
rect -1230 42780 -1206 43052
rect -5202 42760 -1206 42780
rect -5202 42756 -1526 42760
rect 303926 42356 304246 42358
rect 304244 42038 304246 42356
rect -5974 40800 -3762 41120
rect -2674 40722 -2006 40922
rect -1806 40722 -1804 40922
rect -2006 40720 -1804 40722
rect -5202 40052 -1206 40076
rect -5202 39780 -1502 40052
rect -1230 39780 -1206 40052
rect -5202 39760 -1206 39780
rect -5202 39756 -1526 39760
rect 303926 39356 304246 39358
rect 304244 39038 304246 39356
rect -5974 37800 -3762 38120
rect -2674 37722 -2006 37922
rect -1806 37722 -1804 37922
rect -2006 37720 -1804 37722
rect -5202 37052 -1206 37076
rect -5202 36780 -1502 37052
rect -1230 36780 -1206 37052
rect -5202 36760 -1206 36780
rect -5202 36756 -1526 36760
rect 303926 36356 304246 36358
rect 304244 36038 304246 36356
rect -5974 34800 -3762 35120
rect -2674 34722 -2006 34922
rect -1806 34722 -1804 34922
rect -2006 34720 -1804 34722
rect -5202 34052 -1206 34076
rect -5202 33780 -1502 34052
rect -1230 33780 -1206 34052
rect -5202 33760 -1206 33780
rect -5202 33756 -1526 33760
rect 303926 33356 304246 33358
rect 304244 33038 304246 33356
rect -5974 31800 -3762 32120
rect -2674 31722 -2006 31922
rect -1806 31722 -1804 31922
rect -2006 31720 -1804 31722
rect -5202 31052 -1206 31076
rect -5202 30780 -1502 31052
rect -1230 30780 -1206 31052
rect -5202 30760 -1206 30780
rect -5202 30756 -1526 30760
rect 303926 30356 304246 30358
rect 304244 30038 304246 30356
rect -5974 28800 -3762 29120
rect -2674 28722 -2006 28922
rect -1806 28722 -1804 28922
rect -2006 28720 -1804 28722
rect -5202 28052 -1206 28076
rect -5202 27780 -1502 28052
rect -1230 27780 -1206 28052
rect -5202 27760 -1206 27780
rect -5202 27756 -1526 27760
rect 303926 27356 304246 27358
rect 304244 27038 304246 27356
rect -5974 25800 -3762 26120
rect -2674 25722 -2006 25922
rect -1806 25722 -1804 25922
rect -2006 25720 -1804 25722
rect -5202 25052 -1206 25076
rect -5202 24780 -1502 25052
rect -1230 24780 -1206 25052
rect -5202 24760 -1206 24780
rect -5202 24756 -1526 24760
rect 303926 24356 304246 24358
rect 304244 24038 304246 24356
rect -5974 22800 -3762 23120
rect -2674 22722 -2006 22922
rect -1806 22722 -1804 22922
rect -2006 22720 -1804 22722
rect -5202 22052 -1206 22076
rect -5202 21780 -1502 22052
rect -1230 21780 -1206 22052
rect -5202 21760 -1206 21780
rect -5202 21756 -1526 21760
rect 303926 21356 304246 21358
rect 304244 21038 304246 21356
rect -5974 19800 -3762 20120
rect -5202 19052 -1206 19076
rect -5202 18780 -1502 19052
rect -1230 18780 -1206 19052
rect -5202 18760 -1206 18780
rect -780 18794 1738 18904
rect -5202 18756 -1526 18760
rect -5994 17742 -5992 17942
rect -6094 17740 -5992 17742
rect -780 16796 -670 18794
rect 2328 18466 2548 19498
rect 5328 18810 5548 19606
rect 7470 18892 7720 18910
rect 8328 18892 8548 19654
rect 7470 18890 8548 18892
rect 5316 18784 5566 18810
rect 3664 18758 3984 18760
rect 2316 18438 2566 18466
rect 3982 18440 3984 18758
rect 5316 18566 5328 18784
rect 5546 18566 5566 18784
rect 7470 18672 7482 18890
rect 7700 18672 8548 18890
rect 10692 18836 10942 18858
rect 11328 18836 11548 19678
rect 10692 18834 11548 18836
rect 7470 18652 7720 18672
rect 10692 18616 10712 18834
rect 10930 18616 11548 18834
rect 13790 18930 14040 18950
rect 14328 18930 14548 19678
rect 13790 18928 14548 18930
rect 13790 18710 13802 18928
rect 14020 18710 14548 18928
rect 16900 18816 17150 18824
rect 17328 18816 17548 19672
rect 19850 19194 20100 19202
rect 20328 19194 20548 19678
rect 19850 19192 20548 19194
rect 19850 18974 19870 19192
rect 20088 18974 20548 19192
rect 19850 18944 20100 18974
rect 13790 18692 14040 18710
rect 10692 18600 10942 18616
rect 16900 18598 16912 18816
rect 17130 18598 17548 18816
rect 16900 18596 17548 18598
rect 18088 18758 18408 18760
rect 16900 18566 17150 18596
rect 5316 18552 5566 18566
rect 18406 18440 18408 18758
rect 22872 18658 23188 18672
rect 23328 18658 23548 19678
rect 25908 19012 26226 19028
rect 26328 19012 26548 19678
rect 29328 19062 29548 19678
rect 25908 19010 26548 19012
rect 25908 18792 25944 19010
rect 26162 18792 26548 19010
rect 29084 19060 29548 19062
rect 29302 18842 29548 19060
rect 32328 18986 32548 19678
rect 35328 19066 35548 19596
rect 38328 19226 38548 19634
rect 38312 19218 38562 19226
rect 25908 18762 26226 18792
rect 32546 18768 32548 18986
rect 35298 19054 35584 19066
rect 35298 18836 35328 19054
rect 35546 18836 35584 19054
rect 38312 19000 38328 19218
rect 38546 19000 38562 19218
rect 38312 18968 38562 19000
rect 41328 18892 41548 19678
rect 44328 18936 44548 19672
rect 47328 19144 47548 19678
rect 47318 19130 47568 19144
rect 44320 18922 44570 18936
rect 35298 18828 35584 18836
rect 41318 18872 41568 18892
rect 32328 18766 32548 18768
rect 22872 18440 22898 18658
rect 23116 18440 23548 18658
rect 32914 18758 33234 18760
rect 35328 18758 35548 18828
rect 33232 18440 33234 18758
rect 41318 18654 41328 18872
rect 41546 18654 41568 18872
rect 44320 18704 44328 18922
rect 44546 18704 44570 18922
rect 47318 18912 47328 19130
rect 47546 18912 47568 19130
rect 47318 18886 47568 18912
rect 50328 19022 50548 19654
rect 53328 19064 53548 19678
rect 56328 19162 56548 19666
rect 53328 19042 53770 19064
rect 50328 19010 50750 19022
rect 50328 18792 50516 19010
rect 50734 18792 50750 19010
rect 53328 18824 53538 19042
rect 53756 18824 53770 19042
rect 56328 18944 56616 19162
rect 56328 18942 56834 18944
rect 53328 18822 53770 18824
rect 53520 18806 53770 18822
rect 59328 18866 59548 19678
rect 50500 18764 50750 18792
rect 44320 18678 44570 18704
rect 41318 18634 41568 18654
rect 59328 18648 59630 18866
rect 59848 18648 59850 18866
rect 59328 18646 59850 18648
rect 62328 18790 62548 19678
rect 65328 18882 65548 19644
rect 68328 18952 68548 19638
rect 65328 18880 65962 18882
rect 62328 18572 62632 18790
rect 62850 18572 62852 18790
rect 62328 18570 62852 18572
rect 64256 18758 64576 18760
rect 64574 18440 64576 18758
rect 65328 18662 65742 18880
rect 65960 18662 65962 18880
rect 68546 18734 68548 18952
rect 71328 19060 71548 19630
rect 71328 18842 71928 19060
rect 72146 18842 72148 19060
rect 71328 18840 72148 18842
rect 74328 19030 74548 19676
rect 74328 18812 75078 19030
rect 75296 18812 75298 19030
rect 74328 18810 75298 18812
rect 68328 18732 68548 18734
rect 2316 18220 2328 18438
rect 2546 18220 2566 18438
rect 22872 18438 23548 18440
rect 22872 18406 23188 18438
rect 2316 18208 2566 18220
rect 77328 18306 77548 19678
rect 80328 18906 80548 19676
rect 80328 18904 81410 18906
rect 80328 18686 81190 18904
rect 81408 18686 81410 18904
rect 83328 18404 83548 19662
rect 83328 18402 84494 18404
rect 77328 18088 78098 18306
rect 78316 18088 78318 18306
rect 83328 18184 84274 18402
rect 84492 18184 84494 18402
rect 86328 18314 86548 19678
rect 89328 18838 89548 19632
rect 89328 18836 90632 18838
rect 89328 18618 90412 18836
rect 90630 18618 90632 18836
rect 92328 18794 92548 19624
rect 95328 18876 95548 19632
rect 95328 18874 96672 18876
rect 92328 18792 93776 18794
rect 92328 18574 93556 18792
rect 93774 18574 93776 18792
rect 95328 18656 96454 18874
rect 98328 18502 98548 19638
rect 101328 18740 101548 19610
rect 104328 18756 104548 19632
rect 107328 19032 107548 19624
rect 107328 18814 108902 19032
rect 107328 18812 109120 18814
rect 110328 18936 110548 19646
rect 113328 18984 113548 19658
rect 110328 18934 112168 18936
rect 104328 18754 105894 18756
rect 101328 18522 102712 18740
rect 104328 18536 105676 18754
rect 110328 18716 111948 18934
rect 112166 18716 112168 18934
rect 113328 18766 114954 18984
rect 113328 18764 115172 18766
rect 116328 18978 116548 19612
rect 116328 18976 118188 18978
rect 116328 18758 117968 18976
rect 118186 18758 118188 18976
rect 119328 18864 119548 19678
rect 119328 18646 121150 18864
rect 121368 18646 121370 18864
rect 122328 18852 122548 19658
rect 125328 18942 125548 19678
rect 122328 18850 124338 18852
rect 119328 18644 121370 18646
rect 121678 18758 121998 18760
rect 101328 18520 102930 18522
rect 98328 18500 99816 18502
rect 86328 18096 87336 18314
rect 98328 18282 99598 18500
rect 121996 18440 121998 18758
rect 122328 18632 124118 18850
rect 124336 18632 124338 18850
rect 125328 18724 127242 18942
rect 125328 18722 127460 18724
rect 128328 18814 128548 19644
rect 131328 18866 131548 19674
rect 128328 18812 130470 18814
rect 128328 18594 130250 18812
rect 130468 18594 130470 18812
rect 131328 18648 133412 18866
rect 133630 18648 133632 18866
rect 131328 18646 133632 18648
rect 86328 18094 87554 18096
rect 134328 18242 134548 19658
rect 137328 18600 137548 19614
rect 140328 18668 140548 19678
rect 143328 18844 143548 19674
rect 146328 18844 146548 19666
rect 143328 18842 145798 18844
rect 137328 18382 139552 18600
rect 139770 18382 139772 18600
rect 140328 18450 142600 18668
rect 143328 18624 145578 18842
rect 145796 18624 145798 18842
rect 146328 18842 148974 18844
rect 146328 18624 148754 18842
rect 148972 18624 148974 18842
rect 149328 18774 149548 19658
rect 152328 18858 152548 19658
rect 155328 18998 155548 19658
rect 155328 18996 158062 18998
rect 149328 18556 151772 18774
rect 151990 18556 151992 18774
rect 152328 18640 154792 18858
rect 155010 18640 155012 18858
rect 155328 18778 157844 18996
rect 152328 18638 155012 18640
rect 158328 18758 158548 19678
rect 161328 18890 161548 19666
rect 164328 19028 164548 19666
rect 167328 19136 167548 19658
rect 149328 18554 151992 18556
rect 158328 18540 160886 18758
rect 161104 18540 161152 18758
rect 161328 18670 163556 18890
rect 164328 18808 166148 19028
rect 167328 18916 169082 19136
rect 158328 18538 161152 18540
rect 140328 18448 142818 18450
rect 163238 18458 163458 18670
rect 137328 18380 139772 18382
rect 134328 18240 136686 18242
rect 163456 18240 163458 18458
rect 77328 18086 78318 18088
rect 134328 18022 136468 18240
rect 165928 18174 166148 18808
rect 167548 18758 167868 18760
rect 167866 18440 167868 18758
rect 166146 17956 166148 18174
rect 165928 17954 166148 17956
rect 168862 17420 169082 18916
rect 170328 18490 170548 19642
rect 173328 19136 173548 19678
rect 173328 19134 174586 19136
rect 173328 18916 174366 19134
rect 174584 18916 174586 19134
rect 176328 18812 176548 19628
rect 176546 18594 176548 18812
rect 176328 18592 176548 18594
rect 170328 18488 173302 18490
rect 170328 18270 173082 18488
rect 173300 18270 173302 18488
rect 179328 17860 179548 19678
rect 182328 18782 182548 19658
rect 180548 18758 180868 18760
rect 180866 18440 180868 18758
rect 182328 18562 184230 18782
rect 179328 17858 182692 17860
rect 179328 17640 182474 17858
rect 168862 17202 168864 17420
rect 184010 17152 184230 18562
rect 185328 18036 185548 19678
rect 185546 17818 185548 18036
rect 185328 17816 185548 17818
rect 188328 17658 188548 19658
rect 189548 18758 189868 18760
rect 189866 18440 189868 18758
rect 191328 18626 191548 19634
rect 191328 18406 193684 18626
rect 188546 17440 188548 17658
rect 184228 16934 184230 17152
rect 184010 16932 184230 16934
rect 193464 17018 193684 18406
rect 194328 17930 194548 19624
rect 197328 17956 197548 19660
rect 200328 18804 200548 19624
rect 198548 18758 198868 18760
rect 198866 18440 198868 18758
rect 200328 18584 202222 18804
rect 194328 17928 197012 17930
rect 194328 17710 196794 17928
rect 197328 17738 200916 17956
rect 197328 17736 201134 17738
rect 193464 16800 193466 17018
rect 202002 16894 202222 18584
rect 203328 17752 203548 19670
rect 204548 18758 204868 18760
rect 204866 18440 204868 18758
rect 206328 18454 206548 19678
rect 206546 18236 206548 18454
rect 209328 18098 209548 19652
rect 212328 18884 212548 19634
rect 211548 18758 211868 18760
rect 211866 18440 211868 18758
rect 212328 18664 214124 18884
rect 209328 17880 213156 18098
rect 209328 17878 213374 17880
rect 203328 17750 207218 17752
rect 203328 17532 207000 17750
rect 213904 17268 214124 18664
rect 215328 18562 215548 19666
rect 218328 18894 218548 19678
rect 218328 18674 220908 18894
rect 215546 18344 215548 18562
rect 214122 17050 214124 17268
rect 220688 17228 220908 18674
rect 221328 17710 221548 19666
rect 223548 18758 223868 18760
rect 223866 18440 223868 18758
rect 224328 18428 224548 19656
rect 227328 18940 227548 19674
rect 227328 18938 229878 18940
rect 227328 18720 229658 18938
rect 229876 18720 229878 18938
rect 224328 18210 227194 18428
rect 227412 18210 227414 18428
rect 224328 18208 227414 18210
rect 230328 18304 230548 19648
rect 232548 18758 232868 18760
rect 232866 18440 232868 18758
rect 233328 18688 233548 19678
rect 233546 18470 233548 18688
rect 230328 18302 234870 18304
rect 230328 18084 234650 18302
rect 234868 18084 234870 18302
rect 236328 18016 236548 19498
rect 238548 18758 238868 18760
rect 238866 18440 238868 18758
rect 239328 18534 239548 19610
rect 242328 18570 242548 19678
rect 239328 18316 241672 18534
rect 241890 18316 241892 18534
rect 242546 18352 242548 18570
rect 245328 18598 245548 19678
rect 248328 19090 248548 19654
rect 248328 18870 249886 19090
rect 245328 18378 248930 18598
rect 242328 18350 242548 18352
rect 239328 18314 241892 18316
rect 236328 18014 241136 18016
rect 236328 17796 240916 18014
rect 241134 17796 241136 18014
rect 221546 17492 221548 17710
rect 220906 17010 220908 17228
rect 220688 17008 220908 17010
rect 248710 17076 248930 18378
rect 249666 17860 249886 18870
rect 250548 18758 250868 18760
rect 250866 18440 250868 18758
rect 251328 18510 251548 19678
rect 254328 18700 254548 19678
rect 251328 18508 254144 18510
rect 251328 18290 253926 18508
rect 254546 18482 254548 18700
rect 254328 18480 254548 18482
rect 257328 18576 257548 19670
rect 260328 19116 260548 19678
rect 260328 18896 261264 19116
rect 257328 18356 260272 18576
rect 249666 17642 249668 17860
rect 249666 17640 249886 17642
rect -4334 16686 -670 16796
rect -4334 13976 -4224 16686
rect 202002 16676 202004 16894
rect 248710 16858 248712 17076
rect 260052 17246 260272 18356
rect 261044 18124 261264 18896
rect 261262 17906 261264 18124
rect 263328 17964 263548 19678
rect 263948 18758 264268 18760
rect 264266 18440 264268 18758
rect 266328 18560 266548 19620
rect 266328 18342 269032 18560
rect 269250 18342 269252 18560
rect 266328 18340 269252 18342
rect 269328 18268 269548 19594
rect 269948 18758 270268 18760
rect 270266 18440 270268 18758
rect 269546 18050 269548 18268
rect 269328 18048 269548 18050
rect 263328 17962 266146 17964
rect 263328 17744 265870 17962
rect 266088 17744 266146 17962
rect 272328 17582 272548 19648
rect 272948 18758 273268 18760
rect 273266 18440 273268 18758
rect 275328 18206 275548 19648
rect 275948 18758 276268 18760
rect 276266 18440 276268 18758
rect 278328 18698 278548 19670
rect 278328 18480 279676 18698
rect 279894 18480 279896 18698
rect 278328 18478 279896 18480
rect 275328 17988 278878 18206
rect 279096 17988 279098 18206
rect 275328 17986 279098 17988
rect 272328 17364 277694 17582
rect 272328 17362 277912 17364
rect 281328 17512 281548 19678
rect 281948 18758 282268 18760
rect 282266 18440 282268 18758
rect 284328 18136 284548 19678
rect 285948 18758 286268 18760
rect 286266 18440 286268 18758
rect 284546 17918 284548 18136
rect 287328 18228 287548 19670
rect 290328 18954 290548 19678
rect 290546 18736 290548 18954
rect 287328 18226 292626 18228
rect 287328 18008 292408 18226
rect 293328 17724 293548 19642
rect 293948 18758 294268 18760
rect 294266 18440 294268 18758
rect 296328 18328 296548 19654
rect 299328 19100 299548 19678
rect 299328 19098 305604 19100
rect 299328 18880 305386 19098
rect 296948 18758 297268 18760
rect 297266 18440 297268 18758
rect 299948 18758 300268 18760
rect 300266 18440 300268 18758
rect 302948 18758 303268 18760
rect 303266 18440 303268 18758
rect 296328 18108 300470 18328
rect 293328 17722 299478 17724
rect 281328 17294 286930 17512
rect 293328 17504 299258 17722
rect 299476 17504 299478 17722
rect 281328 17292 287148 17294
rect 260052 17028 260054 17246
rect 260052 17026 260272 17028
rect 300250 17104 300470 18108
rect 300250 16886 300252 17104
rect 303866 17264 304186 17288
rect 303866 16992 303890 17264
rect 304162 16992 304186 17264
rect 202002 16674 202222 16676
rect 302940 16410 303274 16412
rect 18082 15706 18414 15708
rect 167542 15706 167874 15708
rect 3658 15688 3990 15690
rect 121672 15704 122004 15706
rect 64250 15690 64582 15692
rect 32908 15682 33240 15684
rect 180542 15706 180874 15708
rect 189542 15706 189874 15708
rect 198542 15706 198874 15708
rect 204542 15706 204874 15708
rect 211542 15706 211874 15708
rect 223542 15706 223874 15708
rect 232542 15706 232874 15708
rect 238542 15706 238874 15708
rect 250542 15706 250874 15708
rect 263942 15706 264274 15708
rect 269942 15706 270274 15708
rect 272942 15706 273274 15708
rect 275942 15706 276274 15708
rect 281942 15706 282274 15708
rect 285942 15706 286274 15708
rect 293942 15706 294274 15708
rect 296942 15706 297274 15708
rect 299942 15706 300274 15708
rect 302942 15706 303274 15708
rect 303866 15692 304186 16992
rect 303682 15396 303866 15668
<< via4 >>
rect -5522 321756 -5202 322076
rect -1502 321780 -1230 322052
rect 302448 324538 302768 324598
rect 302448 324338 302502 324538
rect 302502 324338 302712 324538
rect 302712 324338 302768 324538
rect 302448 324278 302768 324338
rect 303950 321062 304222 321334
rect -6294 319800 -5974 320120
rect -3762 319800 -3442 320120
rect -2994 319662 -2674 319982
rect -5522 318756 -5202 319076
rect -1502 318780 -1230 319052
rect 303950 318062 304222 318334
rect -6294 316800 -5974 317120
rect -3762 316800 -3442 317120
rect -2994 316662 -2674 316982
rect -5522 315756 -5202 316076
rect -1502 315780 -1230 316052
rect 303950 315062 304222 315334
rect -6294 313800 -5974 314120
rect -3762 313800 -3442 314120
rect -2994 313662 -2674 313982
rect -5522 312756 -5202 313076
rect -1502 312780 -1230 313052
rect 303950 312062 304222 312334
rect -6294 310800 -5974 311120
rect -3762 310800 -3442 311120
rect -2994 310662 -2674 310982
rect -5522 309756 -5202 310076
rect -1502 309780 -1230 310052
rect 303950 309062 304222 309334
rect -6294 307800 -5974 308120
rect -3762 307800 -3442 308120
rect -2994 307662 -2674 307982
rect -5522 306756 -5202 307076
rect -1502 306780 -1230 307052
rect 303950 306062 304222 306334
rect -6294 304800 -5974 305120
rect -3762 304800 -3442 305120
rect -2994 304662 -2674 304982
rect -5522 303756 -5202 304076
rect -1502 303780 -1230 304052
rect 303950 303062 304222 303334
rect -6294 301800 -5974 302120
rect -3762 301800 -3442 302120
rect -2994 301662 -2674 301982
rect -5522 300756 -5202 301076
rect -1502 300780 -1230 301052
rect 303950 300062 304222 300334
rect -6294 298800 -5974 299120
rect -3762 298800 -3442 299120
rect -2994 298662 -2674 298982
rect -5522 297756 -5202 298076
rect -1502 297780 -1230 298052
rect 303950 297062 304222 297334
rect -6294 295800 -5974 296120
rect -3762 295800 -3442 296120
rect -2994 295662 -2674 295982
rect -5522 294756 -5202 295076
rect -1502 294780 -1230 295052
rect 303950 294062 304222 294334
rect -6294 292800 -5974 293120
rect -3762 292800 -3442 293120
rect -2994 292662 -2674 292982
rect -5522 291756 -5202 292076
rect -1502 291780 -1230 292052
rect 303950 291062 304222 291334
rect -6294 289800 -5974 290120
rect -3762 289800 -3442 290120
rect -2994 289662 -2674 289982
rect -5522 288756 -5202 289076
rect -1502 288780 -1230 289052
rect 303950 288062 304222 288334
rect -6294 286800 -5974 287120
rect -3762 286800 -3442 287120
rect -2994 286662 -2674 286982
rect -5522 285756 -5202 286076
rect -1502 285780 -1230 286052
rect 303950 285062 304222 285334
rect -6294 283800 -5974 284120
rect -3762 283800 -3442 284120
rect -2994 283662 -2674 283982
rect -5522 282756 -5202 283076
rect -1502 282780 -1230 283052
rect 303950 282062 304222 282334
rect -6294 280800 -5974 281120
rect -3762 280800 -3442 281120
rect -2994 280662 -2674 280982
rect -5522 279756 -5202 280076
rect -1502 279780 -1230 280052
rect 303950 279062 304222 279334
rect -6294 277800 -5974 278120
rect -3762 277800 -3442 278120
rect -2994 277662 -2674 277982
rect -5522 276756 -5202 277076
rect -1502 276780 -1230 277052
rect 303950 276062 304222 276334
rect -6294 274800 -5974 275120
rect -3762 274800 -3442 275120
rect -2994 274662 -2674 274982
rect -5522 273756 -5202 274076
rect -1502 273780 -1230 274052
rect 303950 273062 304222 273334
rect -6294 271800 -5974 272120
rect -3762 271800 -3442 272120
rect -2994 271662 -2674 271982
rect -5522 270756 -5202 271076
rect -1502 270780 -1230 271052
rect 303950 270062 304222 270334
rect -6294 268800 -5974 269120
rect -3762 268800 -3442 269120
rect -2994 268662 -2674 268982
rect -5522 267756 -5202 268076
rect -1502 267780 -1230 268052
rect 303950 267062 304222 267334
rect -6294 265800 -5974 266120
rect -3762 265800 -3442 266120
rect -2994 265662 -2674 265982
rect -5522 264756 -5202 265076
rect -1502 264780 -1230 265052
rect 303950 264062 304222 264334
rect -6294 262800 -5974 263120
rect -3762 262800 -3442 263120
rect -2994 262662 -2674 262982
rect -5522 261756 -5202 262076
rect -1502 261780 -1230 262052
rect 303950 261062 304222 261334
rect -6294 259800 -5974 260120
rect -3762 259800 -3442 260120
rect -2994 259662 -2674 259982
rect -5522 258756 -5202 259076
rect -1502 258780 -1230 259052
rect 303950 258062 304222 258334
rect -6294 256800 -5974 257120
rect -3762 256800 -3442 257120
rect -2994 256662 -2674 256982
rect -5522 255756 -5202 256076
rect -1502 255780 -1230 256052
rect 303950 255062 304222 255334
rect -6294 253800 -5974 254120
rect -3762 253800 -3442 254120
rect -2994 253662 -2674 253982
rect -5522 252756 -5202 253076
rect -1502 252780 -1230 253052
rect 303950 252062 304222 252334
rect -6294 250800 -5974 251120
rect -3762 250800 -3442 251120
rect -2994 250662 -2674 250982
rect -5522 249756 -5202 250076
rect -1502 249780 -1230 250052
rect 303950 249062 304222 249334
rect -6294 247800 -5974 248120
rect -3762 247800 -3442 248120
rect -2994 247662 -2674 247982
rect 303950 246062 304222 246334
rect -6294 244800 -5974 245120
rect -3762 244800 -3442 245120
rect -2994 244662 -2674 244982
rect -5522 243756 -5202 244076
rect -1502 243780 -1230 244052
rect 303950 243062 304222 243334
rect -6294 241800 -5974 242120
rect -3762 241800 -3442 242120
rect -2994 241662 -2674 241982
rect -5522 240756 -5202 241076
rect -1502 240780 -1230 241052
rect 303950 240062 304222 240334
rect -6294 238800 -5974 239120
rect -3762 238800 -3442 239120
rect -2994 238662 -2674 238982
rect -5522 237756 -5202 238076
rect -1502 237780 -1230 238052
rect 303950 237062 304222 237334
rect -6294 235800 -5974 236120
rect -3762 235800 -3442 236120
rect -2994 235662 -2674 235982
rect -5522 234756 -5202 235076
rect -1502 234780 -1230 235052
rect 303950 234062 304222 234334
rect -6294 232800 -5974 233120
rect -3762 232800 -3442 233120
rect -2994 232662 -2674 232982
rect -5522 231756 -5202 232076
rect -1502 231780 -1230 232052
rect 303950 231062 304222 231334
rect -6294 229800 -5974 230120
rect -3762 229800 -3442 230120
rect -2994 229662 -2674 229982
rect -5522 228756 -5202 229076
rect -1502 228780 -1230 229052
rect 303950 228062 304222 228334
rect -6294 226800 -5974 227120
rect -3762 226800 -3442 227120
rect -2994 226662 -2674 226982
rect -5522 225756 -5202 226076
rect -1502 225780 -1230 226052
rect 303950 225062 304222 225334
rect -6294 223800 -5974 224120
rect -3762 223800 -3442 224120
rect -2994 223662 -2674 223982
rect -5522 222756 -5202 223076
rect -1502 222780 -1230 223052
rect 303950 222062 304222 222334
rect -6294 220800 -5974 221120
rect -3762 220800 -3442 221120
rect -2994 220662 -2674 220982
rect -5522 219756 -5202 220076
rect -1502 219780 -1230 220052
rect 303950 219062 304222 219334
rect -6294 217800 -5974 218120
rect -3762 217800 -3442 218120
rect -2994 217662 -2674 217982
rect -5522 216756 -5202 217076
rect -1502 216780 -1230 217052
rect 303950 216062 304222 216334
rect -6294 214800 -5974 215120
rect -3762 214800 -3442 215120
rect -2994 214662 -2674 214982
rect -5522 213756 -5202 214076
rect -1502 213780 -1230 214052
rect 303950 213062 304222 213334
rect -6294 211800 -5974 212120
rect -3762 211800 -3442 212120
rect -2994 211662 -2674 211982
rect -5522 210756 -5202 211076
rect -1502 210780 -1230 211052
rect 303950 210062 304222 210334
rect -2994 208662 -2674 208982
rect -5522 207756 -5202 208076
rect -1502 207780 -1230 208052
rect 303950 207062 304222 207334
rect -6294 205800 -5974 206120
rect -3762 205800 -3442 206120
rect -2994 205662 -2674 205982
rect -5522 204756 -5202 205076
rect -1502 204780 -1230 205052
rect 303950 204062 304222 204334
rect -6294 202800 -5974 203120
rect -3762 202800 -3442 203120
rect -2994 202662 -2674 202982
rect -5522 201756 -5202 202076
rect -1502 201780 -1230 202052
rect 303950 201062 304222 201334
rect -6294 199800 -5974 200120
rect -3762 199800 -3442 200120
rect -2994 199662 -2674 199982
rect -5522 198756 -5202 199076
rect -1502 198780 -1230 199052
rect 303950 198062 304222 198334
rect -6294 196800 -5974 197120
rect -3762 196800 -3442 197120
rect -2994 196662 -2674 196982
rect -5522 195756 -5202 196076
rect -1502 195780 -1230 196052
rect 303950 195062 304222 195334
rect -6294 193800 -5974 194120
rect -3762 193800 -3442 194120
rect -2994 193662 -2674 193982
rect -5522 192756 -5202 193076
rect -1502 192780 -1230 193052
rect 303950 192062 304222 192334
rect -6294 190800 -5974 191120
rect -3762 190800 -3442 191120
rect -2994 190662 -2674 190982
rect -5522 189756 -5202 190076
rect -1502 189780 -1230 190052
rect 303950 189062 304222 189334
rect -6294 187800 -5974 188120
rect -3762 187800 -3442 188120
rect -2994 187662 -2674 187982
rect -5522 186756 -5202 187076
rect -1502 186780 -1230 187052
rect 303950 186062 304222 186334
rect -6294 184800 -5974 185120
rect -3762 184800 -3442 185120
rect -2994 184662 -2674 184982
rect -5522 183756 -5202 184076
rect -1502 183780 -1230 184052
rect 303950 183062 304222 183334
rect -6294 181800 -5974 182120
rect -3762 181800 -3442 182120
rect -2994 181662 -2674 181982
rect -5522 180756 -5202 181076
rect -1502 180780 -1230 181052
rect 303950 180062 304222 180334
rect -6294 178800 -5974 179120
rect -3762 178800 -3442 179120
rect -2994 178662 -2674 178982
rect -5522 177756 -5202 178076
rect -1502 177780 -1230 178052
rect 303950 177062 304222 177334
rect -6294 175800 -5974 176120
rect -3762 175800 -3442 176120
rect -2994 175662 -2674 175982
rect -5522 174756 -5202 175076
rect -1502 174780 -1230 175052
rect 303950 174062 304222 174334
rect -6294 172800 -5974 173120
rect -3762 172800 -3442 173120
rect -2994 172662 -2674 172982
rect -5522 171756 -5202 172076
rect -1502 171780 -1230 172052
rect 303950 171062 304222 171334
rect -6294 169800 -5974 170120
rect -3762 169800 -3442 170120
rect -2994 169662 -2674 169982
rect -5522 168756 -5202 169076
rect -1502 168780 -1230 169052
rect 303950 168062 304222 168334
rect -6294 166800 -5974 167120
rect -3762 166800 -3442 167120
rect -2994 166662 -2674 166982
rect -5522 165756 -5202 166076
rect -1502 165780 -1230 166052
rect 303950 165062 304222 165334
rect -6294 163800 -5974 164120
rect -3762 163800 -3442 164120
rect -2994 163662 -2674 163982
rect -5522 162756 -5202 163076
rect -1502 162780 -1230 163052
rect 303950 162062 304222 162334
rect -6294 160800 -5974 161120
rect -3762 160800 -3442 161120
rect -2994 160662 -2674 160982
rect -5522 159756 -5202 160076
rect -1502 159780 -1230 160052
rect 303950 159062 304222 159334
rect -6294 157800 -5974 158120
rect -3762 157800 -3442 158120
rect -2994 157662 -2674 157982
rect -5522 156756 -5202 157076
rect -1502 156780 -1230 157052
rect 303950 156062 304222 156334
rect -6294 154800 -5974 155120
rect -3762 154800 -3442 155120
rect -2994 154662 -2674 154982
rect -5522 153756 -5202 154076
rect -1502 153780 -1230 154052
rect 303950 153062 304222 153334
rect -6294 151800 -5974 152120
rect -3762 151800 -3442 152120
rect -2994 151662 -2674 151982
rect -5522 150756 -5202 151076
rect -1502 150780 -1230 151052
rect 303950 150062 304222 150334
rect -6294 148800 -5974 149120
rect -3762 148800 -3442 149120
rect -2994 148662 -2674 148982
rect -5522 147756 -5202 148076
rect -1502 147780 -1230 148052
rect 303950 147062 304222 147334
rect -6294 145800 -5974 146120
rect -3762 145800 -3442 146120
rect -2994 145662 -2674 145982
rect -5522 144756 -5202 145076
rect -1502 144780 -1230 145052
rect 303950 144062 304222 144334
rect -6294 142800 -5974 143120
rect -3762 142800 -3442 143120
rect -2994 142662 -2674 142982
rect -5522 141756 -5202 142076
rect -1502 141780 -1230 142052
rect 303950 141062 304222 141334
rect -6294 139800 -5974 140120
rect -3762 139800 -3442 140120
rect -2994 139662 -2674 139982
rect -5522 138756 -5202 139076
rect -1502 138780 -1230 139052
rect 303950 138062 304222 138334
rect -6294 136800 -5974 137120
rect -3762 136800 -3442 137120
rect -2994 136662 -2674 136982
rect -5522 135756 -5202 136076
rect -1502 135780 -1230 136052
rect 303950 135062 304222 135334
rect -6294 133800 -5974 134120
rect -3762 133800 -3442 134120
rect -2994 133662 -2674 133982
rect -5522 132756 -5202 133076
rect -1502 132780 -1230 133052
rect 303950 132062 304222 132334
rect -6294 130800 -5974 131120
rect -3762 130800 -3442 131120
rect -2994 130662 -2674 130982
rect -5522 129756 -5202 130076
rect -1502 129780 -1230 130052
rect 303950 129062 304222 129334
rect -6294 127800 -5974 128120
rect -3762 127800 -3442 128120
rect -2994 127662 -2674 127982
rect -5522 126756 -5202 127076
rect -1502 126780 -1230 127052
rect 303950 126062 304222 126334
rect -6294 124800 -5974 125120
rect -3762 124800 -3442 125120
rect -2994 124662 -2674 124982
rect -5522 123756 -5202 124076
rect -1502 123780 -1230 124052
rect 303950 123062 304222 123334
rect -6294 121800 -5974 122120
rect -3762 121800 -3442 122120
rect -2994 121662 -2674 121982
rect -5522 120756 -5202 121076
rect -1502 120780 -1230 121052
rect 303950 120062 304222 120334
rect -6294 118800 -5974 119120
rect -3762 118800 -3442 119120
rect -2994 118662 -2674 118982
rect -5522 117756 -5202 118076
rect -1502 117780 -1230 118052
rect 303950 117062 304222 117334
rect -6294 115800 -5974 116120
rect -3762 115800 -3442 116120
rect -2994 115662 -2674 115982
rect -5522 114756 -5202 115076
rect -1502 114780 -1230 115052
rect 303950 114062 304222 114334
rect -6294 112800 -5974 113120
rect -3762 112800 -3442 113120
rect -2994 112662 -2674 112982
rect -5522 111756 -5202 112076
rect -1502 111780 -1230 112052
rect 303950 111062 304222 111334
rect -6294 109800 -5974 110120
rect -3762 109800 -3442 110120
rect -2994 109662 -2674 109982
rect -5522 108756 -5202 109076
rect -1502 108780 -1230 109052
rect 303950 108062 304222 108334
rect -6294 106800 -5974 107120
rect -3762 106800 -3442 107120
rect -2994 106662 -2674 106982
rect -5522 105756 -5202 106076
rect -1502 105780 -1230 106052
rect 303950 105062 304222 105334
rect -6294 103800 -5974 104120
rect -3762 103800 -3442 104120
rect -2994 103662 -2674 103982
rect -5522 102756 -5202 103076
rect -1502 102780 -1230 103052
rect 303950 102062 304222 102334
rect -6294 100800 -5974 101120
rect -3762 100800 -3442 101120
rect -2994 100662 -2674 100982
rect -5522 99756 -5202 100076
rect -1502 99780 -1230 100052
rect 303950 99062 304222 99334
rect -6294 97800 -5974 98120
rect -3762 97800 -3442 98120
rect -2994 97662 -2674 97982
rect -5522 96756 -5202 97076
rect -1502 96780 -1230 97052
rect 303950 96062 304222 96334
rect -6294 94800 -5974 95120
rect -3762 94800 -3442 95120
rect -2994 94662 -2674 94982
rect 303950 93062 304222 93334
rect -6294 91800 -5974 92120
rect -3762 91800 -3442 92120
rect -2994 91662 -2674 91982
rect -5522 90756 -5202 91076
rect -1502 90780 -1230 91052
rect 303950 90062 304222 90334
rect -6294 88800 -5974 89120
rect -3762 88800 -3442 89120
rect -2994 88662 -2674 88982
rect -5522 87756 -5202 88076
rect -1502 87780 -1230 88052
rect 303950 87062 304222 87334
rect -6294 85800 -5974 86120
rect -3762 85800 -3442 86120
rect -2994 85662 -2674 85982
rect -5522 84756 -5202 85076
rect -1502 84780 -1230 85052
rect 303950 84062 304222 84334
rect -6294 82800 -5974 83120
rect -3762 82800 -3442 83120
rect -2994 82662 -2674 82982
rect -5522 81756 -5202 82076
rect -1502 81780 -1230 82052
rect 303950 81062 304222 81334
rect -6294 79800 -5974 80120
rect -3762 79800 -3442 80120
rect -2994 79662 -2674 79982
rect -5522 78756 -5202 79076
rect -1502 78780 -1230 79052
rect 303950 78062 304222 78334
rect -6294 76800 -5974 77120
rect -3762 76800 -3442 77120
rect -2994 76662 -2674 76982
rect -5522 75756 -5202 76076
rect -1502 75780 -1230 76052
rect 303950 75062 304222 75334
rect -6294 73800 -5974 74120
rect -3762 73800 -3442 74120
rect -2994 73662 -2674 73982
rect -5522 72756 -5202 73076
rect -1502 72780 -1230 73052
rect 303950 72062 304222 72334
rect -6294 70800 -5974 71120
rect -3762 70800 -3442 71120
rect -2994 70662 -2674 70982
rect -5522 69756 -5202 70076
rect -1502 69780 -1230 70052
rect 303950 69062 304222 69334
rect -6294 67800 -5974 68120
rect -3762 67800 -3442 68120
rect -2994 67662 -2674 67982
rect -5522 66756 -5202 67076
rect -1502 66780 -1230 67052
rect 303950 66062 304222 66334
rect -6294 64800 -5974 65120
rect -3762 64800 -3442 65120
rect -2994 64662 -2674 64982
rect -5522 63756 -5202 64076
rect -1502 63780 -1230 64052
rect 303950 63062 304222 63334
rect -6294 61800 -5974 62120
rect -3762 61800 -3442 62120
rect -2994 61662 -2674 61982
rect -5522 60756 -5202 61076
rect -1502 60780 -1230 61052
rect 303950 60062 304222 60334
rect -6294 58800 -5974 59120
rect -3762 58800 -3442 59120
rect -2994 58662 -2674 58982
rect -5522 57756 -5202 58076
rect -1502 57780 -1230 58052
rect 303950 57062 304222 57334
rect -2994 55662 -2674 55982
rect -5522 54756 -5202 55076
rect -1502 54780 -1230 55052
rect 303950 54062 304222 54334
rect -6294 52800 -5974 53120
rect -3762 52800 -3442 53120
rect -2994 52662 -2674 52982
rect -5522 51756 -5202 52076
rect -1502 51780 -1230 52052
rect 303950 51062 304222 51334
rect -6294 49800 -5974 50120
rect -3762 49800 -3442 50120
rect -2994 49662 -2674 49982
rect -5522 48756 -5202 49076
rect -1502 48780 -1230 49052
rect 303950 48062 304222 48334
rect -6294 46800 -5974 47120
rect -3762 46800 -3442 47120
rect -2994 46662 -2674 46982
rect -5522 45756 -5202 46076
rect -1502 45780 -1230 46052
rect 303950 45062 304222 45334
rect -6294 43800 -5974 44120
rect -3762 43800 -3442 44120
rect -2994 43662 -2674 43982
rect -5522 42756 -5202 43076
rect -1502 42780 -1230 43052
rect 303950 42062 304222 42334
rect -6294 40800 -5974 41120
rect -3762 40800 -3442 41120
rect -2994 40662 -2674 40982
rect -5522 39756 -5202 40076
rect -1502 39780 -1230 40052
rect 303950 39062 304222 39334
rect -6294 37800 -5974 38120
rect -3762 37800 -3442 38120
rect -2994 37662 -2674 37982
rect -5522 36756 -5202 37076
rect -1502 36780 -1230 37052
rect 303950 36062 304222 36334
rect -6294 34800 -5974 35120
rect -3762 34800 -3442 35120
rect -2994 34662 -2674 34982
rect -5522 33756 -5202 34076
rect -1502 33780 -1230 34052
rect 303950 33062 304222 33334
rect -6294 31800 -5974 32120
rect -3762 31800 -3442 32120
rect -2994 31662 -2674 31982
rect -5522 30756 -5202 31076
rect -1502 30780 -1230 31052
rect 303950 30062 304222 30334
rect -6294 28800 -5974 29120
rect -3762 28800 -3442 29120
rect -2994 28662 -2674 28982
rect -5522 27756 -5202 28076
rect -1502 27780 -1230 28052
rect 303950 27062 304222 27334
rect -6294 25800 -5974 26120
rect -3762 25800 -3442 26120
rect -2994 25662 -2674 25982
rect -5522 24756 -5202 25076
rect -1502 24780 -1230 25052
rect 303950 24062 304222 24334
rect -6294 22800 -5974 23120
rect -3762 22800 -3442 23120
rect -2994 22662 -2674 22982
rect -5522 21756 -5202 22076
rect -1502 21780 -1230 22052
rect 303950 21062 304222 21334
rect -6294 19800 -5974 20120
rect -3762 19800 -3442 20120
rect -5522 18756 -5202 19076
rect -1502 18780 -1230 19052
rect -6414 17942 -6094 18002
rect -6414 17742 -6204 17942
rect -6204 17742 -6094 17942
rect -6414 17682 -6094 17742
rect 3688 18464 3960 18736
rect 18112 18464 18384 18736
rect 32938 18464 33210 18736
rect 64280 18464 64552 18736
rect 121702 18464 121974 18736
rect 167572 18464 167844 18736
rect 180572 18464 180844 18736
rect 189572 18464 189844 18736
rect 198572 18464 198844 18736
rect 204572 18464 204844 18736
rect 211572 18464 211844 18736
rect 223572 18464 223844 18736
rect 232572 18464 232844 18736
rect 238572 18464 238844 18736
rect 250572 18464 250844 18736
rect 263972 18464 264244 18736
rect 269972 18464 270244 18736
rect 272972 18464 273244 18736
rect 275972 18464 276244 18736
rect 281972 18464 282244 18736
rect 285972 18464 286244 18736
rect 293972 18464 294244 18736
rect 296972 18464 297244 18736
rect 299972 18464 300244 18736
rect 302972 18464 303244 18736
rect 303890 16992 304162 17264
rect 302940 16088 302942 16410
rect 302942 16088 303274 16410
rect 48 15582 368 15642
rect 48 15382 102 15582
rect 102 15382 312 15582
rect 312 15382 368 15582
rect 48 15322 368 15382
rect 3658 15368 3988 15688
rect 3988 15368 3990 15688
rect 18082 15386 18412 15706
rect 18412 15386 18414 15706
rect 32908 15362 33238 15682
rect 33238 15362 33240 15682
rect 64250 15370 64580 15690
rect 64580 15370 64582 15690
rect 121672 15384 122002 15704
rect 122002 15384 122004 15704
rect 167542 15386 167872 15706
rect 167872 15386 167874 15706
rect 180542 15386 180872 15706
rect 180872 15386 180874 15706
rect 189542 15386 189872 15706
rect 189872 15386 189874 15706
rect 198542 15386 198872 15706
rect 198872 15386 198874 15706
rect 204542 15386 204872 15706
rect 204872 15386 204874 15706
rect 211542 15386 211872 15706
rect 211872 15386 211874 15706
rect 223542 15386 223872 15706
rect 223872 15386 223874 15706
rect 232542 15386 232872 15706
rect 232872 15386 232874 15706
rect 238542 15386 238872 15706
rect 238872 15386 238874 15706
rect 250542 15386 250872 15706
rect 250872 15386 250874 15706
rect 263942 15386 264272 15706
rect 264272 15386 264274 15706
rect 269942 15386 270272 15706
rect 270272 15386 270274 15706
rect 272942 15386 273272 15706
rect 273272 15386 273274 15706
rect 275942 15386 276272 15706
rect 276272 15386 276274 15706
rect 281942 15386 282272 15706
rect 282272 15386 282274 15706
rect 285942 15386 286272 15706
rect 286272 15386 286274 15706
rect 293942 15386 294272 15706
rect 294272 15386 294274 15706
rect 296942 15386 297272 15706
rect 297272 15386 297274 15706
rect 299942 15386 300272 15706
rect 300272 15386 300274 15706
rect 302942 15386 303272 15706
rect 303272 15386 303274 15706
rect 303866 15372 304186 15692
<< metal5 >>
rect -2946 326542 -2626 326564
rect -1526 326542 -1206 326564
rect -2946 326222 305854 326542
rect -5546 322076 -5178 322100
rect -5546 321756 -5522 322076
rect -5202 321756 -5178 322076
rect -5546 321732 -5178 321756
rect -6318 320120 -5950 320144
rect -6318 319800 -6294 320120
rect -5974 319800 -5950 320120
rect -6318 319776 -5950 319800
rect -3786 320120 -3418 320144
rect -2946 320120 -2626 326222
rect -1526 326068 -1206 326222
rect -1526 324636 -1206 324684
rect 302448 324636 302768 324994
rect -1928 324598 304434 324636
rect -1928 324316 302448 324598
rect -3786 319800 -3762 320120
rect -3442 319982 -2626 320120
rect -3442 319800 -2994 319982
rect -3786 319776 -3418 319800
rect -3018 319662 -2994 319800
rect -2674 319662 -2626 319982
rect -3018 319638 -2626 319662
rect -5546 319076 -5178 319100
rect -5546 318756 -5522 319076
rect -5202 318756 -5178 319076
rect -5546 318732 -5178 318756
rect -6318 317120 -5950 317144
rect -6318 316800 -6294 317120
rect -5974 316800 -5950 317120
rect -6318 316776 -5950 316800
rect -3786 317120 -3418 317144
rect -2946 317120 -2626 319638
rect -3786 316800 -3762 317120
rect -3442 316982 -2626 317120
rect -3442 316800 -2994 316982
rect -3786 316776 -3418 316800
rect -3018 316662 -2994 316800
rect -2674 316662 -2626 316982
rect -1526 322052 -1206 324316
rect 302424 324278 302448 324316
rect 302768 324316 304434 324598
rect 302768 324278 302792 324316
rect 302424 324254 302792 324278
rect -1526 321780 -1502 322052
rect -1230 321780 -1206 322052
rect -1526 319052 -1206 321780
rect 303926 321334 304246 324316
rect 303926 321062 303950 321334
rect 304222 321062 304246 321334
rect 288 320218 854 320538
rect -1526 318780 -1502 319052
rect -1230 318780 -1206 319052
rect -1526 316960 -1206 318780
rect -3018 316638 -2626 316662
rect -1528 316640 -1206 316960
rect -5546 316076 -5178 316100
rect -5546 315756 -5522 316076
rect -5202 315756 -5178 316076
rect -5546 315732 -5178 315756
rect -6318 314120 -5950 314144
rect -6318 313800 -6294 314120
rect -5974 313800 -5950 314120
rect -6318 313776 -5950 313800
rect -3786 314120 -3418 314144
rect -2946 314120 -2626 316638
rect -3786 313800 -3762 314120
rect -3442 313982 -2626 314120
rect -3442 313800 -2994 313982
rect -3786 313776 -3418 313800
rect -3018 313662 -2994 313800
rect -2674 313662 -2626 313982
rect -1526 316052 -1206 316640
rect -1526 315780 -1502 316052
rect -1230 315780 -1206 316052
rect -1526 313960 -1206 315780
rect -3018 313638 -2626 313662
rect -1528 313640 -1206 313960
rect -5546 313076 -5178 313100
rect -5546 312756 -5522 313076
rect -5202 312756 -5178 313076
rect -5546 312732 -5178 312756
rect -6318 311120 -5950 311144
rect -6318 310800 -6294 311120
rect -5974 310800 -5950 311120
rect -6318 310776 -5950 310800
rect -3786 311120 -3418 311144
rect -2946 311120 -2626 313638
rect -3786 310800 -3762 311120
rect -3442 310982 -2626 311120
rect -3442 310800 -2994 310982
rect -3786 310776 -3418 310800
rect -3018 310662 -2994 310800
rect -2674 310662 -2626 310982
rect -1526 313052 -1206 313640
rect -1526 312780 -1502 313052
rect -1230 312780 -1206 313052
rect -1526 310960 -1206 312780
rect -3018 310638 -2626 310662
rect -1528 310640 -1206 310960
rect -5546 310076 -5178 310100
rect -5546 309756 -5522 310076
rect -5202 309756 -5178 310076
rect -5546 309732 -5178 309756
rect -6318 308120 -5950 308144
rect -6318 307800 -6294 308120
rect -5974 307800 -5950 308120
rect -6318 307776 -5950 307800
rect -3786 308120 -3418 308144
rect -2946 308120 -2626 310638
rect -3786 307800 -3762 308120
rect -3442 307982 -2626 308120
rect -3442 307800 -2994 307982
rect -3786 307776 -3418 307800
rect -3018 307662 -2994 307800
rect -2674 307662 -2626 307982
rect -1526 310052 -1206 310640
rect -1526 309780 -1502 310052
rect -1230 309780 -1206 310052
rect -1526 307960 -1206 309780
rect -3018 307638 -2626 307662
rect -1528 307640 -1206 307960
rect -5546 307076 -5178 307100
rect -5546 306756 -5522 307076
rect -5202 306756 -5178 307076
rect -5546 306732 -5178 306756
rect -6318 305120 -5950 305144
rect -6318 304800 -6294 305120
rect -5974 304800 -5950 305120
rect -6318 304776 -5950 304800
rect -3786 305120 -3418 305144
rect -2946 305120 -2626 307638
rect -3786 304800 -3762 305120
rect -3442 304982 -2626 305120
rect -3442 304800 -2994 304982
rect -3786 304776 -3418 304800
rect -3018 304662 -2994 304800
rect -2674 304662 -2626 304982
rect -1526 307052 -1206 307640
rect -1526 306780 -1502 307052
rect -1230 306780 -1206 307052
rect -1526 304960 -1206 306780
rect -3018 304638 -2626 304662
rect -1528 304640 -1206 304960
rect -5546 304076 -5178 304100
rect -5546 303756 -5522 304076
rect -5202 303756 -5178 304076
rect -5546 303732 -5178 303756
rect -6318 302120 -5950 302144
rect -6318 301800 -6294 302120
rect -5974 301800 -5950 302120
rect -6318 301776 -5950 301800
rect -3786 302120 -3418 302144
rect -2946 302120 -2626 304638
rect -3786 301800 -3762 302120
rect -3442 301982 -2626 302120
rect -3442 301800 -2994 301982
rect -3786 301776 -3418 301800
rect -3018 301662 -2994 301800
rect -2674 301662 -2626 301982
rect -1526 304052 -1206 304640
rect -1526 303780 -1502 304052
rect -1230 303780 -1206 304052
rect -1526 301960 -1206 303780
rect -3018 301638 -2626 301662
rect -1528 301640 -1206 301960
rect -5546 301076 -5178 301100
rect -5546 300756 -5522 301076
rect -5202 300756 -5178 301076
rect -5546 300732 -5178 300756
rect -6318 299120 -5950 299144
rect -6318 298800 -6294 299120
rect -5974 298800 -5950 299120
rect -6318 298776 -5950 298800
rect -3786 299120 -3418 299144
rect -2946 299120 -2626 301638
rect -3786 298800 -3762 299120
rect -3442 298982 -2626 299120
rect -3442 298800 -2994 298982
rect -3786 298776 -3418 298800
rect -3018 298662 -2994 298800
rect -2674 298662 -2626 298982
rect -1526 301052 -1206 301640
rect -1526 300780 -1502 301052
rect -1230 300780 -1206 301052
rect -1526 298960 -1206 300780
rect -3018 298638 -2626 298662
rect -1528 298640 -1206 298960
rect -5546 298076 -5178 298100
rect -5546 297756 -5522 298076
rect -5202 297756 -5178 298076
rect -5546 297732 -5178 297756
rect -6318 296120 -5950 296144
rect -6318 295800 -6294 296120
rect -5974 295800 -5950 296120
rect -6318 295776 -5950 295800
rect -3786 296120 -3418 296144
rect -2946 296120 -2626 298638
rect -3786 295800 -3762 296120
rect -3442 295982 -2626 296120
rect -3442 295800 -2994 295982
rect -3786 295776 -3418 295800
rect -3018 295662 -2994 295800
rect -2674 295662 -2626 295982
rect -1526 298052 -1206 298640
rect -1526 297780 -1502 298052
rect -1230 297780 -1206 298052
rect -1526 295960 -1206 297780
rect -3018 295638 -2626 295662
rect -1528 295640 -1206 295960
rect -5546 295076 -5178 295100
rect -5546 294756 -5522 295076
rect -5202 294756 -5178 295076
rect -5546 294732 -5178 294756
rect -6318 293120 -5950 293144
rect -6318 292800 -6294 293120
rect -5974 292800 -5950 293120
rect -6318 292776 -5950 292800
rect -3786 293120 -3418 293144
rect -2946 293120 -2626 295638
rect -3786 292800 -3762 293120
rect -3442 292982 -2626 293120
rect -3442 292800 -2994 292982
rect -3786 292776 -3418 292800
rect -3018 292662 -2994 292800
rect -2674 292662 -2626 292982
rect -1526 295052 -1206 295640
rect -1526 294780 -1502 295052
rect -1230 294780 -1206 295052
rect -1526 292960 -1206 294780
rect -3018 292638 -2626 292662
rect -1528 292640 -1206 292960
rect -5546 292076 -5178 292100
rect -5546 291756 -5522 292076
rect -5202 291756 -5178 292076
rect -5546 291732 -5178 291756
rect -6318 290120 -5950 290144
rect -6318 289800 -6294 290120
rect -5974 289800 -5950 290120
rect -6318 289776 -5950 289800
rect -3786 290120 -3418 290144
rect -2946 290120 -2626 292638
rect -3786 289800 -3762 290120
rect -3442 289982 -2626 290120
rect -3442 289800 -2994 289982
rect -3786 289776 -3418 289800
rect -3018 289662 -2994 289800
rect -2674 289662 -2626 289982
rect -1526 292052 -1206 292640
rect -1526 291780 -1502 292052
rect -1230 291780 -1206 292052
rect -1526 289960 -1206 291780
rect -3018 289638 -2626 289662
rect -1528 289640 -1206 289960
rect -5546 289076 -5178 289100
rect -5546 288756 -5522 289076
rect -5202 288756 -5178 289076
rect -5546 288732 -5178 288756
rect -6318 287120 -5950 287144
rect -6318 286800 -6294 287120
rect -5974 286800 -5950 287120
rect -6318 286776 -5950 286800
rect -3786 287120 -3418 287144
rect -2946 287120 -2626 289638
rect -3786 286800 -3762 287120
rect -3442 286982 -2626 287120
rect -3442 286800 -2994 286982
rect -3786 286776 -3418 286800
rect -3018 286662 -2994 286800
rect -2674 286662 -2626 286982
rect -1526 289052 -1206 289640
rect -1526 288780 -1502 289052
rect -1230 288780 -1206 289052
rect -1526 286960 -1206 288780
rect -3018 286638 -2626 286662
rect -1528 286640 -1206 286960
rect -5546 286076 -5178 286100
rect -5546 285756 -5522 286076
rect -5202 285756 -5178 286076
rect -5546 285732 -5178 285756
rect -6318 284120 -5950 284144
rect -6318 283800 -6294 284120
rect -5974 283800 -5950 284120
rect -6318 283776 -5950 283800
rect -3786 284120 -3418 284144
rect -2946 284120 -2626 286638
rect -3786 283800 -3762 284120
rect -3442 283982 -2626 284120
rect -3442 283800 -2994 283982
rect -3786 283776 -3418 283800
rect -3018 283662 -2994 283800
rect -2674 283662 -2626 283982
rect -1526 286052 -1206 286640
rect -1526 285780 -1502 286052
rect -1230 285780 -1206 286052
rect -1526 283960 -1206 285780
rect -3018 283638 -2626 283662
rect -1528 283640 -1206 283960
rect -5546 283076 -5178 283100
rect -5546 282756 -5522 283076
rect -5202 282756 -5178 283076
rect -5546 282732 -5178 282756
rect -6318 281120 -5950 281144
rect -6318 280800 -6294 281120
rect -5974 280800 -5950 281120
rect -6318 280776 -5950 280800
rect -3786 281120 -3418 281144
rect -2946 281120 -2626 283638
rect -3786 280800 -3762 281120
rect -3442 280982 -2626 281120
rect -3442 280800 -2994 280982
rect -3786 280776 -3418 280800
rect -3018 280662 -2994 280800
rect -2674 280662 -2626 280982
rect -1526 283052 -1206 283640
rect -1526 282780 -1502 283052
rect -1230 282780 -1206 283052
rect -1526 280960 -1206 282780
rect -3018 280638 -2626 280662
rect -1528 280640 -1206 280960
rect -5546 280076 -5178 280100
rect -5546 279756 -5522 280076
rect -5202 279756 -5178 280076
rect -5546 279732 -5178 279756
rect -6318 278120 -5950 278144
rect -6318 277800 -6294 278120
rect -5974 277800 -5950 278120
rect -6318 277776 -5950 277800
rect -3786 278120 -3418 278144
rect -2946 278120 -2626 280638
rect -3786 277800 -3762 278120
rect -3442 277982 -2626 278120
rect -3442 277800 -2994 277982
rect -3786 277776 -3418 277800
rect -3018 277662 -2994 277800
rect -2674 277662 -2626 277982
rect -1526 280052 -1206 280640
rect -1526 279780 -1502 280052
rect -1230 279780 -1206 280052
rect -1526 277960 -1206 279780
rect -3018 277638 -2626 277662
rect -1528 277640 -1206 277960
rect -5546 277076 -5178 277100
rect -5546 276756 -5522 277076
rect -5202 276756 -5178 277076
rect -5546 276732 -5178 276756
rect -6318 275120 -5950 275144
rect -6318 274800 -6294 275120
rect -5974 274800 -5950 275120
rect -6318 274776 -5950 274800
rect -3786 275120 -3418 275144
rect -2946 275120 -2626 277638
rect -3786 274800 -3762 275120
rect -3442 274982 -2626 275120
rect -3442 274800 -2994 274982
rect -3786 274776 -3418 274800
rect -3018 274662 -2994 274800
rect -2674 274662 -2626 274982
rect -1526 277052 -1206 277640
rect -1526 276780 -1502 277052
rect -1230 276780 -1206 277052
rect -1526 274960 -1206 276780
rect -3018 274638 -2626 274662
rect -1528 274640 -1206 274960
rect -5546 274076 -5178 274100
rect -5546 273756 -5522 274076
rect -5202 273756 -5178 274076
rect -5546 273732 -5178 273756
rect -6318 272120 -5950 272144
rect -6318 271800 -6294 272120
rect -5974 271800 -5950 272120
rect -6318 271776 -5950 271800
rect -3786 272120 -3418 272144
rect -2946 272120 -2626 274638
rect -3786 271800 -3762 272120
rect -3442 271982 -2626 272120
rect -3442 271800 -2994 271982
rect -3786 271776 -3418 271800
rect -3018 271662 -2994 271800
rect -2674 271662 -2626 271982
rect -1526 274052 -1206 274640
rect -1526 273780 -1502 274052
rect -1230 273780 -1206 274052
rect -1526 271960 -1206 273780
rect -3018 271638 -2626 271662
rect -1528 271640 -1206 271960
rect -5546 271076 -5178 271100
rect -5546 270756 -5522 271076
rect -5202 270756 -5178 271076
rect -5546 270732 -5178 270756
rect -6318 269120 -5950 269144
rect -6318 268800 -6294 269120
rect -5974 268800 -5950 269120
rect -6318 268776 -5950 268800
rect -3786 269120 -3418 269144
rect -2946 269120 -2626 271638
rect -3786 268800 -3762 269120
rect -3442 268982 -2626 269120
rect -3442 268800 -2994 268982
rect -3786 268776 -3418 268800
rect -3018 268662 -2994 268800
rect -2674 268662 -2626 268982
rect -1526 271052 -1206 271640
rect -1526 270780 -1502 271052
rect -1230 270780 -1206 271052
rect -1526 268960 -1206 270780
rect -3018 268638 -2626 268662
rect -1528 268640 -1206 268960
rect -5546 268076 -5178 268100
rect -5546 267756 -5522 268076
rect -5202 267756 -5178 268076
rect -5546 267732 -5178 267756
rect -6318 266120 -5950 266144
rect -6318 265800 -6294 266120
rect -5974 265800 -5950 266120
rect -6318 265776 -5950 265800
rect -3786 266120 -3418 266144
rect -2946 266120 -2626 268638
rect -3786 265800 -3762 266120
rect -3442 265982 -2626 266120
rect -3442 265800 -2994 265982
rect -3786 265776 -3418 265800
rect -3018 265662 -2994 265800
rect -2674 265662 -2626 265982
rect -1526 268052 -1206 268640
rect -1526 267780 -1502 268052
rect -1230 267780 -1206 268052
rect -1526 265960 -1206 267780
rect -3018 265638 -2626 265662
rect -1528 265640 -1206 265960
rect -5546 265076 -5178 265100
rect -5546 264756 -5522 265076
rect -5202 264756 -5178 265076
rect -5546 264732 -5178 264756
rect -6318 263120 -5950 263144
rect -6318 262800 -6294 263120
rect -5974 262800 -5950 263120
rect -6318 262776 -5950 262800
rect -3786 263120 -3418 263144
rect -2946 263120 -2626 265638
rect -3786 262800 -3762 263120
rect -3442 262982 -2626 263120
rect -3442 262800 -2994 262982
rect -3786 262776 -3418 262800
rect -3018 262662 -2994 262800
rect -2674 262662 -2626 262982
rect -1526 265052 -1206 265640
rect -1526 264780 -1502 265052
rect -1230 264780 -1206 265052
rect -1526 262960 -1206 264780
rect -3018 262638 -2626 262662
rect -1528 262640 -1206 262960
rect -5546 262076 -5178 262100
rect -5546 261756 -5522 262076
rect -5202 261756 -5178 262076
rect -5546 261732 -5178 261756
rect -6318 260120 -5950 260144
rect -6318 259800 -6294 260120
rect -5974 259800 -5950 260120
rect -6318 259776 -5950 259800
rect -3786 260120 -3418 260144
rect -2946 260120 -2626 262638
rect -3786 259800 -3762 260120
rect -3442 259982 -2626 260120
rect -3442 259800 -2994 259982
rect -3786 259776 -3418 259800
rect -3018 259662 -2994 259800
rect -2674 259662 -2626 259982
rect -1526 262052 -1206 262640
rect -1526 261780 -1502 262052
rect -1230 261780 -1206 262052
rect -1526 259960 -1206 261780
rect -3018 259638 -2626 259662
rect -1528 259640 -1206 259960
rect -5546 259076 -5178 259100
rect -5546 258756 -5522 259076
rect -5202 258756 -5178 259076
rect -5546 258732 -5178 258756
rect -6318 257120 -5950 257144
rect -6318 256800 -6294 257120
rect -5974 256800 -5950 257120
rect -6318 256776 -5950 256800
rect -3786 257120 -3418 257144
rect -2946 257120 -2626 259638
rect -3786 256800 -3762 257120
rect -3442 256982 -2626 257120
rect -3442 256800 -2994 256982
rect -3786 256776 -3418 256800
rect -3018 256662 -2994 256800
rect -2674 256662 -2626 256982
rect -1526 259052 -1206 259640
rect -1526 258780 -1502 259052
rect -1230 258780 -1206 259052
rect -1526 256960 -1206 258780
rect -3018 256638 -2626 256662
rect -1528 256640 -1206 256960
rect -5546 256076 -5178 256100
rect -5546 255756 -5522 256076
rect -5202 255756 -5178 256076
rect -5546 255732 -5178 255756
rect -6318 254120 -5950 254144
rect -6318 253800 -6294 254120
rect -5974 253800 -5950 254120
rect -6318 253776 -5950 253800
rect -3786 254120 -3418 254144
rect -2946 254120 -2626 256638
rect -3786 253800 -3762 254120
rect -3442 253982 -2626 254120
rect -3442 253800 -2994 253982
rect -3786 253776 -3418 253800
rect -3018 253662 -2994 253800
rect -2674 253662 -2626 253982
rect -1526 256052 -1206 256640
rect -1526 255780 -1502 256052
rect -1230 255780 -1206 256052
rect -1526 253960 -1206 255780
rect -3018 253638 -2626 253662
rect -1528 253640 -1206 253960
rect -5546 253076 -5178 253100
rect -5546 252756 -5522 253076
rect -5202 252756 -5178 253076
rect -5546 252732 -5178 252756
rect -6318 251120 -5950 251144
rect -6318 250800 -6294 251120
rect -5974 250800 -5950 251120
rect -6318 250776 -5950 250800
rect -3786 251120 -3418 251144
rect -2946 251120 -2626 253638
rect -3786 250800 -3762 251120
rect -3442 250982 -2626 251120
rect -3442 250800 -2994 250982
rect -3786 250776 -3418 250800
rect -3018 250662 -2994 250800
rect -2674 250662 -2626 250982
rect -1526 253052 -1206 253640
rect -1526 252780 -1502 253052
rect -1230 252780 -1206 253052
rect -1526 250960 -1206 252780
rect -3018 250638 -2626 250662
rect -1528 250640 -1206 250960
rect -5546 250076 -5178 250100
rect -5546 249756 -5522 250076
rect -5202 249756 -5178 250076
rect -5546 249732 -5178 249756
rect -6318 248120 -5950 248144
rect -6318 247800 -6294 248120
rect -5974 247800 -5950 248120
rect -6318 247776 -5950 247800
rect -3786 248120 -3418 248144
rect -2946 248120 -2626 250638
rect -3786 247800 -3762 248120
rect -3442 247982 -2626 248120
rect -3442 247800 -2994 247982
rect -3786 247776 -3418 247800
rect -3018 247662 -2994 247800
rect -2674 247662 -2626 247982
rect -1526 250052 -1206 250640
rect -1526 249780 -1502 250052
rect -1230 249780 -1206 250052
rect -1526 247960 -1206 249780
rect -3018 247638 -2626 247662
rect -1528 247640 -1206 247960
rect -6318 245120 -5950 245144
rect -6318 244800 -6294 245120
rect -5974 244800 -5950 245120
rect -6318 244776 -5950 244800
rect -3786 245120 -3418 245144
rect -2946 245120 -2626 247638
rect -3786 244800 -3762 245120
rect -3442 244982 -2626 245120
rect -3442 244800 -2994 244982
rect -3786 244776 -3418 244800
rect -3018 244662 -2994 244800
rect -2674 244662 -2626 244982
rect -1526 244960 -1206 247640
rect -3018 244638 -2626 244662
rect -1528 244640 -1206 244960
rect -5546 244076 -5178 244100
rect -5546 243756 -5522 244076
rect -5202 243756 -5178 244076
rect -5546 243732 -5178 243756
rect -6318 242120 -5950 242144
rect -6318 241800 -6294 242120
rect -5974 241800 -5950 242120
rect -6318 241776 -5950 241800
rect -3786 242120 -3418 242144
rect -2946 242120 -2626 244638
rect -3786 241800 -3762 242120
rect -3442 241982 -2626 242120
rect -3442 241800 -2994 241982
rect -3786 241776 -3418 241800
rect -3018 241662 -2994 241800
rect -2674 241662 -2626 241982
rect -1526 244052 -1206 244640
rect -1526 243780 -1502 244052
rect -1230 243780 -1206 244052
rect -1526 241960 -1206 243780
rect -3018 241638 -2626 241662
rect -1528 241640 -1206 241960
rect -5546 241076 -5178 241100
rect -5546 240756 -5522 241076
rect -5202 240756 -5178 241076
rect -5546 240732 -5178 240756
rect -6318 239120 -5950 239144
rect -6318 238800 -6294 239120
rect -5974 238800 -5950 239120
rect -6318 238776 -5950 238800
rect -3786 239120 -3418 239144
rect -2946 239120 -2626 241638
rect -3786 238800 -3762 239120
rect -3442 238982 -2626 239120
rect -3442 238800 -2994 238982
rect -3786 238776 -3418 238800
rect -3018 238662 -2994 238800
rect -2674 238662 -2626 238982
rect -1526 241052 -1206 241640
rect -1526 240780 -1502 241052
rect -1230 240780 -1206 241052
rect -1526 238960 -1206 240780
rect -3018 238638 -2626 238662
rect -1528 238640 -1206 238960
rect -5546 238076 -5178 238100
rect -5546 237756 -5522 238076
rect -5202 237756 -5178 238076
rect -5546 237732 -5178 237756
rect -6318 236120 -5950 236144
rect -6318 235800 -6294 236120
rect -5974 235800 -5950 236120
rect -6318 235776 -5950 235800
rect -3786 236120 -3418 236144
rect -2946 236120 -2626 238638
rect -3786 235800 -3762 236120
rect -3442 235982 -2626 236120
rect -3442 235800 -2994 235982
rect -3786 235776 -3418 235800
rect -3018 235662 -2994 235800
rect -2674 235662 -2626 235982
rect -1526 238052 -1206 238640
rect -1526 237780 -1502 238052
rect -1230 237780 -1206 238052
rect -1526 235960 -1206 237780
rect -3018 235638 -2626 235662
rect -1528 235640 -1206 235960
rect -5546 235076 -5178 235100
rect -5546 234756 -5522 235076
rect -5202 234756 -5178 235076
rect -5546 234732 -5178 234756
rect -6318 233120 -5950 233144
rect -6318 232800 -6294 233120
rect -5974 232800 -5950 233120
rect -6318 232776 -5950 232800
rect -3786 233120 -3418 233144
rect -2946 233120 -2626 235638
rect -3786 232800 -3762 233120
rect -3442 232982 -2626 233120
rect -3442 232800 -2994 232982
rect -3786 232776 -3418 232800
rect -3018 232662 -2994 232800
rect -2674 232662 -2626 232982
rect -1526 235052 -1206 235640
rect -1526 234780 -1502 235052
rect -1230 234780 -1206 235052
rect -1526 232960 -1206 234780
rect -3018 232638 -2626 232662
rect -1528 232640 -1206 232960
rect -5546 232076 -5178 232100
rect -5546 231756 -5522 232076
rect -5202 231756 -5178 232076
rect -5546 231732 -5178 231756
rect -6318 230120 -5950 230144
rect -6318 229800 -6294 230120
rect -5974 229800 -5950 230120
rect -6318 229776 -5950 229800
rect -3786 230120 -3418 230144
rect -2946 230120 -2626 232638
rect -3786 229800 -3762 230120
rect -3442 229982 -2626 230120
rect -3442 229800 -2994 229982
rect -3786 229776 -3418 229800
rect -3018 229662 -2994 229800
rect -2674 229662 -2626 229982
rect -1526 232052 -1206 232640
rect -1526 231780 -1502 232052
rect -1230 231780 -1206 232052
rect -1526 229960 -1206 231780
rect -3018 229638 -2626 229662
rect -1528 229640 -1206 229960
rect -5546 229076 -5178 229100
rect -5546 228756 -5522 229076
rect -5202 228756 -5178 229076
rect -5546 228732 -5178 228756
rect -6318 227120 -5950 227144
rect -6318 226800 -6294 227120
rect -5974 226800 -5950 227120
rect -6318 226776 -5950 226800
rect -3786 227120 -3418 227144
rect -2946 227120 -2626 229638
rect -3786 226800 -3762 227120
rect -3442 226982 -2626 227120
rect -3442 226800 -2994 226982
rect -3786 226776 -3418 226800
rect -3018 226662 -2994 226800
rect -2674 226662 -2626 226982
rect -1526 229052 -1206 229640
rect -1526 228780 -1502 229052
rect -1230 228780 -1206 229052
rect -1526 226960 -1206 228780
rect -3018 226638 -2626 226662
rect -1528 226640 -1206 226960
rect -5546 226076 -5178 226100
rect -5546 225756 -5522 226076
rect -5202 225756 -5178 226076
rect -5546 225732 -5178 225756
rect -6318 224120 -5950 224144
rect -6318 223800 -6294 224120
rect -5974 223800 -5950 224120
rect -6318 223776 -5950 223800
rect -3786 224120 -3418 224144
rect -2946 224120 -2626 226638
rect -3786 223800 -3762 224120
rect -3442 223982 -2626 224120
rect -3442 223800 -2994 223982
rect -3786 223776 -3418 223800
rect -3018 223662 -2994 223800
rect -2674 223662 -2626 223982
rect -1526 226052 -1206 226640
rect -1526 225780 -1502 226052
rect -1230 225780 -1206 226052
rect -1526 223960 -1206 225780
rect -3018 223638 -2626 223662
rect -1528 223640 -1206 223960
rect -5546 223076 -5178 223100
rect -5546 222756 -5522 223076
rect -5202 222756 -5178 223076
rect -5546 222732 -5178 222756
rect -6318 221120 -5950 221144
rect -6318 220800 -6294 221120
rect -5974 220800 -5950 221120
rect -6318 220776 -5950 220800
rect -3786 221120 -3418 221144
rect -2946 221120 -2626 223638
rect -3786 220800 -3762 221120
rect -3442 220982 -2626 221120
rect -3442 220800 -2994 220982
rect -3786 220776 -3418 220800
rect -3018 220662 -2994 220800
rect -2674 220662 -2626 220982
rect -1526 223052 -1206 223640
rect -1526 222780 -1502 223052
rect -1230 222780 -1206 223052
rect -1526 220960 -1206 222780
rect -3018 220638 -2626 220662
rect -1528 220640 -1206 220960
rect -5546 220076 -5178 220100
rect -5546 219756 -5522 220076
rect -5202 219756 -5178 220076
rect -5546 219732 -5178 219756
rect -6318 218120 -5950 218144
rect -6318 217800 -6294 218120
rect -5974 217800 -5950 218120
rect -6318 217776 -5950 217800
rect -3786 218120 -3418 218144
rect -2946 218120 -2626 220638
rect -3786 217800 -3762 218120
rect -3442 217982 -2626 218120
rect -3442 217800 -2994 217982
rect -3786 217776 -3418 217800
rect -3018 217662 -2994 217800
rect -2674 217662 -2626 217982
rect -1526 220052 -1206 220640
rect -1526 219780 -1502 220052
rect -1230 219780 -1206 220052
rect -1526 217960 -1206 219780
rect -3018 217638 -2626 217662
rect -1528 217640 -1206 217960
rect -5546 217076 -5178 217100
rect -5546 216756 -5522 217076
rect -5202 216756 -5178 217076
rect -5546 216732 -5178 216756
rect -6318 215120 -5950 215144
rect -6318 214800 -6294 215120
rect -5974 214800 -5950 215120
rect -6318 214776 -5950 214800
rect -3786 215120 -3418 215144
rect -2946 215120 -2626 217638
rect -3786 214800 -3762 215120
rect -3442 214982 -2626 215120
rect -3442 214800 -2994 214982
rect -3786 214776 -3418 214800
rect -3018 214662 -2994 214800
rect -2674 214662 -2626 214982
rect -1526 217052 -1206 217640
rect -1526 216780 -1502 217052
rect -1230 216780 -1206 217052
rect -1526 214960 -1206 216780
rect -3018 214638 -2626 214662
rect -1528 214640 -1206 214960
rect -5546 214076 -5178 214100
rect -5546 213756 -5522 214076
rect -5202 213756 -5178 214076
rect -5546 213732 -5178 213756
rect -6318 212120 -5950 212144
rect -6318 211800 -6294 212120
rect -5974 211800 -5950 212120
rect -6318 211776 -5950 211800
rect -3786 212120 -3418 212144
rect -2946 212120 -2626 214638
rect -3786 211800 -3762 212120
rect -3442 211982 -2626 212120
rect -3442 211800 -2994 211982
rect -3786 211776 -3418 211800
rect -3018 211662 -2994 211800
rect -2674 211662 -2626 211982
rect -1526 214052 -1206 214640
rect -1526 213780 -1502 214052
rect -1230 213780 -1206 214052
rect -1526 211960 -1206 213780
rect -3018 211638 -2626 211662
rect -1528 211640 -1206 211960
rect -5546 211076 -5178 211100
rect -5546 210756 -5522 211076
rect -5202 210756 -5178 211076
rect -5546 210732 -5178 210756
rect -2946 209120 -2626 211638
rect -3120 208982 -2626 209120
rect -3120 208800 -2994 208982
rect -3018 208662 -2994 208800
rect -2674 208662 -2626 208982
rect -1526 211052 -1206 211640
rect -1526 210780 -1502 211052
rect -1230 210780 -1206 211052
rect -1526 208960 -1206 210780
rect -3018 208638 -2626 208662
rect -1528 208640 -1206 208960
rect -5546 208076 -5178 208100
rect -5546 207756 -5522 208076
rect -5202 207756 -5178 208076
rect -5546 207732 -5178 207756
rect -6318 206120 -5950 206144
rect -6318 205800 -6294 206120
rect -5974 205800 -5950 206120
rect -6318 205776 -5950 205800
rect -3786 206120 -3418 206144
rect -2946 206120 -2626 208638
rect -3786 205800 -3762 206120
rect -3442 205982 -2626 206120
rect -3442 205800 -2994 205982
rect -3786 205776 -3418 205800
rect -3018 205662 -2994 205800
rect -2674 205662 -2626 205982
rect -1526 208052 -1206 208640
rect -1526 207780 -1502 208052
rect -1230 207780 -1206 208052
rect -1526 205960 -1206 207780
rect -3018 205638 -2626 205662
rect -1528 205640 -1206 205960
rect -5546 205076 -5178 205100
rect -5546 204756 -5522 205076
rect -5202 204756 -5178 205076
rect -5546 204732 -5178 204756
rect -6318 203120 -5950 203144
rect -6318 202800 -6294 203120
rect -5974 202800 -5950 203120
rect -6318 202776 -5950 202800
rect -3786 203120 -3418 203144
rect -2946 203120 -2626 205638
rect -3786 202800 -3762 203120
rect -3442 202982 -2626 203120
rect -3442 202800 -2994 202982
rect -3786 202776 -3418 202800
rect -3018 202662 -2994 202800
rect -2674 202662 -2626 202982
rect -1526 205052 -1206 205640
rect -1526 204780 -1502 205052
rect -1230 204780 -1206 205052
rect -1526 202960 -1206 204780
rect -3018 202638 -2626 202662
rect -1528 202640 -1206 202960
rect -5546 202076 -5178 202100
rect -5546 201756 -5522 202076
rect -5202 201756 -5178 202076
rect -5546 201732 -5178 201756
rect -6318 200120 -5950 200144
rect -6318 199800 -6294 200120
rect -5974 199800 -5950 200120
rect -6318 199776 -5950 199800
rect -3786 200120 -3418 200144
rect -2946 200120 -2626 202638
rect -3786 199800 -3762 200120
rect -3442 199982 -2626 200120
rect -3442 199800 -2994 199982
rect -3786 199776 -3418 199800
rect -3018 199662 -2994 199800
rect -2674 199662 -2626 199982
rect -1526 202052 -1206 202640
rect -1526 201780 -1502 202052
rect -1230 201780 -1206 202052
rect -1526 199960 -1206 201780
rect -3018 199638 -2626 199662
rect -1528 199640 -1206 199960
rect -5546 199076 -5178 199100
rect -5546 198756 -5522 199076
rect -5202 198756 -5178 199076
rect -5546 198732 -5178 198756
rect -6318 197120 -5950 197144
rect -6318 196800 -6294 197120
rect -5974 196800 -5950 197120
rect -6318 196776 -5950 196800
rect -3786 197120 -3418 197144
rect -2946 197120 -2626 199638
rect -3786 196800 -3762 197120
rect -3442 196982 -2626 197120
rect -3442 196800 -2994 196982
rect -3786 196776 -3418 196800
rect -3018 196662 -2994 196800
rect -2674 196662 -2626 196982
rect -1526 199052 -1206 199640
rect -1526 198780 -1502 199052
rect -1230 198780 -1206 199052
rect -1526 196960 -1206 198780
rect -3018 196638 -2626 196662
rect -1528 196640 -1206 196960
rect -5546 196076 -5178 196100
rect -5546 195756 -5522 196076
rect -5202 195756 -5178 196076
rect -5546 195732 -5178 195756
rect -6318 194120 -5950 194144
rect -6318 193800 -6294 194120
rect -5974 193800 -5950 194120
rect -6318 193776 -5950 193800
rect -3786 194120 -3418 194144
rect -2946 194120 -2626 196638
rect -3786 193800 -3762 194120
rect -3442 193982 -2626 194120
rect -3442 193800 -2994 193982
rect -3786 193776 -3418 193800
rect -3018 193662 -2994 193800
rect -2674 193662 -2626 193982
rect -1526 196052 -1206 196640
rect -1526 195780 -1502 196052
rect -1230 195780 -1206 196052
rect -1526 193960 -1206 195780
rect -3018 193638 -2626 193662
rect -1528 193640 -1206 193960
rect -5546 193076 -5178 193100
rect -5546 192756 -5522 193076
rect -5202 192756 -5178 193076
rect -5546 192732 -5178 192756
rect -6318 191120 -5950 191144
rect -6318 190800 -6294 191120
rect -5974 190800 -5950 191120
rect -6318 190776 -5950 190800
rect -3786 191120 -3418 191144
rect -2946 191120 -2626 193638
rect -3786 190800 -3762 191120
rect -3442 190982 -2626 191120
rect -3442 190800 -2994 190982
rect -3786 190776 -3418 190800
rect -3018 190662 -2994 190800
rect -2674 190662 -2626 190982
rect -1526 193052 -1206 193640
rect -1526 192780 -1502 193052
rect -1230 192780 -1206 193052
rect -1526 190960 -1206 192780
rect -3018 190638 -2626 190662
rect -1528 190640 -1206 190960
rect -5546 190076 -5178 190100
rect -5546 189756 -5522 190076
rect -5202 189756 -5178 190076
rect -5546 189732 -5178 189756
rect -6318 188120 -5950 188144
rect -6318 187800 -6294 188120
rect -5974 187800 -5950 188120
rect -6318 187776 -5950 187800
rect -3786 188120 -3418 188144
rect -2946 188120 -2626 190638
rect -3786 187800 -3762 188120
rect -3442 187982 -2626 188120
rect -3442 187800 -2994 187982
rect -3786 187776 -3418 187800
rect -3018 187662 -2994 187800
rect -2674 187662 -2626 187982
rect -1526 190052 -1206 190640
rect -1526 189780 -1502 190052
rect -1230 189780 -1206 190052
rect -1526 187960 -1206 189780
rect -3018 187638 -2626 187662
rect -1528 187640 -1206 187960
rect -5546 187076 -5178 187100
rect -5546 186756 -5522 187076
rect -5202 186756 -5178 187076
rect -5546 186732 -5178 186756
rect -6318 185120 -5950 185144
rect -6318 184800 -6294 185120
rect -5974 184800 -5950 185120
rect -6318 184776 -5950 184800
rect -3786 185120 -3418 185144
rect -2946 185120 -2626 187638
rect -3786 184800 -3762 185120
rect -3442 184982 -2626 185120
rect -3442 184800 -2994 184982
rect -3786 184776 -3418 184800
rect -3018 184662 -2994 184800
rect -2674 184662 -2626 184982
rect -1526 187052 -1206 187640
rect -1526 186780 -1502 187052
rect -1230 186780 -1206 187052
rect -1526 184960 -1206 186780
rect -3018 184638 -2626 184662
rect -1528 184640 -1206 184960
rect -5546 184076 -5178 184100
rect -5546 183756 -5522 184076
rect -5202 183756 -5178 184076
rect -5546 183732 -5178 183756
rect -6318 182120 -5950 182144
rect -6318 181800 -6294 182120
rect -5974 181800 -5950 182120
rect -6318 181776 -5950 181800
rect -3786 182120 -3418 182144
rect -2946 182120 -2626 184638
rect -3786 181800 -3762 182120
rect -3442 181982 -2626 182120
rect -3442 181800 -2994 181982
rect -3786 181776 -3418 181800
rect -3018 181662 -2994 181800
rect -2674 181662 -2626 181982
rect -1526 184052 -1206 184640
rect -1526 183780 -1502 184052
rect -1230 183780 -1206 184052
rect -1526 181960 -1206 183780
rect -3018 181638 -2626 181662
rect -1528 181640 -1206 181960
rect -5546 181076 -5178 181100
rect -5546 180756 -5522 181076
rect -5202 180756 -5178 181076
rect -5546 180732 -5178 180756
rect -6318 179120 -5950 179144
rect -6318 178800 -6294 179120
rect -5974 178800 -5950 179120
rect -6318 178776 -5950 178800
rect -3786 179120 -3418 179144
rect -2946 179120 -2626 181638
rect -3786 178800 -3762 179120
rect -3442 178982 -2626 179120
rect -3442 178800 -2994 178982
rect -3786 178776 -3418 178800
rect -3018 178662 -2994 178800
rect -2674 178662 -2626 178982
rect -1526 181052 -1206 181640
rect -1526 180780 -1502 181052
rect -1230 180780 -1206 181052
rect -1526 178960 -1206 180780
rect -3018 178638 -2626 178662
rect -1528 178640 -1206 178960
rect -5546 178076 -5178 178100
rect -5546 177756 -5522 178076
rect -5202 177756 -5178 178076
rect -5546 177732 -5178 177756
rect -6318 176120 -5950 176144
rect -6318 175800 -6294 176120
rect -5974 175800 -5950 176120
rect -6318 175776 -5950 175800
rect -3786 176120 -3418 176144
rect -2946 176120 -2626 178638
rect -3786 175800 -3762 176120
rect -3442 175982 -2626 176120
rect -3442 175800 -2994 175982
rect -3786 175776 -3418 175800
rect -3018 175662 -2994 175800
rect -2674 175662 -2626 175982
rect -1526 178052 -1206 178640
rect -1526 177780 -1502 178052
rect -1230 177780 -1206 178052
rect -1526 175960 -1206 177780
rect -3018 175638 -2626 175662
rect -1528 175640 -1206 175960
rect -5546 175076 -5178 175100
rect -5546 174756 -5522 175076
rect -5202 174756 -5178 175076
rect -5546 174732 -5178 174756
rect -6318 173120 -5950 173144
rect -6318 172800 -6294 173120
rect -5974 172800 -5950 173120
rect -6318 172776 -5950 172800
rect -3786 173120 -3418 173144
rect -2946 173120 -2626 175638
rect -3786 172800 -3762 173120
rect -3442 172982 -2626 173120
rect -3442 172800 -2994 172982
rect -3786 172776 -3418 172800
rect -3018 172662 -2994 172800
rect -2674 172662 -2626 172982
rect -1526 175052 -1206 175640
rect -1526 174780 -1502 175052
rect -1230 174780 -1206 175052
rect -1526 172960 -1206 174780
rect -3018 172638 -2626 172662
rect -1528 172640 -1206 172960
rect -5546 172076 -5178 172100
rect -5546 171756 -5522 172076
rect -5202 171756 -5178 172076
rect -5546 171732 -5178 171756
rect -6318 170120 -5950 170144
rect -6318 169800 -6294 170120
rect -5974 169800 -5950 170120
rect -6318 169776 -5950 169800
rect -3786 170120 -3418 170144
rect -2946 170120 -2626 172638
rect -3786 169800 -3762 170120
rect -3442 169982 -2626 170120
rect -3442 169800 -2994 169982
rect -3786 169776 -3418 169800
rect -3018 169662 -2994 169800
rect -2674 169662 -2626 169982
rect -1526 172052 -1206 172640
rect -1526 171780 -1502 172052
rect -1230 171780 -1206 172052
rect -1526 169960 -1206 171780
rect -3018 169638 -2626 169662
rect -1528 169640 -1206 169960
rect -5546 169076 -5178 169100
rect -5546 168756 -5522 169076
rect -5202 168756 -5178 169076
rect -5546 168732 -5178 168756
rect -6318 167120 -5950 167144
rect -6318 166800 -6294 167120
rect -5974 166800 -5950 167120
rect -6318 166776 -5950 166800
rect -3786 167120 -3418 167144
rect -2946 167120 -2626 169638
rect -3786 166800 -3762 167120
rect -3442 166982 -2626 167120
rect -3442 166800 -2994 166982
rect -3786 166776 -3418 166800
rect -3018 166662 -2994 166800
rect -2674 166662 -2626 166982
rect -1526 169052 -1206 169640
rect -1526 168780 -1502 169052
rect -1230 168780 -1206 169052
rect -1526 166960 -1206 168780
rect -3018 166638 -2626 166662
rect -1528 166640 -1206 166960
rect -5546 166076 -5178 166100
rect -5546 165756 -5522 166076
rect -5202 165756 -5178 166076
rect -5546 165732 -5178 165756
rect -6318 164120 -5950 164144
rect -6318 163800 -6294 164120
rect -5974 163800 -5950 164120
rect -6318 163776 -5950 163800
rect -3786 164120 -3418 164144
rect -2946 164120 -2626 166638
rect -3786 163800 -3762 164120
rect -3442 163982 -2626 164120
rect -3442 163800 -2994 163982
rect -3786 163776 -3418 163800
rect -3018 163662 -2994 163800
rect -2674 163662 -2626 163982
rect -1526 166052 -1206 166640
rect -1526 165780 -1502 166052
rect -1230 165780 -1206 166052
rect -1526 163960 -1206 165780
rect -3018 163638 -2626 163662
rect -1528 163640 -1206 163960
rect -5546 163076 -5178 163100
rect -5546 162756 -5522 163076
rect -5202 162756 -5178 163076
rect -5546 162732 -5178 162756
rect -6318 161120 -5950 161144
rect -6318 160800 -6294 161120
rect -5974 160800 -5950 161120
rect -6318 160776 -5950 160800
rect -3786 161120 -3418 161144
rect -2946 161120 -2626 163638
rect -3786 160800 -3762 161120
rect -3442 160982 -2626 161120
rect -3442 160800 -2994 160982
rect -3786 160776 -3418 160800
rect -3018 160662 -2994 160800
rect -2674 160662 -2626 160982
rect -1526 163052 -1206 163640
rect -1526 162780 -1502 163052
rect -1230 162780 -1206 163052
rect -1526 160960 -1206 162780
rect -3018 160638 -2626 160662
rect -1528 160640 -1206 160960
rect -5546 160076 -5178 160100
rect -5546 159756 -5522 160076
rect -5202 159756 -5178 160076
rect -5546 159732 -5178 159756
rect -6318 158120 -5950 158144
rect -6318 157800 -6294 158120
rect -5974 157800 -5950 158120
rect -6318 157776 -5950 157800
rect -3786 158120 -3418 158144
rect -2946 158120 -2626 160638
rect -3786 157800 -3762 158120
rect -3442 157982 -2626 158120
rect -3442 157800 -2994 157982
rect -3786 157776 -3418 157800
rect -3018 157662 -2994 157800
rect -2674 157662 -2626 157982
rect -1526 160052 -1206 160640
rect -1526 159780 -1502 160052
rect -1230 159780 -1206 160052
rect -1526 157960 -1206 159780
rect -3018 157638 -2626 157662
rect -1528 157640 -1206 157960
rect -5546 157076 -5178 157100
rect -5546 156756 -5522 157076
rect -5202 156756 -5178 157076
rect -5546 156732 -5178 156756
rect -6318 155120 -5950 155144
rect -6318 154800 -6294 155120
rect -5974 154800 -5950 155120
rect -6318 154776 -5950 154800
rect -3786 155120 -3418 155144
rect -2946 155120 -2626 157638
rect -3786 154800 -3762 155120
rect -3442 154982 -2626 155120
rect -3442 154800 -2994 154982
rect -3786 154776 -3418 154800
rect -3018 154662 -2994 154800
rect -2674 154662 -2626 154982
rect -1526 157052 -1206 157640
rect -1526 156780 -1502 157052
rect -1230 156780 -1206 157052
rect -1526 154960 -1206 156780
rect -3018 154638 -2626 154662
rect -1528 154640 -1206 154960
rect -5546 154076 -5178 154100
rect -5546 153756 -5522 154076
rect -5202 153756 -5178 154076
rect -5546 153732 -5178 153756
rect -6318 152120 -5950 152144
rect -6318 151800 -6294 152120
rect -5974 151800 -5950 152120
rect -6318 151776 -5950 151800
rect -3786 152120 -3418 152144
rect -2946 152120 -2626 154638
rect -3786 151800 -3762 152120
rect -3442 151982 -2626 152120
rect -3442 151800 -2994 151982
rect -3786 151776 -3418 151800
rect -3018 151662 -2994 151800
rect -2674 151662 -2626 151982
rect -1526 154052 -1206 154640
rect -1526 153780 -1502 154052
rect -1230 153780 -1206 154052
rect -1526 151960 -1206 153780
rect -3018 151638 -2626 151662
rect -1528 151640 -1206 151960
rect -5546 151076 -5178 151100
rect -5546 150756 -5522 151076
rect -5202 150756 -5178 151076
rect -5546 150732 -5178 150756
rect -6318 149120 -5950 149144
rect -6318 148800 -6294 149120
rect -5974 148800 -5950 149120
rect -6318 148776 -5950 148800
rect -3786 149120 -3418 149144
rect -2946 149120 -2626 151638
rect -3786 148800 -3762 149120
rect -3442 148982 -2626 149120
rect -3442 148800 -2994 148982
rect -3786 148776 -3418 148800
rect -3018 148662 -2994 148800
rect -2674 148662 -2626 148982
rect -1526 151052 -1206 151640
rect -1526 150780 -1502 151052
rect -1230 150780 -1206 151052
rect -1526 148960 -1206 150780
rect -3018 148638 -2626 148662
rect -1528 148640 -1206 148960
rect -5546 148076 -5178 148100
rect -5546 147756 -5522 148076
rect -5202 147756 -5178 148076
rect -5546 147732 -5178 147756
rect -6318 146120 -5950 146144
rect -6318 145800 -6294 146120
rect -5974 145800 -5950 146120
rect -6318 145776 -5950 145800
rect -3786 146120 -3418 146144
rect -2946 146120 -2626 148638
rect -3786 145800 -3762 146120
rect -3442 145982 -2626 146120
rect -3442 145800 -2994 145982
rect -3786 145776 -3418 145800
rect -3018 145662 -2994 145800
rect -2674 145662 -2626 145982
rect -1526 148052 -1206 148640
rect -1526 147780 -1502 148052
rect -1230 147780 -1206 148052
rect -1526 145960 -1206 147780
rect -3018 145638 -2626 145662
rect -1528 145640 -1206 145960
rect -5546 145076 -5178 145100
rect -5546 144756 -5522 145076
rect -5202 144756 -5178 145076
rect -5546 144732 -5178 144756
rect -6318 143120 -5950 143144
rect -6318 142800 -6294 143120
rect -5974 142800 -5950 143120
rect -6318 142776 -5950 142800
rect -3786 143120 -3418 143144
rect -2946 143120 -2626 145638
rect -3786 142800 -3762 143120
rect -3442 142982 -2626 143120
rect -3442 142800 -2994 142982
rect -3786 142776 -3418 142800
rect -3018 142662 -2994 142800
rect -2674 142662 -2626 142982
rect -1526 145052 -1206 145640
rect -1526 144780 -1502 145052
rect -1230 144780 -1206 145052
rect -1526 142960 -1206 144780
rect -3018 142638 -2626 142662
rect -1528 142640 -1206 142960
rect -5546 142076 -5178 142100
rect -5546 141756 -5522 142076
rect -5202 141756 -5178 142076
rect -5546 141732 -5178 141756
rect -6318 140120 -5950 140144
rect -6318 139800 -6294 140120
rect -5974 139800 -5950 140120
rect -6318 139776 -5950 139800
rect -3786 140120 -3418 140144
rect -2946 140120 -2626 142638
rect -3786 139800 -3762 140120
rect -3442 139982 -2626 140120
rect -3442 139800 -2994 139982
rect -3786 139776 -3418 139800
rect -3018 139662 -2994 139800
rect -2674 139662 -2626 139982
rect -1526 142052 -1206 142640
rect -1526 141780 -1502 142052
rect -1230 141780 -1206 142052
rect -1526 139960 -1206 141780
rect -3018 139638 -2626 139662
rect -1528 139640 -1206 139960
rect -5546 139076 -5178 139100
rect -5546 138756 -5522 139076
rect -5202 138756 -5178 139076
rect -5546 138732 -5178 138756
rect -6318 137120 -5950 137144
rect -6318 136800 -6294 137120
rect -5974 136800 -5950 137120
rect -6318 136776 -5950 136800
rect -3786 137120 -3418 137144
rect -2946 137120 -2626 139638
rect -3786 136800 -3762 137120
rect -3442 136982 -2626 137120
rect -3442 136800 -2994 136982
rect -3786 136776 -3418 136800
rect -3018 136662 -2994 136800
rect -2674 136662 -2626 136982
rect -1526 139052 -1206 139640
rect -1526 138780 -1502 139052
rect -1230 138780 -1206 139052
rect -1526 136960 -1206 138780
rect -3018 136638 -2626 136662
rect -1528 136640 -1206 136960
rect -5546 136076 -5178 136100
rect -5546 135756 -5522 136076
rect -5202 135756 -5178 136076
rect -5546 135732 -5178 135756
rect -6318 134120 -5950 134144
rect -6318 133800 -6294 134120
rect -5974 133800 -5950 134120
rect -6318 133776 -5950 133800
rect -3786 134120 -3418 134144
rect -2946 134120 -2626 136638
rect -3786 133800 -3762 134120
rect -3442 133982 -2626 134120
rect -3442 133800 -2994 133982
rect -3786 133776 -3418 133800
rect -3018 133662 -2994 133800
rect -2674 133662 -2626 133982
rect -1526 136052 -1206 136640
rect -1526 135780 -1502 136052
rect -1230 135780 -1206 136052
rect -1526 133960 -1206 135780
rect -3018 133638 -2626 133662
rect -1528 133640 -1206 133960
rect -5546 133076 -5178 133100
rect -5546 132756 -5522 133076
rect -5202 132756 -5178 133076
rect -5546 132732 -5178 132756
rect -6318 131120 -5950 131144
rect -6318 130800 -6294 131120
rect -5974 130800 -5950 131120
rect -6318 130776 -5950 130800
rect -3786 131120 -3418 131144
rect -2946 131120 -2626 133638
rect -3786 130800 -3762 131120
rect -3442 130982 -2626 131120
rect -3442 130800 -2994 130982
rect -3786 130776 -3418 130800
rect -3018 130662 -2994 130800
rect -2674 130662 -2626 130982
rect -1526 133052 -1206 133640
rect -1526 132780 -1502 133052
rect -1230 132780 -1206 133052
rect -1526 130960 -1206 132780
rect -3018 130638 -2626 130662
rect -1528 130640 -1206 130960
rect -5546 130076 -5178 130100
rect -5546 129756 -5522 130076
rect -5202 129756 -5178 130076
rect -5546 129732 -5178 129756
rect -6318 128120 -5950 128144
rect -6318 127800 -6294 128120
rect -5974 127800 -5950 128120
rect -6318 127776 -5950 127800
rect -3786 128120 -3418 128144
rect -2946 128120 -2626 130638
rect -3786 127800 -3762 128120
rect -3442 127982 -2626 128120
rect -3442 127800 -2994 127982
rect -3786 127776 -3418 127800
rect -3018 127662 -2994 127800
rect -2674 127662 -2626 127982
rect -1526 130052 -1206 130640
rect -1526 129780 -1502 130052
rect -1230 129780 -1206 130052
rect -1526 127960 -1206 129780
rect -3018 127638 -2626 127662
rect -1528 127640 -1206 127960
rect -5546 127076 -5178 127100
rect -5546 126756 -5522 127076
rect -5202 126756 -5178 127076
rect -5546 126732 -5178 126756
rect -6318 125120 -5950 125144
rect -6318 124800 -6294 125120
rect -5974 124800 -5950 125120
rect -6318 124776 -5950 124800
rect -3786 125120 -3418 125144
rect -2946 125120 -2626 127638
rect -3786 124800 -3762 125120
rect -3442 124982 -2626 125120
rect -3442 124800 -2994 124982
rect -3786 124776 -3418 124800
rect -3018 124662 -2994 124800
rect -2674 124662 -2626 124982
rect -1526 127052 -1206 127640
rect -1526 126780 -1502 127052
rect -1230 126780 -1206 127052
rect -1526 124960 -1206 126780
rect -3018 124638 -2626 124662
rect -1528 124640 -1206 124960
rect -5546 124076 -5178 124100
rect -5546 123756 -5522 124076
rect -5202 123756 -5178 124076
rect -5546 123732 -5178 123756
rect -6318 122120 -5950 122144
rect -6318 121800 -6294 122120
rect -5974 121800 -5950 122120
rect -6318 121776 -5950 121800
rect -3786 122120 -3418 122144
rect -2946 122120 -2626 124638
rect -3786 121800 -3762 122120
rect -3442 121982 -2626 122120
rect -3442 121800 -2994 121982
rect -3786 121776 -3418 121800
rect -3018 121662 -2994 121800
rect -2674 121662 -2626 121982
rect -1526 124052 -1206 124640
rect -1526 123780 -1502 124052
rect -1230 123780 -1206 124052
rect -1526 121960 -1206 123780
rect -3018 121638 -2626 121662
rect -1528 121640 -1206 121960
rect -5546 121076 -5178 121100
rect -5546 120756 -5522 121076
rect -5202 120756 -5178 121076
rect -5546 120732 -5178 120756
rect -6318 119120 -5950 119144
rect -6318 118800 -6294 119120
rect -5974 118800 -5950 119120
rect -6318 118776 -5950 118800
rect -3786 119120 -3418 119144
rect -2946 119120 -2626 121638
rect -3786 118800 -3762 119120
rect -3442 118982 -2626 119120
rect -3442 118800 -2994 118982
rect -3786 118776 -3418 118800
rect -3018 118662 -2994 118800
rect -2674 118662 -2626 118982
rect -1526 121052 -1206 121640
rect -1526 120780 -1502 121052
rect -1230 120780 -1206 121052
rect -1526 118960 -1206 120780
rect -3018 118638 -2626 118662
rect -1528 118640 -1206 118960
rect -5546 118076 -5178 118100
rect -5546 117756 -5522 118076
rect -5202 117756 -5178 118076
rect -5546 117732 -5178 117756
rect -6318 116120 -5950 116144
rect -6318 115800 -6294 116120
rect -5974 115800 -5950 116120
rect -6318 115776 -5950 115800
rect -3786 116120 -3418 116144
rect -2946 116120 -2626 118638
rect -3786 115800 -3762 116120
rect -3442 115982 -2626 116120
rect -3442 115800 -2994 115982
rect -3786 115776 -3418 115800
rect -3018 115662 -2994 115800
rect -2674 115662 -2626 115982
rect -1526 118052 -1206 118640
rect -1526 117780 -1502 118052
rect -1230 117780 -1206 118052
rect -1526 115960 -1206 117780
rect -3018 115638 -2626 115662
rect -1528 115640 -1206 115960
rect -5546 115076 -5178 115100
rect -5546 114756 -5522 115076
rect -5202 114756 -5178 115076
rect -5546 114732 -5178 114756
rect -6318 113120 -5950 113144
rect -6318 112800 -6294 113120
rect -5974 112800 -5950 113120
rect -6318 112776 -5950 112800
rect -3786 113120 -3418 113144
rect -2946 113120 -2626 115638
rect -3786 112800 -3762 113120
rect -3442 112982 -2626 113120
rect -3442 112800 -2994 112982
rect -3786 112776 -3418 112800
rect -3018 112662 -2994 112800
rect -2674 112662 -2626 112982
rect -1526 115052 -1206 115640
rect -1526 114780 -1502 115052
rect -1230 114780 -1206 115052
rect -1526 112960 -1206 114780
rect -3018 112638 -2626 112662
rect -1528 112640 -1206 112960
rect -5546 112076 -5178 112100
rect -5546 111756 -5522 112076
rect -5202 111756 -5178 112076
rect -5546 111732 -5178 111756
rect -6318 110120 -5950 110144
rect -6318 109800 -6294 110120
rect -5974 109800 -5950 110120
rect -6318 109776 -5950 109800
rect -3786 110120 -3418 110144
rect -2946 110120 -2626 112638
rect -3786 109800 -3762 110120
rect -3442 109982 -2626 110120
rect -3442 109800 -2994 109982
rect -3786 109776 -3418 109800
rect -3018 109662 -2994 109800
rect -2674 109662 -2626 109982
rect -1526 112052 -1206 112640
rect -1526 111780 -1502 112052
rect -1230 111780 -1206 112052
rect -1526 109960 -1206 111780
rect -3018 109638 -2626 109662
rect -1528 109640 -1206 109960
rect -5546 109076 -5178 109100
rect -5546 108756 -5522 109076
rect -5202 108756 -5178 109076
rect -5546 108732 -5178 108756
rect -6318 107120 -5950 107144
rect -6318 106800 -6294 107120
rect -5974 106800 -5950 107120
rect -6318 106776 -5950 106800
rect -3786 107120 -3418 107144
rect -2946 107120 -2626 109638
rect -3786 106800 -3762 107120
rect -3442 106982 -2626 107120
rect -3442 106800 -2994 106982
rect -3786 106776 -3418 106800
rect -3018 106662 -2994 106800
rect -2674 106662 -2626 106982
rect -1526 109052 -1206 109640
rect -1526 108780 -1502 109052
rect -1230 108780 -1206 109052
rect -1526 106960 -1206 108780
rect -3018 106638 -2626 106662
rect -1528 106640 -1206 106960
rect -5546 106076 -5178 106100
rect -5546 105756 -5522 106076
rect -5202 105756 -5178 106076
rect -5546 105732 -5178 105756
rect -6318 104120 -5950 104144
rect -6318 103800 -6294 104120
rect -5974 103800 -5950 104120
rect -6318 103776 -5950 103800
rect -3786 104120 -3418 104144
rect -2946 104120 -2626 106638
rect -3786 103800 -3762 104120
rect -3442 103982 -2626 104120
rect -3442 103800 -2994 103982
rect -3786 103776 -3418 103800
rect -3018 103662 -2994 103800
rect -2674 103662 -2626 103982
rect -1526 106052 -1206 106640
rect -1526 105780 -1502 106052
rect -1230 105780 -1206 106052
rect -1526 103960 -1206 105780
rect -3018 103638 -2626 103662
rect -1528 103640 -1206 103960
rect -5546 103076 -5178 103100
rect -5546 102756 -5522 103076
rect -5202 102756 -5178 103076
rect -5546 102732 -5178 102756
rect -6318 101120 -5950 101144
rect -6318 100800 -6294 101120
rect -5974 100800 -5950 101120
rect -6318 100776 -5950 100800
rect -3786 101120 -3418 101144
rect -2946 101120 -2626 103638
rect -3786 100800 -3762 101120
rect -3442 100982 -2626 101120
rect -3442 100800 -2994 100982
rect -3786 100776 -3418 100800
rect -3018 100662 -2994 100800
rect -2674 100662 -2626 100982
rect -1526 103052 -1206 103640
rect -1526 102780 -1502 103052
rect -1230 102780 -1206 103052
rect -1526 100960 -1206 102780
rect -3018 100638 -2626 100662
rect -1528 100640 -1206 100960
rect -5546 100076 -5178 100100
rect -5546 99756 -5522 100076
rect -5202 99756 -5178 100076
rect -5546 99732 -5178 99756
rect -6318 98120 -5950 98144
rect -6318 97800 -6294 98120
rect -5974 97800 -5950 98120
rect -6318 97776 -5950 97800
rect -3786 98120 -3418 98144
rect -2946 98120 -2626 100638
rect -3786 97800 -3762 98120
rect -3442 97982 -2626 98120
rect -3442 97800 -2994 97982
rect -3786 97776 -3418 97800
rect -3018 97662 -2994 97800
rect -2674 97662 -2626 97982
rect -1526 100052 -1206 100640
rect -1526 99780 -1502 100052
rect -1230 99780 -1206 100052
rect -1526 97960 -1206 99780
rect -3018 97638 -2626 97662
rect -1528 97640 -1206 97960
rect -5546 97076 -5178 97100
rect -5546 96756 -5522 97076
rect -5202 96756 -5178 97076
rect -5546 96732 -5178 96756
rect -6318 95120 -5950 95144
rect -6318 94800 -6294 95120
rect -5974 94800 -5950 95120
rect -6318 94776 -5950 94800
rect -3786 95120 -3418 95144
rect -2946 95120 -2626 97638
rect -3786 94800 -3762 95120
rect -3442 94982 -2626 95120
rect -3442 94800 -2994 94982
rect -3786 94776 -3418 94800
rect -3018 94662 -2994 94800
rect -2674 94662 -2626 94982
rect -1526 97052 -1206 97640
rect -1526 96780 -1502 97052
rect -1230 96780 -1206 97052
rect -1526 94960 -1206 96780
rect -3018 94638 -2626 94662
rect -1528 94640 -1206 94960
rect -6318 92120 -5950 92144
rect -6318 91800 -6294 92120
rect -5974 91800 -5950 92120
rect -6318 91776 -5950 91800
rect -3786 92120 -3418 92144
rect -2946 92120 -2626 94638
rect -3786 91800 -3762 92120
rect -3442 91982 -2626 92120
rect -3442 91800 -2994 91982
rect -3786 91776 -3418 91800
rect -3018 91662 -2994 91800
rect -2674 91662 -2626 91982
rect -1526 91960 -1206 94640
rect -3018 91638 -2626 91662
rect -1528 91640 -1206 91960
rect -5546 91076 -5178 91100
rect -5546 90756 -5522 91076
rect -5202 90756 -5178 91076
rect -5546 90732 -5178 90756
rect -6318 89120 -5950 89144
rect -6318 88800 -6294 89120
rect -5974 88800 -5950 89120
rect -6318 88776 -5950 88800
rect -3786 89120 -3418 89144
rect -2946 89120 -2626 91638
rect -3786 88800 -3762 89120
rect -3442 88982 -2626 89120
rect -3442 88800 -2994 88982
rect -3786 88776 -3418 88800
rect -3018 88662 -2994 88800
rect -2674 88662 -2626 88982
rect -1526 91052 -1206 91640
rect -1526 90780 -1502 91052
rect -1230 90780 -1206 91052
rect -1526 88960 -1206 90780
rect -3018 88638 -2626 88662
rect -1528 88640 -1206 88960
rect -5546 88076 -5178 88100
rect -5546 87756 -5522 88076
rect -5202 87756 -5178 88076
rect -5546 87732 -5178 87756
rect -6318 86120 -5950 86144
rect -6318 85800 -6294 86120
rect -5974 85800 -5950 86120
rect -6318 85776 -5950 85800
rect -3786 86120 -3418 86144
rect -2946 86120 -2626 88638
rect -3786 85800 -3762 86120
rect -3442 85982 -2626 86120
rect -3442 85800 -2994 85982
rect -3786 85776 -3418 85800
rect -3018 85662 -2994 85800
rect -2674 85662 -2626 85982
rect -1526 88052 -1206 88640
rect -1526 87780 -1502 88052
rect -1230 87780 -1206 88052
rect -1526 85960 -1206 87780
rect -3018 85638 -2626 85662
rect -1528 85640 -1206 85960
rect -5546 85076 -5178 85100
rect -5546 84756 -5522 85076
rect -5202 84756 -5178 85076
rect -5546 84732 -5178 84756
rect -6318 83120 -5950 83144
rect -6318 82800 -6294 83120
rect -5974 82800 -5950 83120
rect -6318 82776 -5950 82800
rect -3786 83120 -3418 83144
rect -2946 83120 -2626 85638
rect -3786 82800 -3762 83120
rect -3442 82982 -2626 83120
rect -3442 82800 -2994 82982
rect -3786 82776 -3418 82800
rect -3018 82662 -2994 82800
rect -2674 82662 -2626 82982
rect -1526 85052 -1206 85640
rect -1526 84780 -1502 85052
rect -1230 84780 -1206 85052
rect -1526 82960 -1206 84780
rect -3018 82638 -2626 82662
rect -1528 82640 -1206 82960
rect -5546 82076 -5178 82100
rect -5546 81756 -5522 82076
rect -5202 81756 -5178 82076
rect -5546 81732 -5178 81756
rect -6318 80120 -5950 80144
rect -6318 79800 -6294 80120
rect -5974 79800 -5950 80120
rect -6318 79776 -5950 79800
rect -3786 80120 -3418 80144
rect -2946 80120 -2626 82638
rect -3786 79800 -3762 80120
rect -3442 79982 -2626 80120
rect -3442 79800 -2994 79982
rect -3786 79776 -3418 79800
rect -3018 79662 -2994 79800
rect -2674 79662 -2626 79982
rect -1526 82052 -1206 82640
rect -1526 81780 -1502 82052
rect -1230 81780 -1206 82052
rect -1526 79960 -1206 81780
rect -3018 79638 -2626 79662
rect -1528 79640 -1206 79960
rect -5546 79076 -5178 79100
rect -5546 78756 -5522 79076
rect -5202 78756 -5178 79076
rect -5546 78732 -5178 78756
rect -6318 77120 -5950 77144
rect -6318 76800 -6294 77120
rect -5974 76800 -5950 77120
rect -6318 76776 -5950 76800
rect -3786 77120 -3418 77144
rect -2946 77120 -2626 79638
rect -3786 76800 -3762 77120
rect -3442 76982 -2626 77120
rect -3442 76800 -2994 76982
rect -3786 76776 -3418 76800
rect -3018 76662 -2994 76800
rect -2674 76662 -2626 76982
rect -1526 79052 -1206 79640
rect -1526 78780 -1502 79052
rect -1230 78780 -1206 79052
rect -1526 76960 -1206 78780
rect -3018 76638 -2626 76662
rect -1528 76640 -1206 76960
rect -5546 76076 -5178 76100
rect -5546 75756 -5522 76076
rect -5202 75756 -5178 76076
rect -5546 75732 -5178 75756
rect -6318 74120 -5950 74144
rect -6318 73800 -6294 74120
rect -5974 73800 -5950 74120
rect -6318 73776 -5950 73800
rect -3786 74120 -3418 74144
rect -2946 74120 -2626 76638
rect -3786 73800 -3762 74120
rect -3442 73982 -2626 74120
rect -3442 73800 -2994 73982
rect -3786 73776 -3418 73800
rect -3018 73662 -2994 73800
rect -2674 73662 -2626 73982
rect -1526 76052 -1206 76640
rect -1526 75780 -1502 76052
rect -1230 75780 -1206 76052
rect -1526 73960 -1206 75780
rect -3018 73638 -2626 73662
rect -1528 73640 -1206 73960
rect -5546 73076 -5178 73100
rect -5546 72756 -5522 73076
rect -5202 72756 -5178 73076
rect -5546 72732 -5178 72756
rect -6318 71120 -5950 71144
rect -6318 70800 -6294 71120
rect -5974 70800 -5950 71120
rect -6318 70776 -5950 70800
rect -3786 71120 -3418 71144
rect -2946 71120 -2626 73638
rect -3786 70800 -3762 71120
rect -3442 70982 -2626 71120
rect -3442 70800 -2994 70982
rect -3786 70776 -3418 70800
rect -3018 70662 -2994 70800
rect -2674 70662 -2626 70982
rect -1526 73052 -1206 73640
rect -1526 72780 -1502 73052
rect -1230 72780 -1206 73052
rect -1526 70960 -1206 72780
rect -3018 70638 -2626 70662
rect -1528 70640 -1206 70960
rect -5546 70076 -5178 70100
rect -5546 69756 -5522 70076
rect -5202 69756 -5178 70076
rect -5546 69732 -5178 69756
rect -6318 68120 -5950 68144
rect -6318 67800 -6294 68120
rect -5974 67800 -5950 68120
rect -6318 67776 -5950 67800
rect -3786 68120 -3418 68144
rect -2946 68120 -2626 70638
rect -3786 67800 -3762 68120
rect -3442 67982 -2626 68120
rect -3442 67800 -2994 67982
rect -3786 67776 -3418 67800
rect -3018 67662 -2994 67800
rect -2674 67662 -2626 67982
rect -1526 70052 -1206 70640
rect -1526 69780 -1502 70052
rect -1230 69780 -1206 70052
rect -1526 67960 -1206 69780
rect -3018 67638 -2626 67662
rect -1528 67640 -1206 67960
rect -5546 67076 -5178 67100
rect -5546 66756 -5522 67076
rect -5202 66756 -5178 67076
rect -5546 66732 -5178 66756
rect -6318 65120 -5950 65144
rect -6318 64800 -6294 65120
rect -5974 64800 -5950 65120
rect -6318 64776 -5950 64800
rect -3786 65120 -3418 65144
rect -2946 65120 -2626 67638
rect -3786 64800 -3762 65120
rect -3442 64982 -2626 65120
rect -3442 64800 -2994 64982
rect -3786 64776 -3418 64800
rect -3018 64662 -2994 64800
rect -2674 64662 -2626 64982
rect -1526 67052 -1206 67640
rect -1526 66780 -1502 67052
rect -1230 66780 -1206 67052
rect -1526 64960 -1206 66780
rect -3018 64638 -2626 64662
rect -1528 64640 -1206 64960
rect -5546 64076 -5178 64100
rect -5546 63756 -5522 64076
rect -5202 63756 -5178 64076
rect -5546 63732 -5178 63756
rect -6318 62120 -5950 62144
rect -6318 61800 -6294 62120
rect -5974 61800 -5950 62120
rect -6318 61776 -5950 61800
rect -3786 62120 -3418 62144
rect -2946 62120 -2626 64638
rect -3786 61800 -3762 62120
rect -3442 61982 -2626 62120
rect -3442 61800 -2994 61982
rect -3786 61776 -3418 61800
rect -3018 61662 -2994 61800
rect -2674 61662 -2626 61982
rect -1526 64052 -1206 64640
rect -1526 63780 -1502 64052
rect -1230 63780 -1206 64052
rect -1526 61960 -1206 63780
rect -3018 61638 -2626 61662
rect -1528 61640 -1206 61960
rect -5546 61076 -5178 61100
rect -5546 60756 -5522 61076
rect -5202 60756 -5178 61076
rect -5546 60732 -5178 60756
rect -6318 59120 -5950 59144
rect -6318 58800 -6294 59120
rect -5974 58800 -5950 59120
rect -6318 58776 -5950 58800
rect -3786 59120 -3418 59144
rect -2946 59120 -2626 61638
rect -3786 58800 -3762 59120
rect -3442 58982 -2626 59120
rect -3442 58800 -2994 58982
rect -3786 58776 -3418 58800
rect -3018 58662 -2994 58800
rect -2674 58662 -2626 58982
rect -1526 61052 -1206 61640
rect -1526 60780 -1502 61052
rect -1230 60780 -1206 61052
rect -1526 58960 -1206 60780
rect -3018 58638 -2626 58662
rect -1528 58640 -1206 58960
rect -5546 58076 -5178 58100
rect -5546 57756 -5522 58076
rect -5202 57756 -5178 58076
rect -5546 57732 -5178 57756
rect -2946 56120 -2626 58638
rect -3120 55982 -2626 56120
rect -3120 55800 -2994 55982
rect -3018 55662 -2994 55800
rect -2674 55662 -2626 55982
rect -1526 58052 -1206 58640
rect -1526 57780 -1502 58052
rect -1230 57780 -1206 58052
rect -1526 55960 -1206 57780
rect -3018 55638 -2626 55662
rect -1528 55640 -1206 55960
rect -5546 55076 -5178 55100
rect -5546 54756 -5522 55076
rect -5202 54756 -5178 55076
rect -5546 54732 -5178 54756
rect -6318 53120 -5950 53144
rect -6318 52800 -6294 53120
rect -5974 52800 -5950 53120
rect -6318 52776 -5950 52800
rect -3786 53120 -3418 53144
rect -2946 53120 -2626 55638
rect -3786 52800 -3762 53120
rect -3442 52982 -2626 53120
rect -3442 52800 -2994 52982
rect -3786 52776 -3418 52800
rect -3018 52662 -2994 52800
rect -2674 52662 -2626 52982
rect -1526 55052 -1206 55640
rect -1526 54780 -1502 55052
rect -1230 54780 -1206 55052
rect -1526 52960 -1206 54780
rect -3018 52638 -2626 52662
rect -1528 52640 -1206 52960
rect -5546 52076 -5178 52100
rect -5546 51756 -5522 52076
rect -5202 51756 -5178 52076
rect -5546 51732 -5178 51756
rect -6318 50120 -5950 50144
rect -6318 49800 -6294 50120
rect -5974 49800 -5950 50120
rect -6318 49776 -5950 49800
rect -3786 50120 -3418 50144
rect -2946 50120 -2626 52638
rect -3786 49800 -3762 50120
rect -3442 49982 -2626 50120
rect -3442 49800 -2994 49982
rect -3786 49776 -3418 49800
rect -3018 49662 -2994 49800
rect -2674 49662 -2626 49982
rect -1526 52052 -1206 52640
rect -1526 51780 -1502 52052
rect -1230 51780 -1206 52052
rect -1526 49960 -1206 51780
rect -3018 49638 -2626 49662
rect -1528 49640 -1206 49960
rect -5546 49076 -5178 49100
rect -5546 48756 -5522 49076
rect -5202 48756 -5178 49076
rect -5546 48732 -5178 48756
rect -6318 47120 -5950 47144
rect -6318 46800 -6294 47120
rect -5974 46800 -5950 47120
rect -6318 46776 -5950 46800
rect -3786 47120 -3418 47144
rect -2946 47120 -2626 49638
rect -3786 46800 -3762 47120
rect -3442 46982 -2626 47120
rect -3442 46800 -2994 46982
rect -3786 46776 -3418 46800
rect -3018 46662 -2994 46800
rect -2674 46662 -2626 46982
rect -1526 49052 -1206 49640
rect -1526 48780 -1502 49052
rect -1230 48780 -1206 49052
rect -1526 46960 -1206 48780
rect -3018 46638 -2626 46662
rect -1528 46640 -1206 46960
rect -5546 46076 -5178 46100
rect -5546 45756 -5522 46076
rect -5202 45756 -5178 46076
rect -5546 45732 -5178 45756
rect -6318 44120 -5950 44144
rect -6318 43800 -6294 44120
rect -5974 43800 -5950 44120
rect -6318 43776 -5950 43800
rect -3786 44120 -3418 44144
rect -2946 44120 -2626 46638
rect -3786 43800 -3762 44120
rect -3442 43982 -2626 44120
rect -3442 43800 -2994 43982
rect -3786 43776 -3418 43800
rect -3018 43662 -2994 43800
rect -2674 43662 -2626 43982
rect -1526 46052 -1206 46640
rect -1526 45780 -1502 46052
rect -1230 45780 -1206 46052
rect -1526 43960 -1206 45780
rect -3018 43638 -2626 43662
rect -1528 43640 -1206 43960
rect -5546 43076 -5178 43100
rect -5546 42756 -5522 43076
rect -5202 42756 -5178 43076
rect -5546 42732 -5178 42756
rect -6318 41120 -5950 41144
rect -6318 40800 -6294 41120
rect -5974 40800 -5950 41120
rect -6318 40776 -5950 40800
rect -3786 41120 -3418 41144
rect -2946 41120 -2626 43638
rect -3786 40800 -3762 41120
rect -3442 40982 -2626 41120
rect -3442 40800 -2994 40982
rect -3786 40776 -3418 40800
rect -3018 40662 -2994 40800
rect -2674 40662 -2626 40982
rect -1526 43052 -1206 43640
rect -1526 42780 -1502 43052
rect -1230 42780 -1206 43052
rect -1526 40960 -1206 42780
rect -3018 40638 -2626 40662
rect -1528 40640 -1206 40960
rect -5546 40076 -5178 40100
rect -5546 39756 -5522 40076
rect -5202 39756 -5178 40076
rect -5546 39732 -5178 39756
rect -6318 38120 -5950 38144
rect -6318 37800 -6294 38120
rect -5974 37800 -5950 38120
rect -6318 37776 -5950 37800
rect -3786 38120 -3418 38144
rect -2946 38120 -2626 40638
rect -3786 37800 -3762 38120
rect -3442 37982 -2626 38120
rect -3442 37800 -2994 37982
rect -3786 37776 -3418 37800
rect -3018 37662 -2994 37800
rect -2674 37662 -2626 37982
rect -1526 40052 -1206 40640
rect -1526 39780 -1502 40052
rect -1230 39780 -1206 40052
rect -1526 37960 -1206 39780
rect -3018 37638 -2626 37662
rect -1528 37640 -1206 37960
rect -5546 37076 -5178 37100
rect -5546 36756 -5522 37076
rect -5202 36756 -5178 37076
rect -5546 36732 -5178 36756
rect -6318 35120 -5950 35144
rect -6318 34800 -6294 35120
rect -5974 34800 -5950 35120
rect -6318 34776 -5950 34800
rect -3786 35120 -3418 35144
rect -2946 35120 -2626 37638
rect -3786 34800 -3762 35120
rect -3442 34982 -2626 35120
rect -3442 34800 -2994 34982
rect -3786 34776 -3418 34800
rect -3018 34662 -2994 34800
rect -2674 34662 -2626 34982
rect -1526 37052 -1206 37640
rect -1526 36780 -1502 37052
rect -1230 36780 -1206 37052
rect -1526 34960 -1206 36780
rect -3018 34638 -2626 34662
rect -1528 34640 -1206 34960
rect -5546 34076 -5178 34100
rect -5546 33756 -5522 34076
rect -5202 33756 -5178 34076
rect -5546 33732 -5178 33756
rect -6318 32120 -5950 32144
rect -6318 31800 -6294 32120
rect -5974 31800 -5950 32120
rect -6318 31776 -5950 31800
rect -3786 32120 -3418 32144
rect -2946 32120 -2626 34638
rect -3786 31800 -3762 32120
rect -3442 31982 -2626 32120
rect -3442 31800 -2994 31982
rect -3786 31776 -3418 31800
rect -3018 31662 -2994 31800
rect -2674 31662 -2626 31982
rect -1526 34052 -1206 34640
rect -1526 33780 -1502 34052
rect -1230 33780 -1206 34052
rect -1526 31960 -1206 33780
rect -3018 31638 -2626 31662
rect -1528 31640 -1206 31960
rect -5546 31076 -5178 31100
rect -5546 30756 -5522 31076
rect -5202 30756 -5178 31076
rect -5546 30732 -5178 30756
rect -6318 29120 -5950 29144
rect -6318 28800 -6294 29120
rect -5974 28800 -5950 29120
rect -6318 28776 -5950 28800
rect -3786 29120 -3418 29144
rect -2946 29120 -2626 31638
rect -3786 28800 -3762 29120
rect -3442 28982 -2626 29120
rect -3442 28800 -2994 28982
rect -3786 28776 -3418 28800
rect -3018 28662 -2994 28800
rect -2674 28662 -2626 28982
rect -1526 31052 -1206 31640
rect -1526 30780 -1502 31052
rect -1230 30780 -1206 31052
rect -1526 28960 -1206 30780
rect -3018 28638 -2626 28662
rect -1528 28640 -1206 28960
rect -5546 28076 -5178 28100
rect -5546 27756 -5522 28076
rect -5202 27756 -5178 28076
rect -5546 27732 -5178 27756
rect -6318 26120 -5950 26144
rect -6318 25800 -6294 26120
rect -5974 25800 -5950 26120
rect -6318 25776 -5950 25800
rect -3786 26120 -3418 26144
rect -2946 26120 -2626 28638
rect -3786 25800 -3762 26120
rect -3442 25982 -2626 26120
rect -3442 25800 -2994 25982
rect -3786 25776 -3418 25800
rect -3018 25662 -2994 25800
rect -2674 25662 -2626 25982
rect -1526 28052 -1206 28640
rect -1526 27780 -1502 28052
rect -1230 27780 -1206 28052
rect -1526 25960 -1206 27780
rect -3018 25638 -2626 25662
rect -1528 25640 -1206 25960
rect -5546 25076 -5178 25100
rect -5546 24756 -5522 25076
rect -5202 24756 -5178 25076
rect -5546 24732 -5178 24756
rect -6318 23120 -5950 23144
rect -6318 22800 -6294 23120
rect -5974 22800 -5950 23120
rect -6318 22776 -5950 22800
rect -3786 23120 -3418 23144
rect -2946 23120 -2626 25638
rect -3786 22800 -3762 23120
rect -3442 22982 -2626 23120
rect -3442 22800 -2994 22982
rect -3786 22776 -3418 22800
rect -3018 22662 -2994 22800
rect -2674 22662 -2626 22982
rect -1526 25052 -1206 25640
rect -1526 24780 -1502 25052
rect -1230 24780 -1206 25052
rect -1526 22960 -1206 24780
rect -3018 22638 -2626 22662
rect -1528 22640 -1206 22960
rect -5546 22076 -5178 22100
rect -5546 21756 -5522 22076
rect -5202 21756 -5178 22076
rect -5546 21732 -5178 21756
rect -6318 20120 -5950 20144
rect -6318 19800 -6294 20120
rect -5974 19800 -5950 20120
rect -6318 19776 -5950 19800
rect -3786 20120 -3418 20144
rect -2946 20120 -2626 22638
rect -3786 19800 -3762 20120
rect -3442 19800 -2626 20120
rect -1526 22052 -1206 22640
rect -1526 21780 -1502 22052
rect -1230 21780 -1206 22052
rect -1526 19960 -1206 21780
rect -3786 19776 -3418 19800
rect -5546 19076 -5178 19100
rect -5546 18756 -5522 19076
rect -5202 18756 -5178 19076
rect -5546 18732 -5178 18756
rect -6414 18026 -6094 18186
rect -6438 18002 -6070 18026
rect -6438 17682 -6414 18002
rect -6094 17682 -6070 18002
rect -6438 17658 -6070 17682
rect -6414 17374 -6094 17658
rect -2946 17288 -2626 19800
rect -1528 19640 -1206 19960
rect -1526 19052 -1206 19640
rect -1526 18780 -1502 19052
rect -1230 18780 -1206 19052
rect 303926 318334 304246 321062
rect 303926 318062 303950 318334
rect 304222 318062 304246 318334
rect 303926 315334 304246 318062
rect 303926 315062 303950 315334
rect 304222 315062 304246 315334
rect 303926 312334 304246 315062
rect 303926 312062 303950 312334
rect 304222 312062 304246 312334
rect 303926 309334 304246 312062
rect 303926 309062 303950 309334
rect 304222 309062 304246 309334
rect 303926 306334 304246 309062
rect 303926 306062 303950 306334
rect 304222 306062 304246 306334
rect 303926 303334 304246 306062
rect 303926 303062 303950 303334
rect 304222 303062 304246 303334
rect 303926 300334 304246 303062
rect 303926 300062 303950 300334
rect 304222 300062 304246 300334
rect 303926 297334 304246 300062
rect 303926 297062 303950 297334
rect 304222 297062 304246 297334
rect 303926 294334 304246 297062
rect 303926 294062 303950 294334
rect 304222 294062 304246 294334
rect 303926 291334 304246 294062
rect 303926 291062 303950 291334
rect 304222 291062 304246 291334
rect 303926 288334 304246 291062
rect 303926 288062 303950 288334
rect 304222 288062 304246 288334
rect 303926 285334 304246 288062
rect 303926 285062 303950 285334
rect 304222 285062 304246 285334
rect 303926 282334 304246 285062
rect 303926 282062 303950 282334
rect 304222 282062 304246 282334
rect 303926 279334 304246 282062
rect 303926 279062 303950 279334
rect 304222 279062 304246 279334
rect 303926 276334 304246 279062
rect 303926 276062 303950 276334
rect 304222 276062 304246 276334
rect 303926 273334 304246 276062
rect 303926 273062 303950 273334
rect 304222 273062 304246 273334
rect 303926 270334 304246 273062
rect 303926 270062 303950 270334
rect 304222 270062 304246 270334
rect 303926 267334 304246 270062
rect 303926 267062 303950 267334
rect 304222 267062 304246 267334
rect 303926 264334 304246 267062
rect 303926 264062 303950 264334
rect 304222 264062 304246 264334
rect 303926 261334 304246 264062
rect 303926 261062 303950 261334
rect 304222 261062 304246 261334
rect 303926 258334 304246 261062
rect 303926 258062 303950 258334
rect 304222 258062 304246 258334
rect 303926 255334 304246 258062
rect 303926 255062 303950 255334
rect 304222 255062 304246 255334
rect 303926 252334 304246 255062
rect 303926 252062 303950 252334
rect 304222 252062 304246 252334
rect 303926 249334 304246 252062
rect 303926 249062 303950 249334
rect 304222 249062 304246 249334
rect 303926 246334 304246 249062
rect 303926 246062 303950 246334
rect 304222 246062 304246 246334
rect 303926 243334 304246 246062
rect 303926 243062 303950 243334
rect 304222 243062 304246 243334
rect 303926 240334 304246 243062
rect 303926 240062 303950 240334
rect 304222 240062 304246 240334
rect 303926 237334 304246 240062
rect 303926 237062 303950 237334
rect 304222 237062 304246 237334
rect 303926 234334 304246 237062
rect 303926 234062 303950 234334
rect 304222 234062 304246 234334
rect 303926 231334 304246 234062
rect 303926 231062 303950 231334
rect 304222 231062 304246 231334
rect 303926 228334 304246 231062
rect 303926 228062 303950 228334
rect 304222 228062 304246 228334
rect 303926 225334 304246 228062
rect 303926 225062 303950 225334
rect 304222 225062 304246 225334
rect 303926 222334 304246 225062
rect 303926 222062 303950 222334
rect 304222 222062 304246 222334
rect 303926 219334 304246 222062
rect 303926 219062 303950 219334
rect 304222 219062 304246 219334
rect 303926 216334 304246 219062
rect 303926 216062 303950 216334
rect 304222 216062 304246 216334
rect 303926 213334 304246 216062
rect 303926 213062 303950 213334
rect 304222 213062 304246 213334
rect 303926 210334 304246 213062
rect 303926 210062 303950 210334
rect 304222 210062 304246 210334
rect 303926 207334 304246 210062
rect 303926 207062 303950 207334
rect 304222 207062 304246 207334
rect 303926 204334 304246 207062
rect 303926 204062 303950 204334
rect 304222 204062 304246 204334
rect 303926 201334 304246 204062
rect 303926 201062 303950 201334
rect 304222 201062 304246 201334
rect 303926 198334 304246 201062
rect 303926 198062 303950 198334
rect 304222 198062 304246 198334
rect 303926 195334 304246 198062
rect 303926 195062 303950 195334
rect 304222 195062 304246 195334
rect 303926 192334 304246 195062
rect 303926 192062 303950 192334
rect 304222 192062 304246 192334
rect 303926 189334 304246 192062
rect 303926 189062 303950 189334
rect 304222 189062 304246 189334
rect 303926 186334 304246 189062
rect 303926 186062 303950 186334
rect 304222 186062 304246 186334
rect 303926 183334 304246 186062
rect 303926 183062 303950 183334
rect 304222 183062 304246 183334
rect 303926 180334 304246 183062
rect 303926 180062 303950 180334
rect 304222 180062 304246 180334
rect 303926 177334 304246 180062
rect 303926 177062 303950 177334
rect 304222 177062 304246 177334
rect 303926 174334 304246 177062
rect 303926 174062 303950 174334
rect 304222 174062 304246 174334
rect 303926 171334 304246 174062
rect 303926 171062 303950 171334
rect 304222 171062 304246 171334
rect 303926 168334 304246 171062
rect 303926 168062 303950 168334
rect 304222 168062 304246 168334
rect 303926 165334 304246 168062
rect 303926 165062 303950 165334
rect 304222 165062 304246 165334
rect 303926 162334 304246 165062
rect 303926 162062 303950 162334
rect 304222 162062 304246 162334
rect 303926 159334 304246 162062
rect 303926 159062 303950 159334
rect 304222 159062 304246 159334
rect 303926 156334 304246 159062
rect 303926 156062 303950 156334
rect 304222 156062 304246 156334
rect 303926 153334 304246 156062
rect 303926 153062 303950 153334
rect 304222 153062 304246 153334
rect 303926 150334 304246 153062
rect 303926 150062 303950 150334
rect 304222 150062 304246 150334
rect 303926 147334 304246 150062
rect 303926 147062 303950 147334
rect 304222 147062 304246 147334
rect 303926 144334 304246 147062
rect 303926 144062 303950 144334
rect 304222 144062 304246 144334
rect 303926 141334 304246 144062
rect 303926 141062 303950 141334
rect 304222 141062 304246 141334
rect 303926 138334 304246 141062
rect 303926 138062 303950 138334
rect 304222 138062 304246 138334
rect 303926 135334 304246 138062
rect 303926 135062 303950 135334
rect 304222 135062 304246 135334
rect 303926 132334 304246 135062
rect 303926 132062 303950 132334
rect 304222 132062 304246 132334
rect 303926 129334 304246 132062
rect 303926 129062 303950 129334
rect 304222 129062 304246 129334
rect 303926 126334 304246 129062
rect 303926 126062 303950 126334
rect 304222 126062 304246 126334
rect 303926 123334 304246 126062
rect 303926 123062 303950 123334
rect 304222 123062 304246 123334
rect 303926 120334 304246 123062
rect 303926 120062 303950 120334
rect 304222 120062 304246 120334
rect 303926 117334 304246 120062
rect 303926 117062 303950 117334
rect 304222 117062 304246 117334
rect 303926 114334 304246 117062
rect 303926 114062 303950 114334
rect 304222 114062 304246 114334
rect 303926 111334 304246 114062
rect 303926 111062 303950 111334
rect 304222 111062 304246 111334
rect 303926 108334 304246 111062
rect 303926 108062 303950 108334
rect 304222 108062 304246 108334
rect 303926 105334 304246 108062
rect 303926 105062 303950 105334
rect 304222 105062 304246 105334
rect 303926 102334 304246 105062
rect 303926 102062 303950 102334
rect 304222 102062 304246 102334
rect 303926 99334 304246 102062
rect 303926 99062 303950 99334
rect 304222 99062 304246 99334
rect 303926 96334 304246 99062
rect 303926 96062 303950 96334
rect 304222 96062 304246 96334
rect 303926 93334 304246 96062
rect 303926 93062 303950 93334
rect 304222 93062 304246 93334
rect 303926 90334 304246 93062
rect 303926 90062 303950 90334
rect 304222 90062 304246 90334
rect 303926 87334 304246 90062
rect 303926 87062 303950 87334
rect 304222 87062 304246 87334
rect 303926 84334 304246 87062
rect 303926 84062 303950 84334
rect 304222 84062 304246 84334
rect 303926 81334 304246 84062
rect 303926 81062 303950 81334
rect 304222 81062 304246 81334
rect 303926 78334 304246 81062
rect 303926 78062 303950 78334
rect 304222 78062 304246 78334
rect 303926 75334 304246 78062
rect 303926 75062 303950 75334
rect 304222 75062 304246 75334
rect 303926 72334 304246 75062
rect 303926 72062 303950 72334
rect 304222 72062 304246 72334
rect 303926 69334 304246 72062
rect 303926 69062 303950 69334
rect 304222 69062 304246 69334
rect 303926 66334 304246 69062
rect 303926 66062 303950 66334
rect 304222 66062 304246 66334
rect 303926 63334 304246 66062
rect 303926 63062 303950 63334
rect 304222 63062 304246 63334
rect 303926 60334 304246 63062
rect 303926 60062 303950 60334
rect 304222 60062 304246 60334
rect 303926 57334 304246 60062
rect 303926 57062 303950 57334
rect 304222 57062 304246 57334
rect 303926 54334 304246 57062
rect 303926 54062 303950 54334
rect 304222 54062 304246 54334
rect 303926 51334 304246 54062
rect 303926 51062 303950 51334
rect 304222 51062 304246 51334
rect 303926 48334 304246 51062
rect 303926 48062 303950 48334
rect 304222 48062 304246 48334
rect 303926 45334 304246 48062
rect 303926 45062 303950 45334
rect 304222 45062 304246 45334
rect 303926 42334 304246 45062
rect 303926 42062 303950 42334
rect 304222 42062 304246 42334
rect 303926 39334 304246 42062
rect 303926 39062 303950 39334
rect 304222 39062 304246 39334
rect 303926 36334 304246 39062
rect 303926 36062 303950 36334
rect 304222 36062 304246 36334
rect 303926 33334 304246 36062
rect 303926 33062 303950 33334
rect 304222 33062 304246 33334
rect 303926 30334 304246 33062
rect 303926 30062 303950 30334
rect 304222 30062 304246 30334
rect 303926 27334 304246 30062
rect 303926 27062 303950 27334
rect 304222 27062 304246 27334
rect 303926 24334 304246 27062
rect 303926 24062 303950 24334
rect 304222 24062 304246 24334
rect 303926 21334 304246 24062
rect 303926 21062 303950 21334
rect 304222 21062 304246 21334
rect -1526 18760 -1206 18780
rect 289572 18760 289952 18790
rect 303926 18760 304246 21062
rect -1578 18736 304262 18760
rect -1578 18464 3688 18736
rect 3960 18464 18112 18736
rect 18384 18464 32938 18736
rect 33210 18464 64280 18736
rect 64552 18464 121702 18736
rect 121974 18464 167572 18736
rect 167844 18464 180572 18736
rect 180844 18464 189572 18736
rect 189844 18464 198572 18736
rect 198844 18464 204572 18736
rect 204844 18464 211572 18736
rect 211844 18464 223572 18736
rect 223844 18464 232572 18736
rect 232844 18464 238572 18736
rect 238844 18464 250572 18736
rect 250844 18464 263972 18736
rect 264244 18464 269972 18736
rect 270244 18464 272972 18736
rect 273244 18464 275972 18736
rect 276244 18464 281972 18736
rect 282244 18464 285972 18736
rect 286244 18464 293972 18736
rect 294244 18464 296972 18736
rect 297244 18464 299972 18736
rect 300244 18464 302972 18736
rect 303244 18464 304262 18736
rect -1578 18440 304262 18464
rect 289572 18422 289952 18440
rect 303926 18104 304246 18440
rect 305436 17288 305756 326222
rect -2982 17264 305756 17288
rect -2982 16992 303890 17264
rect 304162 16992 305756 17264
rect -2982 16968 305756 16992
rect -2946 16904 -2626 16968
rect 644 16874 964 16968
rect 3644 16874 3964 16968
rect 6644 16874 6964 16968
rect 9644 16874 9964 16968
rect 12644 16874 12964 16968
rect 15644 16874 15964 16968
rect 18644 16874 18964 16968
rect 21644 16874 21964 16968
rect 24644 16874 24964 16968
rect 27644 16874 27964 16968
rect 30644 16874 30964 16968
rect 33644 16874 33964 16968
rect 36644 16874 36964 16968
rect 39644 16874 39964 16968
rect 42644 16874 42964 16968
rect 45644 16874 45964 16968
rect 48644 16874 48964 16968
rect 51644 16874 51964 16968
rect 54644 16874 54964 16968
rect 57644 16874 57964 16968
rect 60644 16874 60964 16968
rect 63644 16874 63964 16968
rect 66644 16874 66964 16968
rect 69644 16874 69964 16968
rect 72644 16874 72964 16968
rect 75644 16874 75964 16968
rect 78644 16874 78964 16968
rect 81644 16874 81964 16968
rect 84644 16874 84964 16968
rect 87644 16874 87964 16968
rect 90644 16874 90964 16968
rect 93644 16874 93964 16968
rect 96644 16874 96964 16968
rect 99644 16874 99964 16968
rect 102644 16874 102964 16968
rect 105644 16874 105964 16968
rect 108644 16874 108964 16968
rect 111644 16874 111964 16968
rect 114644 16874 114964 16968
rect 117644 16874 117964 16968
rect 120644 16874 120964 16968
rect 123644 16874 123964 16968
rect 126644 16874 126964 16968
rect 129644 16874 129964 16968
rect 132644 16874 132964 16968
rect 135644 16874 135964 16968
rect 138644 16874 138964 16968
rect 141644 16874 141964 16968
rect 144644 16874 144964 16968
rect 147644 16874 147964 16968
rect 150644 16874 150964 16968
rect 153644 16874 153964 16968
rect 156644 16874 156964 16968
rect 159644 16874 159964 16968
rect 162644 16874 162964 16968
rect 165644 16874 165964 16968
rect 168644 16874 168964 16968
rect 171644 16874 171964 16968
rect 174644 16874 174964 16968
rect 177644 16874 177964 16968
rect 180644 16874 180964 16968
rect 183644 16874 183964 16968
rect 186644 16874 186964 16968
rect 189644 16874 189964 16968
rect 192644 16874 192964 16968
rect 195644 16874 195964 16968
rect 198644 16874 198964 16968
rect 201644 16874 201964 16968
rect 204644 16874 204964 16968
rect 207644 16874 207964 16968
rect 210644 16874 210964 16968
rect 213644 16874 213964 16968
rect 216644 16874 216964 16968
rect 219644 16874 219964 16968
rect 222644 16874 222964 16968
rect 225644 16874 225964 16968
rect 228644 16874 228964 16968
rect 231644 16874 231964 16968
rect 234644 16874 234964 16968
rect 237644 16874 237964 16968
rect 240644 16874 240964 16968
rect 243644 16874 243964 16968
rect 246644 16874 246964 16968
rect 249644 16874 249964 16968
rect 252644 16874 252964 16968
rect 255644 16874 255964 16968
rect 258644 16874 258964 16968
rect 261644 16874 261964 16968
rect 264644 16874 264964 16968
rect 270644 16874 270964 16968
rect 273644 16874 273964 16968
rect 276644 16874 276964 16968
rect 279644 16874 279964 16968
rect 282644 16874 282964 16968
rect 285644 16874 285964 16968
rect 288644 16874 288964 16968
rect 291644 16874 291964 16968
rect 294644 16874 294964 16968
rect 297644 16874 297964 16968
rect 300644 16874 300964 16968
rect 302916 16410 303298 16434
rect 302916 16088 302940 16410
rect 303274 16088 303298 16410
rect 302916 16064 303298 16088
rect 306874 16048 307194 16842
rect 3634 15688 4014 15712
rect 24 15642 392 15666
rect 24 15322 48 15642
rect 368 15322 836 15642
rect 3634 15368 3658 15688
rect 3990 15368 4014 15688
rect 3634 15344 4014 15368
rect 18058 15706 18438 15730
rect 18058 15386 18082 15706
rect 18414 15386 18438 15706
rect 18058 15362 18438 15386
rect 32884 15682 33264 15706
rect 32884 15362 32908 15682
rect 33240 15362 33264 15682
rect 32884 15338 33264 15362
rect 64226 15690 64606 15714
rect 64226 15370 64250 15690
rect 64582 15370 64606 15690
rect 64226 15346 64606 15370
rect 121648 15704 122028 15728
rect 121648 15384 121672 15704
rect 122004 15384 122028 15704
rect 121648 15360 122028 15384
rect 167518 15706 167898 15730
rect 167518 15386 167542 15706
rect 167874 15386 167898 15706
rect 167518 15362 167898 15386
rect 180518 15706 180898 15730
rect 180518 15386 180542 15706
rect 180874 15386 180898 15706
rect 180518 15362 180898 15386
rect 189518 15706 189898 15730
rect 189518 15386 189542 15706
rect 189874 15386 189898 15706
rect 189518 15362 189898 15386
rect 198518 15706 198898 15730
rect 198518 15386 198542 15706
rect 198874 15386 198898 15706
rect 198518 15362 198898 15386
rect 204518 15706 204898 15730
rect 204518 15386 204542 15706
rect 204874 15386 204898 15706
rect 204518 15362 204898 15386
rect 211518 15706 211898 15730
rect 211518 15386 211542 15706
rect 211874 15386 211898 15706
rect 211518 15362 211898 15386
rect 223518 15706 223898 15730
rect 223518 15386 223542 15706
rect 223874 15386 223898 15706
rect 223518 15362 223898 15386
rect 232518 15706 232898 15730
rect 232518 15386 232542 15706
rect 232874 15386 232898 15706
rect 232518 15362 232898 15386
rect 238518 15706 238898 15730
rect 238518 15386 238542 15706
rect 238874 15386 238898 15706
rect 238518 15362 238898 15386
rect 250518 15706 250898 15730
rect 250518 15386 250542 15706
rect 250874 15386 250898 15706
rect 250518 15362 250898 15386
rect 263918 15706 264298 15730
rect 263918 15386 263942 15706
rect 264274 15386 264298 15706
rect 263918 15362 264298 15386
rect 269918 15706 270298 15730
rect 269918 15386 269942 15706
rect 270274 15386 270298 15706
rect 269918 15362 270298 15386
rect 272918 15706 273298 15730
rect 272918 15386 272942 15706
rect 273274 15386 273298 15706
rect 272918 15362 273298 15386
rect 275918 15706 276298 15730
rect 275918 15386 275942 15706
rect 276274 15386 276298 15706
rect 275918 15362 276298 15386
rect 281918 15706 282298 15730
rect 281918 15386 281942 15706
rect 282274 15386 282298 15706
rect 281918 15362 282298 15386
rect 285918 15706 286298 15730
rect 285918 15386 285942 15706
rect 286274 15386 286298 15706
rect 285918 15362 286298 15386
rect 293918 15706 294298 15730
rect 293918 15386 293942 15706
rect 294274 15386 294298 15706
rect 293918 15362 294298 15386
rect 296918 15706 297298 15730
rect 296918 15386 296942 15706
rect 297274 15386 297298 15706
rect 296918 15362 297298 15386
rect 299918 15706 300298 15730
rect 299918 15386 299942 15706
rect 300274 15386 300298 15706
rect 299918 15362 300298 15386
rect 302918 15706 303298 15730
rect 302918 15386 302942 15706
rect 303274 15386 303298 15706
rect 302918 15362 303298 15386
rect 303842 15692 304210 15716
rect 303842 15372 303866 15692
rect 304186 15372 304210 15692
rect 303842 15348 304210 15372
rect 24 15298 392 15322
use pixel_array100x100  pixel_array100x100_0
timestamp 1757995770
transform 1 0 2108 0 1 317378
box -3000 -298600 300740 5000
use shift_register  shift_register_0
timestamp 1757709129
transform 0 1 -21072 -1 0 323984
box -1076 -4 307988 16000
use shift_registerC  shift_registerC_0
timestamp 1757709129
transform 1 0 58 0 1 590
box -1076 -4 307988 16000
<< labels >>
rlabel metal5 -2842 18750 -2834 18760 1 VDD
port 1 n
rlabel metal5 -1354 19538 -1354 19538 1 GND
port 2 n
rlabel space 306642 6498 306642 6498 1 COL_ENA
port 3 n
rlabel metal3 306826 6496 306826 6496 1 COL_ENA
port 3 n
rlabel metal3 306748 10568 306748 10568 1 COL_RST
port 4 n
rlabel metal3 306704 14532 306704 14532 1 COL_DIN
port 5 n
rlabel metal3 306718 2558 306718 2558 1 COL_CLK
port 6 n
rlabel metal3 196 8622 316 8742 1 COL_DOUT
port 7 n
rlabel metal4 -4276 14472 -4276 14472 1 CSA_VREF
port 8 n
rlabel metal2 304782 19400 304782 19400 1 ARRAY_OUT
port 9 n
rlabel metal2 1414 325058 1414 325058 1 NB1
port 10 n
rlabel metal2 2166 325646 2166 325646 1 NB2
port 11 n
rlabel metal4 -7482 325904 -7482 325904 1 VBIAS
port 12 n
rlabel metal2 -7646 325424 -7614 325458 1 VREF
port 13 n
rlabel metal3 942 325236 942 325236 1 SF_IB
port 14 n
rlabel metal3 -7150 17524 -7150 17524 1 ROW_DIN
port 16 n
rlabel metal3 -11058 17572 -11058 17572 1 ROW_RST
port 17 n
rlabel metal3 -15162 17518 -15162 17518 1 ROW_ENA
port 18 n
rlabel metal3 -19086 17484 -19086 17484 1 ROW_CLK
port 19 n
rlabel metal5 666 320402 666 320402 1 gring
port 20 n
<< end >>
