** sch_path: /home/hni/TopmetalSe-Respin/xschem/array3.sch
.subckt array3 VDD GND SF_IB gring VBIAS ARRAY_OUT ROW_SEL[0] ROW_SEL[1] ROW_SEL[2] VREF PIX_IN[0] PIX_IN[1] PIX_IN[2] PIX_IN[3]
+ PIX_IN[4] PIX_IN[5] PIX_IN[6] PIX_IN[7] PIX_IN[8] NB2 NB1 CSA_VREF COL_SEL[0] COL_SEL[1] COL_SEL[2]
*.PININFO VDD:I GND:I SF_IB:I gring:I VBIAS:I ARRAY_OUT:O ROW_SEL[0:2]:I VREF:I PIX_IN[0:8]:I NB2:I NB1:I CSA_VREF:I
*+ COL_SEL[0:2]:I
xPix0 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[0] VREF PIX_IN[0] NB2 NB1 CSA_VREF pixel
xPix1 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[0] VREF PIX_IN[1] NB2 NB1 CSA_VREF pixel
xPix2 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[0] VREF PIX_IN[2] NB2 NB1 CSA_VREF pixel
xPix3 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[1] VREF PIX_IN[3] NB2 NB1 CSA_VREF pixel
xPix4 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[1] VREF PIX_IN[4] NB2 NB1 CSA_VREF pixel
xPix5 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[1] VREF PIX_IN[5] NB2 NB1 CSA_VREF pixel
xPix6 VDD GND SF_IB gring VBIAS COL_OUT[0] ROW_SEL[2] VREF PIX_IN[6] NB2 NB1 CSA_VREF pixel
xPix7 VDD GND SF_IB gring VBIAS COL_OUT[1] ROW_SEL[2] VREF PIX_IN[7] NB2 NB1 CSA_VREF pixel
xPix8 VDD GND SF_IB gring VBIAS COL_OUT[2] ROW_SEL[2] VREF PIX_IN[8] NB2 NB1 CSA_VREF pixel
XM0 COL_OUT[0] COL_SEL[0] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 m=1
XM1 COL_OUT[1] COL_SEL[1] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 m=1
XM2 COL_OUT[2] COL_SEL[2] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=1 m=1
.ends

* expanding   symbol:  pixel/pixel.sym # of pins=12
** sym_path: /home/hni/TopmetalSe-Respin/xschem/pixel/pixel.sym
** sch_path: /home/hni/TopmetalSe-Respin/xschem/pixel/pixel.sch
.subckt pixel VDD GND SF_IB gring VBIAS pix_out ROW_SEL VREF AMP_IN NB2 NB1 CSA_VREF
*.PININFO pix_out:O SF_IB:I ROW_SEL:I VREF:I AMP_IN:I NB1:I CSA_VREF:I VBIAS:I NB2:I VDD:I GND:I gring:I
XM2 net2 ROW_SEL pix_out GND sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 m=1
XM3 GND AMP_OUT net1 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XM5 net1 SF_IB VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XM7 VDD net1 net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM1 VDD net6 AMP_OUT GND sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM8 net5 net5 net7 VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM10 net8 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM11 net7 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM15 AMP_OUT NB2 GND GND sky130_fd_pr__nfet_01v8_lvt L=1.15 W=1 nf=1 m=1
XM16 net4 NB1 GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=1.2 nf=1 m=1
XC3 AMP_IN AMP_OUT sky130_fd_pr__cap_mim_m3_1 W=2 L=2 m=1
XM4 net3 VREF net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7 nf=1 m=1
XM6 AMP_IN CSA_VREF AMP_OUT VDD sky130_fd_pr__pfet_01v8_lvt L=7.95 W=0.42 nf=1 m=1
XM9 net6 net5 net8 VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM12 net5 VBIAS net3 GND sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 m=1
XM13 net9 AMP_IN net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7 nf=1 m=1
XM14 net6 VBIAS net9 GND sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 m=1
XMD_4 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.6 nf=1 m=1
XMD_1 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
XMD_2 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt L=3.35 W=2 nf=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
