magic
tech sky130A
magscale 1 2
timestamp 1758314889
<< metal1 >>
rect 302440 324532 302792 324614
rect 302440 324332 302508 324532
rect 302708 324332 302792 324532
rect 302440 324258 302792 324332
rect 302508 321358 302708 324258
rect 303888 321358 304300 322140
rect 302508 321038 303926 321358
rect 304246 321038 304300 321358
rect 108 319922 308 320310
rect 302508 320098 302708 321038
rect 102 319722 108 319922
rect 308 319722 314 319922
rect 102 319700 314 319722
rect 108 319450 308 319700
rect 303888 318358 304300 321038
rect 302536 318038 303926 318358
rect 304246 318038 304300 318358
rect 108 316942 308 317310
rect 76 316922 354 316942
rect 76 316722 108 316922
rect 308 316722 354 316922
rect 76 316670 354 316722
rect 108 316450 308 316670
rect 303888 315358 304300 318038
rect 302536 315038 303926 315358
rect 304246 315038 304300 315358
rect 108 313960 308 314310
rect 82 313922 350 313960
rect 82 313722 108 313922
rect 308 313722 350 313922
rect 82 313682 350 313722
rect 108 313450 308 313682
rect 303888 312358 304300 315038
rect 302536 312038 303926 312358
rect 304246 312038 304300 312358
rect 108 310934 308 311310
rect 76 310922 334 310934
rect 76 310722 108 310922
rect 308 310722 334 310922
rect 76 310692 334 310722
rect 108 310450 308 310692
rect 303888 309358 304300 312038
rect 302536 309038 303926 309358
rect 304246 309038 304300 309358
rect 108 307922 308 308310
rect 102 307722 108 307922
rect 308 307722 314 307922
rect 102 307700 314 307722
rect 108 307450 308 307700
rect 303888 306358 304300 309038
rect 302536 306038 303926 306358
rect 304246 306038 304300 306358
rect 108 304922 308 305310
rect 102 304722 108 304922
rect 308 304722 314 304922
rect 102 304700 314 304722
rect 108 304450 308 304700
rect 303888 303358 304300 306038
rect 302536 303038 303926 303358
rect 304246 303038 304300 303358
rect 108 301922 308 302310
rect 102 301722 108 301922
rect 308 301722 314 301922
rect 102 301700 314 301722
rect 108 301450 308 301700
rect 303888 300358 304300 303038
rect 302536 300038 303926 300358
rect 304246 300038 304300 300358
rect 108 298922 308 299310
rect 102 298722 108 298922
rect 308 298722 314 298922
rect 102 298700 314 298722
rect 108 298450 308 298700
rect 303888 297358 304300 300038
rect 302536 297038 303926 297358
rect 304246 297038 304300 297358
rect 108 295922 308 296310
rect 102 295722 108 295922
rect 308 295722 314 295922
rect 102 295700 314 295722
rect 108 295450 308 295700
rect 303888 294358 304300 297038
rect 302536 294038 303926 294358
rect 304246 294038 304300 294358
rect 108 292922 308 293310
rect 102 292722 108 292922
rect 308 292722 314 292922
rect 102 292700 314 292722
rect 108 292450 308 292700
rect 303888 291358 304300 294038
rect 302536 291038 303926 291358
rect 304246 291038 304300 291358
rect 108 289922 308 290310
rect 102 289722 108 289922
rect 308 289722 314 289922
rect 102 289700 314 289722
rect 108 289450 308 289700
rect 303888 288358 304300 291038
rect 302536 288038 303926 288358
rect 304246 288038 304300 288358
rect 108 286922 308 287310
rect 102 286722 108 286922
rect 308 286722 314 286922
rect 102 286700 314 286722
rect 108 286450 308 286700
rect 303888 285358 304300 288038
rect 302536 285038 303926 285358
rect 304246 285038 304300 285358
rect 108 283922 308 284310
rect 102 283722 108 283922
rect 308 283722 314 283922
rect 102 283700 314 283722
rect 108 283450 308 283700
rect 303888 282358 304300 285038
rect 302536 282038 303926 282358
rect 304246 282038 304300 282358
rect 108 280922 308 281310
rect 102 280722 108 280922
rect 308 280722 314 280922
rect 102 280700 314 280722
rect 108 280450 308 280700
rect 303888 279358 304300 282038
rect 302536 279038 303926 279358
rect 304246 279038 304300 279358
rect 108 277922 308 278310
rect 102 277722 108 277922
rect 308 277722 314 277922
rect 102 277700 314 277722
rect 108 277450 308 277700
rect 303888 276358 304300 279038
rect 302536 276038 303926 276358
rect 304246 276038 304300 276358
rect 108 274922 308 275310
rect 102 274722 108 274922
rect 308 274722 314 274922
rect 102 274700 314 274722
rect 108 274450 308 274700
rect 303888 273358 304300 276038
rect 302536 273038 303926 273358
rect 304246 273038 304300 273358
rect 108 271922 308 272310
rect 102 271722 108 271922
rect 308 271722 314 271922
rect 102 271700 314 271722
rect 108 271450 308 271700
rect 303888 270358 304300 273038
rect 302536 270038 303926 270358
rect 304246 270038 304300 270358
rect 108 268922 308 269310
rect 102 268722 108 268922
rect 308 268722 314 268922
rect 102 268700 314 268722
rect 108 268450 308 268700
rect 303888 267358 304300 270038
rect 302536 267038 303926 267358
rect 304246 267038 304300 267358
rect 108 265922 308 266310
rect 102 265722 108 265922
rect 308 265722 314 265922
rect 102 265700 314 265722
rect 108 265450 308 265700
rect 303888 264358 304300 267038
rect 302536 264038 303926 264358
rect 304246 264038 304300 264358
rect 108 262922 308 263310
rect 102 262722 108 262922
rect 308 262722 314 262922
rect 102 262700 314 262722
rect 108 262450 308 262700
rect 303888 261358 304300 264038
rect 302536 261038 303926 261358
rect 304246 261038 304300 261358
rect 108 259922 308 260310
rect 102 259722 108 259922
rect 308 259722 314 259922
rect 102 259700 314 259722
rect 108 259450 308 259700
rect 303888 258358 304300 261038
rect 302536 258038 303926 258358
rect 304246 258038 304300 258358
rect 108 256922 308 257310
rect 102 256722 108 256922
rect 308 256722 314 256922
rect 102 256700 314 256722
rect 108 256450 308 256700
rect 303888 255358 304300 258038
rect 302536 255038 303926 255358
rect 304246 255038 304300 255358
rect 108 253922 308 254310
rect 102 253722 108 253922
rect 308 253722 314 253922
rect 102 253700 314 253722
rect 108 253450 308 253700
rect 303888 252358 304300 255038
rect 302536 252038 303926 252358
rect 304246 252038 304300 252358
rect 108 250922 308 251310
rect 102 250722 108 250922
rect 308 250722 314 250922
rect 102 250700 314 250722
rect 108 250450 308 250700
rect 303888 249358 304300 252038
rect 302536 249038 303926 249358
rect 304246 249038 304300 249358
rect 108 247922 308 248310
rect 102 247722 108 247922
rect 308 247722 314 247922
rect 102 247700 314 247722
rect 108 247450 308 247700
rect 303888 246358 304300 249038
rect 302536 246038 303926 246358
rect 304246 246038 304300 246358
rect 108 244922 308 245310
rect 102 244722 108 244922
rect 308 244722 314 244922
rect 102 244700 314 244722
rect 108 244450 308 244700
rect 303888 243358 304300 246038
rect 302536 243038 303926 243358
rect 304246 243038 304300 243358
rect 108 241922 308 242310
rect 102 241722 108 241922
rect 308 241722 314 241922
rect 102 241700 314 241722
rect 108 241450 308 241700
rect 303888 240358 304300 243038
rect 302536 240038 303926 240358
rect 304246 240038 304300 240358
rect 108 238922 308 239310
rect 102 238722 108 238922
rect 308 238722 314 238922
rect 102 238700 314 238722
rect 108 238450 308 238700
rect 303888 237358 304300 240038
rect 302536 237038 303926 237358
rect 304246 237038 304300 237358
rect 108 235922 308 236310
rect 102 235722 108 235922
rect 308 235722 314 235922
rect 102 235700 314 235722
rect 108 235450 308 235700
rect 303888 234358 304300 237038
rect 302536 234038 303926 234358
rect 304246 234038 304300 234358
rect 108 232922 308 233310
rect 102 232722 108 232922
rect 308 232722 314 232922
rect 102 232700 314 232722
rect 108 232450 308 232700
rect 303888 231358 304300 234038
rect 302536 231038 303926 231358
rect 304246 231038 304300 231358
rect 108 229922 308 230310
rect 102 229722 108 229922
rect 308 229722 314 229922
rect 102 229700 314 229722
rect 108 229450 308 229700
rect 303888 228358 304300 231038
rect 302536 228038 303926 228358
rect 304246 228038 304300 228358
rect 108 226922 308 227310
rect 102 226722 108 226922
rect 308 226722 314 226922
rect 102 226700 314 226722
rect 108 226450 308 226700
rect 303888 225358 304300 228038
rect 302536 225038 303926 225358
rect 304246 225038 304300 225358
rect 108 223922 308 224310
rect 102 223722 108 223922
rect 308 223722 314 223922
rect 102 223700 314 223722
rect 108 223450 308 223700
rect 303888 222358 304300 225038
rect 302536 222038 303926 222358
rect 304246 222038 304300 222358
rect 108 220922 308 221310
rect 102 220722 108 220922
rect 308 220722 314 220922
rect 102 220700 314 220722
rect 108 220450 308 220700
rect 303888 219358 304300 222038
rect 302536 219038 303926 219358
rect 304246 219038 304300 219358
rect 108 217922 308 218310
rect 102 217722 108 217922
rect 308 217722 314 217922
rect 102 217700 314 217722
rect 108 217450 308 217700
rect 303888 216358 304300 219038
rect 302536 216038 303926 216358
rect 304246 216038 304300 216358
rect 108 214922 308 215310
rect 102 214722 108 214922
rect 308 214722 314 214922
rect 102 214700 314 214722
rect 108 214450 308 214700
rect 303888 213358 304300 216038
rect 302536 213038 303926 213358
rect 304246 213038 304300 213358
rect 108 211922 308 212310
rect 102 211722 108 211922
rect 308 211722 314 211922
rect 102 211700 314 211722
rect 108 211450 308 211700
rect 303888 210358 304300 213038
rect 302536 210038 303926 210358
rect 304246 210038 304300 210358
rect 108 208922 308 209310
rect 102 208722 108 208922
rect 308 208722 314 208922
rect 102 208700 314 208722
rect 108 208450 308 208700
rect 303888 207358 304300 210038
rect 302536 207038 303926 207358
rect 304246 207038 304300 207358
rect 108 205922 308 206310
rect 102 205722 108 205922
rect 308 205722 314 205922
rect 102 205700 314 205722
rect 108 205450 308 205700
rect 303888 204358 304300 207038
rect 302536 204038 303926 204358
rect 304246 204038 304300 204358
rect 108 202922 308 203310
rect 102 202722 108 202922
rect 308 202722 314 202922
rect 102 202700 314 202722
rect 108 202450 308 202700
rect 303888 201358 304300 204038
rect 302536 201038 303926 201358
rect 304246 201038 304300 201358
rect 108 199922 308 200310
rect 102 199722 108 199922
rect 308 199722 314 199922
rect 102 199700 314 199722
rect 108 199450 308 199700
rect 303888 198358 304300 201038
rect 302536 198038 303926 198358
rect 304246 198038 304300 198358
rect 108 196922 308 197310
rect 102 196722 108 196922
rect 308 196722 314 196922
rect 102 196700 314 196722
rect 108 196450 308 196700
rect 303888 195358 304300 198038
rect 302536 195038 303926 195358
rect 304246 195038 304300 195358
rect 108 193922 308 194310
rect 102 193722 108 193922
rect 308 193722 314 193922
rect 102 193700 314 193722
rect 108 193450 308 193700
rect 303888 192358 304300 195038
rect 302536 192038 303926 192358
rect 304246 192038 304300 192358
rect 108 190922 308 191310
rect 102 190722 108 190922
rect 308 190722 314 190922
rect 102 190700 314 190722
rect 108 190450 308 190700
rect 303888 189358 304300 192038
rect 302536 189038 303926 189358
rect 304246 189038 304300 189358
rect 108 187922 308 188310
rect 102 187722 108 187922
rect 308 187722 314 187922
rect 102 187700 314 187722
rect 108 187450 308 187700
rect 303888 186358 304300 189038
rect 302536 186038 303926 186358
rect 304246 186038 304300 186358
rect 108 184922 308 185310
rect 102 184722 108 184922
rect 308 184722 314 184922
rect 102 184700 314 184722
rect 108 184450 308 184700
rect 303888 183358 304300 186038
rect 302536 183038 303926 183358
rect 304246 183038 304300 183358
rect 108 181922 308 182310
rect 102 181722 108 181922
rect 308 181722 314 181922
rect 102 181700 314 181722
rect 108 181450 308 181700
rect 303888 180358 304300 183038
rect 302536 180038 303926 180358
rect 304246 180038 304300 180358
rect 108 178922 308 179310
rect 102 178722 108 178922
rect 308 178722 314 178922
rect 102 178700 314 178722
rect 108 178450 308 178700
rect 303888 177358 304300 180038
rect 302536 177038 303926 177358
rect 304246 177038 304300 177358
rect 108 175922 308 176310
rect 102 175722 108 175922
rect 308 175722 314 175922
rect 102 175700 314 175722
rect 108 175450 308 175700
rect 303888 174358 304300 177038
rect 302536 174038 303926 174358
rect 304246 174038 304300 174358
rect 108 172922 308 173310
rect 102 172722 108 172922
rect 308 172722 314 172922
rect 102 172700 314 172722
rect 108 172450 308 172700
rect 303888 171358 304300 174038
rect 302536 171038 303926 171358
rect 304246 171038 304300 171358
rect 108 169922 308 170310
rect 102 169722 108 169922
rect 308 169722 314 169922
rect 102 169700 314 169722
rect 108 169450 308 169700
rect 303888 168358 304300 171038
rect 302536 168038 303926 168358
rect 304246 168038 304300 168358
rect 108 166922 308 167310
rect 102 166722 108 166922
rect 308 166722 314 166922
rect 102 166700 314 166722
rect 108 166450 308 166700
rect 303888 165358 304300 168038
rect 302536 165038 303926 165358
rect 304246 165038 304300 165358
rect 108 163922 308 164310
rect 102 163722 108 163922
rect 308 163722 314 163922
rect 102 163700 314 163722
rect 108 163450 308 163700
rect 303888 162358 304300 165038
rect 302536 162038 303926 162358
rect 304246 162038 304300 162358
rect 108 160922 308 161310
rect 102 160722 108 160922
rect 308 160722 314 160922
rect 102 160700 314 160722
rect 108 160450 308 160700
rect 303888 159358 304300 162038
rect 302536 159038 303926 159358
rect 304246 159038 304300 159358
rect 108 157922 308 158310
rect 102 157722 108 157922
rect 308 157722 314 157922
rect 102 157700 314 157722
rect 108 157450 308 157700
rect 303888 156358 304300 159038
rect 302536 156038 303926 156358
rect 304246 156038 304300 156358
rect 108 154922 308 155310
rect 102 154722 108 154922
rect 308 154722 314 154922
rect 102 154700 314 154722
rect 108 154450 308 154700
rect 303888 153358 304300 156038
rect 302536 153038 303926 153358
rect 304246 153038 304300 153358
rect 108 151922 308 152310
rect 102 151722 108 151922
rect 308 151722 314 151922
rect 102 151700 314 151722
rect 108 151450 308 151700
rect 303888 150358 304300 153038
rect 302536 150038 303926 150358
rect 304246 150038 304300 150358
rect 108 148922 308 149310
rect 102 148722 108 148922
rect 308 148722 314 148922
rect 102 148700 314 148722
rect 108 148450 308 148700
rect 303888 147358 304300 150038
rect 302536 147038 303926 147358
rect 304246 147038 304300 147358
rect 108 145922 308 146310
rect 102 145722 108 145922
rect 308 145722 314 145922
rect 102 145700 314 145722
rect 108 145450 308 145700
rect 303888 144358 304300 147038
rect 302536 144038 303926 144358
rect 304246 144038 304300 144358
rect 108 142922 308 143310
rect 102 142722 108 142922
rect 308 142722 314 142922
rect 102 142700 314 142722
rect 108 142450 308 142700
rect 303888 141358 304300 144038
rect 302536 141038 303926 141358
rect 304246 141038 304300 141358
rect 108 139922 308 140310
rect 102 139722 108 139922
rect 308 139722 314 139922
rect 102 139700 314 139722
rect 108 139450 308 139700
rect 303888 138358 304300 141038
rect 302536 138038 303926 138358
rect 304246 138038 304300 138358
rect 108 136922 308 137310
rect 102 136722 108 136922
rect 308 136722 314 136922
rect 102 136700 314 136722
rect 108 136450 308 136700
rect 303888 135358 304300 138038
rect 302536 135038 303926 135358
rect 304246 135038 304300 135358
rect 108 133922 308 134310
rect 102 133722 108 133922
rect 308 133722 314 133922
rect 102 133700 314 133722
rect 108 133450 308 133700
rect 303888 132358 304300 135038
rect 302536 132038 303926 132358
rect 304246 132038 304300 132358
rect 108 130922 308 131310
rect 102 130722 108 130922
rect 308 130722 314 130922
rect 102 130700 314 130722
rect 108 130450 308 130700
rect 303888 129358 304300 132038
rect 302536 129038 303926 129358
rect 304246 129038 304300 129358
rect 108 127922 308 128310
rect 102 127722 108 127922
rect 308 127722 314 127922
rect 102 127700 314 127722
rect 108 127450 308 127700
rect 303888 126358 304300 129038
rect 302536 126038 303926 126358
rect 304246 126038 304300 126358
rect 108 124922 308 125310
rect 102 124722 108 124922
rect 308 124722 314 124922
rect 102 124700 314 124722
rect 108 124450 308 124700
rect 303888 123358 304300 126038
rect 302536 123038 303926 123358
rect 304246 123038 304300 123358
rect 108 121922 308 122310
rect 102 121722 108 121922
rect 308 121722 314 121922
rect 102 121700 314 121722
rect 108 121450 308 121700
rect 303888 120358 304300 123038
rect 302536 120038 303926 120358
rect 304246 120038 304300 120358
rect 108 118922 308 119310
rect 102 118722 108 118922
rect 308 118722 314 118922
rect 102 118700 314 118722
rect 108 118450 308 118700
rect 303888 117358 304300 120038
rect 302536 117038 303926 117358
rect 304246 117038 304300 117358
rect 108 115922 308 116310
rect 102 115722 108 115922
rect 308 115722 314 115922
rect 102 115700 314 115722
rect 108 115450 308 115700
rect 303888 114358 304300 117038
rect 302536 114038 303926 114358
rect 304246 114038 304300 114358
rect 108 112922 308 113310
rect 102 112722 108 112922
rect 308 112722 314 112922
rect 102 112700 314 112722
rect 108 112450 308 112700
rect 303888 111358 304300 114038
rect 302536 111038 303926 111358
rect 304246 111038 304300 111358
rect 108 109922 308 110310
rect 102 109722 108 109922
rect 308 109722 314 109922
rect 102 109700 314 109722
rect 108 109450 308 109700
rect 303888 108358 304300 111038
rect 302536 108038 303926 108358
rect 304246 108038 304300 108358
rect 108 106922 308 107310
rect 102 106722 108 106922
rect 308 106722 314 106922
rect 102 106700 314 106722
rect 108 106450 308 106700
rect 303888 105358 304300 108038
rect 302536 105038 303926 105358
rect 304246 105038 304300 105358
rect 108 103922 308 104310
rect 102 103722 108 103922
rect 308 103722 314 103922
rect 102 103700 314 103722
rect 108 103450 308 103700
rect 303888 102358 304300 105038
rect 302536 102038 303926 102358
rect 304246 102038 304300 102358
rect 108 100922 308 101310
rect 102 100722 108 100922
rect 308 100722 314 100922
rect 102 100700 314 100722
rect 108 100450 308 100700
rect 303888 99358 304300 102038
rect 302536 99038 303926 99358
rect 304246 99038 304300 99358
rect 108 97922 308 98310
rect 102 97722 108 97922
rect 308 97722 314 97922
rect 102 97700 314 97722
rect 108 97450 308 97700
rect 303888 96358 304300 99038
rect 302536 96038 303926 96358
rect 304246 96038 304300 96358
rect 108 94922 308 95310
rect 102 94722 108 94922
rect 308 94722 314 94922
rect 102 94700 314 94722
rect 108 94450 308 94700
rect 303888 93358 304300 96038
rect 302536 93038 303926 93358
rect 304246 93038 304300 93358
rect 108 91922 308 92310
rect 102 91722 108 91922
rect 308 91722 314 91922
rect 102 91700 314 91722
rect 108 91450 308 91700
rect 303888 90358 304300 93038
rect 302536 90038 303926 90358
rect 304246 90038 304300 90358
rect 108 88922 308 89310
rect 102 88722 108 88922
rect 308 88722 314 88922
rect 102 88700 314 88722
rect 108 88450 308 88700
rect 303888 87358 304300 90038
rect 302536 87038 303926 87358
rect 304246 87038 304300 87358
rect 108 85922 308 86310
rect 102 85722 108 85922
rect 308 85722 314 85922
rect 102 85700 314 85722
rect 108 85450 308 85700
rect 303888 84358 304300 87038
rect 302536 84038 303926 84358
rect 304246 84038 304300 84358
rect 108 82922 308 83310
rect 102 82722 108 82922
rect 308 82722 314 82922
rect 102 82700 314 82722
rect 108 82450 308 82700
rect 303888 81358 304300 84038
rect 302536 81038 303926 81358
rect 304246 81038 304300 81358
rect 108 79922 308 80310
rect 102 79722 108 79922
rect 308 79722 314 79922
rect 102 79700 314 79722
rect 108 79450 308 79700
rect 303888 78358 304300 81038
rect 302536 78038 303926 78358
rect 304246 78038 304300 78358
rect 108 76922 308 77310
rect 102 76722 108 76922
rect 308 76722 314 76922
rect 102 76700 314 76722
rect 108 76450 308 76700
rect 303888 75358 304300 78038
rect 302536 75038 303926 75358
rect 304246 75038 304300 75358
rect 108 73922 308 74310
rect 102 73722 108 73922
rect 308 73722 314 73922
rect 102 73700 314 73722
rect 108 73450 308 73700
rect 303888 72358 304300 75038
rect 302536 72038 303926 72358
rect 304246 72038 304300 72358
rect 108 70922 308 71310
rect 102 70722 108 70922
rect 308 70722 314 70922
rect 102 70700 314 70722
rect 108 70450 308 70700
rect 303888 69358 304300 72038
rect 302536 69038 303926 69358
rect 304246 69038 304300 69358
rect 108 67922 308 68310
rect 102 67722 108 67922
rect 308 67722 314 67922
rect 102 67700 314 67722
rect 108 67450 308 67700
rect 303888 66358 304300 69038
rect 302536 66038 303926 66358
rect 304246 66038 304300 66358
rect 108 64922 308 65310
rect 102 64722 108 64922
rect 308 64722 314 64922
rect 102 64700 314 64722
rect 108 64450 308 64700
rect 303888 63358 304300 66038
rect 302536 63038 303926 63358
rect 304246 63038 304300 63358
rect 108 61922 308 62310
rect 102 61722 108 61922
rect 308 61722 314 61922
rect 102 61700 314 61722
rect 108 61450 308 61700
rect 303888 60358 304300 63038
rect 302536 60038 303926 60358
rect 304246 60038 304300 60358
rect 108 58922 308 59310
rect 102 58722 108 58922
rect 308 58722 314 58922
rect 102 58700 314 58722
rect 108 58450 308 58700
rect 303888 57358 304300 60038
rect 302536 57038 303926 57358
rect 304246 57038 304300 57358
rect 108 55922 308 56310
rect 102 55722 108 55922
rect 308 55722 314 55922
rect 102 55700 314 55722
rect 108 55450 308 55700
rect 303888 54358 304300 57038
rect 302536 54038 303926 54358
rect 304246 54038 304300 54358
rect 108 52922 308 53310
rect 102 52722 108 52922
rect 308 52722 314 52922
rect 102 52700 314 52722
rect 108 52450 308 52700
rect 303888 51358 304300 54038
rect 302536 51038 303926 51358
rect 304246 51038 304300 51358
rect 108 49922 308 50310
rect 102 49722 108 49922
rect 308 49722 314 49922
rect 102 49700 314 49722
rect 108 49450 308 49700
rect 303888 48358 304300 51038
rect 302536 48038 303926 48358
rect 304246 48038 304300 48358
rect 108 46922 308 47310
rect 102 46722 108 46922
rect 308 46722 314 46922
rect 102 46700 314 46722
rect 108 46450 308 46700
rect 303888 45358 304300 48038
rect 302536 45038 303926 45358
rect 304246 45038 304300 45358
rect 108 43922 308 44310
rect 102 43722 108 43922
rect 308 43722 314 43922
rect 102 43700 314 43722
rect 108 43450 308 43700
rect 303888 42358 304300 45038
rect 302536 42038 303926 42358
rect 304246 42038 304300 42358
rect 108 40922 308 41310
rect 102 40722 108 40922
rect 308 40722 314 40922
rect 102 40700 314 40722
rect 108 40450 308 40700
rect 303888 39358 304300 42038
rect 302536 39038 303926 39358
rect 304246 39038 304300 39358
rect 108 37922 308 38310
rect 102 37722 108 37922
rect 308 37722 314 37922
rect 102 37700 314 37722
rect 108 37450 308 37700
rect 303888 36358 304300 39038
rect 302536 36038 303926 36358
rect 304246 36038 304300 36358
rect 108 34922 308 35310
rect 102 34722 108 34922
rect 308 34722 314 34922
rect 102 34700 314 34722
rect 108 34450 308 34700
rect 303888 33358 304300 36038
rect 302536 33038 303926 33358
rect 304246 33038 304300 33358
rect 108 31938 308 32310
rect 72 31922 352 31938
rect 72 31722 108 31922
rect 308 31722 352 31922
rect 72 31684 352 31722
rect 108 31450 308 31684
rect 303888 30358 304300 33038
rect 302536 30038 303926 30358
rect 304246 30038 304300 30358
rect 108 28944 308 29310
rect 82 28922 354 28944
rect 82 28722 108 28922
rect 308 28722 354 28922
rect 82 28692 354 28722
rect 108 28450 308 28692
rect 303888 27358 304300 30038
rect 302536 27038 303926 27358
rect 304246 27038 304300 27358
rect 108 25946 308 26310
rect 70 25922 330 25946
rect 70 25722 108 25922
rect 308 25722 330 25922
rect 70 25684 330 25722
rect 108 25450 308 25684
rect 303888 24358 304300 27038
rect 302536 24038 303926 24358
rect 304246 24038 304300 24358
rect 108 22932 308 23310
rect 90 22922 338 22932
rect 90 22722 108 22922
rect 308 22722 338 22922
rect 90 22704 338 22722
rect 102 22700 314 22704
rect 108 22450 308 22700
rect 303888 21372 304300 24038
rect 303888 21358 304304 21372
rect 302536 21038 303926 21358
rect 304246 21038 304304 21358
rect 303888 21004 304304 21038
rect 303888 20952 304300 21004
rect 108 19900 308 20808
rect 302508 20408 302828 20608
rect 102 19700 314 19900
rect -6210 17946 -5984 17960
rect 108 17946 308 19700
rect -6210 17746 -6198 17946
rect -5998 17746 308 17946
rect 198548 17938 198868 18170
rect 211548 17938 211868 18300
rect 232548 17938 232868 18370
rect 238548 17938 238868 18116
rect 250548 17938 250868 18332
rect 263948 17938 264268 18238
rect 269948 17938 270268 18366
rect 272948 17938 273268 18360
rect 275948 17938 276268 18326
rect 281948 17938 282268 18316
rect 285948 17938 286268 18280
rect 293948 17938 294268 18336
rect 296948 17938 297268 18364
rect 299948 17938 300268 18392
rect 302948 18264 303268 18390
rect 302946 18258 303268 18264
rect -6210 17734 -5984 17746
rect 108 15664 308 17746
rect 302946 16448 303268 17936
rect 302888 16416 303316 16448
rect 302888 16094 302946 16416
rect 303268 16094 303316 16416
rect 302888 16036 303316 16094
rect 26 15588 390 15664
rect 26 15388 108 15588
rect 308 15388 390 15588
rect 26 15298 390 15388
<< via1 >>
rect 302508 324332 302708 324532
rect 303926 321038 304246 321358
rect 108 319722 308 319922
rect 303926 318038 304246 318358
rect 108 316722 308 316922
rect 303926 315038 304246 315358
rect 108 313722 308 313922
rect 303926 312038 304246 312358
rect 108 310722 308 310922
rect 303926 309038 304246 309358
rect 108 307722 308 307922
rect 303926 306038 304246 306358
rect 108 304722 308 304922
rect 303926 303038 304246 303358
rect 108 301722 308 301922
rect 303926 300038 304246 300358
rect 108 298722 308 298922
rect 303926 297038 304246 297358
rect 108 295722 308 295922
rect 303926 294038 304246 294358
rect 108 292722 308 292922
rect 303926 291038 304246 291358
rect 108 289722 308 289922
rect 303926 288038 304246 288358
rect 108 286722 308 286922
rect 303926 285038 304246 285358
rect 108 283722 308 283922
rect 303926 282038 304246 282358
rect 108 280722 308 280922
rect 303926 279038 304246 279358
rect 108 277722 308 277922
rect 303926 276038 304246 276358
rect 108 274722 308 274922
rect 303926 273038 304246 273358
rect 108 271722 308 271922
rect 303926 270038 304246 270358
rect 108 268722 308 268922
rect 303926 267038 304246 267358
rect 108 265722 308 265922
rect 303926 264038 304246 264358
rect 108 262722 308 262922
rect 303926 261038 304246 261358
rect 108 259722 308 259922
rect 303926 258038 304246 258358
rect 108 256722 308 256922
rect 303926 255038 304246 255358
rect 108 253722 308 253922
rect 303926 252038 304246 252358
rect 108 250722 308 250922
rect 303926 249038 304246 249358
rect 108 247722 308 247922
rect 303926 246038 304246 246358
rect 108 244722 308 244922
rect 303926 243038 304246 243358
rect 108 241722 308 241922
rect 303926 240038 304246 240358
rect 108 238722 308 238922
rect 303926 237038 304246 237358
rect 108 235722 308 235922
rect 303926 234038 304246 234358
rect 108 232722 308 232922
rect 303926 231038 304246 231358
rect 108 229722 308 229922
rect 303926 228038 304246 228358
rect 108 226722 308 226922
rect 303926 225038 304246 225358
rect 108 223722 308 223922
rect 303926 222038 304246 222358
rect 108 220722 308 220922
rect 303926 219038 304246 219358
rect 108 217722 308 217922
rect 303926 216038 304246 216358
rect 108 214722 308 214922
rect 303926 213038 304246 213358
rect 108 211722 308 211922
rect 303926 210038 304246 210358
rect 108 208722 308 208922
rect 303926 207038 304246 207358
rect 108 205722 308 205922
rect 303926 204038 304246 204358
rect 108 202722 308 202922
rect 303926 201038 304246 201358
rect 108 199722 308 199922
rect 303926 198038 304246 198358
rect 108 196722 308 196922
rect 303926 195038 304246 195358
rect 108 193722 308 193922
rect 303926 192038 304246 192358
rect 108 190722 308 190922
rect 303926 189038 304246 189358
rect 108 187722 308 187922
rect 303926 186038 304246 186358
rect 108 184722 308 184922
rect 303926 183038 304246 183358
rect 108 181722 308 181922
rect 303926 180038 304246 180358
rect 108 178722 308 178922
rect 303926 177038 304246 177358
rect 108 175722 308 175922
rect 303926 174038 304246 174358
rect 108 172722 308 172922
rect 303926 171038 304246 171358
rect 108 169722 308 169922
rect 303926 168038 304246 168358
rect 108 166722 308 166922
rect 303926 165038 304246 165358
rect 108 163722 308 163922
rect 303926 162038 304246 162358
rect 108 160722 308 160922
rect 303926 159038 304246 159358
rect 108 157722 308 157922
rect 303926 156038 304246 156358
rect 108 154722 308 154922
rect 303926 153038 304246 153358
rect 108 151722 308 151922
rect 303926 150038 304246 150358
rect 108 148722 308 148922
rect 303926 147038 304246 147358
rect 108 145722 308 145922
rect 303926 144038 304246 144358
rect 108 142722 308 142922
rect 303926 141038 304246 141358
rect 108 139722 308 139922
rect 303926 138038 304246 138358
rect 108 136722 308 136922
rect 303926 135038 304246 135358
rect 108 133722 308 133922
rect 303926 132038 304246 132358
rect 108 130722 308 130922
rect 303926 129038 304246 129358
rect 108 127722 308 127922
rect 303926 126038 304246 126358
rect 108 124722 308 124922
rect 303926 123038 304246 123358
rect 108 121722 308 121922
rect 303926 120038 304246 120358
rect 108 118722 308 118922
rect 303926 117038 304246 117358
rect 108 115722 308 115922
rect 303926 114038 304246 114358
rect 108 112722 308 112922
rect 303926 111038 304246 111358
rect 108 109722 308 109922
rect 303926 108038 304246 108358
rect 108 106722 308 106922
rect 303926 105038 304246 105358
rect 108 103722 308 103922
rect 303926 102038 304246 102358
rect 108 100722 308 100922
rect 303926 99038 304246 99358
rect 108 97722 308 97922
rect 303926 96038 304246 96358
rect 108 94722 308 94922
rect 303926 93038 304246 93358
rect 108 91722 308 91922
rect 303926 90038 304246 90358
rect 108 88722 308 88922
rect 303926 87038 304246 87358
rect 108 85722 308 85922
rect 303926 84038 304246 84358
rect 108 82722 308 82922
rect 303926 81038 304246 81358
rect 108 79722 308 79922
rect 303926 78038 304246 78358
rect 108 76722 308 76922
rect 303926 75038 304246 75358
rect 108 73722 308 73922
rect 303926 72038 304246 72358
rect 108 70722 308 70922
rect 303926 69038 304246 69358
rect 108 67722 308 67922
rect 303926 66038 304246 66358
rect 108 64722 308 64922
rect 303926 63038 304246 63358
rect 108 61722 308 61922
rect 303926 60038 304246 60358
rect 108 58722 308 58922
rect 303926 57038 304246 57358
rect 108 55722 308 55922
rect 303926 54038 304246 54358
rect 108 52722 308 52922
rect 303926 51038 304246 51358
rect 108 49722 308 49922
rect 303926 48038 304246 48358
rect 108 46722 308 46922
rect 303926 45038 304246 45358
rect 108 43722 308 43922
rect 303926 42038 304246 42358
rect 108 40722 308 40922
rect 303926 39038 304246 39358
rect 108 37722 308 37922
rect 303926 36038 304246 36358
rect 108 34722 308 34922
rect 303926 33038 304246 33358
rect 108 31722 308 31922
rect 303926 30038 304246 30358
rect 108 28722 308 28922
rect 303926 27038 304246 27358
rect 108 25722 308 25922
rect 303926 24038 304246 24358
rect 108 22722 308 22922
rect 303926 21038 304246 21358
rect -6198 17746 -5998 17946
rect 302946 17936 303268 18258
rect 302946 16094 303268 16416
rect 108 15388 308 15588
<< metal2 >>
rect -8166 325380 -1626 325490
rect -5180 322442 -2032 322532
rect -5132 319402 -2402 319458
rect -5168 316366 -2742 316422
rect -5148 313238 -3102 313294
rect -3534 310258 -3444 310274
rect -5148 310202 -3444 310258
rect -5138 307166 -3932 307222
rect -5158 304038 -4342 304094
rect -4398 302338 -4342 304038
rect -3988 303948 -3932 307166
rect -3534 306948 -3444 310202
rect -3158 309948 -3102 313238
rect -2798 312948 -2742 316366
rect -2458 315930 -2402 319402
rect -2122 318948 -2032 322442
rect -1736 320838 -1626 325380
rect 1358 321238 1468 327120
rect 2118 321418 2228 326996
rect 302440 324532 302792 324614
rect 302440 324332 302508 324532
rect 302708 324332 302792 324532
rect 302440 324258 302792 324332
rect 303888 321358 304300 322140
rect 303888 321038 303926 321358
rect 304246 321038 304300 321358
rect -1736 320728 -782 320838
rect 94 319922 358 319948
rect 94 319722 108 319922
rect 308 319722 358 319922
rect 94 319698 358 319722
rect -2122 318858 -802 318948
rect 303888 318358 304300 321038
rect 303888 318038 303926 318358
rect 304246 318038 304300 318358
rect 76 316922 354 316942
rect 76 316722 108 316922
rect 308 316722 354 316922
rect 76 316670 354 316722
rect -2458 315874 -578 315930
rect 303888 315358 304300 318038
rect 303888 315038 303926 315358
rect 304246 315038 304300 315358
rect 82 313922 350 313960
rect 82 313722 108 313922
rect 308 313722 350 313922
rect 82 313682 350 313722
rect -2798 312892 -622 312948
rect 303888 312358 304300 315038
rect 303888 312038 303926 312358
rect 304246 312038 304300 312358
rect 76 310922 334 310934
rect 76 310722 108 310922
rect 308 310722 334 310922
rect 76 310692 334 310722
rect -3164 309858 -754 309948
rect 303888 309358 304300 312038
rect 303888 309038 303926 309358
rect 304246 309038 304300 309358
rect 80 307922 328 307932
rect 80 307722 108 307922
rect 308 307722 328 307922
rect 80 307694 328 307722
rect -3534 306858 -802 306948
rect 303888 306358 304300 309038
rect 303888 306038 303926 306358
rect 304246 306038 304300 306358
rect 88 304922 358 304948
rect 88 304722 108 304922
rect 308 304722 358 304922
rect 88 304698 358 304722
rect -4004 303858 -774 303948
rect 303888 303358 304300 306038
rect 303888 303038 303926 303358
rect 304246 303038 304300 303358
rect -4398 302282 -692 302338
rect -1484 301058 -1004 301064
rect -5128 301002 -1004 301058
rect -1484 300974 -1004 301002
rect -5148 297966 -1542 298022
rect -1634 294948 -1544 297966
rect -1094 297948 -1004 300974
rect -834 300858 -744 302282
rect 98 301922 332 301954
rect 98 301722 108 301922
rect 308 301722 332 301922
rect 98 301688 332 301722
rect 303888 300358 304300 303038
rect 303888 300038 303926 300358
rect 304246 300038 304300 300358
rect 82 298922 322 298930
rect 82 298722 108 298922
rect 308 298722 322 298922
rect 82 298698 322 298722
rect -1094 297858 -744 297948
rect 303888 297358 304300 300038
rect 303888 297038 303926 297358
rect 304246 297038 304300 297358
rect 96 295922 318 295934
rect 96 295722 108 295922
rect 308 295722 318 295922
rect 96 295702 318 295722
rect -5148 294838 -2152 294894
rect -1634 294858 -724 294948
rect -3094 291858 -3004 292054
rect -2208 291918 -2152 294838
rect 303888 294358 304300 297038
rect 303888 294038 303926 294358
rect 304246 294038 304300 294358
rect 84 292922 336 292942
rect 84 292722 108 292922
rect 308 292722 336 292922
rect 84 292698 336 292722
rect -2208 291862 -452 291918
rect -5148 291802 -3004 291858
rect -3094 288948 -3004 291802
rect 303888 291358 304300 294038
rect 303888 291038 303926 291358
rect 304246 291038 304300 291358
rect 84 289922 336 289942
rect 84 289722 108 289922
rect 308 289722 336 289922
rect 84 289698 336 289722
rect -3094 288858 -784 288948
rect -3914 288730 -3824 288814
rect -5148 288674 -3824 288730
rect -3914 285948 -3824 288674
rect 303888 288358 304300 291038
rect 303888 288038 303926 288358
rect 304246 288038 304300 288358
rect 84 286922 336 286942
rect 84 286722 108 286922
rect 308 286722 336 286922
rect 84 286698 336 286722
rect -3914 285858 -764 285948
rect -5138 285638 -4232 285694
rect -4288 284088 -4232 285638
rect 303888 285358 304300 288038
rect 303888 285038 303926 285358
rect 304246 285038 304300 285358
rect -1104 284088 -1014 284104
rect -4288 284032 -962 284088
rect -1104 282948 -1014 284032
rect 84 283922 336 283942
rect 84 283722 108 283922
rect 308 283722 336 283922
rect 84 283698 336 283722
rect -1104 282858 -802 282948
rect -2204 282658 -2114 282764
rect -5158 282602 -2114 282658
rect -2204 279948 -2114 282602
rect 303888 282358 304300 285038
rect 303888 282038 303926 282358
rect 304246 282038 304300 282358
rect 84 280922 336 280942
rect 84 280722 108 280922
rect 308 280722 336 280922
rect 84 280698 336 280722
rect -2204 279858 -802 279948
rect -5218 279474 -1962 279530
rect -2054 276948 -1964 279474
rect 303888 279358 304300 282038
rect 303888 279038 303926 279358
rect 304246 279038 304300 279358
rect 84 277922 336 277942
rect 84 277722 108 277922
rect 308 277722 336 277922
rect 84 277698 336 277722
rect -2054 276858 -784 276948
rect -892 276494 -802 276524
rect -5188 276438 -802 276494
rect -892 273858 -802 276438
rect 303888 276358 304300 279038
rect 303888 276038 303926 276358
rect 304246 276038 304300 276358
rect 84 274922 336 274942
rect 84 274722 108 274922
rect 308 274722 336 274922
rect 84 274698 336 274722
rect -3964 273458 -3874 273584
rect -5228 273402 -3874 273458
rect -3964 270948 -3874 273402
rect 303888 273358 304300 276038
rect 303888 273038 303926 273358
rect 304246 273038 304300 273358
rect 84 271922 336 271942
rect 84 271722 108 271922
rect 308 271722 336 271922
rect 84 271698 336 271722
rect -3964 270858 -802 270948
rect 303888 270358 304300 273038
rect -5168 270274 -4582 270330
rect -4638 267948 -4582 270274
rect 303888 270038 303926 270358
rect 304246 270038 304300 270358
rect 84 268922 336 268942
rect 84 268722 108 268922
rect 308 268722 336 268922
rect 84 268698 336 268722
rect -4638 267882 -802 267948
rect -4614 267858 -802 267882
rect -4284 267294 -4194 267424
rect -5148 267238 -4194 267294
rect -4284 264948 -4194 267238
rect 303888 267358 304300 270038
rect 303888 267038 303926 267358
rect 304246 267038 304300 267358
rect 84 265922 336 265942
rect 84 265722 108 265922
rect 308 265722 336 265922
rect 84 265698 336 265722
rect -4284 264858 -802 264948
rect 303888 264358 304300 267038
rect -5148 264110 -1932 264166
rect -1988 261948 -1932 264110
rect 303888 264038 303926 264358
rect 304246 264038 304300 264358
rect 84 262922 336 262942
rect 84 262722 108 262922
rect 308 262722 336 262922
rect 84 262698 336 262722
rect -1988 261858 -802 261948
rect -1988 261812 -1932 261858
rect 303888 261358 304300 264038
rect -5178 261074 -1092 261130
rect -1148 258948 -1092 261074
rect 303888 261038 303926 261358
rect 304246 261038 304300 261358
rect 84 259922 336 259942
rect 84 259722 108 259922
rect 308 259722 336 259922
rect 84 259698 336 259722
rect -1148 258858 -774 258948
rect -1148 258822 -1092 258858
rect 303888 258358 304300 261038
rect -5218 258038 -1112 258094
rect -1168 255948 -1112 258038
rect 303888 258038 303926 258358
rect 304246 258038 304300 258358
rect 84 256922 336 256942
rect 84 256722 108 256922
rect 308 256722 336 256922
rect 84 256698 336 256722
rect -1168 255858 -802 255948
rect -1168 255842 -1112 255858
rect 303888 255358 304300 258038
rect 303888 255038 303926 255358
rect 304246 255038 304300 255358
rect -5168 254910 -1172 254966
rect -1228 252948 -1172 254910
rect 84 253922 336 253942
rect 84 253722 108 253922
rect 308 253722 336 253922
rect 84 253698 336 253722
rect -1228 252858 -802 252948
rect -1228 252852 -1172 252858
rect 303888 252358 304300 255038
rect 303888 252038 303926 252358
rect 304246 252038 304300 252358
rect -5208 251874 -1402 251930
rect -1458 249948 -1402 251874
rect 84 250922 336 250942
rect 84 250722 108 250922
rect 308 250722 336 250922
rect 84 250698 336 250722
rect -1458 249892 -794 249948
rect -1434 249858 -794 249892
rect 303888 249358 304300 252038
rect -884 248894 -794 249084
rect 303888 249038 303926 249358
rect 304246 249038 304300 249358
rect -5128 248838 -792 248894
rect -884 246858 -794 248838
rect 84 247922 336 247942
rect 84 247722 108 247922
rect 308 247722 336 247922
rect 84 247698 336 247722
rect 303888 246358 304300 249038
rect 303888 246038 303926 246358
rect 304246 246038 304300 246358
rect -892 245766 -802 245884
rect -5268 245710 -802 245766
rect -892 243858 -802 245710
rect 84 244922 336 244942
rect 84 244722 108 244922
rect 308 244722 336 244922
rect 84 244698 336 244722
rect 303888 243358 304300 246038
rect 303888 243038 303926 243358
rect 304246 243038 304300 243358
rect -5228 242674 -832 242730
rect -888 240852 -832 242674
rect 84 241922 336 241942
rect 84 241722 108 241922
rect 308 241722 336 241922
rect 84 241698 336 241722
rect 303888 240358 304300 243038
rect 303888 240038 303926 240358
rect 304246 240038 304300 240358
rect -5158 239638 -812 239694
rect -868 237892 -812 239638
rect 84 238922 336 238942
rect 84 238722 108 238922
rect 308 238722 336 238922
rect 84 238698 336 238722
rect 303888 237358 304300 240038
rect 303888 237038 303926 237358
rect 304246 237038 304300 237358
rect -892 236566 -802 236724
rect -5188 236510 -802 236566
rect -892 234858 -802 236510
rect 84 235922 336 235942
rect 84 235722 108 235922
rect 308 235722 336 235922
rect 84 235698 336 235722
rect 303888 234358 304300 237038
rect 303888 234038 303926 234358
rect 304246 234038 304300 234358
rect -5168 233474 -892 233530
rect -948 231852 -892 233474
rect 84 232922 336 232942
rect 84 232722 108 232922
rect 308 232722 336 232922
rect 84 232698 336 232722
rect 303888 231358 304300 234038
rect 303888 231038 303926 231358
rect 304246 231038 304300 231358
rect -5168 228948 -5112 230402
rect 84 229922 336 229942
rect 84 229722 108 229922
rect 308 229722 336 229922
rect 84 229698 336 229722
rect -5168 228892 -784 228948
rect -5154 228858 -784 228892
rect 303888 228358 304300 231038
rect 303888 228038 303926 228358
rect 304246 228038 304300 228358
rect -5138 227310 -612 227366
rect -834 225858 -744 227310
rect 84 226922 336 226942
rect 84 226722 108 226922
rect 308 226722 336 226922
rect 84 226698 336 226722
rect 303888 225358 304300 228038
rect 303888 225038 303926 225358
rect 304246 225038 304300 225358
rect -5194 224264 -802 224354
rect -892 222858 -802 224264
rect 84 223922 336 223942
rect 84 223722 108 223922
rect 308 223722 336 223922
rect 84 223698 336 223722
rect 303888 222358 304300 225038
rect 303888 222038 303926 222358
rect 304246 222038 304300 222358
rect -5148 221146 -808 221202
rect -864 219882 -808 221146
rect 84 220922 336 220942
rect 84 220722 108 220922
rect 308 220722 336 220922
rect 84 220698 336 220722
rect 303888 219358 304300 222038
rect 303888 219038 303926 219358
rect 304246 219038 304300 219358
rect -808 218178 -752 218202
rect -5128 218122 -752 218178
rect -808 216872 -752 218122
rect 84 217922 336 217942
rect 84 217722 108 217922
rect 308 217722 336 217922
rect 84 217698 336 217722
rect 303888 216358 304300 219038
rect 303888 216038 303926 216358
rect 304246 216038 304300 216358
rect -5128 215082 -752 215138
rect -808 213858 -752 215082
rect 84 214922 336 214942
rect 84 214722 108 214922
rect 308 214722 336 214922
rect 84 214698 336 214722
rect 303888 213358 304300 216038
rect 303888 213038 303926 213358
rect 304246 213038 304300 213358
rect -5134 211914 -802 212004
rect -892 210858 -802 211914
rect 84 211922 336 211942
rect 84 211722 108 211922
rect 308 211722 336 211922
rect 84 211698 336 211722
rect 303888 210358 304300 213038
rect 303888 210038 303926 210358
rect 304246 210038 304300 210358
rect -5128 208910 -732 208966
rect -892 207872 -732 208910
rect 84 208922 336 208942
rect 84 208722 108 208922
rect 308 208722 336 208922
rect 84 208698 336 208722
rect -892 207858 -764 207872
rect 303888 207358 304300 210038
rect 303888 207038 303926 207358
rect 304246 207038 304300 207358
rect 84 205922 336 205942
rect -5168 205782 -802 205838
rect -858 204842 -802 205782
rect 84 205722 108 205922
rect 308 205722 336 205922
rect 84 205698 336 205722
rect 303888 204358 304300 207038
rect 303888 204038 303926 204358
rect 304246 204038 304300 204358
rect 84 202922 336 202942
rect -5158 202746 -762 202802
rect -884 201858 -794 202746
rect 84 202722 108 202922
rect 308 202722 336 202922
rect 84 202698 336 202722
rect 303888 201358 304300 204038
rect 303888 201038 303926 201358
rect 304246 201038 304300 201358
rect 84 199922 336 199942
rect -5208 199710 -722 199766
rect -778 198852 -722 199710
rect 84 199722 108 199922
rect 308 199722 336 199922
rect 84 199698 336 199722
rect 303888 198358 304300 201038
rect 303888 198038 303926 198358
rect 304246 198038 304300 198358
rect 84 196922 336 196942
rect 84 196722 108 196922
rect 308 196722 336 196922
rect 84 196698 336 196722
rect -5144 196582 -1202 196638
rect -1258 195948 -1202 196582
rect -1258 195858 -792 195948
rect -1258 195804 -1202 195858
rect 303888 195358 304300 198038
rect 303888 195038 303926 195358
rect 304246 195038 304300 195358
rect 84 193922 336 193942
rect 84 193722 108 193922
rect 308 193722 336 193922
rect 84 193698 336 193722
rect -5144 193552 -4890 193642
rect -4980 192948 -4890 193552
rect -4980 192858 -782 192948
rect 303888 192358 304300 195038
rect 303888 192038 303926 192358
rect 304246 192038 304300 192358
rect 84 190922 336 190942
rect 84 190722 108 190922
rect 308 190722 336 190922
rect 84 190698 336 190722
rect -5134 190510 -736 190566
rect -792 189806 -736 190510
rect 303888 189358 304300 192038
rect 303888 189038 303926 189358
rect 304246 189038 304300 189358
rect 84 187922 336 187942
rect 84 187722 108 187922
rect 308 187722 336 187922
rect 84 187698 336 187722
rect -5140 186948 -5050 187460
rect -5140 186858 -792 186948
rect 303888 186358 304300 189038
rect 303888 186038 303926 186358
rect 304246 186038 304300 186358
rect 84 184922 336 184942
rect 84 184722 108 184922
rect 308 184722 336 184922
rect 84 184698 336 184722
rect -5140 183948 -5050 184424
rect -5140 183858 -578 183948
rect 303888 183358 304300 186038
rect 303888 183038 303926 183358
rect 304246 183038 304300 183358
rect 84 181922 336 181942
rect 84 181722 108 181922
rect 308 181722 336 181922
rect 84 181698 336 181722
rect -5184 180948 -5094 181338
rect -5184 180858 -802 180948
rect 303888 180358 304300 183038
rect 303888 180038 303926 180358
rect 304246 180038 304300 180358
rect 84 178922 336 178942
rect 84 178722 108 178922
rect 308 178722 336 178922
rect 84 178698 336 178722
rect -5168 177948 -5078 178234
rect -5168 177858 -572 177948
rect 303888 177358 304300 180038
rect 303888 177038 303926 177358
rect 304246 177038 304300 177358
rect 84 175922 336 175942
rect 84 175722 108 175922
rect 308 175722 336 175922
rect 84 175698 336 175722
rect -5128 174948 -5072 175202
rect -5128 174858 -690 174948
rect -5128 174790 -5072 174858
rect 303888 174358 304300 177038
rect 303888 174038 303926 174358
rect 304246 174038 304300 174358
rect 84 172922 336 172942
rect 84 172722 108 172922
rect 308 172722 336 172922
rect 84 172698 336 172722
rect -5208 171948 -5118 172064
rect -5208 171858 -782 171948
rect 303888 171358 304300 174038
rect 303888 171038 303926 171358
rect 304246 171038 304300 171358
rect 84 169922 336 169942
rect 84 169722 108 169922
rect 308 169722 336 169922
rect 84 169698 336 169722
rect -5156 168948 -5066 169080
rect -5156 168858 -802 168948
rect 303888 168358 304300 171038
rect 303888 168038 303926 168358
rect 304246 168038 304300 168358
rect 84 166922 336 166942
rect 84 166722 108 166922
rect 308 166722 336 166922
rect 84 166698 336 166722
rect -5144 165948 -5054 166032
rect -5144 165858 -730 165948
rect 303888 165358 304300 168038
rect 303888 165038 303926 165358
rect 304246 165038 304300 165358
rect 84 163922 336 163942
rect 84 163722 108 163922
rect 308 163722 336 163922
rect 84 163698 336 163722
rect -5144 162858 -770 162948
rect 303888 162358 304300 165038
rect 303888 162038 303926 162358
rect 304246 162038 304300 162358
rect 84 160922 336 160942
rect 84 160722 108 160922
rect 308 160722 336 160922
rect 84 160698 336 160722
rect -5922 159858 -798 159948
rect -5922 159778 -816 159858
rect 303888 159358 304300 162038
rect 303888 159038 303926 159358
rect 304246 159038 304300 159358
rect 84 157922 336 157942
rect 84 157722 108 157922
rect 308 157722 336 157922
rect 84 157698 336 157722
rect -826 156900 -736 156948
rect -5162 156856 -736 156900
rect -5168 156742 -736 156856
rect 303888 156358 304300 159038
rect 303888 156038 303926 156358
rect 304246 156038 304300 156358
rect 84 154922 336 154942
rect 84 154722 108 154922
rect 308 154722 336 154922
rect 84 154698 336 154722
rect -882 153678 -792 153948
rect -5134 153588 -792 153678
rect 303888 153358 304300 156038
rect 303888 153038 303926 153358
rect 304246 153038 304300 153358
rect 84 151922 336 151942
rect 84 151722 108 151922
rect 308 151722 336 151922
rect 84 151698 336 151722
rect -5242 150584 -5010 150658
rect -892 150584 -802 150948
rect -5242 150568 -802 150584
rect -5100 150494 -802 150568
rect 303888 150358 304300 153038
rect 303888 150038 303926 150358
rect 304246 150038 304300 150358
rect 84 148922 336 148942
rect 84 148722 108 148922
rect 308 148722 336 148922
rect 84 148698 336 148722
rect -5122 147428 -5032 147554
rect -882 147428 -792 147948
rect -5122 147338 -792 147428
rect 303888 147358 304300 150038
rect 303888 147038 303926 147358
rect 304246 147038 304300 147358
rect 84 145922 336 145942
rect 84 145722 108 145922
rect 308 145722 336 145922
rect 84 145698 336 145722
rect -882 144568 -792 144948
rect -5178 144478 -792 144568
rect -5178 144416 -838 144478
rect 303888 144358 304300 147038
rect 303888 144038 303926 144358
rect 304246 144038 304300 144358
rect 84 142922 336 142942
rect 84 142722 108 142922
rect 308 142722 336 142922
rect 84 142698 336 142722
rect -866 141504 -776 141948
rect -5140 141414 -776 141504
rect -5140 141352 -816 141414
rect 303888 141358 304300 144038
rect 303888 141038 303926 141358
rect 304246 141038 304300 141358
rect 84 139922 336 139942
rect 84 139722 108 139922
rect 308 139722 336 139922
rect 84 139698 336 139722
rect -860 138338 -770 138948
rect -5178 138248 -770 138338
rect 303888 138358 304300 141038
rect 303888 138038 303926 138358
rect 304246 138038 304300 138358
rect 84 136922 336 136942
rect 84 136722 108 136922
rect 308 136722 336 136922
rect 84 136698 336 136722
rect -892 135340 -802 135948
rect -5190 135250 -802 135340
rect 303888 135358 304300 138038
rect -5134 135182 -804 135250
rect 303888 135038 303926 135358
rect 304246 135038 304300 135358
rect 84 133922 336 133942
rect 84 133722 108 133922
rect 308 133722 336 133922
rect 84 133698 336 133722
rect -848 132368 -758 132948
rect -5174 132278 -758 132368
rect 303888 132358 304300 135038
rect -5174 132186 -5084 132278
rect 303888 132038 303926 132358
rect 304246 132038 304300 132358
rect 84 130922 336 130942
rect 84 130722 108 130922
rect 308 130722 336 130922
rect 84 130698 336 130722
rect -880 129084 -790 129948
rect -5186 128936 -790 129084
rect 303888 129358 304300 132038
rect 303888 129038 303926 129358
rect 304246 129038 304300 129358
rect 84 127922 336 127942
rect 84 127722 108 127922
rect 308 127722 336 127922
rect 84 127698 336 127722
rect -852 126084 -762 126948
rect -5198 125938 -762 126084
rect 303888 126358 304300 129038
rect 303888 126038 303926 126358
rect 304246 126038 304300 126358
rect 84 124922 336 124942
rect 84 124722 108 124922
rect 308 124722 336 124922
rect 84 124698 336 124722
rect -892 122976 -802 123948
rect -5140 122790 -802 122976
rect 303888 123358 304300 126038
rect 303888 123038 303926 123358
rect 304246 123038 304300 123358
rect 84 121922 336 121942
rect 84 121722 108 121922
rect 308 121722 336 121922
rect 84 121698 336 121722
rect -5128 120948 -5072 121158
rect -5140 120858 -762 120948
rect -5128 119854 -5072 120858
rect 303888 120358 304300 123038
rect 303888 120038 303926 120358
rect 304246 120038 304300 120358
rect 84 118922 336 118942
rect 84 118722 108 118922
rect 308 118722 336 118922
rect 84 118698 336 118722
rect -5186 117858 -802 117948
rect -5186 116774 -5096 117858
rect 303888 117358 304300 120038
rect 303888 117038 303926 117358
rect 304246 117038 304300 117358
rect 84 115922 336 115942
rect 84 115722 108 115922
rect 308 115722 336 115922
rect 84 115698 336 115722
rect -5158 114858 -614 114948
rect -5158 113650 -5068 114858
rect 303888 114358 304300 117038
rect 303888 114038 303926 114358
rect 304246 114038 304300 114358
rect 84 112922 336 112942
rect 84 112722 108 112922
rect 308 112722 336 112922
rect 84 112698 336 112722
rect -5192 111858 -768 111948
rect -5192 110632 -5102 111858
rect 303888 111358 304300 114038
rect 303888 111038 303926 111358
rect 304246 111038 304300 111358
rect 84 109922 336 109942
rect 84 109722 108 109922
rect 308 109722 336 109922
rect 84 109698 336 109722
rect -5124 108858 -802 108948
rect -5124 107622 -5034 108858
rect 303888 108358 304300 111038
rect 303888 108038 303926 108358
rect 304246 108038 304300 108358
rect 84 106922 336 106942
rect 84 106722 108 106922
rect 308 106722 336 106922
rect 84 106698 336 106722
rect -836 104588 -746 105948
rect -5164 104498 -746 104588
rect 303888 105358 304300 108038
rect 303888 105038 303926 105358
rect 304246 105038 304300 105358
rect -5164 104490 -768 104498
rect 84 103922 336 103942
rect 84 103722 108 103922
rect 308 103722 336 103922
rect 84 103698 336 103722
rect -892 101548 -802 102948
rect -5174 101458 -802 101548
rect -892 101258 -802 101458
rect 303888 102358 304300 105038
rect 303888 102038 303926 102358
rect 304246 102038 304300 102358
rect 84 100922 336 100942
rect 84 100722 108 100922
rect 308 100722 336 100922
rect 84 100698 336 100722
rect -892 98428 -802 99948
rect -5208 98338 -802 98428
rect -892 98076 -802 98338
rect 303888 99358 304300 102038
rect 303888 99038 303926 99358
rect 304246 99038 304300 99358
rect 84 97922 336 97942
rect 84 97722 108 97922
rect 308 97722 336 97922
rect 84 97698 336 97722
rect -880 95396 -790 96948
rect -5180 95306 -790 95396
rect -880 95008 -790 95306
rect 303888 96358 304300 99038
rect 303888 96038 303926 96358
rect 304246 96038 304300 96358
rect 84 94922 336 94942
rect 84 94722 108 94922
rect 308 94722 336 94922
rect 84 94698 336 94722
rect -870 92316 -780 93948
rect -5232 92226 -780 92316
rect -870 91912 -780 92226
rect 303888 93358 304300 96038
rect 303888 93038 303926 93358
rect 304246 93038 304300 93358
rect 84 91922 336 91942
rect 84 91722 108 91922
rect 308 91722 336 91922
rect 84 91698 336 91722
rect -852 89208 -762 90948
rect -5192 89118 -762 89208
rect -852 89016 -762 89118
rect 303888 90358 304300 93038
rect 303888 90038 303926 90358
rect 304246 90038 304300 90358
rect 84 88922 336 88942
rect 84 88722 108 88922
rect 308 88722 336 88922
rect 84 88698 336 88722
rect -836 86198 -746 87948
rect -5128 86108 -746 86198
rect -836 85976 -746 86108
rect 303888 87358 304300 90038
rect 303888 87038 303926 87358
rect 304246 87038 304300 87358
rect 84 85922 336 85942
rect 84 85722 108 85922
rect 308 85722 336 85922
rect 84 85698 336 85722
rect -796 83152 -706 84948
rect -5220 83062 -706 83152
rect -796 82720 -706 83062
rect 303888 84358 304300 87038
rect 303888 84038 303926 84358
rect 304246 84038 304300 84358
rect 84 82922 336 82942
rect 84 82722 108 82922
rect 308 82722 336 82922
rect 84 82698 336 82722
rect -880 80022 -790 81948
rect -5202 79932 -790 80022
rect 303888 81358 304300 84038
rect 303888 81038 303926 81358
rect 304246 81038 304300 81358
rect -880 79526 -790 79932
rect 84 79922 336 79942
rect 84 79722 108 79922
rect 308 79722 336 79922
rect 84 79698 336 79722
rect -858 76948 -768 78948
rect -5208 76858 -768 76948
rect 303888 78358 304300 81038
rect 303888 78038 303926 78358
rect 304246 78038 304300 78358
rect -858 76390 -768 76858
rect 84 76922 336 76942
rect 84 76722 108 76922
rect 308 76722 336 76922
rect 84 76698 336 76722
rect -5164 73772 -5074 74058
rect -790 73772 -700 75948
rect 303888 75358 304300 78038
rect 303888 75038 303926 75358
rect 304246 75038 304300 75358
rect -5164 73682 -700 73772
rect 84 73922 336 73942
rect 84 73722 108 73922
rect 308 73722 336 73922
rect 84 73698 336 73722
rect -790 73476 -700 73682
rect -830 70796 -740 72948
rect 303888 72358 304300 75038
rect 303888 72038 303926 72358
rect 304246 72038 304300 72358
rect -5152 70706 -740 70796
rect -830 70580 -740 70706
rect 84 70922 336 70942
rect 84 70722 108 70922
rect 308 70722 336 70922
rect 84 70698 336 70722
rect -5168 67654 -5078 67774
rect -892 67654 -802 69948
rect 303888 69358 304300 72038
rect 303888 69038 303926 69358
rect 304246 69038 304300 69358
rect 84 67922 336 67942
rect 84 67722 108 67922
rect 308 67722 336 67922
rect 84 67698 336 67722
rect -5168 67564 -802 67654
rect -892 67370 -802 67564
rect -608 64618 -552 66924
rect 303888 66358 304300 69038
rect 303888 66038 303926 66358
rect 304246 66038 304300 66358
rect 84 64922 336 64942
rect 84 64722 108 64922
rect 308 64722 336 64922
rect 84 64698 336 64722
rect -5226 64562 -552 64618
rect -5208 63858 -642 63948
rect -5208 61354 -5118 63858
rect 303888 63358 304300 66038
rect 303888 63038 303926 63358
rect 304246 63038 304300 63358
rect 84 61922 336 61942
rect 84 61722 108 61922
rect 308 61722 336 61922
rect 84 61698 336 61722
rect -5242 60858 -700 60948
rect -5242 58378 -5152 60858
rect 303888 60358 304300 63038
rect 303888 60038 303926 60358
rect 304246 60038 304300 60358
rect 84 58922 336 58942
rect 84 58722 108 58922
rect 308 58722 336 58922
rect 84 58698 336 58722
rect -5214 57858 -774 57948
rect -5214 55224 -5124 57858
rect 303888 57358 304300 60038
rect 303888 57038 303926 57358
rect 304246 57038 304300 57358
rect 84 55922 336 55942
rect 84 55722 108 55922
rect 308 55722 336 55922
rect 84 55698 336 55722
rect -5242 54858 -774 54948
rect -5242 52316 -5152 54858
rect 303888 54358 304300 57038
rect 303888 54038 303926 54358
rect 304246 54038 304300 54358
rect 84 52922 336 52942
rect 84 52722 108 52922
rect 308 52722 336 52922
rect 84 52698 336 52722
rect -322 49346 -266 52178
rect 303888 51358 304300 54038
rect 303888 51038 303926 51358
rect 304246 51038 304300 51358
rect 84 49922 336 49942
rect 84 49722 108 49922
rect 308 49722 336 49922
rect 84 49698 336 49722
rect -5146 49290 -266 49346
rect -5226 48858 -488 48948
rect -5226 45970 -5136 48858
rect 303888 48358 304300 51038
rect 303888 48038 303926 48358
rect 304246 48038 304300 48358
rect 84 46922 336 46942
rect 84 46722 108 46922
rect 308 46722 336 46922
rect 84 46698 336 46722
rect -3540 45858 -802 45948
rect -3540 43182 -3450 45858
rect 303888 45358 304300 48038
rect 303888 45038 303926 45358
rect 304246 45038 304300 45358
rect 84 43922 336 43942
rect 84 43722 108 43922
rect 308 43722 336 43922
rect 84 43698 336 43722
rect -5188 43126 -3342 43182
rect -3540 42490 -3450 43126
rect -2360 42948 -2304 43190
rect -2458 42858 -802 42948
rect -2360 40054 -2304 42858
rect 303888 42358 304300 45038
rect 303888 42038 303926 42358
rect 304246 42038 304300 42358
rect 84 40922 336 40942
rect 84 40722 108 40922
rect 308 40722 336 40922
rect 84 40698 336 40722
rect -5256 39998 -2304 40054
rect -750 38442 -660 39948
rect 303888 39358 304300 42038
rect 303888 39038 303926 39358
rect 304246 39038 304300 39358
rect -1990 38386 -496 38442
rect -1990 37018 -1934 38386
rect -750 38280 -660 38386
rect 84 37922 336 37942
rect 84 37722 108 37922
rect 308 37722 336 37922
rect 84 37698 336 37722
rect -5130 36962 -1934 37018
rect -462 35564 -372 36948
rect -2434 35508 -372 35564
rect -2434 33982 -2378 35508
rect -462 35254 -372 35508
rect 303888 36358 304300 39038
rect 303888 36038 303926 36358
rect 304246 36038 304300 36358
rect 84 34922 336 34942
rect 84 34722 108 34922
rect 308 34722 336 34922
rect 84 34698 336 34722
rect -5144 33926 -2378 33982
rect -772 32850 -716 34558
rect -3298 32794 -716 32850
rect 303888 33358 304300 36038
rect 303888 33038 303926 33358
rect 304246 33038 304300 33358
rect -3298 30854 -3242 32794
rect 84 31938 336 31942
rect 72 31922 352 31938
rect 72 31722 108 31922
rect 308 31722 352 31922
rect 72 31684 352 31722
rect -5174 30798 -3242 30854
rect -720 29740 -630 30948
rect 303888 30358 304300 33038
rect 303888 30038 303926 30358
rect 304246 30038 304300 30358
rect -2904 29684 -584 29740
rect -2904 27818 -2848 29684
rect -720 29384 -584 29684
rect -720 29260 -630 29384
rect 82 28922 354 28944
rect 82 28722 108 28922
rect 308 28722 354 28922
rect 82 28692 354 28722
rect -5174 27762 -2848 27818
rect -756 26900 -666 27948
rect 303888 27358 304300 30038
rect 303888 27038 303926 27358
rect 304246 27038 304300 27358
rect -2592 26844 -628 26900
rect -2592 24782 -2536 26844
rect -756 26590 -666 26844
rect 70 25942 330 25946
rect 70 25922 336 25942
rect 70 25722 108 25922
rect 308 25722 336 25922
rect 70 25698 336 25722
rect 70 25684 330 25698
rect -5188 24726 -2536 24782
rect -764 23910 -674 24948
rect 303888 24358 304300 27038
rect 303888 24038 303926 24358
rect 304246 24038 304300 24358
rect -5244 23854 -458 23910
rect -5244 21598 -5188 23854
rect -764 23518 -674 23854
rect 84 22932 336 22942
rect 84 22922 338 22932
rect 84 22722 108 22922
rect 308 22722 338 22922
rect 84 22704 338 22722
rect 84 22698 336 22704
rect -4016 21858 -736 21948
rect -4016 18618 -3926 21858
rect 303888 21372 304300 24038
rect 303888 21358 304304 21372
rect 303888 21038 303926 21358
rect 304246 21038 304304 21358
rect 303888 21004 304304 21038
rect 303888 20952 304300 21004
rect 302848 19472 303028 19478
rect 302848 19292 307364 19472
rect 302848 19278 303028 19292
rect 38312 19214 38562 19226
rect 19850 19188 20100 19202
rect 19850 18978 19874 19188
rect 20084 18978 20100 19188
rect 29066 19062 29328 19096
rect 13790 18930 14040 18950
rect 19850 18944 20100 18978
rect 25908 19006 26226 19028
rect 13650 18924 14040 18930
rect 7470 18886 7720 18910
rect 5316 18784 5566 18810
rect 4518 18780 5566 18784
rect -5180 18510 -3804 18618
rect 4518 18570 5332 18780
rect 5542 18570 5566 18780
rect 7470 18676 7486 18886
rect 7696 18676 7720 18886
rect 7470 18652 7720 18676
rect 10692 18830 10942 18858
rect 4518 18564 5566 18570
rect -5180 18496 -3926 18510
rect 2316 18440 2566 18466
rect 1498 18434 2566 18440
rect 1498 18224 2332 18434
rect 2542 18224 2566 18434
rect 1498 18220 2566 18224
rect -6210 17946 -5984 17960
rect -6210 17746 -6198 17946
rect -5998 17746 -5984 17946
rect -6210 17734 -5984 17746
rect 1498 16556 1718 18220
rect 2316 18208 2566 18220
rect 4518 16430 4738 18564
rect 5316 18552 5566 18564
rect 7482 16456 7702 18652
rect 10692 18620 10716 18830
rect 10926 18620 10942 18830
rect 10692 18600 10942 18620
rect 13650 18714 13806 18924
rect 14016 18714 14040 18924
rect 13650 18692 14040 18714
rect 16900 18812 17150 18824
rect 10710 16526 10930 18600
rect 13650 16450 13870 18692
rect 16900 18602 16916 18812
rect 17126 18602 17150 18812
rect 16900 18566 17150 18602
rect 16910 16694 17130 18566
rect 16746 16474 17130 16694
rect 19868 16482 20088 18944
rect 25908 18796 25948 19006
rect 26158 18796 26226 19006
rect 29066 18842 29084 19062
rect 29304 18842 29328 19062
rect 35298 19050 35584 19066
rect 32330 18986 32556 18990
rect 29066 18824 29328 18842
rect 32124 18982 32556 18986
rect 25908 18762 26226 18796
rect 22880 18672 23142 18674
rect 22872 18654 23188 18672
rect 22872 18444 22902 18654
rect 23112 18444 23188 18654
rect 22872 18406 23188 18444
rect 22896 16456 23116 18406
rect 25942 16450 26162 18762
rect 29084 16482 29304 18824
rect 32124 18772 32332 18982
rect 32542 18772 32556 18982
rect 35298 18840 35332 19050
rect 35542 18840 35584 19050
rect 38312 19004 38332 19214
rect 38542 19004 38562 19214
rect 56594 19158 56844 19178
rect 38312 18968 38562 19004
rect 47292 19126 47590 19154
rect 35298 18828 35584 18840
rect 32124 18754 32556 18772
rect 32124 16526 32344 18754
rect 35328 17248 35548 18828
rect 35196 17028 35548 17248
rect 35196 16482 35416 17028
rect 38328 16512 38548 18968
rect 44320 18918 44570 18936
rect 41318 18868 41568 18892
rect 41318 18658 41332 18868
rect 41542 18658 41568 18868
rect 44320 18708 44332 18918
rect 44542 18708 44570 18918
rect 47292 18916 47332 19126
rect 47542 18916 47590 19126
rect 53520 19038 53770 19064
rect 47292 18900 47590 18916
rect 50500 19006 50750 19022
rect 47318 18886 47568 18900
rect 44320 18678 44570 18708
rect 41318 18634 41568 18658
rect 41328 16456 41548 18634
rect 44328 16424 44548 18678
rect 47328 17632 47548 18886
rect 50500 18796 50520 19006
rect 50730 18796 50750 19006
rect 53520 18828 53542 19038
rect 53752 18828 53770 19038
rect 56594 18948 56620 19158
rect 56830 18948 56844 19158
rect 174332 19130 174626 19162
rect 75052 19026 75346 19044
rect 56594 18920 56844 18948
rect 68518 18952 68808 18988
rect 68518 18948 69258 18952
rect 53520 18806 53770 18828
rect 50500 18764 50750 18796
rect 47328 17412 47734 17632
rect 47514 16506 47734 17412
rect 50516 16474 50736 18764
rect 53536 17810 53756 18806
rect 53536 17590 53888 17810
rect 53668 16506 53888 17590
rect 56614 16444 56834 18920
rect 59608 18866 59858 18886
rect 65736 18876 66010 18892
rect 59608 18862 60000 18866
rect 59608 18652 59634 18862
rect 59844 18652 60000 18862
rect 59608 18628 60000 18652
rect 59780 16494 60000 18628
rect 62572 18790 62974 18834
rect 62572 18786 62996 18790
rect 62572 18576 62636 18786
rect 62846 18576 62996 18786
rect 65736 18666 65746 18876
rect 65956 18666 66010 18876
rect 68518 18738 68554 18948
rect 68764 18738 69258 18948
rect 75052 18816 75082 19026
rect 75292 18816 75346 19026
rect 108892 19028 109134 19040
rect 96442 18870 96684 18884
rect 75052 18782 75346 18816
rect 90400 18832 90652 18856
rect 68518 18732 69258 18738
rect 68518 18722 68808 18732
rect 65736 18610 66010 18666
rect 62572 18542 62996 18576
rect 62776 16468 62996 18542
rect 65946 16498 66002 18610
rect 69038 16506 69258 18732
rect 71910 18520 72162 18536
rect 71910 18310 71932 18520
rect 72142 18310 72162 18520
rect 71910 18292 72162 18310
rect 71928 17006 72148 18292
rect 71928 16786 72278 17006
rect 72058 16506 72278 16786
rect 75078 16416 75298 18782
rect 81172 18706 81430 18720
rect 81172 18496 81194 18706
rect 81404 18496 81430 18706
rect 90400 18622 90416 18832
rect 90626 18622 90652 18832
rect 90400 18608 90652 18622
rect 93536 18788 93788 18810
rect 81172 18482 81430 18496
rect 78074 18076 78350 18088
rect 78074 17866 78102 18076
rect 78312 17866 78350 18076
rect 78074 17848 78350 17866
rect 78098 17154 78318 17848
rect 78098 16934 78452 17154
rect 78232 16492 78452 16934
rect 81190 16478 81410 18482
rect 87330 18310 87580 18326
rect 87330 18100 87340 18310
rect 87550 18100 87580 18310
rect 87330 18086 87580 18100
rect 84246 17980 84526 18028
rect 84246 17770 84278 17980
rect 84488 17770 84526 17980
rect 84246 17732 84526 17770
rect 84274 16492 84494 17732
rect 87334 16380 87554 18086
rect 90412 16440 90632 18608
rect 93536 18578 93560 18788
rect 93770 18578 93788 18788
rect 96442 18660 96458 18870
rect 96668 18660 96684 18870
rect 108892 18818 108906 19028
rect 109116 18818 109134 19028
rect 114930 18980 115200 19008
rect 108892 18808 109134 18818
rect 111936 18930 112184 18948
rect 96442 18650 96684 18660
rect 102658 18736 102952 18774
rect 93536 18562 93788 18578
rect 93556 16448 93776 18562
rect 96452 17026 96672 18650
rect 102658 18526 102716 18736
rect 102926 18526 102952 18736
rect 99582 18496 99842 18518
rect 99582 18286 99602 18496
rect 99812 18286 99842 18496
rect 102658 18468 102952 18526
rect 105620 18750 105914 18790
rect 105620 18540 105680 18750
rect 105890 18540 105914 18750
rect 105620 18484 105914 18540
rect 99582 18248 99842 18286
rect 96452 16806 96814 17026
rect 96594 16478 96814 16806
rect 99596 16514 99816 18248
rect 102710 16410 102930 18468
rect 105674 16996 105894 18484
rect 105674 16776 106014 16996
rect 105794 16462 106014 16776
rect 108900 16454 109120 18808
rect 111936 18720 111952 18930
rect 112162 18720 112184 18930
rect 114930 18770 114958 18980
rect 115168 18770 115200 18980
rect 114930 18744 115200 18770
rect 117942 18972 118250 18998
rect 117942 18762 117972 18972
rect 118182 18762 118250 18972
rect 157794 18992 158088 19008
rect 127190 18938 127500 18970
rect 111936 18712 112184 18720
rect 111948 16514 112168 18712
rect 114952 16452 115172 18744
rect 117942 18686 118250 18762
rect 121128 18860 121382 18878
rect 117968 17904 118188 18686
rect 121128 18650 121154 18860
rect 121364 18650 121382 18860
rect 121128 18614 121382 18650
rect 124096 18852 124354 18864
rect 124096 18632 124118 18852
rect 124338 18632 124354 18852
rect 127190 18728 127246 18938
rect 127456 18728 127500 18938
rect 133376 18866 133686 18894
rect 127190 18678 127500 18728
rect 130210 18808 130520 18858
rect 124096 18624 124354 18632
rect 117968 17684 118368 17904
rect 118148 16482 118368 17684
rect 121150 16460 121370 18614
rect 124118 16552 124338 18624
rect 127240 16460 127460 18678
rect 130210 18598 130254 18808
rect 130464 18598 130520 18808
rect 133376 18646 133412 18866
rect 133632 18646 133686 18866
rect 145538 18838 145832 18860
rect 133376 18602 133686 18646
rect 142542 18664 142852 18692
rect 130210 18566 130520 18598
rect 130250 16476 130470 18566
rect 133412 16460 133632 18602
rect 139492 18596 139802 18606
rect 139492 18386 139556 18596
rect 139766 18386 139802 18596
rect 142542 18454 142604 18664
rect 142814 18454 142852 18664
rect 145538 18628 145582 18838
rect 145792 18628 145832 18838
rect 145538 18580 145832 18628
rect 148714 18838 149008 18874
rect 148714 18628 148758 18838
rect 148968 18628 149008 18838
rect 154754 18854 155048 18876
rect 148714 18594 149008 18628
rect 151732 18770 152026 18802
rect 142542 18400 142852 18454
rect 139492 18314 139802 18386
rect 136442 18236 136752 18286
rect 136442 18026 136472 18236
rect 136682 18026 136752 18236
rect 136442 17994 136752 18026
rect 136466 16400 136686 17994
rect 139552 16484 139772 18314
rect 142598 16468 142818 18400
rect 145578 16946 145798 18580
rect 145578 16726 145918 16946
rect 145698 16452 145918 16726
rect 148754 16406 148974 18594
rect 151732 18560 151776 18770
rect 151986 18560 152026 18770
rect 154754 18644 154796 18854
rect 155006 18644 155048 18854
rect 157794 18782 157848 18992
rect 158058 18782 158088 18992
rect 174332 18920 174370 19130
rect 174580 18920 174626 19130
rect 305362 19094 305616 19106
rect 290286 18956 290586 18982
rect 174332 18882 174626 18920
rect 229636 18934 229916 18952
rect 157794 18728 158088 18782
rect 160862 18754 161156 18778
rect 154754 18596 155048 18644
rect 151732 18522 152026 18560
rect 151772 16372 151992 18522
rect 154792 17614 155012 18596
rect 154792 17394 155166 17614
rect 154946 16464 155166 17394
rect 157842 17038 158062 18728
rect 160862 18544 160890 18754
rect 161100 18544 161156 18754
rect 160862 18498 161156 18544
rect 173066 18508 173336 18534
rect 160886 17192 161106 18498
rect 163202 18460 163496 18486
rect 173060 18484 173354 18508
rect 163202 18454 164318 18460
rect 163202 18244 163242 18454
rect 163452 18244 164318 18454
rect 163202 18240 164318 18244
rect 163202 18206 163496 18240
rect 164098 17688 164318 18240
rect 173060 18274 173086 18484
rect 173296 18274 173354 18484
rect 173060 18228 173354 18274
rect 165896 18174 166190 18202
rect 165896 18170 167322 18174
rect 165896 17960 165932 18170
rect 166142 17960 167322 18170
rect 165896 17954 167322 17960
rect 165896 17922 166190 17954
rect 164052 17332 164318 17688
rect 157842 16818 158224 17038
rect 160886 16972 161244 17192
rect 158004 16494 158224 16818
rect 161024 16540 161244 16972
rect 164052 16440 164272 17332
rect 167102 16440 167322 17954
rect 173082 17606 173302 18228
rect 168824 17422 169118 17446
rect 168824 17416 170482 17422
rect 168824 17206 168868 17416
rect 169078 17206 170482 17416
rect 173082 17386 173510 17606
rect 168824 17202 170482 17206
rect 168824 17166 169118 17202
rect 170262 16502 170482 17202
rect 173290 16464 173510 17386
rect 174366 17560 174586 18882
rect 176292 18812 176586 18846
rect 176292 18808 179212 18812
rect 176292 18598 176332 18808
rect 176542 18598 179212 18808
rect 229636 18724 229662 18934
rect 229872 18724 229916 18934
rect 290286 18950 293618 18956
rect 290286 18740 290332 18950
rect 290542 18740 293618 18950
rect 305362 18884 305390 19094
rect 305600 18884 305616 19094
rect 305362 18850 305616 18884
rect 290286 18736 293618 18740
rect 229636 18700 229916 18724
rect 176292 18592 179212 18598
rect 176292 18566 176586 18592
rect 174366 17340 176668 17560
rect 176448 16456 176668 17340
rect 178992 17290 179212 18592
rect 215300 18564 215570 18576
rect 215300 18558 219616 18564
rect 206300 18456 206560 18470
rect 206300 18450 208700 18456
rect 206300 18240 206332 18450
rect 206542 18240 208700 18450
rect 215300 18348 215332 18558
rect 215542 18348 219616 18558
rect 215300 18344 219616 18348
rect 215300 18338 215570 18344
rect 206300 18236 208700 18240
rect 206300 18216 206560 18236
rect 185290 18036 185584 18060
rect 185290 18032 188126 18036
rect 182444 17854 182738 17894
rect 182444 17644 182478 17854
rect 182688 17644 182738 17854
rect 185290 17822 185332 18032
rect 185542 17822 188126 18032
rect 185290 17816 188126 17822
rect 185290 17780 185584 17816
rect 182444 17614 182738 17644
rect 178992 17070 179704 17290
rect 179484 16494 179704 17070
rect 182472 16480 182692 17614
rect 183972 17152 184266 17190
rect 183972 17148 185874 17152
rect 183972 16938 184014 17148
rect 184224 16938 185874 17148
rect 183972 16932 185874 16938
rect 183972 16910 184266 16932
rect 185654 16456 185874 16932
rect 187906 16884 188126 17816
rect 196770 17924 197064 17956
rect 196770 17714 196798 17924
rect 197008 17714 197064 17924
rect 188280 17660 188574 17686
rect 196770 17676 197064 17714
rect 200892 17952 201204 18006
rect 200892 17742 200920 17952
rect 201130 17742 201204 17952
rect 200892 17700 201204 17742
rect 206974 17746 207242 17790
rect 188280 17654 191876 17660
rect 188280 17444 188332 17654
rect 188542 17444 191876 17654
rect 188280 17440 191876 17444
rect 188280 17406 188574 17440
rect 187906 16664 188840 16884
rect 188620 16448 188840 16664
rect 191656 16486 191876 17440
rect 193426 17020 193720 17048
rect 196792 17020 197012 17676
rect 193426 17014 195050 17020
rect 193426 16804 193470 17014
rect 193680 16804 195050 17014
rect 193426 16800 195050 16804
rect 196792 16800 198136 17020
rect 193426 16768 193720 16800
rect 194830 16452 195050 16800
rect 197916 16380 198136 16800
rect 200914 16470 201134 17700
rect 206974 17536 207004 17746
rect 207214 17536 207242 17746
rect 206974 17516 207242 17536
rect 201984 16894 202244 16902
rect 201984 16890 204256 16894
rect 201984 16680 202008 16890
rect 202218 16680 204256 16890
rect 201984 16674 204256 16680
rect 201984 16656 202244 16674
rect 204036 16514 204256 16674
rect 206998 16522 207218 17516
rect 208480 17090 208700 18236
rect 213128 18094 213386 18108
rect 213128 17884 213160 18094
rect 213370 17884 213386 18094
rect 213128 17848 213386 17884
rect 208480 16870 210430 17090
rect 210210 16506 210430 16870
rect 213154 16434 213374 17848
rect 213898 17276 214144 17278
rect 213876 17270 214144 17276
rect 213876 17264 216496 17270
rect 213876 17054 213908 17264
rect 214118 17054 216496 17264
rect 213876 17050 216496 17054
rect 213876 17032 214144 17050
rect 213876 17030 214122 17032
rect 216276 16372 216496 17050
rect 219396 16434 219616 18344
rect 227174 18424 227460 18436
rect 227174 18214 227198 18424
rect 227408 18214 227460 18424
rect 227174 18192 227460 18214
rect 221292 17712 221614 17730
rect 221292 17706 225720 17712
rect 221292 17496 221332 17706
rect 221542 17496 225720 17706
rect 221292 17492 225720 17496
rect 221292 17460 221614 17492
rect 220666 17228 220962 17238
rect 220666 17224 222682 17228
rect 220666 17014 220692 17224
rect 220902 17014 222682 17224
rect 220666 17008 222682 17014
rect 220666 17000 220962 17008
rect 222462 16426 222682 17008
rect 225500 16498 225720 17492
rect 227194 17524 227414 18192
rect 227194 17304 228838 17524
rect 228618 16480 228838 17304
rect 229658 17434 229878 18700
rect 233310 18690 233574 18702
rect 254314 18700 254612 18736
rect 254314 18696 257536 18700
rect 233310 18684 237602 18690
rect 233310 18474 233332 18684
rect 233542 18680 237602 18684
rect 233542 18474 237948 18680
rect 242314 18570 242552 18578
rect 242314 18566 245088 18570
rect 233310 18470 237948 18474
rect 233310 18442 233574 18470
rect 237356 18460 237948 18470
rect 234638 18304 234884 18322
rect 234638 18298 235040 18304
rect 234638 18088 234654 18298
rect 234864 18088 235040 18298
rect 234638 18062 235040 18088
rect 229658 17214 231876 17434
rect 231656 16542 231876 17214
rect 234820 16506 235040 18062
rect 237728 17960 237948 18460
rect 241664 18530 241902 18544
rect 241664 18320 241676 18530
rect 241886 18320 241902 18530
rect 242314 18356 242332 18566
rect 242542 18356 245088 18566
rect 242314 18350 245088 18356
rect 242314 18346 242552 18350
rect 241664 18312 241902 18320
rect 237706 17778 237948 17960
rect 240890 18010 241174 18054
rect 240890 17800 240920 18010
rect 241130 17800 241174 18010
rect 237706 16426 237926 17778
rect 240890 17770 241174 17800
rect 240916 16484 241136 17770
rect 241672 17214 241892 18312
rect 241672 16994 244150 17214
rect 243930 16320 244150 16994
rect 244868 16986 245088 18350
rect 253898 18504 254148 18520
rect 253898 18294 253930 18504
rect 254140 18294 254148 18504
rect 254314 18486 254332 18696
rect 254542 18486 257536 18696
rect 279642 18694 279942 18730
rect 290286 18696 290586 18736
rect 254314 18480 257536 18486
rect 254314 18462 254612 18480
rect 253898 18276 254148 18294
rect 249644 17860 249924 17882
rect 249644 17856 253346 17860
rect 249644 17646 249672 17856
rect 249882 17646 253346 17856
rect 249644 17640 253346 17646
rect 249644 17622 249924 17640
rect 248702 17078 248952 17090
rect 248702 17072 250268 17078
rect 244868 16766 247272 16986
rect 248702 16862 248716 17072
rect 248926 16862 250268 17072
rect 248702 16858 250268 16862
rect 248702 16846 248952 16858
rect 247052 16520 247272 16766
rect 250048 16420 250268 16858
rect 253126 16520 253346 17640
rect 253924 17354 254144 18276
rect 257316 17358 257536 18480
rect 269016 18556 269288 18572
rect 269016 18346 269036 18556
rect 269246 18346 269288 18556
rect 279642 18484 279680 18694
rect 279890 18484 279942 18694
rect 279642 18444 279942 18484
rect 269016 18314 269288 18346
rect 261022 18126 261294 18136
rect 261022 18120 265648 18126
rect 261022 17910 261048 18120
rect 261258 17910 265648 18120
rect 261022 17906 265648 17910
rect 261022 17878 261294 17906
rect 259366 17358 259586 17386
rect 253924 17134 256416 17354
rect 257316 17138 259608 17358
rect 260030 17246 260302 17258
rect 260030 17242 262606 17246
rect 256196 16438 256416 17134
rect 259366 16506 259586 17138
rect 260030 17032 260058 17242
rect 260268 17032 262606 17242
rect 260030 17026 262606 17032
rect 260030 17000 260302 17026
rect 262386 16480 262606 17026
rect 265428 16438 265648 17906
rect 265852 17964 266124 17980
rect 265852 17958 267378 17964
rect 265852 17748 265874 17958
rect 266084 17748 267378 17958
rect 265852 17744 267378 17748
rect 265852 17722 266124 17744
rect 267158 17370 267378 17744
rect 267158 17150 268752 17370
rect 267158 17148 267378 17150
rect 268532 16388 268752 17150
rect 269032 17090 269252 18314
rect 269322 18268 269594 18292
rect 269322 18264 274812 18268
rect 269322 18054 269332 18264
rect 269542 18054 274812 18264
rect 269322 18048 274812 18054
rect 269322 18034 269594 18048
rect 269032 16870 271810 17090
rect 271590 16406 271810 16870
rect 274592 16502 274812 18048
rect 278800 18202 279208 18308
rect 278800 17992 278882 18202
rect 279092 17992 279208 18202
rect 278800 17946 279208 17992
rect 277670 17578 277952 17624
rect 277670 17368 277698 17578
rect 277908 17368 277952 17578
rect 277670 17336 277952 17368
rect 277692 16482 277912 17336
rect 278878 17146 279098 17946
rect 279676 17916 279896 18444
rect 292376 18222 292676 18260
rect 284308 18138 284608 18176
rect 284308 18132 287822 18138
rect 284308 17922 284332 18132
rect 284542 17922 287822 18132
rect 292376 18012 292412 18222
rect 292622 18012 292676 18222
rect 292376 17974 292676 18012
rect 284308 17918 287822 17922
rect 279676 17696 284112 17916
rect 284308 17890 284608 17918
rect 278878 16926 280970 17146
rect 280750 16364 280970 16926
rect 283892 16454 284112 17696
rect 286910 17508 287210 17550
rect 286910 17298 286934 17508
rect 287144 17298 287210 17508
rect 286910 17264 287210 17298
rect 286928 16446 287148 17264
rect 287602 16980 287822 17918
rect 287602 16760 290186 16980
rect 289966 16488 290186 16760
rect 292406 16924 292626 17974
rect 293398 17354 293618 18736
rect 302946 18469 303268 18478
rect 302940 17936 302946 18258
rect 303268 17936 303274 18258
rect 299228 17718 299528 17758
rect 299228 17508 299262 17718
rect 299472 17508 299528 17718
rect 299228 17472 299528 17508
rect 293398 17134 296406 17354
rect 292406 16704 293306 16924
rect 293086 16446 293306 16704
rect 296186 16460 296406 17134
rect 299258 16890 299478 17472
rect 299146 16670 299478 16890
rect 300208 17106 300508 17140
rect 300208 17100 302500 17106
rect 300208 16890 300256 17100
rect 300466 16890 302500 17100
rect 300208 16886 302500 16890
rect 300208 16854 300508 16886
rect 299146 16398 299366 16670
rect 302280 16510 302500 16886
rect 305384 16504 305604 18850
rect 302888 16416 303316 16448
rect 302888 16094 302946 16416
rect 303268 16094 303316 16416
rect 302888 16036 303316 16094
rect 26 15588 390 15664
rect 26 15388 108 15588
rect 308 15388 390 15588
rect 26 15298 390 15388
<< via2 >>
rect 302508 324332 302708 324532
rect 303930 321042 304240 321352
rect 108 319722 308 319922
rect 303930 318042 304240 318352
rect 108 316722 308 316922
rect 303930 315042 304240 315352
rect 108 313722 308 313922
rect 303930 312042 304240 312352
rect 108 310722 308 310922
rect 303930 309042 304240 309352
rect 108 307722 308 307922
rect 303930 306042 304240 306352
rect 108 304722 308 304922
rect 303930 303042 304240 303352
rect 108 301722 308 301922
rect 303930 300042 304240 300352
rect 108 298722 308 298922
rect 303930 297042 304240 297352
rect 108 295722 308 295922
rect 303930 294042 304240 294352
rect 108 292722 308 292922
rect 303930 291042 304240 291352
rect 108 289722 308 289922
rect 303930 288042 304240 288352
rect 108 286722 308 286922
rect 303930 285042 304240 285352
rect 108 283722 308 283922
rect 303930 282042 304240 282352
rect 108 280722 308 280922
rect 303930 279042 304240 279352
rect 108 277722 308 277922
rect 303930 276042 304240 276352
rect 108 274722 308 274922
rect 303930 273042 304240 273352
rect 108 271722 308 271922
rect 303930 270042 304240 270352
rect 108 268722 308 268922
rect 303930 267042 304240 267352
rect 108 265722 308 265922
rect 303930 264042 304240 264352
rect 108 262722 308 262922
rect 303930 261042 304240 261352
rect 108 259722 308 259922
rect 303930 258042 304240 258352
rect 108 256722 308 256922
rect 303930 255042 304240 255352
rect 108 253722 308 253922
rect 303930 252042 304240 252352
rect 108 250722 308 250922
rect 303930 249042 304240 249352
rect 108 247722 308 247922
rect 303930 246042 304240 246352
rect 108 244722 308 244922
rect 303930 243042 304240 243352
rect 108 241722 308 241922
rect 303930 240042 304240 240352
rect 108 238722 308 238922
rect 303930 237042 304240 237352
rect 108 235722 308 235922
rect 303930 234042 304240 234352
rect 108 232722 308 232922
rect 303930 231042 304240 231352
rect 108 229722 308 229922
rect 303930 228042 304240 228352
rect 108 226722 308 226922
rect 303930 225042 304240 225352
rect 108 223722 308 223922
rect 303930 222042 304240 222352
rect 108 220722 308 220922
rect 303930 219042 304240 219352
rect 108 217722 308 217922
rect 303930 216042 304240 216352
rect 108 214722 308 214922
rect 303930 213042 304240 213352
rect 108 211722 308 211922
rect 303930 210042 304240 210352
rect 108 208722 308 208922
rect 303930 207042 304240 207352
rect 108 205722 308 205922
rect 303930 204042 304240 204352
rect 108 202722 308 202922
rect 303930 201042 304240 201352
rect 108 199722 308 199922
rect 303930 198042 304240 198352
rect 108 196722 308 196922
rect 303930 195042 304240 195352
rect 108 193722 308 193922
rect 303930 192042 304240 192352
rect 108 190722 308 190922
rect 303930 189042 304240 189352
rect 108 187722 308 187922
rect 303930 186042 304240 186352
rect 108 184722 308 184922
rect 303930 183042 304240 183352
rect 108 181722 308 181922
rect 303930 180042 304240 180352
rect 108 178722 308 178922
rect 303930 177042 304240 177352
rect 108 175722 308 175922
rect 303930 174042 304240 174352
rect 108 172722 308 172922
rect 303930 171042 304240 171352
rect 108 169722 308 169922
rect 303930 168042 304240 168352
rect 108 166722 308 166922
rect 303930 165042 304240 165352
rect 108 163722 308 163922
rect 303930 162042 304240 162352
rect 108 160722 308 160922
rect 303930 159042 304240 159352
rect 108 157722 308 157922
rect 303930 156042 304240 156352
rect 108 154722 308 154922
rect 303930 153042 304240 153352
rect 108 151722 308 151922
rect 303930 150042 304240 150352
rect 108 148722 308 148922
rect 303930 147042 304240 147352
rect 108 145722 308 145922
rect 303930 144042 304240 144352
rect 108 142722 308 142922
rect 303930 141042 304240 141352
rect 108 139722 308 139922
rect 303930 138042 304240 138352
rect 108 136722 308 136922
rect 303930 135042 304240 135352
rect 108 133722 308 133922
rect 303930 132042 304240 132352
rect 108 130722 308 130922
rect 303930 129042 304240 129352
rect 108 127722 308 127922
rect 303930 126042 304240 126352
rect 108 124722 308 124922
rect 303930 123042 304240 123352
rect 108 121722 308 121922
rect 303930 120042 304240 120352
rect 108 118722 308 118922
rect 303930 117042 304240 117352
rect 108 115722 308 115922
rect 303930 114042 304240 114352
rect 108 112722 308 112922
rect 303930 111042 304240 111352
rect 108 109722 308 109922
rect 303930 108042 304240 108352
rect 108 106722 308 106922
rect 303930 105042 304240 105352
rect 108 103722 308 103922
rect 303930 102042 304240 102352
rect 108 100722 308 100922
rect 303930 99042 304240 99352
rect 108 97722 308 97922
rect 303930 96042 304240 96352
rect 108 94722 308 94922
rect 303930 93042 304240 93352
rect 108 91722 308 91922
rect 303930 90042 304240 90352
rect 108 88722 308 88922
rect 303930 87042 304240 87352
rect 108 85722 308 85922
rect 303930 84042 304240 84352
rect 108 82722 308 82922
rect 303930 81042 304240 81352
rect 108 79722 308 79922
rect 303930 78042 304240 78352
rect 108 76722 308 76922
rect 303930 75042 304240 75352
rect 108 73722 308 73922
rect 303930 72042 304240 72352
rect 108 70722 308 70922
rect 303930 69042 304240 69352
rect 108 67722 308 67922
rect 303930 66042 304240 66352
rect 108 64722 308 64922
rect 303930 63042 304240 63352
rect 108 61722 308 61922
rect 303930 60042 304240 60352
rect 108 58722 308 58922
rect 303930 57042 304240 57352
rect 108 55722 308 55922
rect 303930 54042 304240 54352
rect 108 52722 308 52922
rect 303930 51042 304240 51352
rect 108 49722 308 49922
rect 303930 48042 304240 48352
rect 108 46722 308 46922
rect 303930 45042 304240 45352
rect 108 43722 308 43922
rect 303930 42042 304240 42352
rect 108 40722 308 40922
rect 303930 39042 304240 39352
rect 108 37722 308 37922
rect 303930 36042 304240 36352
rect 108 34722 308 34922
rect 303930 33042 304240 33352
rect 108 31722 308 31922
rect 303930 30042 304240 30352
rect 108 28722 308 28922
rect 303930 27042 304240 27352
rect 108 25722 308 25922
rect 303930 24042 304240 24352
rect 108 22722 308 22922
rect 303930 21042 304240 21352
rect 19874 18978 20084 19188
rect 5332 18570 5542 18780
rect 7486 18676 7696 18886
rect 2332 18224 2542 18434
rect -6198 17746 -5998 17946
rect 10716 18620 10926 18830
rect 13806 18714 14016 18924
rect 16916 18602 17126 18812
rect 25948 18796 26158 19006
rect 29084 18842 29304 19062
rect 22902 18444 23112 18654
rect 32332 18772 32542 18982
rect 35332 18840 35542 19050
rect 38332 19004 38542 19214
rect 41332 18658 41542 18868
rect 44332 18708 44542 18918
rect 47332 18916 47542 19126
rect 50520 18796 50730 19006
rect 53542 18828 53752 19038
rect 56620 18948 56830 19158
rect 59634 18652 59844 18862
rect 62636 18576 62846 18786
rect 65746 18666 65956 18876
rect 68554 18738 68764 18948
rect 75082 18816 75292 19026
rect 71932 18310 72142 18520
rect 81194 18496 81404 18706
rect 90416 18622 90626 18832
rect 78102 17866 78312 18076
rect 87340 18100 87550 18310
rect 84278 17770 84488 17980
rect 93560 18578 93770 18788
rect 96458 18660 96668 18870
rect 108906 18818 109116 19028
rect 102716 18526 102926 18736
rect 99602 18286 99812 18496
rect 105680 18540 105890 18750
rect 111952 18720 112162 18930
rect 114958 18770 115168 18980
rect 117972 18762 118182 18972
rect 121154 18650 121364 18860
rect 124118 18632 124338 18852
rect 127246 18728 127456 18938
rect 130254 18598 130464 18808
rect 133412 18646 133632 18866
rect 139556 18386 139766 18596
rect 142604 18454 142814 18664
rect 145582 18628 145792 18838
rect 148758 18628 148968 18838
rect 136472 18026 136682 18236
rect 151776 18560 151986 18770
rect 154796 18644 155006 18854
rect 157848 18782 158058 18992
rect 174370 18920 174580 19130
rect 160890 18544 161100 18754
rect 163242 18244 163452 18454
rect 173086 18274 173296 18484
rect 165932 17960 166142 18170
rect 168868 17206 169078 17416
rect 176332 18598 176542 18808
rect 229662 18724 229872 18934
rect 290332 18740 290542 18950
rect 305390 18884 305600 19094
rect 206332 18240 206542 18450
rect 215332 18348 215542 18558
rect 182478 17644 182688 17854
rect 185332 17822 185542 18032
rect 184014 16938 184224 17148
rect 196798 17714 197008 17924
rect 200920 17742 201130 17952
rect 188332 17444 188542 17654
rect 193470 16804 193680 17014
rect 207004 17536 207214 17746
rect 202008 16680 202218 16890
rect 213160 17884 213370 18094
rect 213908 17054 214118 17264
rect 227198 18214 227408 18424
rect 221332 17496 221542 17706
rect 220692 17014 220902 17224
rect 233332 18474 233542 18684
rect 234654 18088 234864 18298
rect 241676 18320 241886 18530
rect 242332 18356 242542 18566
rect 240920 17800 241130 18010
rect 253930 18294 254140 18504
rect 254332 18486 254542 18696
rect 249672 17646 249882 17856
rect 248716 16862 248926 17072
rect 269036 18346 269246 18556
rect 279680 18484 279890 18694
rect 261048 17910 261258 18120
rect 260058 17032 260268 17242
rect 265874 17748 266084 17958
rect 269332 18054 269542 18264
rect 278882 17992 279092 18202
rect 277698 17368 277908 17578
rect 284332 17922 284542 18132
rect 292412 18012 292622 18222
rect 286934 17298 287144 17508
rect 302946 18258 303268 18469
rect 302946 18147 303268 18258
rect 299262 17508 299472 17718
rect 300256 16890 300466 17100
rect 302946 16094 303268 16416
rect 108 15388 308 15588
<< metal3 >>
rect -13040 323508 -12920 323868
rect 908 322280 998 327366
rect 302440 324538 302792 324614
rect 302440 324338 302502 324538
rect 302712 324338 302792 324538
rect 302440 324332 302508 324338
rect 302708 324332 302792 324338
rect 302440 324258 302792 324332
rect 303888 321356 304300 322140
rect 303888 321038 303926 321356
rect 304244 321038 304300 321356
rect -2066 319922 -1726 319998
rect 60 319922 352 319968
rect -2066 319723 -2006 319922
rect -2066 319722 -2005 319723
rect -1806 319722 108 319922
rect 308 319722 400 319922
rect -2066 319684 -1726 319722
rect 60 319702 352 319722
rect 303888 318356 304300 321038
rect 303888 318038 303926 318356
rect 304244 318038 304300 318356
rect -2038 316922 -1776 317004
rect 76 316922 354 316942
rect -2038 316722 -2006 316922
rect -1806 316722 108 316922
rect 308 316722 354 316922
rect -2038 316694 -1776 316722
rect 76 316670 354 316722
rect 303888 315356 304300 318038
rect 303888 315038 303926 315356
rect 304244 315038 304300 315356
rect 82 313922 350 313960
rect -2012 313722 -2006 313922
rect -1806 313722 108 313922
rect 308 313722 350 313922
rect 82 313682 350 313722
rect 303888 312356 304300 315038
rect 303888 312038 303926 312356
rect 304244 312038 304300 312356
rect -2026 310922 -1780 310940
rect 76 310922 334 310934
rect -2026 310722 -2006 310922
rect -1806 310722 108 310922
rect 308 310722 334 310922
rect -2026 310708 -1780 310722
rect 76 310692 334 310722
rect 303888 309356 304300 312038
rect 303888 309038 303926 309356
rect 304244 309038 304300 309356
rect 80 307922 328 307932
rect -2012 307722 -2006 307922
rect -1806 307722 108 307922
rect 308 307722 328 307922
rect 80 307694 328 307722
rect 303888 306356 304300 309038
rect 303888 306038 303926 306356
rect 304244 306038 304300 306356
rect 88 304922 358 304948
rect -2012 304722 -2006 304922
rect -1806 304722 108 304922
rect 308 304722 358 304922
rect 88 304698 358 304722
rect 303888 303356 304300 306038
rect 303888 303038 303926 303356
rect 304244 303038 304300 303356
rect -2018 301922 -1790 301926
rect 98 301922 332 301954
rect -2018 301722 -2006 301922
rect -1806 301722 108 301922
rect 308 301722 332 301922
rect -2018 301712 -1790 301722
rect 98 301688 332 301722
rect 303888 300356 304300 303038
rect 303888 300038 303926 300356
rect 304244 300038 304300 300356
rect 82 298922 322 298930
rect -2012 298722 -2006 298922
rect -1806 298722 108 298922
rect 308 298722 322 298922
rect 82 298698 322 298722
rect 303888 297356 304300 300038
rect 303888 297038 303926 297356
rect 304244 297038 304300 297356
rect 96 295922 318 295934
rect -2012 295722 -2006 295922
rect -1806 295722 108 295922
rect 308 295722 318 295922
rect 96 295702 318 295722
rect 303888 294356 304300 297038
rect 303888 294038 303926 294356
rect 304244 294038 304300 294356
rect 84 292922 336 292942
rect -2012 292722 -2006 292922
rect -1806 292722 108 292922
rect 308 292722 336 292922
rect 84 292698 336 292722
rect 303888 291356 304300 294038
rect 303888 291038 303926 291356
rect 304244 291038 304300 291356
rect 84 289922 336 289942
rect -2012 289722 -2006 289922
rect -1806 289722 108 289922
rect 308 289722 336 289922
rect 84 289698 336 289722
rect 303888 288356 304300 291038
rect 303888 288038 303926 288356
rect 304244 288038 304300 288356
rect 84 286930 336 286942
rect -2016 286922 -1786 286930
rect 82 286922 336 286930
rect -2016 286722 -2006 286922
rect -1806 286722 108 286922
rect 308 286722 336 286922
rect -2016 286708 -1786 286722
rect 82 286698 336 286722
rect 303888 285356 304300 288038
rect 303888 285038 303926 285356
rect 304244 285038 304300 285356
rect 84 283930 336 283942
rect -2016 283922 -1786 283930
rect 82 283922 336 283930
rect -2016 283722 -2006 283922
rect -1806 283722 108 283922
rect 308 283722 336 283922
rect -2016 283708 -1786 283722
rect 82 283698 336 283722
rect 303888 282356 304300 285038
rect 303888 282038 303926 282356
rect 304244 282038 304300 282356
rect 84 280930 336 280942
rect -2016 280922 -1786 280930
rect 82 280922 336 280930
rect -2016 280722 -2006 280922
rect -1806 280722 108 280922
rect 308 280722 336 280922
rect -2016 280708 -1786 280722
rect 82 280698 336 280722
rect 303888 279356 304300 282038
rect 303888 279038 303926 279356
rect 304244 279038 304300 279356
rect -2016 277922 -1786 277930
rect 84 277922 336 277942
rect -2016 277722 -2006 277922
rect -1806 277722 108 277922
rect 308 277722 336 277922
rect -2016 277708 -1786 277722
rect 84 277698 336 277722
rect 303888 276356 304300 279038
rect 303888 276038 303926 276356
rect 304244 276038 304300 276356
rect -2016 274922 -1786 274930
rect 84 274922 336 274942
rect -2016 274722 -2006 274922
rect -1806 274722 108 274922
rect 308 274722 336 274922
rect -2016 274708 -1786 274722
rect 84 274698 336 274722
rect 303888 273356 304300 276038
rect 303888 273038 303926 273356
rect 304244 273038 304300 273356
rect -2016 271922 -1786 271930
rect 84 271922 336 271942
rect -2016 271722 -2006 271922
rect -1806 271722 108 271922
rect 308 271722 336 271922
rect -2016 271708 -1786 271722
rect 84 271698 336 271722
rect 303888 270356 304300 273038
rect 303888 270038 303926 270356
rect 304244 270038 304300 270356
rect -2016 268922 -1786 268930
rect 84 268922 336 268942
rect -2016 268722 -2006 268922
rect -1806 268722 108 268922
rect 308 268722 336 268922
rect -2016 268708 -1786 268722
rect 84 268698 336 268722
rect 303888 267356 304300 270038
rect 303888 267038 303926 267356
rect 304244 267038 304300 267356
rect -2016 265922 -1786 265930
rect 84 265922 336 265942
rect -2016 265722 -2006 265922
rect -1806 265722 108 265922
rect 308 265722 336 265922
rect -2016 265708 -1786 265722
rect 84 265698 336 265722
rect 303888 264356 304300 267038
rect 303888 264038 303926 264356
rect 304244 264038 304300 264356
rect -2016 262922 -1786 262930
rect 84 262922 336 262942
rect -2016 262722 -2006 262922
rect -1806 262722 108 262922
rect 308 262722 336 262922
rect -2016 262708 -1786 262722
rect 84 262698 336 262722
rect 303888 261356 304300 264038
rect 303888 261038 303926 261356
rect 304244 261038 304300 261356
rect -2016 259922 -1786 259930
rect 84 259922 336 259942
rect -2016 259722 -2006 259922
rect -1806 259722 108 259922
rect 308 259722 336 259922
rect -2016 259708 -1786 259722
rect 84 259698 336 259722
rect 303888 258356 304300 261038
rect 303888 258038 303926 258356
rect 304244 258038 304300 258356
rect -2016 256922 -1786 256930
rect 84 256922 336 256942
rect -2016 256722 -2006 256922
rect -1806 256722 108 256922
rect 308 256722 336 256922
rect -2016 256708 -1786 256722
rect 84 256698 336 256722
rect 303888 255356 304300 258038
rect 303888 255038 303926 255356
rect 304244 255038 304300 255356
rect -2016 253922 -1786 253930
rect 84 253922 336 253942
rect -2016 253722 -2006 253922
rect -1806 253722 108 253922
rect 308 253722 336 253922
rect -2016 253708 -1786 253722
rect 84 253698 336 253722
rect 303888 252356 304300 255038
rect 303888 252038 303926 252356
rect 304244 252038 304300 252356
rect -2016 250922 -1786 250930
rect 84 250922 336 250942
rect -2016 250722 -2006 250922
rect -1806 250722 108 250922
rect 308 250722 336 250922
rect -2016 250708 -1786 250722
rect 84 250698 336 250722
rect 303888 249356 304300 252038
rect 303888 249038 303926 249356
rect 304244 249038 304300 249356
rect -2016 247922 -1786 247930
rect 84 247922 336 247942
rect -2016 247722 -2006 247922
rect -1806 247722 108 247922
rect 308 247722 336 247922
rect -2016 247708 -1786 247722
rect 84 247698 336 247722
rect 303888 246356 304300 249038
rect 303888 246038 303926 246356
rect 304244 246038 304300 246356
rect -2016 244922 -1786 244930
rect 84 244922 336 244942
rect -2016 244722 -2006 244922
rect -1806 244722 108 244922
rect 308 244722 336 244922
rect -2016 244708 -1786 244722
rect 84 244698 336 244722
rect 303888 243356 304300 246038
rect 303888 243038 303926 243356
rect 304244 243038 304300 243356
rect -2016 241922 -1786 241930
rect 84 241922 336 241942
rect -2016 241722 -2006 241922
rect -1806 241722 108 241922
rect 308 241722 336 241922
rect -2016 241708 -1786 241722
rect 84 241698 336 241722
rect 303888 240356 304300 243038
rect 303888 240038 303926 240356
rect 304244 240038 304300 240356
rect -2016 238922 -1786 238930
rect 84 238922 336 238942
rect -2016 238722 -2006 238922
rect -1806 238722 108 238922
rect 308 238722 336 238922
rect -2016 238708 -1786 238722
rect 84 238698 336 238722
rect 303888 237356 304300 240038
rect 303888 237038 303926 237356
rect 304244 237038 304300 237356
rect -2016 235922 -1786 235930
rect 84 235922 336 235942
rect -2016 235722 -2006 235922
rect -1806 235722 108 235922
rect 308 235722 336 235922
rect -2016 235708 -1786 235722
rect 84 235698 336 235722
rect 303888 234356 304300 237038
rect 303888 234038 303926 234356
rect 304244 234038 304300 234356
rect -2016 232922 -1786 232930
rect 84 232922 336 232942
rect -2016 232722 -2006 232922
rect -1806 232722 108 232922
rect 308 232722 336 232922
rect -2016 232708 -1786 232722
rect 84 232698 336 232722
rect 303888 231356 304300 234038
rect 303888 231038 303926 231356
rect 304244 231038 304300 231356
rect -2016 229922 -1786 229930
rect 84 229922 336 229942
rect -2016 229722 -2006 229922
rect -1806 229722 108 229922
rect 308 229722 336 229922
rect -2016 229708 -1786 229722
rect 84 229698 336 229722
rect 303888 228356 304300 231038
rect 303888 228038 303926 228356
rect 304244 228038 304300 228356
rect -2016 226922 -1786 226930
rect 84 226922 336 226942
rect -2016 226722 -2006 226922
rect -1806 226722 108 226922
rect 308 226722 336 226922
rect -2016 226708 -1786 226722
rect 84 226698 336 226722
rect 303888 225356 304300 228038
rect 303888 225038 303926 225356
rect 304244 225038 304300 225356
rect -2016 223922 -1786 223930
rect 84 223922 336 223942
rect -2016 223722 -2006 223922
rect -1806 223722 108 223922
rect 308 223722 336 223922
rect -2016 223708 -1786 223722
rect 84 223698 336 223722
rect 303888 222356 304300 225038
rect 303888 222038 303926 222356
rect 304244 222038 304300 222356
rect -2016 220922 -1786 220930
rect 84 220922 336 220942
rect -2016 220722 -2006 220922
rect -1806 220722 108 220922
rect 308 220722 336 220922
rect -2016 220708 -1786 220722
rect 84 220698 336 220722
rect 303888 219356 304300 222038
rect 303888 219038 303926 219356
rect 304244 219038 304300 219356
rect -2016 217922 -1786 217930
rect 84 217922 336 217942
rect -2016 217722 -2006 217922
rect -1806 217722 108 217922
rect 308 217722 336 217922
rect -2016 217708 -1786 217722
rect 84 217698 336 217722
rect 303888 216356 304300 219038
rect 303888 216038 303926 216356
rect 304244 216038 304300 216356
rect -2016 214922 -1786 214930
rect 84 214922 336 214942
rect -2016 214722 -2006 214922
rect -1806 214722 108 214922
rect 308 214722 336 214922
rect -2016 214708 -1786 214722
rect 84 214698 336 214722
rect 303888 213356 304300 216038
rect 303888 213038 303926 213356
rect 304244 213038 304300 213356
rect -2016 211922 -1786 211930
rect 84 211922 336 211942
rect -2016 211722 -2006 211922
rect -1806 211722 108 211922
rect 308 211722 336 211922
rect -2016 211708 -1786 211722
rect 84 211698 336 211722
rect 303888 210356 304300 213038
rect 303888 210038 303926 210356
rect 304244 210038 304300 210356
rect -2016 208922 -1786 208930
rect 84 208922 336 208942
rect -2016 208722 -2006 208922
rect -1806 208722 108 208922
rect 308 208722 336 208922
rect -2016 208708 -1786 208722
rect 84 208698 336 208722
rect 303888 207356 304300 210038
rect 303888 207038 303926 207356
rect 304244 207038 304300 207356
rect -2016 205922 -1786 205930
rect 84 205922 336 205942
rect -2016 205722 -2006 205922
rect -1806 205722 108 205922
rect 308 205722 336 205922
rect -2016 205708 -1786 205722
rect 84 205698 336 205722
rect 303888 204356 304300 207038
rect 303888 204038 303926 204356
rect 304244 204038 304300 204356
rect -2016 202922 -1786 202930
rect 84 202922 336 202942
rect -2016 202722 -2006 202922
rect -1806 202722 108 202922
rect 308 202722 336 202922
rect -2016 202708 -1786 202722
rect 84 202698 336 202722
rect 303888 201356 304300 204038
rect 303888 201038 303926 201356
rect 304244 201038 304300 201356
rect -2016 199922 -1786 199930
rect 84 199922 336 199942
rect -2016 199722 -2006 199922
rect -1806 199722 108 199922
rect 308 199722 336 199922
rect -2016 199708 -1786 199722
rect 84 199698 336 199722
rect 303888 198356 304300 201038
rect 303888 198038 303926 198356
rect 304244 198038 304300 198356
rect -2016 196922 -1786 196930
rect 84 196922 336 196942
rect -2016 196722 -2006 196922
rect -1806 196722 108 196922
rect 308 196722 336 196922
rect -2016 196708 -1786 196722
rect 84 196698 336 196722
rect 303888 195356 304300 198038
rect 303888 195038 303926 195356
rect 304244 195038 304300 195356
rect -2016 193922 -1786 193930
rect 84 193922 336 193942
rect -2016 193722 -2006 193922
rect -1806 193722 108 193922
rect 308 193722 336 193922
rect -2016 193708 -1786 193722
rect 84 193698 336 193722
rect 303888 192356 304300 195038
rect 303888 192038 303926 192356
rect 304244 192038 304300 192356
rect -2016 190922 -1786 190930
rect 84 190922 336 190942
rect -2016 190722 -2006 190922
rect -1806 190722 108 190922
rect 308 190722 336 190922
rect -2016 190708 -1786 190722
rect 84 190698 336 190722
rect 303888 189356 304300 192038
rect 303888 189038 303926 189356
rect 304244 189038 304300 189356
rect -2016 187922 -1786 187930
rect 84 187922 336 187942
rect -2016 187722 -2006 187922
rect -1806 187722 108 187922
rect 308 187722 336 187922
rect -2016 187708 -1786 187722
rect 84 187698 336 187722
rect 303888 186356 304300 189038
rect 303888 186038 303926 186356
rect 304244 186038 304300 186356
rect -2016 184922 -1786 184930
rect 84 184922 336 184942
rect -2016 184722 -2006 184922
rect -1806 184722 108 184922
rect 308 184722 336 184922
rect -2016 184708 -1786 184722
rect 84 184698 336 184722
rect 303888 183356 304300 186038
rect 303888 183038 303926 183356
rect 304244 183038 304300 183356
rect -2016 181922 -1786 181930
rect 84 181922 336 181942
rect -2016 181722 -2006 181922
rect -1806 181722 108 181922
rect 308 181722 336 181922
rect -2016 181708 -1786 181722
rect 84 181698 336 181722
rect 303888 180356 304300 183038
rect 303888 180038 303926 180356
rect 304244 180038 304300 180356
rect -2016 178922 -1786 178930
rect 84 178922 336 178942
rect -2016 178722 -2006 178922
rect -1806 178722 108 178922
rect 308 178722 336 178922
rect -2016 178708 -1786 178722
rect 84 178698 336 178722
rect 303888 177356 304300 180038
rect 303888 177038 303926 177356
rect 304244 177038 304300 177356
rect -2016 175922 -1786 175930
rect 84 175922 336 175942
rect -2016 175722 -2006 175922
rect -1806 175722 108 175922
rect 308 175722 336 175922
rect -2016 175708 -1786 175722
rect 84 175698 336 175722
rect 303888 174356 304300 177038
rect 303888 174038 303926 174356
rect 304244 174038 304300 174356
rect -2016 172922 -1786 172930
rect 84 172922 336 172942
rect -2016 172722 -2006 172922
rect -1806 172722 108 172922
rect 308 172722 336 172922
rect -2016 172708 -1786 172722
rect 84 172698 336 172722
rect 303888 171356 304300 174038
rect 303888 171038 303926 171356
rect 304244 171038 304300 171356
rect -2016 169922 -1786 169930
rect 84 169922 336 169942
rect -2016 169722 -2006 169922
rect -1806 169722 108 169922
rect 308 169722 336 169922
rect -2016 169708 -1786 169722
rect 84 169698 336 169722
rect 303888 168356 304300 171038
rect 303888 168038 303926 168356
rect 304244 168038 304300 168356
rect -2016 166922 -1786 166930
rect 84 166922 336 166942
rect -2016 166722 -2006 166922
rect -1806 166722 108 166922
rect 308 166722 336 166922
rect -2016 166708 -1786 166722
rect 84 166698 336 166722
rect 303888 165356 304300 168038
rect 303888 165038 303926 165356
rect 304244 165038 304300 165356
rect -2016 163922 -1786 163930
rect 84 163922 336 163942
rect -2016 163722 -2006 163922
rect -1806 163722 108 163922
rect 308 163722 336 163922
rect -2016 163708 -1786 163722
rect 84 163698 336 163722
rect 303888 162356 304300 165038
rect 303888 162038 303926 162356
rect 304244 162038 304300 162356
rect -2016 160922 -1786 160930
rect 84 160922 336 160942
rect -2016 160722 -2006 160922
rect -1806 160722 108 160922
rect 308 160722 336 160922
rect -2016 160708 -1786 160722
rect 84 160698 336 160722
rect 303888 159356 304300 162038
rect 303888 159038 303926 159356
rect 304244 159038 304300 159356
rect -2016 157922 -1786 157930
rect 84 157922 336 157942
rect -2016 157722 -2006 157922
rect -1806 157722 108 157922
rect 308 157722 336 157922
rect -2016 157708 -1786 157722
rect 84 157698 336 157722
rect 303888 156356 304300 159038
rect 303888 156038 303926 156356
rect 304244 156038 304300 156356
rect -2016 154922 -1786 154930
rect 84 154922 336 154942
rect -2016 154722 -2006 154922
rect -1806 154722 108 154922
rect 308 154722 336 154922
rect -2016 154708 -1786 154722
rect 84 154698 336 154722
rect 303888 153356 304300 156038
rect 303888 153038 303926 153356
rect 304244 153038 304300 153356
rect -2016 151922 -1786 151930
rect 84 151922 336 151942
rect -2016 151722 -2006 151922
rect -1806 151722 108 151922
rect 308 151722 336 151922
rect -2016 151708 -1786 151722
rect 84 151698 336 151722
rect 303888 150356 304300 153038
rect 303888 150038 303926 150356
rect 304244 150038 304300 150356
rect -2016 148922 -1786 148930
rect 84 148922 336 148942
rect -2016 148722 -2006 148922
rect -1806 148722 108 148922
rect 308 148722 336 148922
rect -2016 148708 -1786 148722
rect 84 148698 336 148722
rect 303888 147356 304300 150038
rect 303888 147038 303926 147356
rect 304244 147038 304300 147356
rect -2016 145922 -1786 145930
rect 84 145922 336 145942
rect -2016 145722 -2006 145922
rect -1806 145722 108 145922
rect 308 145722 336 145922
rect -2016 145708 -1786 145722
rect 84 145698 336 145722
rect 303888 144356 304300 147038
rect 303888 144038 303926 144356
rect 304244 144038 304300 144356
rect -2016 142922 -1786 142930
rect 84 142922 336 142942
rect -2016 142722 -2006 142922
rect -1806 142722 108 142922
rect 308 142722 336 142922
rect -2016 142708 -1786 142722
rect 84 142698 336 142722
rect 303888 141356 304300 144038
rect 303888 141038 303926 141356
rect 304244 141038 304300 141356
rect -2016 139922 -1786 139930
rect 84 139922 336 139942
rect -2016 139722 -2006 139922
rect -1806 139722 108 139922
rect 308 139722 336 139922
rect -2016 139708 -1786 139722
rect 84 139698 336 139722
rect 303888 138356 304300 141038
rect 303888 138038 303926 138356
rect 304244 138038 304300 138356
rect -2016 136922 -1786 136930
rect 84 136922 336 136942
rect -2016 136722 -2006 136922
rect -1806 136722 108 136922
rect 308 136722 336 136922
rect -2016 136708 -1786 136722
rect 84 136698 336 136722
rect 303888 135356 304300 138038
rect 303888 135038 303926 135356
rect 304244 135038 304300 135356
rect -2016 133922 -1786 133930
rect 84 133922 336 133942
rect -2016 133722 -2006 133922
rect -1806 133722 108 133922
rect 308 133722 336 133922
rect -2016 133708 -1786 133722
rect 84 133698 336 133722
rect 303888 132356 304300 135038
rect 303888 132038 303926 132356
rect 304244 132038 304300 132356
rect -2016 130922 -1786 130930
rect 84 130922 336 130942
rect -2016 130722 -2006 130922
rect -1806 130722 108 130922
rect 308 130722 336 130922
rect -2016 130708 -1786 130722
rect 84 130698 336 130722
rect 303888 129356 304300 132038
rect 303888 129038 303926 129356
rect 304244 129038 304300 129356
rect -2016 127922 -1786 127930
rect 84 127922 336 127942
rect -2016 127722 -2006 127922
rect -1806 127722 108 127922
rect 308 127722 336 127922
rect -2016 127708 -1786 127722
rect 84 127698 336 127722
rect 303888 126356 304300 129038
rect 303888 126038 303926 126356
rect 304244 126038 304300 126356
rect -2016 124922 -1786 124930
rect 84 124922 336 124942
rect -2016 124722 -2006 124922
rect -1806 124722 108 124922
rect 308 124722 336 124922
rect -2016 124708 -1786 124722
rect 84 124698 336 124722
rect 303888 123356 304300 126038
rect 303888 123038 303926 123356
rect 304244 123038 304300 123356
rect -2016 121922 -1786 121930
rect 84 121922 336 121942
rect -2016 121722 -2006 121922
rect -1806 121722 108 121922
rect 308 121722 336 121922
rect -2016 121708 -1786 121722
rect 84 121698 336 121722
rect 303888 120356 304300 123038
rect 303888 120038 303926 120356
rect 304244 120038 304300 120356
rect -2016 118922 -1786 118930
rect 84 118922 336 118942
rect -2016 118722 -2006 118922
rect -1806 118722 108 118922
rect 308 118722 336 118922
rect -2016 118708 -1786 118722
rect 84 118698 336 118722
rect 303888 117356 304300 120038
rect 303888 117038 303926 117356
rect 304244 117038 304300 117356
rect -2016 115922 -1786 115930
rect 84 115922 336 115942
rect -2016 115722 -2006 115922
rect -1806 115722 108 115922
rect 308 115722 336 115922
rect -2016 115708 -1786 115722
rect 84 115698 336 115722
rect 303888 114356 304300 117038
rect 303888 114038 303926 114356
rect 304244 114038 304300 114356
rect -2016 112922 -1786 112930
rect 84 112922 336 112942
rect -2016 112722 -2006 112922
rect -1806 112722 108 112922
rect 308 112722 336 112922
rect -2016 112708 -1786 112722
rect 84 112698 336 112722
rect 303888 111356 304300 114038
rect 303888 111038 303926 111356
rect 304244 111038 304300 111356
rect -2016 109922 -1786 109930
rect 84 109922 336 109942
rect -2016 109722 -2006 109922
rect -1806 109722 108 109922
rect 308 109722 336 109922
rect -2016 109708 -1786 109722
rect 84 109698 336 109722
rect 303888 108356 304300 111038
rect 303888 108038 303926 108356
rect 304244 108038 304300 108356
rect -2016 106922 -1786 106930
rect 84 106922 336 106942
rect -2016 106722 -2006 106922
rect -1806 106722 108 106922
rect 308 106722 336 106922
rect -2016 106708 -1786 106722
rect 84 106698 336 106722
rect 303888 105356 304300 108038
rect 303888 105038 303926 105356
rect 304244 105038 304300 105356
rect -2016 103922 -1786 103930
rect 84 103922 336 103942
rect -2016 103722 -2006 103922
rect -1806 103722 108 103922
rect 308 103722 336 103922
rect -2016 103708 -1786 103722
rect 84 103698 336 103722
rect 303888 102356 304300 105038
rect 303888 102038 303926 102356
rect 304244 102038 304300 102356
rect -2016 100922 -1786 100930
rect 84 100922 336 100942
rect -2016 100722 -2006 100922
rect -1806 100722 108 100922
rect 308 100722 336 100922
rect -2016 100708 -1786 100722
rect 84 100698 336 100722
rect 303888 99356 304300 102038
rect 303888 99038 303926 99356
rect 304244 99038 304300 99356
rect -2016 97922 -1786 97930
rect 84 97922 336 97942
rect -2016 97722 -2006 97922
rect -1806 97722 108 97922
rect 308 97722 336 97922
rect -2016 97708 -1786 97722
rect 84 97698 336 97722
rect 303888 96356 304300 99038
rect 303888 96038 303926 96356
rect 304244 96038 304300 96356
rect -2016 94922 -1786 94930
rect 84 94922 336 94942
rect -2016 94722 -2006 94922
rect -1806 94722 108 94922
rect 308 94722 336 94922
rect -2016 94708 -1786 94722
rect 84 94698 336 94722
rect 303888 93356 304300 96038
rect 303888 93038 303926 93356
rect 304244 93038 304300 93356
rect -2016 91922 -1786 91930
rect 84 91922 336 91942
rect -2016 91722 -2006 91922
rect -1806 91722 108 91922
rect 308 91722 336 91922
rect -2016 91708 -1786 91722
rect 84 91698 336 91722
rect 303888 90356 304300 93038
rect 303888 90038 303926 90356
rect 304244 90038 304300 90356
rect -2016 88922 -1786 88930
rect 84 88922 336 88942
rect -2016 88722 -2006 88922
rect -1806 88722 108 88922
rect 308 88722 336 88922
rect -2016 88708 -1786 88722
rect 84 88698 336 88722
rect 303888 87356 304300 90038
rect 303888 87038 303926 87356
rect 304244 87038 304300 87356
rect -2016 85922 -1786 85930
rect 84 85922 336 85942
rect -2016 85722 -2006 85922
rect -1806 85722 108 85922
rect 308 85722 336 85922
rect -2016 85708 -1786 85722
rect 84 85698 336 85722
rect 303888 84356 304300 87038
rect 303888 84038 303926 84356
rect 304244 84038 304300 84356
rect -2016 82922 -1786 82930
rect 84 82922 336 82942
rect -2016 82722 -2006 82922
rect -1806 82722 108 82922
rect 308 82722 336 82922
rect -2016 82708 -1786 82722
rect 84 82698 336 82722
rect 303888 81356 304300 84038
rect 303888 81038 303926 81356
rect 304244 81038 304300 81356
rect -2016 79922 -1786 79930
rect 84 79922 336 79942
rect -2016 79722 -2006 79922
rect -1806 79722 108 79922
rect 308 79722 336 79922
rect -2016 79708 -1786 79722
rect 84 79698 336 79722
rect 303888 78356 304300 81038
rect 303888 78038 303926 78356
rect 304244 78038 304300 78356
rect -2016 76922 -1786 76930
rect 84 76922 336 76942
rect -2016 76722 -2006 76922
rect -1806 76722 108 76922
rect 308 76722 336 76922
rect -2016 76708 -1786 76722
rect 84 76698 336 76722
rect 303888 75356 304300 78038
rect 303888 75038 303926 75356
rect 304244 75038 304300 75356
rect -2016 73922 -1786 73930
rect 84 73922 336 73942
rect -2016 73722 -2006 73922
rect -1806 73722 108 73922
rect 308 73722 336 73922
rect -2016 73708 -1786 73722
rect 84 73698 336 73722
rect 303888 72356 304300 75038
rect 303888 72038 303926 72356
rect 304244 72038 304300 72356
rect -2016 70922 -1786 70930
rect 84 70922 336 70942
rect -2016 70722 -2006 70922
rect -1806 70722 108 70922
rect 308 70722 336 70922
rect -2016 70708 -1786 70722
rect 84 70698 336 70722
rect 303888 69356 304300 72038
rect 303888 69038 303926 69356
rect 304244 69038 304300 69356
rect -2016 67922 -1786 67930
rect 84 67922 336 67942
rect -2016 67722 -2006 67922
rect -1806 67722 108 67922
rect 308 67722 336 67922
rect -2016 67708 -1786 67722
rect 84 67698 336 67722
rect 303888 66356 304300 69038
rect 303888 66038 303926 66356
rect 304244 66038 304300 66356
rect -2016 64922 -1786 64930
rect 84 64922 336 64942
rect -2016 64722 -2006 64922
rect -1806 64722 108 64922
rect 308 64722 336 64922
rect -2016 64708 -1786 64722
rect 84 64698 336 64722
rect 303888 63356 304300 66038
rect 303888 63038 303926 63356
rect 304244 63038 304300 63356
rect -2016 61922 -1786 61930
rect 84 61922 336 61942
rect -2016 61722 -2006 61922
rect -1806 61722 108 61922
rect 308 61722 336 61922
rect -2016 61708 -1786 61722
rect 84 61698 336 61722
rect 303888 60356 304300 63038
rect 303888 60038 303926 60356
rect 304244 60038 304300 60356
rect -2016 58922 -1786 58930
rect 84 58922 336 58942
rect -2016 58722 -2006 58922
rect -1806 58722 108 58922
rect 308 58722 336 58922
rect -2016 58708 -1786 58722
rect 84 58698 336 58722
rect 303888 57356 304300 60038
rect 303888 57038 303926 57356
rect 304244 57038 304300 57356
rect -2016 55922 -1786 55930
rect 84 55922 336 55942
rect -2016 55722 -2006 55922
rect -1806 55722 108 55922
rect 308 55722 336 55922
rect -2016 55708 -1786 55722
rect 84 55698 336 55722
rect 303888 54356 304300 57038
rect 303888 54038 303926 54356
rect 304244 54038 304300 54356
rect -2016 52922 -1786 52930
rect 84 52922 336 52942
rect -2016 52722 -2006 52922
rect -1806 52722 108 52922
rect 308 52722 336 52922
rect -2016 52708 -1786 52722
rect 84 52698 336 52722
rect 303888 51356 304300 54038
rect 303888 51038 303926 51356
rect 304244 51038 304300 51356
rect -2016 49922 -1786 49930
rect 84 49922 336 49942
rect -2016 49722 -2006 49922
rect -1806 49722 108 49922
rect 308 49722 336 49922
rect -2016 49708 -1786 49722
rect 84 49698 336 49722
rect 303888 48356 304300 51038
rect 303888 48038 303926 48356
rect 304244 48038 304300 48356
rect -2016 46922 -1786 46930
rect 84 46922 336 46942
rect -2016 46722 -2006 46922
rect -1806 46722 108 46922
rect 308 46722 336 46922
rect -2016 46708 -1786 46722
rect 84 46698 336 46722
rect 303888 45356 304300 48038
rect 303888 45038 303926 45356
rect 304244 45038 304300 45356
rect -2016 43922 -1786 43930
rect 84 43922 336 43942
rect -2016 43722 -2006 43922
rect -1806 43722 108 43922
rect 308 43722 336 43922
rect -2016 43708 -1786 43722
rect 84 43698 336 43722
rect 303888 42356 304300 45038
rect 303888 42038 303926 42356
rect 304244 42038 304300 42356
rect -2016 40922 -1786 40930
rect 84 40922 336 40942
rect -2016 40722 -2006 40922
rect -1806 40722 108 40922
rect 308 40722 336 40922
rect -2016 40708 -1786 40722
rect 84 40698 336 40722
rect 303888 39356 304300 42038
rect 303888 39038 303926 39356
rect 304244 39038 304300 39356
rect -2044 37922 -1762 37940
rect 84 37922 336 37942
rect -2044 37722 -2006 37922
rect -1806 37722 108 37922
rect 308 37722 336 37922
rect -2044 37700 -1762 37722
rect 84 37698 336 37722
rect 303888 36356 304300 39038
rect 303888 36038 303926 36356
rect 304244 36038 304300 36356
rect -2030 34930 -1788 34970
rect -2030 34922 -1786 34930
rect 84 34922 336 34942
rect -2030 34722 -2006 34922
rect -1806 34722 108 34922
rect 308 34722 336 34922
rect -2030 34708 -1786 34722
rect -2030 34702 -1788 34708
rect -2004 34690 -1788 34702
rect 84 34698 336 34722
rect 303888 33356 304300 36038
rect 303888 33038 303926 33356
rect 304244 33038 304300 33356
rect -2046 31922 -1772 31996
rect 84 31938 336 31942
rect 72 31922 352 31938
rect -2046 31722 -2006 31922
rect -1806 31722 108 31922
rect 308 31722 352 31922
rect -2046 31696 -1772 31722
rect 72 31684 352 31722
rect 303888 30356 304300 33038
rect 303888 30038 303926 30356
rect 304244 30038 304300 30356
rect -2016 28922 -1778 28946
rect 82 28922 354 28944
rect -2016 28722 -2006 28922
rect -1806 28722 108 28922
rect 308 28722 354 28922
rect -2016 28696 -1778 28722
rect 82 28692 354 28722
rect 303888 27356 304300 30038
rect 303888 27038 303926 27356
rect 304244 27038 304300 27356
rect 70 25942 330 25946
rect -2050 25930 -1806 25934
rect -2050 25922 -1786 25930
rect 70 25922 336 25942
rect -2050 25722 -2006 25922
rect -1806 25722 108 25922
rect 308 25722 336 25922
rect -2050 25708 -1786 25722
rect -2050 25692 -1806 25708
rect 70 25698 336 25722
rect 70 25684 330 25698
rect 303888 24356 304300 27038
rect 303888 24038 303926 24356
rect 304244 24038 304300 24356
rect -2026 22930 -1792 22942
rect 84 22932 336 22942
rect -2026 22922 -1786 22930
rect 84 22922 338 22932
rect -2026 22722 -2006 22922
rect -1806 22722 108 22922
rect 308 22722 338 22922
rect -2026 22708 -1786 22722
rect -2026 22706 -1792 22708
rect 84 22704 338 22722
rect 84 22698 336 22704
rect 303888 21372 304300 24038
rect 303888 21356 304304 21372
rect 303888 21038 303926 21356
rect 304244 21038 304304 21356
rect 303888 21004 304304 21038
rect 303888 20952 304300 21004
rect 19796 19192 20146 19256
rect 19796 18974 19870 19192
rect 20088 18974 20146 19192
rect 38280 19218 38600 19236
rect 29054 19062 29324 19088
rect 25938 19014 26174 19020
rect 7442 18890 7772 18958
rect 5280 18784 5646 18878
rect 5280 18566 5328 18784
rect 5546 18566 5646 18784
rect 7442 18672 7482 18890
rect 7700 18672 7772 18890
rect 13800 18928 14038 18946
rect 7442 18632 7772 18672
rect 10640 18834 11000 18876
rect 10640 18616 10712 18834
rect 10930 18616 11000 18834
rect 13800 18710 13802 18928
rect 14020 18710 14038 18928
rect 19796 18896 20146 18974
rect 25934 19012 26174 19014
rect 25934 19010 26178 19012
rect 13800 18698 14038 18710
rect 16870 18816 17188 18856
rect 10640 18576 11000 18616
rect 16870 18598 16912 18816
rect 17130 18598 17188 18816
rect 25934 18792 25944 19010
rect 26162 18792 26178 19010
rect 29054 18842 29084 19062
rect 29304 18842 29324 19062
rect 35314 19054 35564 19058
rect 29054 18808 29324 18842
rect 32314 18986 32562 18994
rect 25934 18788 26178 18792
rect 25934 18782 26170 18788
rect 32314 18768 32328 18986
rect 32546 18768 32562 18986
rect 35314 18836 35328 19054
rect 35546 18836 35564 19054
rect 38280 19000 38328 19218
rect 38546 19000 38600 19218
rect 56590 19162 56858 19182
rect 47292 19130 47590 19154
rect 38280 18958 38600 19000
rect 44294 18922 44700 19020
rect 35314 18822 35564 18836
rect 41310 18872 41582 18898
rect 32314 18756 32562 18768
rect 5280 18454 5646 18566
rect 16870 18554 17188 18598
rect 22880 18658 23142 18674
rect 2324 18438 2554 18442
rect 2322 18220 2328 18438
rect 2546 18220 2554 18438
rect 22880 18440 22898 18658
rect 23116 18440 23142 18658
rect 41310 18654 41328 18872
rect 41546 18654 41582 18872
rect 41310 18618 41582 18654
rect 44294 18704 44328 18922
rect 44546 18704 44700 18922
rect 47292 18912 47328 19130
rect 47546 18912 47590 19130
rect 53518 19042 53776 19056
rect 50516 19014 50734 19016
rect 47292 18900 47590 18912
rect 50508 19010 50744 19014
rect 50508 18792 50516 19010
rect 50734 18792 50744 19010
rect 53518 18824 53538 19042
rect 53756 18824 53776 19042
rect 56590 18944 56616 19162
rect 56834 18944 56858 19162
rect 174332 19134 174626 19162
rect 71914 19060 72174 19076
rect 68290 18968 68580 18992
rect 56590 18922 56858 18944
rect 53518 18808 53776 18824
rect 59606 18866 59858 18888
rect 50508 18788 50744 18792
rect 50516 18786 50734 18788
rect 44294 18596 44700 18704
rect 59606 18648 59630 18866
rect 59848 18648 59858 18866
rect 65716 18880 66082 18964
rect 59606 18634 59858 18648
rect 62572 18790 62974 18834
rect 62572 18572 62632 18790
rect 62850 18572 62974 18790
rect 65716 18662 65742 18880
rect 65960 18662 66082 18880
rect 68290 18952 68784 18968
rect 68290 18734 68328 18952
rect 68546 18948 68784 18952
rect 68546 18738 68554 18948
rect 68764 18738 68784 18948
rect 71914 18842 71928 19060
rect 72146 18842 72174 19060
rect 71914 18828 72174 18842
rect 75054 19030 75306 19042
rect 68546 18734 68784 18738
rect 68290 18726 68784 18734
rect 65716 18648 66082 18662
rect 62572 18542 62974 18572
rect 71928 18536 72148 18828
rect 75054 18812 75078 19030
rect 75296 18812 75306 19030
rect 108892 19032 109134 19040
rect 81190 18904 81410 18906
rect 75054 18798 75306 18812
rect 81184 18720 81190 18904
rect 81172 18686 81190 18720
rect 81408 18720 81414 18904
rect 96442 18874 96684 18884
rect 90400 18836 90652 18856
rect 81408 18686 81430 18720
rect 22880 18422 23142 18440
rect 71910 18520 72162 18536
rect 71910 18310 71932 18520
rect 72142 18310 72162 18520
rect 81172 18496 81194 18686
rect 81404 18496 81430 18686
rect 90400 18618 90412 18836
rect 90630 18618 90652 18836
rect 90400 18608 90652 18618
rect 93536 18792 93788 18810
rect 93536 18574 93556 18792
rect 93774 18574 93788 18792
rect 96442 18656 96454 18874
rect 96672 18656 96684 18874
rect 108892 18814 108902 19032
rect 109120 18814 109134 19032
rect 114930 18984 115200 19008
rect 108892 18808 109134 18814
rect 111936 18934 112184 18948
rect 96442 18650 96684 18656
rect 102658 18740 102952 18774
rect 93536 18562 93788 18574
rect 102658 18522 102712 18740
rect 102930 18522 102952 18740
rect 81172 18482 81430 18496
rect 99582 18500 99842 18518
rect 84274 18404 84492 18408
rect 84274 18402 84494 18404
rect 71910 18292 72162 18310
rect 78098 18306 78316 18312
rect 2324 18204 2554 18220
rect 78316 18088 78318 18306
rect 84492 18184 84494 18402
rect 78074 18076 78350 18088
rect -6210 17946 -5984 17960
rect -6210 17942 -6198 17946
rect -5998 17942 -5984 17946
rect -6210 17742 -6204 17942
rect -5994 17742 -5984 17942
rect 78074 17866 78102 18076
rect 78312 17866 78350 18076
rect 84274 18028 84494 18184
rect 87330 18314 87580 18326
rect 87330 18096 87336 18314
rect 87554 18096 87580 18314
rect 99582 18282 99598 18500
rect 99816 18282 99842 18500
rect 102658 18468 102952 18522
rect 105620 18754 105914 18790
rect 105620 18536 105676 18754
rect 105894 18536 105914 18754
rect 111936 18716 111948 18934
rect 112166 18716 112184 18934
rect 114930 18766 114954 18984
rect 115172 18766 115200 18984
rect 114930 18744 115200 18766
rect 117942 18976 118250 18998
rect 117942 18758 117968 18976
rect 118186 18758 118250 18976
rect 157794 18996 158088 19008
rect 127190 18942 127500 18970
rect 111936 18712 112184 18716
rect 111948 18710 112166 18712
rect 117942 18686 118250 18758
rect 121114 18864 121400 18884
rect 121114 18646 121150 18864
rect 121368 18646 121400 18864
rect 121114 18598 121400 18646
rect 124096 18852 124354 18864
rect 124096 18632 124118 18852
rect 124338 18632 124354 18852
rect 127190 18724 127242 18942
rect 127460 18724 127500 18942
rect 133376 18866 133686 18894
rect 127190 18678 127500 18724
rect 130210 18812 130520 18858
rect 124096 18624 124354 18632
rect 130210 18594 130250 18812
rect 130468 18594 130520 18812
rect 133376 18646 133412 18866
rect 133632 18646 133686 18866
rect 145538 18842 145832 18860
rect 133376 18602 133686 18646
rect 142576 18668 142876 18684
rect 130210 18566 130520 18594
rect 139492 18600 139802 18606
rect 105620 18484 105914 18536
rect 139492 18382 139552 18600
rect 139770 18382 139802 18600
rect 142576 18450 142600 18668
rect 142818 18450 142876 18668
rect 145538 18624 145578 18842
rect 145796 18624 145832 18842
rect 145538 18580 145832 18624
rect 148714 18842 149008 18874
rect 148714 18624 148754 18842
rect 148972 18624 149008 18842
rect 154754 18858 155048 18876
rect 148714 18594 149008 18624
rect 151732 18774 152026 18802
rect 151732 18556 151772 18774
rect 151990 18556 152026 18774
rect 154754 18640 154792 18858
rect 155010 18640 155048 18858
rect 157794 18778 157844 18996
rect 158062 18778 158088 18996
rect 174332 18916 174366 19134
rect 174584 18916 174626 19134
rect 305362 19098 305616 19106
rect 290286 18954 290586 18982
rect 174332 18882 174626 18916
rect 229636 18938 229916 18952
rect 176292 18812 176586 18846
rect 157794 18728 158088 18778
rect 160862 18758 161156 18778
rect 154754 18596 155048 18640
rect 151732 18522 152026 18556
rect 160862 18540 160886 18758
rect 161104 18540 161156 18758
rect 176292 18594 176328 18812
rect 176546 18594 176586 18812
rect 229636 18720 229658 18938
rect 229876 18720 229916 18938
rect 290286 18736 290328 18954
rect 290546 18736 290586 18954
rect 305362 18880 305386 19098
rect 305604 18880 305616 19098
rect 305362 18850 305616 18880
rect 229636 18700 229916 18720
rect 176292 18566 176586 18594
rect 233310 18688 233574 18702
rect 160862 18498 161156 18540
rect 215300 18562 215570 18576
rect 173060 18488 173354 18508
rect 142576 18420 142876 18450
rect 163202 18458 163496 18486
rect 139492 18314 139802 18382
rect 99582 18248 99842 18282
rect 87330 18086 87580 18096
rect 136442 18240 136752 18286
rect 78074 17848 78350 17866
rect 84246 17980 84526 18028
rect 136442 18022 136468 18240
rect 136686 18022 136752 18240
rect 163202 18240 163238 18458
rect 163456 18240 163496 18458
rect 163202 18206 163496 18240
rect 173060 18270 173082 18488
rect 173300 18270 173354 18488
rect 173060 18228 173354 18270
rect 206300 18454 206560 18470
rect 206300 18236 206328 18454
rect 206546 18236 206560 18454
rect 215300 18344 215328 18562
rect 215546 18344 215570 18562
rect 233310 18470 233328 18688
rect 233546 18470 233574 18688
rect 254314 18700 254612 18736
rect 242314 18570 242552 18578
rect 233310 18442 233574 18470
rect 241664 18534 241902 18544
rect 215300 18338 215570 18344
rect 227174 18428 227460 18436
rect 206300 18216 206560 18236
rect 227174 18210 227194 18428
rect 227412 18210 227460 18428
rect 136442 17994 136752 18022
rect 165896 18174 166190 18202
rect 227174 18192 227460 18210
rect 234638 18302 234884 18322
rect 241664 18316 241672 18534
rect 241890 18316 241902 18534
rect 242314 18352 242328 18570
rect 242546 18352 242552 18570
rect 242314 18346 242552 18352
rect 253898 18508 254148 18520
rect 241664 18312 241902 18316
rect 241672 18310 241890 18312
rect -6210 17734 -5984 17742
rect 84246 17770 84278 17980
rect 84488 17770 84526 17980
rect 165896 17956 165928 18174
rect 166146 17956 166190 18174
rect 213128 18098 213386 18108
rect 165896 17922 166190 17956
rect 185290 18036 185584 18060
rect 84246 17732 84526 17770
rect 182444 17858 182738 17894
rect -19160 17346 -19040 17596
rect -15216 17346 -15096 17624
rect -11136 17394 -11016 17688
rect -7192 17338 -7072 17696
rect 182444 17640 182474 17858
rect 182692 17640 182738 17858
rect 185290 17818 185328 18036
rect 185546 17818 185584 18036
rect 200892 17956 201204 18006
rect 185290 17780 185584 17818
rect 196770 17928 197064 17956
rect 196770 17710 196794 17928
rect 197012 17710 197064 17928
rect 182444 17614 182738 17640
rect 188280 17658 188574 17686
rect 196770 17676 197064 17710
rect 200892 17738 200916 17956
rect 201134 17738 201204 17956
rect 213128 17880 213156 18098
rect 213374 17880 213386 18098
rect 234638 18084 234650 18302
rect 234868 18084 234884 18302
rect 253898 18290 253926 18508
rect 254144 18290 254150 18508
rect 254314 18482 254328 18700
rect 254546 18482 254612 18700
rect 279642 18698 279942 18730
rect 254314 18462 254612 18482
rect 268990 18560 269262 18570
rect 268990 18342 269032 18560
rect 269250 18342 269262 18560
rect 279642 18480 279676 18698
rect 279894 18480 279942 18698
rect 290286 18696 290586 18736
rect 302946 18717 303268 18723
rect 279642 18444 279942 18480
rect 268990 18312 269262 18342
rect 253898 18276 254148 18290
rect 269322 18268 269594 18292
rect 234638 18062 234884 18084
rect 261022 18124 261294 18136
rect 213128 17848 213386 17880
rect 240890 18014 241174 18054
rect 240890 17796 240916 18014
rect 241134 17796 241174 18014
rect 261022 17906 261044 18124
rect 261262 17906 261294 18124
rect 269322 18050 269328 18268
rect 269546 18050 269594 18268
rect 269322 18034 269594 18050
rect 278800 18206 279208 18308
rect 278800 17988 278878 18206
rect 279096 17988 279208 18206
rect 292376 18226 292676 18260
rect 261022 17878 261294 17906
rect 265852 17962 266124 17980
rect 200892 17700 201204 17738
rect 206974 17750 207242 17790
rect 240890 17770 241174 17796
rect 249648 17860 249898 17866
rect 168824 17420 169118 17446
rect 168824 17202 168864 17420
rect 169082 17202 169118 17420
rect 188280 17440 188328 17658
rect 188546 17440 188574 17658
rect 206974 17532 207000 17750
rect 207218 17532 207242 17750
rect 206974 17516 207242 17532
rect 221292 17710 221614 17730
rect 221292 17492 221328 17710
rect 221546 17492 221614 17710
rect 249648 17642 249668 17860
rect 249886 17642 249898 17860
rect 265852 17744 265870 17962
rect 266088 17744 266124 17962
rect 278800 17946 279208 17988
rect 284308 18136 284608 18176
rect 284308 17918 284328 18136
rect 284546 17918 284608 18136
rect 292376 18008 292408 18226
rect 292626 18008 292676 18226
rect 302941 18147 302946 18474
rect 303268 18147 303273 18474
rect 302941 18142 303273 18147
rect 292376 17974 292676 18008
rect 284308 17890 284608 17918
rect 265852 17722 266124 17744
rect 299228 17722 299528 17758
rect 249648 17622 249898 17642
rect 221292 17460 221614 17492
rect 277670 17582 277952 17624
rect 188280 17406 188574 17440
rect 277670 17364 277694 17582
rect 277912 17364 277952 17582
rect 277670 17336 277952 17364
rect 286910 17512 287210 17550
rect 286910 17294 286930 17512
rect 287148 17294 287210 17512
rect 299228 17504 299258 17722
rect 299476 17504 299528 17722
rect 299228 17472 299528 17504
rect 168824 17166 169118 17202
rect 213876 17270 214122 17276
rect 213876 17268 214124 17270
rect 183972 17152 184266 17190
rect 183972 16934 184010 17152
rect 184228 16934 184266 17152
rect 213876 17050 213904 17268
rect 214122 17050 214124 17268
rect 286910 17264 287210 17294
rect 260030 17246 260302 17258
rect 220666 17228 220962 17238
rect 213876 17030 214122 17050
rect 193466 17022 193684 17024
rect 183972 16910 184266 16934
rect 193440 17018 193702 17022
rect 193440 16800 193466 17018
rect 193684 16800 193702 17018
rect 220666 17010 220688 17228
rect 220906 17010 220962 17228
rect 220666 17000 220962 17010
rect 248702 17076 248952 17090
rect 193440 16776 193702 16800
rect 201984 16894 202244 16902
rect 201984 16676 202004 16894
rect 202222 16676 202244 16894
rect 248702 16858 248712 17076
rect 248930 16858 248952 17076
rect 260030 17028 260054 17246
rect 260272 17028 260302 17246
rect 260030 17000 260302 17028
rect 300208 17104 300508 17140
rect 248702 16846 248952 16858
rect 300208 16886 300252 17104
rect 300470 16886 300508 17104
rect 300208 16854 300508 16886
rect 201984 16656 202244 16676
rect 302888 16416 303316 16448
rect 302888 16410 302946 16416
rect 303268 16410 303316 16416
rect 302888 16088 302942 16410
rect 303274 16088 303316 16410
rect 302888 16036 303316 16088
rect 26 15588 390 15664
rect 26 15582 108 15588
rect 308 15582 390 15588
rect 26 15382 102 15582
rect 312 15382 390 15582
rect 26 15298 390 15382
rect 306608 14470 306790 14590
rect 306628 10526 306844 10646
rect 114 8622 316 8742
rect 306712 6446 306920 6566
rect 306596 2502 306806 2622
<< via3 >>
rect 302502 324532 302712 324538
rect 302502 324338 302508 324532
rect 302508 324338 302708 324532
rect 302708 324338 302712 324532
rect 303926 321352 304244 321356
rect 303926 321042 303930 321352
rect 303930 321042 304240 321352
rect 304240 321042 304244 321352
rect 303926 321038 304244 321042
rect -2006 319723 -1806 319922
rect -2005 319722 -1806 319723
rect 303926 318352 304244 318356
rect 303926 318042 303930 318352
rect 303930 318042 304240 318352
rect 304240 318042 304244 318352
rect 303926 318038 304244 318042
rect -2006 316722 -1806 316922
rect 303926 315352 304244 315356
rect 303926 315042 303930 315352
rect 303930 315042 304240 315352
rect 304240 315042 304244 315352
rect 303926 315038 304244 315042
rect -2006 313722 -1806 313922
rect 303926 312352 304244 312356
rect 303926 312042 303930 312352
rect 303930 312042 304240 312352
rect 304240 312042 304244 312352
rect 303926 312038 304244 312042
rect -2006 310722 -1806 310922
rect 303926 309352 304244 309356
rect 303926 309042 303930 309352
rect 303930 309042 304240 309352
rect 304240 309042 304244 309352
rect 303926 309038 304244 309042
rect -2006 307722 -1806 307922
rect 303926 306352 304244 306356
rect 303926 306042 303930 306352
rect 303930 306042 304240 306352
rect 304240 306042 304244 306352
rect 303926 306038 304244 306042
rect -2006 304722 -1806 304922
rect 303926 303352 304244 303356
rect 303926 303042 303930 303352
rect 303930 303042 304240 303352
rect 304240 303042 304244 303352
rect 303926 303038 304244 303042
rect -2006 301722 -1806 301922
rect 303926 300352 304244 300356
rect 303926 300042 303930 300352
rect 303930 300042 304240 300352
rect 304240 300042 304244 300352
rect 303926 300038 304244 300042
rect -2006 298722 -1806 298922
rect 303926 297352 304244 297356
rect 303926 297042 303930 297352
rect 303930 297042 304240 297352
rect 304240 297042 304244 297352
rect 303926 297038 304244 297042
rect -2006 295722 -1806 295922
rect 303926 294352 304244 294356
rect 303926 294042 303930 294352
rect 303930 294042 304240 294352
rect 304240 294042 304244 294352
rect 303926 294038 304244 294042
rect -2006 292722 -1806 292922
rect 303926 291352 304244 291356
rect 303926 291042 303930 291352
rect 303930 291042 304240 291352
rect 304240 291042 304244 291352
rect 303926 291038 304244 291042
rect -2006 289722 -1806 289922
rect 303926 288352 304244 288356
rect 303926 288042 303930 288352
rect 303930 288042 304240 288352
rect 304240 288042 304244 288352
rect 303926 288038 304244 288042
rect -2006 286722 -1806 286922
rect 303926 285352 304244 285356
rect 303926 285042 303930 285352
rect 303930 285042 304240 285352
rect 304240 285042 304244 285352
rect 303926 285038 304244 285042
rect -2006 283722 -1806 283922
rect 303926 282352 304244 282356
rect 303926 282042 303930 282352
rect 303930 282042 304240 282352
rect 304240 282042 304244 282352
rect 303926 282038 304244 282042
rect -2006 280722 -1806 280922
rect 303926 279352 304244 279356
rect 303926 279042 303930 279352
rect 303930 279042 304240 279352
rect 304240 279042 304244 279352
rect 303926 279038 304244 279042
rect -2006 277722 -1806 277922
rect 303926 276352 304244 276356
rect 303926 276042 303930 276352
rect 303930 276042 304240 276352
rect 304240 276042 304244 276352
rect 303926 276038 304244 276042
rect -2006 274722 -1806 274922
rect 303926 273352 304244 273356
rect 303926 273042 303930 273352
rect 303930 273042 304240 273352
rect 304240 273042 304244 273352
rect 303926 273038 304244 273042
rect -2006 271722 -1806 271922
rect 303926 270352 304244 270356
rect 303926 270042 303930 270352
rect 303930 270042 304240 270352
rect 304240 270042 304244 270352
rect 303926 270038 304244 270042
rect -2006 268722 -1806 268922
rect 303926 267352 304244 267356
rect 303926 267042 303930 267352
rect 303930 267042 304240 267352
rect 304240 267042 304244 267352
rect 303926 267038 304244 267042
rect -2006 265722 -1806 265922
rect 303926 264352 304244 264356
rect 303926 264042 303930 264352
rect 303930 264042 304240 264352
rect 304240 264042 304244 264352
rect 303926 264038 304244 264042
rect -2006 262722 -1806 262922
rect 303926 261352 304244 261356
rect 303926 261042 303930 261352
rect 303930 261042 304240 261352
rect 304240 261042 304244 261352
rect 303926 261038 304244 261042
rect -2006 259722 -1806 259922
rect 303926 258352 304244 258356
rect 303926 258042 303930 258352
rect 303930 258042 304240 258352
rect 304240 258042 304244 258352
rect 303926 258038 304244 258042
rect -2006 256722 -1806 256922
rect 303926 255352 304244 255356
rect 303926 255042 303930 255352
rect 303930 255042 304240 255352
rect 304240 255042 304244 255352
rect 303926 255038 304244 255042
rect -2006 253722 -1806 253922
rect 303926 252352 304244 252356
rect 303926 252042 303930 252352
rect 303930 252042 304240 252352
rect 304240 252042 304244 252352
rect 303926 252038 304244 252042
rect -2006 250722 -1806 250922
rect 303926 249352 304244 249356
rect 303926 249042 303930 249352
rect 303930 249042 304240 249352
rect 304240 249042 304244 249352
rect 303926 249038 304244 249042
rect -2006 247722 -1806 247922
rect 303926 246352 304244 246356
rect 303926 246042 303930 246352
rect 303930 246042 304240 246352
rect 304240 246042 304244 246352
rect 303926 246038 304244 246042
rect -2006 244722 -1806 244922
rect 303926 243352 304244 243356
rect 303926 243042 303930 243352
rect 303930 243042 304240 243352
rect 304240 243042 304244 243352
rect 303926 243038 304244 243042
rect -2006 241722 -1806 241922
rect 303926 240352 304244 240356
rect 303926 240042 303930 240352
rect 303930 240042 304240 240352
rect 304240 240042 304244 240352
rect 303926 240038 304244 240042
rect -2006 238722 -1806 238922
rect 303926 237352 304244 237356
rect 303926 237042 303930 237352
rect 303930 237042 304240 237352
rect 304240 237042 304244 237352
rect 303926 237038 304244 237042
rect -2006 235722 -1806 235922
rect 303926 234352 304244 234356
rect 303926 234042 303930 234352
rect 303930 234042 304240 234352
rect 304240 234042 304244 234352
rect 303926 234038 304244 234042
rect -2006 232722 -1806 232922
rect 303926 231352 304244 231356
rect 303926 231042 303930 231352
rect 303930 231042 304240 231352
rect 304240 231042 304244 231352
rect 303926 231038 304244 231042
rect -2006 229722 -1806 229922
rect 303926 228352 304244 228356
rect 303926 228042 303930 228352
rect 303930 228042 304240 228352
rect 304240 228042 304244 228352
rect 303926 228038 304244 228042
rect -2006 226722 -1806 226922
rect 303926 225352 304244 225356
rect 303926 225042 303930 225352
rect 303930 225042 304240 225352
rect 304240 225042 304244 225352
rect 303926 225038 304244 225042
rect -2006 223722 -1806 223922
rect 303926 222352 304244 222356
rect 303926 222042 303930 222352
rect 303930 222042 304240 222352
rect 304240 222042 304244 222352
rect 303926 222038 304244 222042
rect -2006 220722 -1806 220922
rect 303926 219352 304244 219356
rect 303926 219042 303930 219352
rect 303930 219042 304240 219352
rect 304240 219042 304244 219352
rect 303926 219038 304244 219042
rect -2006 217722 -1806 217922
rect 303926 216352 304244 216356
rect 303926 216042 303930 216352
rect 303930 216042 304240 216352
rect 304240 216042 304244 216352
rect 303926 216038 304244 216042
rect -2006 214722 -1806 214922
rect 303926 213352 304244 213356
rect 303926 213042 303930 213352
rect 303930 213042 304240 213352
rect 304240 213042 304244 213352
rect 303926 213038 304244 213042
rect -2006 211722 -1806 211922
rect 303926 210352 304244 210356
rect 303926 210042 303930 210352
rect 303930 210042 304240 210352
rect 304240 210042 304244 210352
rect 303926 210038 304244 210042
rect -2006 208722 -1806 208922
rect 303926 207352 304244 207356
rect 303926 207042 303930 207352
rect 303930 207042 304240 207352
rect 304240 207042 304244 207352
rect 303926 207038 304244 207042
rect -2006 205722 -1806 205922
rect 303926 204352 304244 204356
rect 303926 204042 303930 204352
rect 303930 204042 304240 204352
rect 304240 204042 304244 204352
rect 303926 204038 304244 204042
rect -2006 202722 -1806 202922
rect 303926 201352 304244 201356
rect 303926 201042 303930 201352
rect 303930 201042 304240 201352
rect 304240 201042 304244 201352
rect 303926 201038 304244 201042
rect -2006 199722 -1806 199922
rect 303926 198352 304244 198356
rect 303926 198042 303930 198352
rect 303930 198042 304240 198352
rect 304240 198042 304244 198352
rect 303926 198038 304244 198042
rect -2006 196722 -1806 196922
rect 303926 195352 304244 195356
rect 303926 195042 303930 195352
rect 303930 195042 304240 195352
rect 304240 195042 304244 195352
rect 303926 195038 304244 195042
rect -2006 193722 -1806 193922
rect 303926 192352 304244 192356
rect 303926 192042 303930 192352
rect 303930 192042 304240 192352
rect 304240 192042 304244 192352
rect 303926 192038 304244 192042
rect -2006 190722 -1806 190922
rect 303926 189352 304244 189356
rect 303926 189042 303930 189352
rect 303930 189042 304240 189352
rect 304240 189042 304244 189352
rect 303926 189038 304244 189042
rect -2006 187722 -1806 187922
rect 303926 186352 304244 186356
rect 303926 186042 303930 186352
rect 303930 186042 304240 186352
rect 304240 186042 304244 186352
rect 303926 186038 304244 186042
rect -2006 184722 -1806 184922
rect 303926 183352 304244 183356
rect 303926 183042 303930 183352
rect 303930 183042 304240 183352
rect 304240 183042 304244 183352
rect 303926 183038 304244 183042
rect -2006 181722 -1806 181922
rect 303926 180352 304244 180356
rect 303926 180042 303930 180352
rect 303930 180042 304240 180352
rect 304240 180042 304244 180352
rect 303926 180038 304244 180042
rect -2006 178722 -1806 178922
rect 303926 177352 304244 177356
rect 303926 177042 303930 177352
rect 303930 177042 304240 177352
rect 304240 177042 304244 177352
rect 303926 177038 304244 177042
rect -2006 175722 -1806 175922
rect 303926 174352 304244 174356
rect 303926 174042 303930 174352
rect 303930 174042 304240 174352
rect 304240 174042 304244 174352
rect 303926 174038 304244 174042
rect -2006 172722 -1806 172922
rect 303926 171352 304244 171356
rect 303926 171042 303930 171352
rect 303930 171042 304240 171352
rect 304240 171042 304244 171352
rect 303926 171038 304244 171042
rect -2006 169722 -1806 169922
rect 303926 168352 304244 168356
rect 303926 168042 303930 168352
rect 303930 168042 304240 168352
rect 304240 168042 304244 168352
rect 303926 168038 304244 168042
rect -2006 166722 -1806 166922
rect 303926 165352 304244 165356
rect 303926 165042 303930 165352
rect 303930 165042 304240 165352
rect 304240 165042 304244 165352
rect 303926 165038 304244 165042
rect -2006 163722 -1806 163922
rect 303926 162352 304244 162356
rect 303926 162042 303930 162352
rect 303930 162042 304240 162352
rect 304240 162042 304244 162352
rect 303926 162038 304244 162042
rect -2006 160722 -1806 160922
rect 303926 159352 304244 159356
rect 303926 159042 303930 159352
rect 303930 159042 304240 159352
rect 304240 159042 304244 159352
rect 303926 159038 304244 159042
rect -2006 157722 -1806 157922
rect 303926 156352 304244 156356
rect 303926 156042 303930 156352
rect 303930 156042 304240 156352
rect 304240 156042 304244 156352
rect 303926 156038 304244 156042
rect -2006 154722 -1806 154922
rect 303926 153352 304244 153356
rect 303926 153042 303930 153352
rect 303930 153042 304240 153352
rect 304240 153042 304244 153352
rect 303926 153038 304244 153042
rect -2006 151722 -1806 151922
rect 303926 150352 304244 150356
rect 303926 150042 303930 150352
rect 303930 150042 304240 150352
rect 304240 150042 304244 150352
rect 303926 150038 304244 150042
rect -2006 148722 -1806 148922
rect 303926 147352 304244 147356
rect 303926 147042 303930 147352
rect 303930 147042 304240 147352
rect 304240 147042 304244 147352
rect 303926 147038 304244 147042
rect -2006 145722 -1806 145922
rect 303926 144352 304244 144356
rect 303926 144042 303930 144352
rect 303930 144042 304240 144352
rect 304240 144042 304244 144352
rect 303926 144038 304244 144042
rect -2006 142722 -1806 142922
rect 303926 141352 304244 141356
rect 303926 141042 303930 141352
rect 303930 141042 304240 141352
rect 304240 141042 304244 141352
rect 303926 141038 304244 141042
rect -2006 139722 -1806 139922
rect 303926 138352 304244 138356
rect 303926 138042 303930 138352
rect 303930 138042 304240 138352
rect 304240 138042 304244 138352
rect 303926 138038 304244 138042
rect -2006 136722 -1806 136922
rect 303926 135352 304244 135356
rect 303926 135042 303930 135352
rect 303930 135042 304240 135352
rect 304240 135042 304244 135352
rect 303926 135038 304244 135042
rect -2006 133722 -1806 133922
rect 303926 132352 304244 132356
rect 303926 132042 303930 132352
rect 303930 132042 304240 132352
rect 304240 132042 304244 132352
rect 303926 132038 304244 132042
rect -2006 130722 -1806 130922
rect 303926 129352 304244 129356
rect 303926 129042 303930 129352
rect 303930 129042 304240 129352
rect 304240 129042 304244 129352
rect 303926 129038 304244 129042
rect -2006 127722 -1806 127922
rect 303926 126352 304244 126356
rect 303926 126042 303930 126352
rect 303930 126042 304240 126352
rect 304240 126042 304244 126352
rect 303926 126038 304244 126042
rect -2006 124722 -1806 124922
rect 303926 123352 304244 123356
rect 303926 123042 303930 123352
rect 303930 123042 304240 123352
rect 304240 123042 304244 123352
rect 303926 123038 304244 123042
rect -2006 121722 -1806 121922
rect 303926 120352 304244 120356
rect 303926 120042 303930 120352
rect 303930 120042 304240 120352
rect 304240 120042 304244 120352
rect 303926 120038 304244 120042
rect -2006 118722 -1806 118922
rect 303926 117352 304244 117356
rect 303926 117042 303930 117352
rect 303930 117042 304240 117352
rect 304240 117042 304244 117352
rect 303926 117038 304244 117042
rect -2006 115722 -1806 115922
rect 303926 114352 304244 114356
rect 303926 114042 303930 114352
rect 303930 114042 304240 114352
rect 304240 114042 304244 114352
rect 303926 114038 304244 114042
rect -2006 112722 -1806 112922
rect 303926 111352 304244 111356
rect 303926 111042 303930 111352
rect 303930 111042 304240 111352
rect 304240 111042 304244 111352
rect 303926 111038 304244 111042
rect -2006 109722 -1806 109922
rect 303926 108352 304244 108356
rect 303926 108042 303930 108352
rect 303930 108042 304240 108352
rect 304240 108042 304244 108352
rect 303926 108038 304244 108042
rect -2006 106722 -1806 106922
rect 303926 105352 304244 105356
rect 303926 105042 303930 105352
rect 303930 105042 304240 105352
rect 304240 105042 304244 105352
rect 303926 105038 304244 105042
rect -2006 103722 -1806 103922
rect 303926 102352 304244 102356
rect 303926 102042 303930 102352
rect 303930 102042 304240 102352
rect 304240 102042 304244 102352
rect 303926 102038 304244 102042
rect -2006 100722 -1806 100922
rect 303926 99352 304244 99356
rect 303926 99042 303930 99352
rect 303930 99042 304240 99352
rect 304240 99042 304244 99352
rect 303926 99038 304244 99042
rect -2006 97722 -1806 97922
rect 303926 96352 304244 96356
rect 303926 96042 303930 96352
rect 303930 96042 304240 96352
rect 304240 96042 304244 96352
rect 303926 96038 304244 96042
rect -2006 94722 -1806 94922
rect 303926 93352 304244 93356
rect 303926 93042 303930 93352
rect 303930 93042 304240 93352
rect 304240 93042 304244 93352
rect 303926 93038 304244 93042
rect -2006 91722 -1806 91922
rect 303926 90352 304244 90356
rect 303926 90042 303930 90352
rect 303930 90042 304240 90352
rect 304240 90042 304244 90352
rect 303926 90038 304244 90042
rect -2006 88722 -1806 88922
rect 303926 87352 304244 87356
rect 303926 87042 303930 87352
rect 303930 87042 304240 87352
rect 304240 87042 304244 87352
rect 303926 87038 304244 87042
rect -2006 85722 -1806 85922
rect 303926 84352 304244 84356
rect 303926 84042 303930 84352
rect 303930 84042 304240 84352
rect 304240 84042 304244 84352
rect 303926 84038 304244 84042
rect -2006 82722 -1806 82922
rect 303926 81352 304244 81356
rect 303926 81042 303930 81352
rect 303930 81042 304240 81352
rect 304240 81042 304244 81352
rect 303926 81038 304244 81042
rect -2006 79722 -1806 79922
rect 303926 78352 304244 78356
rect 303926 78042 303930 78352
rect 303930 78042 304240 78352
rect 304240 78042 304244 78352
rect 303926 78038 304244 78042
rect -2006 76722 -1806 76922
rect 303926 75352 304244 75356
rect 303926 75042 303930 75352
rect 303930 75042 304240 75352
rect 304240 75042 304244 75352
rect 303926 75038 304244 75042
rect -2006 73722 -1806 73922
rect 303926 72352 304244 72356
rect 303926 72042 303930 72352
rect 303930 72042 304240 72352
rect 304240 72042 304244 72352
rect 303926 72038 304244 72042
rect -2006 70722 -1806 70922
rect 303926 69352 304244 69356
rect 303926 69042 303930 69352
rect 303930 69042 304240 69352
rect 304240 69042 304244 69352
rect 303926 69038 304244 69042
rect -2006 67722 -1806 67922
rect 303926 66352 304244 66356
rect 303926 66042 303930 66352
rect 303930 66042 304240 66352
rect 304240 66042 304244 66352
rect 303926 66038 304244 66042
rect -2006 64722 -1806 64922
rect 303926 63352 304244 63356
rect 303926 63042 303930 63352
rect 303930 63042 304240 63352
rect 304240 63042 304244 63352
rect 303926 63038 304244 63042
rect -2006 61722 -1806 61922
rect 303926 60352 304244 60356
rect 303926 60042 303930 60352
rect 303930 60042 304240 60352
rect 304240 60042 304244 60352
rect 303926 60038 304244 60042
rect -2006 58722 -1806 58922
rect 303926 57352 304244 57356
rect 303926 57042 303930 57352
rect 303930 57042 304240 57352
rect 304240 57042 304244 57352
rect 303926 57038 304244 57042
rect -2006 55722 -1806 55922
rect 303926 54352 304244 54356
rect 303926 54042 303930 54352
rect 303930 54042 304240 54352
rect 304240 54042 304244 54352
rect 303926 54038 304244 54042
rect -2006 52722 -1806 52922
rect 303926 51352 304244 51356
rect 303926 51042 303930 51352
rect 303930 51042 304240 51352
rect 304240 51042 304244 51352
rect 303926 51038 304244 51042
rect -2006 49722 -1806 49922
rect 303926 48352 304244 48356
rect 303926 48042 303930 48352
rect 303930 48042 304240 48352
rect 304240 48042 304244 48352
rect 303926 48038 304244 48042
rect -2006 46722 -1806 46922
rect 303926 45352 304244 45356
rect 303926 45042 303930 45352
rect 303930 45042 304240 45352
rect 304240 45042 304244 45352
rect 303926 45038 304244 45042
rect -2006 43722 -1806 43922
rect 303926 42352 304244 42356
rect 303926 42042 303930 42352
rect 303930 42042 304240 42352
rect 304240 42042 304244 42352
rect 303926 42038 304244 42042
rect -2006 40722 -1806 40922
rect 303926 39352 304244 39356
rect 303926 39042 303930 39352
rect 303930 39042 304240 39352
rect 304240 39042 304244 39352
rect 303926 39038 304244 39042
rect -2006 37722 -1806 37922
rect 303926 36352 304244 36356
rect 303926 36042 303930 36352
rect 303930 36042 304240 36352
rect 304240 36042 304244 36352
rect 303926 36038 304244 36042
rect -2006 34722 -1806 34922
rect 303926 33352 304244 33356
rect 303926 33042 303930 33352
rect 303930 33042 304240 33352
rect 304240 33042 304244 33352
rect 303926 33038 304244 33042
rect -2006 31722 -1806 31922
rect 303926 30352 304244 30356
rect 303926 30042 303930 30352
rect 303930 30042 304240 30352
rect 304240 30042 304244 30352
rect 303926 30038 304244 30042
rect -2006 28722 -1806 28922
rect 303926 27352 304244 27356
rect 303926 27042 303930 27352
rect 303930 27042 304240 27352
rect 304240 27042 304244 27352
rect 303926 27038 304244 27042
rect -2006 25722 -1806 25922
rect 303926 24352 304244 24356
rect 303926 24042 303930 24352
rect 303930 24042 304240 24352
rect 304240 24042 304244 24352
rect 303926 24038 304244 24042
rect -2006 22722 -1806 22922
rect 303926 21352 304244 21356
rect 303926 21042 303930 21352
rect 303930 21042 304240 21352
rect 304240 21042 304244 21352
rect 303926 21038 304244 21042
rect 19870 19188 20088 19192
rect 19870 18978 19874 19188
rect 19874 18978 20084 19188
rect 20084 18978 20088 19188
rect 19870 18974 20088 18978
rect 5328 18780 5546 18784
rect 5328 18570 5332 18780
rect 5332 18570 5542 18780
rect 5542 18570 5546 18780
rect 5328 18566 5546 18570
rect 7482 18886 7700 18890
rect 7482 18676 7486 18886
rect 7486 18676 7696 18886
rect 7696 18676 7700 18886
rect 7482 18672 7700 18676
rect 10712 18830 10930 18834
rect 10712 18620 10716 18830
rect 10716 18620 10926 18830
rect 10926 18620 10930 18830
rect 10712 18616 10930 18620
rect 13802 18924 14020 18928
rect 13802 18714 13806 18924
rect 13806 18714 14016 18924
rect 14016 18714 14020 18924
rect 13802 18710 14020 18714
rect 16912 18812 17130 18816
rect 16912 18602 16916 18812
rect 16916 18602 17126 18812
rect 17126 18602 17130 18812
rect 16912 18598 17130 18602
rect 25944 19006 26162 19010
rect 25944 18796 25948 19006
rect 25948 18796 26158 19006
rect 26158 18796 26162 19006
rect 25944 18792 26162 18796
rect 29084 18842 29302 19060
rect 32328 18982 32546 18986
rect 32328 18772 32332 18982
rect 32332 18772 32542 18982
rect 32542 18772 32546 18982
rect 32328 18768 32546 18772
rect 35328 19050 35546 19054
rect 35328 18840 35332 19050
rect 35332 18840 35542 19050
rect 35542 18840 35546 19050
rect 35328 18836 35546 18840
rect 38328 19214 38546 19218
rect 38328 19004 38332 19214
rect 38332 19004 38542 19214
rect 38542 19004 38546 19214
rect 38328 19000 38546 19004
rect 2328 18434 2546 18438
rect 2328 18224 2332 18434
rect 2332 18224 2542 18434
rect 2542 18224 2546 18434
rect 2328 18220 2546 18224
rect 22898 18654 23116 18658
rect 22898 18444 22902 18654
rect 22902 18444 23112 18654
rect 23112 18444 23116 18654
rect 22898 18440 23116 18444
rect 41328 18868 41546 18872
rect 41328 18658 41332 18868
rect 41332 18658 41542 18868
rect 41542 18658 41546 18868
rect 41328 18654 41546 18658
rect 44328 18918 44546 18922
rect 44328 18708 44332 18918
rect 44332 18708 44542 18918
rect 44542 18708 44546 18918
rect 44328 18704 44546 18708
rect 47328 19126 47546 19130
rect 47328 18916 47332 19126
rect 47332 18916 47542 19126
rect 47542 18916 47546 19126
rect 47328 18912 47546 18916
rect 50516 19006 50734 19010
rect 50516 18796 50520 19006
rect 50520 18796 50730 19006
rect 50730 18796 50734 19006
rect 50516 18792 50734 18796
rect 53538 19038 53756 19042
rect 53538 18828 53542 19038
rect 53542 18828 53752 19038
rect 53752 18828 53756 19038
rect 53538 18824 53756 18828
rect 56616 19158 56834 19162
rect 56616 18948 56620 19158
rect 56620 18948 56830 19158
rect 56830 18948 56834 19158
rect 56616 18944 56834 18948
rect 59630 18862 59848 18866
rect 59630 18652 59634 18862
rect 59634 18652 59844 18862
rect 59844 18652 59848 18862
rect 59630 18648 59848 18652
rect 62632 18786 62850 18790
rect 62632 18576 62636 18786
rect 62636 18576 62846 18786
rect 62846 18576 62850 18786
rect 62632 18572 62850 18576
rect 65742 18876 65960 18880
rect 65742 18666 65746 18876
rect 65746 18666 65956 18876
rect 65956 18666 65960 18876
rect 65742 18662 65960 18666
rect 68328 18734 68546 18952
rect 71928 18842 72146 19060
rect 75078 19026 75296 19030
rect 75078 18816 75082 19026
rect 75082 18816 75292 19026
rect 75292 18816 75296 19026
rect 75078 18812 75296 18816
rect 81190 18706 81408 18904
rect 81190 18686 81194 18706
rect 81194 18686 81404 18706
rect 81404 18686 81408 18706
rect 90412 18832 90630 18836
rect 90412 18622 90416 18832
rect 90416 18622 90626 18832
rect 90626 18622 90630 18832
rect 90412 18618 90630 18622
rect 93556 18788 93774 18792
rect 93556 18578 93560 18788
rect 93560 18578 93770 18788
rect 93770 18578 93774 18788
rect 93556 18574 93774 18578
rect 96454 18870 96672 18874
rect 96454 18660 96458 18870
rect 96458 18660 96668 18870
rect 96668 18660 96672 18870
rect 96454 18656 96672 18660
rect 108902 19028 109120 19032
rect 108902 18818 108906 19028
rect 108906 18818 109116 19028
rect 109116 18818 109120 19028
rect 108902 18814 109120 18818
rect 102712 18736 102930 18740
rect 102712 18526 102716 18736
rect 102716 18526 102926 18736
rect 102926 18526 102930 18736
rect 102712 18522 102930 18526
rect 78098 18088 78316 18306
rect 84274 18184 84492 18402
rect -6204 17746 -6198 17942
rect -6198 17746 -5998 17942
rect -5998 17746 -5994 17942
rect -6204 17742 -5994 17746
rect 87336 18310 87554 18314
rect 87336 18100 87340 18310
rect 87340 18100 87550 18310
rect 87550 18100 87554 18310
rect 87336 18096 87554 18100
rect 99598 18496 99816 18500
rect 99598 18286 99602 18496
rect 99602 18286 99812 18496
rect 99812 18286 99816 18496
rect 99598 18282 99816 18286
rect 105676 18750 105894 18754
rect 105676 18540 105680 18750
rect 105680 18540 105890 18750
rect 105890 18540 105894 18750
rect 105676 18536 105894 18540
rect 111948 18930 112166 18934
rect 111948 18720 111952 18930
rect 111952 18720 112162 18930
rect 112162 18720 112166 18930
rect 111948 18716 112166 18720
rect 114954 18980 115172 18984
rect 114954 18770 114958 18980
rect 114958 18770 115168 18980
rect 115168 18770 115172 18980
rect 114954 18766 115172 18770
rect 117968 18972 118186 18976
rect 117968 18762 117972 18972
rect 117972 18762 118182 18972
rect 118182 18762 118186 18972
rect 117968 18758 118186 18762
rect 121150 18860 121368 18864
rect 121150 18650 121154 18860
rect 121154 18650 121364 18860
rect 121364 18650 121368 18860
rect 121150 18646 121368 18650
rect 124118 18632 124336 18850
rect 127242 18938 127460 18942
rect 127242 18728 127246 18938
rect 127246 18728 127456 18938
rect 127456 18728 127460 18938
rect 127242 18724 127460 18728
rect 130250 18808 130468 18812
rect 130250 18598 130254 18808
rect 130254 18598 130464 18808
rect 130464 18598 130468 18808
rect 130250 18594 130468 18598
rect 133412 18648 133630 18866
rect 139552 18596 139770 18600
rect 139552 18386 139556 18596
rect 139556 18386 139766 18596
rect 139766 18386 139770 18596
rect 139552 18382 139770 18386
rect 142600 18664 142818 18668
rect 142600 18454 142604 18664
rect 142604 18454 142814 18664
rect 142814 18454 142818 18664
rect 142600 18450 142818 18454
rect 145578 18838 145796 18842
rect 145578 18628 145582 18838
rect 145582 18628 145792 18838
rect 145792 18628 145796 18838
rect 145578 18624 145796 18628
rect 148754 18838 148972 18842
rect 148754 18628 148758 18838
rect 148758 18628 148968 18838
rect 148968 18628 148972 18838
rect 148754 18624 148972 18628
rect 151772 18770 151990 18774
rect 151772 18560 151776 18770
rect 151776 18560 151986 18770
rect 151986 18560 151990 18770
rect 151772 18556 151990 18560
rect 154792 18854 155010 18858
rect 154792 18644 154796 18854
rect 154796 18644 155006 18854
rect 155006 18644 155010 18854
rect 154792 18640 155010 18644
rect 157844 18992 158062 18996
rect 157844 18782 157848 18992
rect 157848 18782 158058 18992
rect 158058 18782 158062 18992
rect 157844 18778 158062 18782
rect 174366 19130 174584 19134
rect 174366 18920 174370 19130
rect 174370 18920 174580 19130
rect 174580 18920 174584 19130
rect 174366 18916 174584 18920
rect 160886 18754 161104 18758
rect 160886 18544 160890 18754
rect 160890 18544 161100 18754
rect 161100 18544 161104 18754
rect 160886 18540 161104 18544
rect 176328 18808 176546 18812
rect 176328 18598 176332 18808
rect 176332 18598 176542 18808
rect 176542 18598 176546 18808
rect 176328 18594 176546 18598
rect 229658 18934 229876 18938
rect 229658 18724 229662 18934
rect 229662 18724 229872 18934
rect 229872 18724 229876 18934
rect 229658 18720 229876 18724
rect 290328 18950 290546 18954
rect 290328 18740 290332 18950
rect 290332 18740 290542 18950
rect 290542 18740 290546 18950
rect 290328 18736 290546 18740
rect 305386 19094 305604 19098
rect 305386 18884 305390 19094
rect 305390 18884 305600 19094
rect 305600 18884 305604 19094
rect 305386 18880 305604 18884
rect 136468 18236 136686 18240
rect 136468 18026 136472 18236
rect 136472 18026 136682 18236
rect 136682 18026 136686 18236
rect 136468 18022 136686 18026
rect 163238 18454 163456 18458
rect 163238 18244 163242 18454
rect 163242 18244 163452 18454
rect 163452 18244 163456 18454
rect 163238 18240 163456 18244
rect 173082 18484 173300 18488
rect 173082 18274 173086 18484
rect 173086 18274 173296 18484
rect 173296 18274 173300 18484
rect 173082 18270 173300 18274
rect 206328 18450 206546 18454
rect 206328 18240 206332 18450
rect 206332 18240 206542 18450
rect 206542 18240 206546 18450
rect 206328 18236 206546 18240
rect 215328 18558 215546 18562
rect 215328 18348 215332 18558
rect 215332 18348 215542 18558
rect 215542 18348 215546 18558
rect 215328 18344 215546 18348
rect 233328 18684 233546 18688
rect 233328 18474 233332 18684
rect 233332 18474 233542 18684
rect 233542 18474 233546 18684
rect 233328 18470 233546 18474
rect 227194 18424 227412 18428
rect 227194 18214 227198 18424
rect 227198 18214 227408 18424
rect 227408 18214 227412 18424
rect 227194 18210 227412 18214
rect 241672 18530 241890 18534
rect 241672 18320 241676 18530
rect 241676 18320 241886 18530
rect 241886 18320 241890 18530
rect 241672 18316 241890 18320
rect 242328 18566 242546 18570
rect 242328 18356 242332 18566
rect 242332 18356 242542 18566
rect 242542 18356 242546 18566
rect 242328 18352 242546 18356
rect 165928 18170 166146 18174
rect 165928 17960 165932 18170
rect 165932 17960 166142 18170
rect 166142 17960 166146 18170
rect 165928 17956 166146 17960
rect 182474 17854 182692 17858
rect 182474 17644 182478 17854
rect 182478 17644 182688 17854
rect 182688 17644 182692 17854
rect 182474 17640 182692 17644
rect 185328 18032 185546 18036
rect 185328 17822 185332 18032
rect 185332 17822 185542 18032
rect 185542 17822 185546 18032
rect 185328 17818 185546 17822
rect 196794 17924 197012 17928
rect 196794 17714 196798 17924
rect 196798 17714 197008 17924
rect 197008 17714 197012 17924
rect 196794 17710 197012 17714
rect 200916 17952 201134 17956
rect 200916 17742 200920 17952
rect 200920 17742 201130 17952
rect 201130 17742 201134 17952
rect 200916 17738 201134 17742
rect 213156 18094 213374 18098
rect 213156 17884 213160 18094
rect 213160 17884 213370 18094
rect 213370 17884 213374 18094
rect 213156 17880 213374 17884
rect 234650 18298 234868 18302
rect 234650 18088 234654 18298
rect 234654 18088 234864 18298
rect 234864 18088 234868 18298
rect 234650 18084 234868 18088
rect 253926 18504 254144 18508
rect 253926 18294 253930 18504
rect 253930 18294 254140 18504
rect 254140 18294 254144 18504
rect 253926 18290 254144 18294
rect 254328 18696 254546 18700
rect 254328 18486 254332 18696
rect 254332 18486 254542 18696
rect 254542 18486 254546 18696
rect 254328 18482 254546 18486
rect 269032 18556 269250 18560
rect 269032 18346 269036 18556
rect 269036 18346 269246 18556
rect 269246 18346 269250 18556
rect 269032 18342 269250 18346
rect 279676 18694 279894 18698
rect 279676 18484 279680 18694
rect 279680 18484 279890 18694
rect 279890 18484 279894 18694
rect 279676 18480 279894 18484
rect 240916 18010 241134 18014
rect 240916 17800 240920 18010
rect 240920 17800 241130 18010
rect 241130 17800 241134 18010
rect 240916 17796 241134 17800
rect 261044 18120 261262 18124
rect 261044 17910 261048 18120
rect 261048 17910 261258 18120
rect 261258 17910 261262 18120
rect 261044 17906 261262 17910
rect 269328 18264 269546 18268
rect 269328 18054 269332 18264
rect 269332 18054 269542 18264
rect 269542 18054 269546 18264
rect 269328 18050 269546 18054
rect 278878 18202 279096 18206
rect 278878 17992 278882 18202
rect 278882 17992 279092 18202
rect 279092 17992 279096 18202
rect 278878 17988 279096 17992
rect 168864 17416 169082 17420
rect 168864 17206 168868 17416
rect 168868 17206 169078 17416
rect 169078 17206 169082 17416
rect 168864 17202 169082 17206
rect 188328 17654 188546 17658
rect 188328 17444 188332 17654
rect 188332 17444 188542 17654
rect 188542 17444 188546 17654
rect 188328 17440 188546 17444
rect 207000 17746 207218 17750
rect 207000 17536 207004 17746
rect 207004 17536 207214 17746
rect 207214 17536 207218 17746
rect 207000 17532 207218 17536
rect 221328 17706 221546 17710
rect 221328 17496 221332 17706
rect 221332 17496 221542 17706
rect 221542 17496 221546 17706
rect 221328 17492 221546 17496
rect 249668 17856 249886 17860
rect 249668 17646 249672 17856
rect 249672 17646 249882 17856
rect 249882 17646 249886 17856
rect 249668 17642 249886 17646
rect 265870 17958 266088 17962
rect 265870 17748 265874 17958
rect 265874 17748 266084 17958
rect 266084 17748 266088 17958
rect 265870 17744 266088 17748
rect 284328 18132 284546 18136
rect 284328 17922 284332 18132
rect 284332 17922 284542 18132
rect 284542 17922 284546 18132
rect 284328 17918 284546 17922
rect 292408 18222 292626 18226
rect 292408 18012 292412 18222
rect 292412 18012 292622 18222
rect 292622 18012 292626 18222
rect 292408 18008 292626 18012
rect 302946 18469 303268 18717
rect 302946 18395 303268 18469
rect 277694 17578 277912 17582
rect 277694 17368 277698 17578
rect 277698 17368 277908 17578
rect 277908 17368 277912 17578
rect 277694 17364 277912 17368
rect 286930 17508 287148 17512
rect 286930 17298 286934 17508
rect 286934 17298 287144 17508
rect 287144 17298 287148 17508
rect 286930 17294 287148 17298
rect 299258 17718 299476 17722
rect 299258 17508 299262 17718
rect 299262 17508 299472 17718
rect 299472 17508 299476 17718
rect 299258 17504 299476 17508
rect 184010 17148 184228 17152
rect 184010 16938 184014 17148
rect 184014 16938 184224 17148
rect 184224 16938 184228 17148
rect 184010 16934 184228 16938
rect 213904 17264 214122 17268
rect 213904 17054 213908 17264
rect 213908 17054 214118 17264
rect 214118 17054 214122 17264
rect 213904 17050 214122 17054
rect 193466 17014 193684 17018
rect 193466 16804 193470 17014
rect 193470 16804 193680 17014
rect 193680 16804 193684 17014
rect 193466 16800 193684 16804
rect 220688 17224 220906 17228
rect 220688 17014 220692 17224
rect 220692 17014 220902 17224
rect 220902 17014 220906 17224
rect 220688 17010 220906 17014
rect 202004 16890 202222 16894
rect 202004 16680 202008 16890
rect 202008 16680 202218 16890
rect 202218 16680 202222 16890
rect 202004 16676 202222 16680
rect 248712 17072 248930 17076
rect 248712 16862 248716 17072
rect 248716 16862 248926 17072
rect 248926 16862 248930 17072
rect 248712 16858 248930 16862
rect 260054 17242 260272 17246
rect 260054 17032 260058 17242
rect 260058 17032 260268 17242
rect 260268 17032 260272 17242
rect 260054 17028 260272 17032
rect 300252 17100 300470 17104
rect 300252 16890 300256 17100
rect 300256 16890 300466 17100
rect 300466 16890 300470 17100
rect 300252 16886 300470 16890
rect 302942 16094 302946 16410
rect 302946 16094 303268 16410
rect 303268 16094 303274 16410
rect 302942 16088 303274 16094
rect 102 15388 108 15582
rect 108 15388 308 15582
rect 308 15388 312 15582
rect 102 15382 312 15388
<< metal4 >>
rect -7596 325866 -762 325976
rect -5202 322052 -1206 322076
rect -5202 321780 -1502 322052
rect -1230 321780 -1206 322052
rect -5202 321760 -1206 321780
rect -5202 321756 -1526 321760
rect -872 320928 -762 325866
rect 303888 321356 304300 322140
rect 303888 321038 303926 321356
rect 304244 321038 304300 321356
rect -5974 319800 -3762 320120
rect -2066 319922 -1726 319998
rect -2674 319723 -2006 319922
rect -2674 319722 -2005 319723
rect -1806 319722 -1726 319922
rect -2066 319684 -1726 319722
rect -5202 319052 -1206 319076
rect -5202 318780 -1502 319052
rect -1230 318780 -1206 319052
rect -5202 318760 -1206 318780
rect -5202 318756 -1526 318760
rect 303888 318356 304300 321038
rect 303888 318038 303926 318356
rect 304244 318038 304300 318356
rect -5974 316800 -3762 317120
rect -2038 316922 -1776 317004
rect -2674 316722 -2006 316922
rect -1806 316722 -1776 316922
rect -2038 316694 -1776 316722
rect -5202 316052 -1206 316076
rect -5202 315780 -1502 316052
rect -1230 315780 -1206 316052
rect -5202 315760 -1206 315780
rect -5202 315756 -1526 315760
rect 303888 315356 304300 318038
rect 303888 315038 303926 315356
rect 304244 315038 304300 315356
rect -5974 313800 -3762 314120
rect -2050 313922 -1774 313944
rect -2674 313722 -2006 313922
rect -1806 313722 -1774 313922
rect -2050 313672 -1774 313722
rect -5202 313052 -1206 313076
rect -5202 312780 -1502 313052
rect -1230 312780 -1206 313052
rect -5202 312760 -1206 312780
rect -5202 312756 -1526 312760
rect 303888 312356 304300 315038
rect 303888 312038 303926 312356
rect 304244 312038 304300 312356
rect -5974 310800 -3762 311120
rect -2026 310922 -1780 310940
rect -2674 310722 -2006 310922
rect -1806 310722 -1780 310922
rect -2026 310708 -1780 310722
rect -5202 310052 -1206 310076
rect -5202 309780 -1502 310052
rect -1230 309780 -1206 310052
rect -5202 309760 -1206 309780
rect -5202 309756 -1526 309760
rect 303888 309356 304300 312038
rect 303888 309038 303926 309356
rect 304244 309038 304300 309356
rect -5974 307800 -3762 308120
rect -2010 307922 -1804 307930
rect -2674 307722 -2006 307922
rect -1806 307722 -1804 307922
rect -2010 307714 -1804 307722
rect -5202 307052 -1206 307076
rect -5202 306780 -1502 307052
rect -1230 306780 -1206 307052
rect -5202 306760 -1206 306780
rect -5202 306756 -1526 306760
rect 303888 306356 304300 309038
rect 303888 306038 303926 306356
rect 304244 306038 304300 306356
rect -5974 304800 -3762 305120
rect -2014 304922 -1788 304934
rect -2674 304722 -2006 304922
rect -1806 304722 -1788 304922
rect -2014 304700 -1788 304722
rect -5202 304052 -1206 304076
rect -5202 303780 -1502 304052
rect -1230 303780 -1206 304052
rect -5202 303760 -1206 303780
rect -5202 303756 -1526 303760
rect 303888 303356 304300 306038
rect 303888 303038 303926 303356
rect 304244 303038 304300 303356
rect -5974 301800 -3762 302120
rect -2018 301922 -1790 301926
rect -2674 301722 -2006 301922
rect -1806 301722 -1790 301922
rect -2018 301712 -1790 301722
rect -5202 301052 -1206 301076
rect -5202 300780 -1502 301052
rect -1230 300780 -1206 301052
rect -5202 300760 -1206 300780
rect -5202 300756 -1526 300760
rect 303888 300356 304300 303038
rect 303888 300038 303926 300356
rect 304244 300038 304300 300356
rect -5974 298800 -3762 299120
rect -2018 298922 -1800 298954
rect -2674 298722 -2006 298922
rect -1806 298722 -1800 298922
rect -2018 298688 -1800 298722
rect -5202 298052 -1206 298076
rect -5202 297780 -1502 298052
rect -1230 297780 -1206 298052
rect -5202 297760 -1206 297780
rect -5202 297756 -1526 297760
rect 303888 297356 304300 300038
rect 303888 297038 303926 297356
rect 304244 297038 304300 297356
rect -5974 295800 -3762 296120
rect -2014 295922 -1792 295934
rect -2674 295722 -2006 295922
rect -1806 295722 -1792 295922
rect -2014 295708 -1792 295722
rect -5202 295052 -1206 295076
rect -5202 294780 -1502 295052
rect -1230 294780 -1206 295052
rect -5202 294760 -1206 294780
rect -5202 294756 -1526 294760
rect 303888 294356 304300 297038
rect 303888 294038 303926 294356
rect 304244 294038 304300 294356
rect -5974 292800 -3762 293120
rect -2014 292922 -1800 292932
rect -2674 292722 -2006 292922
rect -1806 292722 -1800 292922
rect -2014 292710 -1800 292722
rect -5202 292052 -1206 292076
rect -5202 291780 -1502 292052
rect -1230 291780 -1206 292052
rect -5202 291760 -1206 291780
rect -5202 291756 -1526 291760
rect 303888 291356 304300 294038
rect 303888 291038 303926 291356
rect 304244 291038 304300 291356
rect -5974 289800 -3762 290120
rect -2024 289922 -1788 289950
rect -2674 289722 -2006 289922
rect -1806 289722 -1788 289922
rect -2024 289694 -1788 289722
rect -5202 289052 -1206 289076
rect -5202 288780 -1502 289052
rect -1230 288780 -1206 289052
rect -5202 288760 -1206 288780
rect -5202 288756 -1526 288760
rect 303888 288356 304300 291038
rect 303888 288038 303926 288356
rect 304244 288038 304300 288356
rect -5974 286800 -3762 287120
rect -2016 286922 -1786 286930
rect -2674 286722 -2006 286922
rect -1806 286722 -1786 286922
rect -2016 286708 -1786 286722
rect -5202 286052 -1206 286076
rect -5202 285780 -1502 286052
rect -1230 285780 -1206 286052
rect -5202 285760 -1206 285780
rect -5202 285756 -1526 285760
rect 303888 285356 304300 288038
rect 303888 285038 303926 285356
rect 304244 285038 304300 285356
rect -5974 283800 -3762 284120
rect -2016 283922 -1786 283930
rect -2674 283722 -2006 283922
rect -1806 283722 -1786 283922
rect -2016 283708 -1786 283722
rect -5202 283052 -1206 283076
rect -5202 282780 -1502 283052
rect -1230 282780 -1206 283052
rect -5202 282760 -1206 282780
rect -5202 282756 -1526 282760
rect 303888 282356 304300 285038
rect 303888 282038 303926 282356
rect 304244 282038 304300 282356
rect -5974 280800 -3762 281120
rect -2016 280922 -1786 280930
rect -2674 280722 -2006 280922
rect -1806 280722 -1786 280922
rect -2016 280708 -1786 280722
rect -5202 280052 -1206 280076
rect -5202 279780 -1502 280052
rect -1230 279780 -1206 280052
rect -5202 279760 -1206 279780
rect -5202 279756 -1526 279760
rect 303888 279356 304300 282038
rect 303888 279038 303926 279356
rect 304244 279038 304300 279356
rect -5974 277800 -3762 278120
rect -2016 277922 -1786 277930
rect -2674 277722 -2006 277922
rect -1806 277722 -1786 277922
rect -2016 277708 -1786 277722
rect -5202 277052 -1206 277076
rect -5202 276780 -1502 277052
rect -1230 276780 -1206 277052
rect -5202 276760 -1206 276780
rect -5202 276756 -1526 276760
rect 303888 276356 304300 279038
rect 303888 276038 303926 276356
rect 304244 276038 304300 276356
rect -5974 274800 -3762 275120
rect -2016 274922 -1786 274930
rect -2674 274722 -2006 274922
rect -1806 274722 -1786 274922
rect -2016 274708 -1786 274722
rect -5202 274052 -1206 274076
rect -5202 273780 -1502 274052
rect -1230 273780 -1206 274052
rect -5202 273760 -1206 273780
rect -5202 273756 -1526 273760
rect 303888 273356 304300 276038
rect 303888 273038 303926 273356
rect 304244 273038 304300 273356
rect -5974 271800 -3762 272120
rect -2016 271922 -1786 271930
rect -2674 271722 -2006 271922
rect -1806 271722 -1786 271922
rect -2016 271708 -1786 271722
rect -5202 271052 -1206 271076
rect -5202 270780 -1502 271052
rect -1230 270780 -1206 271052
rect -5202 270760 -1206 270780
rect -5202 270756 -1526 270760
rect 303888 270356 304300 273038
rect 303888 270038 303926 270356
rect 304244 270038 304300 270356
rect -5974 268800 -3762 269120
rect -2016 268922 -1786 268930
rect -2674 268722 -2006 268922
rect -1806 268722 -1786 268922
rect -2016 268708 -1786 268722
rect -5202 268052 -1206 268076
rect -5202 267780 -1502 268052
rect -1230 267780 -1206 268052
rect -5202 267760 -1206 267780
rect -5202 267756 -1526 267760
rect 303888 267356 304300 270038
rect 303888 267038 303926 267356
rect 304244 267038 304300 267356
rect -5974 265800 -3762 266120
rect -2016 265922 -1786 265930
rect -2674 265722 -2006 265922
rect -1806 265722 -1786 265922
rect -2016 265708 -1786 265722
rect -5202 265052 -1206 265076
rect -5202 264780 -1502 265052
rect -1230 264780 -1206 265052
rect -5202 264760 -1206 264780
rect -5202 264756 -1526 264760
rect 303888 264356 304300 267038
rect 303888 264038 303926 264356
rect 304244 264038 304300 264356
rect -5974 262800 -3762 263120
rect -2016 262922 -1786 262930
rect -2674 262722 -2006 262922
rect -1806 262722 -1786 262922
rect -2016 262708 -1786 262722
rect -5202 262052 -1206 262076
rect -5202 261780 -1502 262052
rect -1230 261780 -1206 262052
rect -5202 261760 -1206 261780
rect -5202 261756 -1526 261760
rect 303888 261356 304300 264038
rect 303888 261038 303926 261356
rect 304244 261038 304300 261356
rect -5974 259800 -3762 260120
rect -2016 259922 -1786 259930
rect -2674 259722 -2006 259922
rect -1806 259722 -1786 259922
rect -2016 259708 -1786 259722
rect -5202 259052 -1206 259076
rect -5202 258780 -1502 259052
rect -1230 258780 -1206 259052
rect -5202 258760 -1206 258780
rect -5202 258756 -1526 258760
rect 303888 258356 304300 261038
rect 303888 258038 303926 258356
rect 304244 258038 304300 258356
rect -5974 256800 -3762 257120
rect -2016 256922 -1786 256930
rect -2674 256722 -2006 256922
rect -1806 256722 -1786 256922
rect -2016 256708 -1786 256722
rect -5202 256052 -1206 256076
rect -5202 255780 -1502 256052
rect -1230 255780 -1206 256052
rect -5202 255760 -1206 255780
rect -5202 255756 -1526 255760
rect 303888 255356 304300 258038
rect 303888 255038 303926 255356
rect 304244 255038 304300 255356
rect -5974 253800 -3762 254120
rect -2016 253922 -1786 253930
rect -2674 253722 -2006 253922
rect -1806 253722 -1786 253922
rect -2016 253708 -1786 253722
rect -5202 253052 -1206 253076
rect -5202 252780 -1502 253052
rect -1230 252780 -1206 253052
rect -5202 252760 -1206 252780
rect -5202 252756 -1526 252760
rect 303888 252356 304300 255038
rect 303888 252038 303926 252356
rect 304244 252038 304300 252356
rect -5974 250800 -3762 251120
rect -2016 250922 -1786 250930
rect -2674 250722 -2006 250922
rect -1806 250722 -1786 250922
rect -2016 250708 -1786 250722
rect -5202 250052 -1206 250076
rect -5202 249780 -1502 250052
rect -1230 249780 -1206 250052
rect -5202 249760 -1206 249780
rect -5202 249756 -1526 249760
rect 303888 249356 304300 252038
rect 303888 249038 303926 249356
rect 304244 249038 304300 249356
rect -5974 247800 -3762 248120
rect -2016 247922 -1786 247930
rect -2674 247722 -2006 247922
rect -1806 247722 -1786 247922
rect -2016 247708 -1786 247722
rect 303888 246356 304300 249038
rect 303888 246038 303926 246356
rect 304244 246038 304300 246356
rect -5974 244800 -3762 245120
rect -2016 244922 -1786 244930
rect -2674 244722 -2006 244922
rect -1806 244722 -1786 244922
rect -2016 244708 -1786 244722
rect -5202 244052 -1206 244076
rect -5202 243780 -1502 244052
rect -1230 243780 -1206 244052
rect -5202 243760 -1206 243780
rect -5202 243756 -1526 243760
rect 303888 243356 304300 246038
rect 303888 243038 303926 243356
rect 304244 243038 304300 243356
rect -5974 241800 -3762 242120
rect -2016 241922 -1786 241930
rect -2674 241722 -2006 241922
rect -1806 241722 -1786 241922
rect -2016 241708 -1786 241722
rect -5202 241052 -1206 241076
rect -5202 240780 -1502 241052
rect -1230 240780 -1206 241052
rect -5202 240760 -1206 240780
rect -5202 240756 -1526 240760
rect 303888 240356 304300 243038
rect 303888 240038 303926 240356
rect 304244 240038 304300 240356
rect -5974 238800 -3762 239120
rect -2016 238922 -1786 238930
rect -2674 238722 -2006 238922
rect -1806 238722 -1786 238922
rect -2016 238708 -1786 238722
rect -5202 238052 -1206 238076
rect -5202 237780 -1502 238052
rect -1230 237780 -1206 238052
rect -5202 237760 -1206 237780
rect -5202 237756 -1526 237760
rect 303888 237356 304300 240038
rect 303888 237038 303926 237356
rect 304244 237038 304300 237356
rect -5974 235800 -3762 236120
rect -2016 235922 -1786 235930
rect -2674 235722 -2006 235922
rect -1806 235722 -1786 235922
rect -2016 235708 -1786 235722
rect -5202 235052 -1206 235076
rect -5202 234780 -1502 235052
rect -1230 234780 -1206 235052
rect -5202 234760 -1206 234780
rect -5202 234756 -1526 234760
rect 303888 234356 304300 237038
rect 303888 234038 303926 234356
rect 304244 234038 304300 234356
rect -5974 232800 -3762 233120
rect -2016 232922 -1786 232930
rect -2674 232722 -2006 232922
rect -1806 232722 -1786 232922
rect -2016 232708 -1786 232722
rect -5202 232052 -1206 232076
rect -5202 231780 -1502 232052
rect -1230 231780 -1206 232052
rect -5202 231760 -1206 231780
rect -5202 231756 -1526 231760
rect 303888 231356 304300 234038
rect 303888 231038 303926 231356
rect 304244 231038 304300 231356
rect -5974 229800 -3762 230120
rect -2016 229922 -1786 229930
rect -2674 229722 -2006 229922
rect -1806 229722 -1786 229922
rect -2016 229708 -1786 229722
rect -5202 229052 -1206 229076
rect -5202 228780 -1502 229052
rect -1230 228780 -1206 229052
rect -5202 228760 -1206 228780
rect -5202 228756 -1526 228760
rect 303888 228356 304300 231038
rect 303888 228038 303926 228356
rect 304244 228038 304300 228356
rect -5974 226800 -3762 227120
rect -2016 226922 -1786 226930
rect -2674 226722 -2006 226922
rect -1806 226722 -1786 226922
rect -2016 226708 -1786 226722
rect -5202 226052 -1206 226076
rect -5202 225780 -1502 226052
rect -1230 225780 -1206 226052
rect -5202 225760 -1206 225780
rect -5202 225756 -1526 225760
rect 303888 225356 304300 228038
rect 303888 225038 303926 225356
rect 304244 225038 304300 225356
rect -5974 223800 -3762 224120
rect -2016 223922 -1786 223930
rect -2674 223722 -2006 223922
rect -1806 223722 -1786 223922
rect -2016 223708 -1786 223722
rect -5202 223052 -1206 223076
rect -5202 222780 -1502 223052
rect -1230 222780 -1206 223052
rect -5202 222760 -1206 222780
rect -5202 222756 -1526 222760
rect 303888 222356 304300 225038
rect 303888 222038 303926 222356
rect 304244 222038 304300 222356
rect -5974 220800 -3762 221120
rect -2016 220922 -1786 220930
rect -2674 220722 -2006 220922
rect -1806 220722 -1786 220922
rect -2016 220708 -1786 220722
rect -5202 220052 -1206 220076
rect -5202 219780 -1502 220052
rect -1230 219780 -1206 220052
rect -5202 219760 -1206 219780
rect -5202 219756 -1526 219760
rect 303888 219356 304300 222038
rect 303888 219038 303926 219356
rect 304244 219038 304300 219356
rect -5974 217800 -3762 218120
rect -2016 217922 -1786 217930
rect -2674 217722 -2006 217922
rect -1806 217722 -1786 217922
rect -2016 217708 -1786 217722
rect -5202 217052 -1206 217076
rect -5202 216780 -1502 217052
rect -1230 216780 -1206 217052
rect -5202 216760 -1206 216780
rect -5202 216756 -1526 216760
rect 303888 216356 304300 219038
rect 303888 216038 303926 216356
rect 304244 216038 304300 216356
rect -5974 214800 -3762 215120
rect -2016 214922 -1786 214930
rect -2674 214722 -2006 214922
rect -1806 214722 -1786 214922
rect -2016 214708 -1786 214722
rect -5202 214052 -1206 214076
rect -5202 213780 -1502 214052
rect -1230 213780 -1206 214052
rect -5202 213760 -1206 213780
rect -5202 213756 -1526 213760
rect 303888 213356 304300 216038
rect 303888 213038 303926 213356
rect 304244 213038 304300 213356
rect -5974 211800 -3762 212120
rect -2016 211922 -1786 211930
rect -2674 211722 -2006 211922
rect -1806 211722 -1786 211922
rect -2016 211708 -1786 211722
rect -5202 211052 -1206 211076
rect -5202 210780 -1502 211052
rect -1230 210780 -1206 211052
rect -5202 210760 -1206 210780
rect -5202 210756 -1526 210760
rect 303888 210356 304300 213038
rect 303888 210038 303926 210356
rect 304244 210038 304300 210356
rect -2016 208922 -1786 208930
rect -2674 208722 -2006 208922
rect -1806 208722 -1786 208922
rect -2016 208708 -1786 208722
rect -5202 208052 -1206 208076
rect -5202 207780 -1502 208052
rect -1230 207780 -1206 208052
rect -5202 207760 -1206 207780
rect -5202 207756 -1526 207760
rect 303888 207356 304300 210038
rect 303888 207038 303926 207356
rect 304244 207038 304300 207356
rect -5974 205800 -3762 206120
rect -2016 205922 -1786 205930
rect -2674 205722 -2006 205922
rect -1806 205722 -1786 205922
rect -2016 205708 -1786 205722
rect -5202 205052 -1206 205076
rect -5202 204780 -1502 205052
rect -1230 204780 -1206 205052
rect -5202 204760 -1206 204780
rect -5202 204756 -1526 204760
rect 303888 204356 304300 207038
rect 303888 204038 303926 204356
rect 304244 204038 304300 204356
rect -5974 202800 -3762 203120
rect -2016 202922 -1786 202930
rect -2674 202722 -2006 202922
rect -1806 202722 -1786 202922
rect -2016 202708 -1786 202722
rect -5202 202052 -1206 202076
rect -5202 201780 -1502 202052
rect -1230 201780 -1206 202052
rect -5202 201760 -1206 201780
rect -5202 201756 -1526 201760
rect 303888 201356 304300 204038
rect 303888 201038 303926 201356
rect 304244 201038 304300 201356
rect -5974 199800 -3762 200120
rect -2016 199922 -1786 199930
rect -2674 199722 -2006 199922
rect -1806 199722 -1786 199922
rect -2016 199708 -1786 199722
rect -5202 199052 -1206 199076
rect -5202 198780 -1502 199052
rect -1230 198780 -1206 199052
rect -5202 198760 -1206 198780
rect -5202 198756 -1526 198760
rect 303888 198356 304300 201038
rect 303888 198038 303926 198356
rect 304244 198038 304300 198356
rect -5974 196800 -3762 197120
rect -2016 196922 -1786 196930
rect -2674 196722 -2006 196922
rect -1806 196722 -1786 196922
rect -2016 196708 -1786 196722
rect -5202 196052 -1206 196076
rect -5202 195780 -1502 196052
rect -1230 195780 -1206 196052
rect -5202 195760 -1206 195780
rect -5202 195756 -1526 195760
rect 303888 195356 304300 198038
rect 303888 195038 303926 195356
rect 304244 195038 304300 195356
rect -5974 193800 -3762 194120
rect -2016 193922 -1786 193930
rect -2674 193722 -2006 193922
rect -1806 193722 -1786 193922
rect -2016 193708 -1786 193722
rect -5202 193052 -1206 193076
rect -5202 192780 -1502 193052
rect -1230 192780 -1206 193052
rect -5202 192760 -1206 192780
rect -5202 192756 -1526 192760
rect 303888 192356 304300 195038
rect 303888 192038 303926 192356
rect 304244 192038 304300 192356
rect -5974 190800 -3762 191120
rect -2016 190922 -1786 190930
rect -2674 190722 -2006 190922
rect -1806 190722 -1786 190922
rect -2016 190708 -1786 190722
rect -5202 190052 -1206 190076
rect -5202 189780 -1502 190052
rect -1230 189780 -1206 190052
rect -5202 189760 -1206 189780
rect -5202 189756 -1526 189760
rect 303888 189356 304300 192038
rect 303888 189038 303926 189356
rect 304244 189038 304300 189356
rect -5974 187800 -3762 188120
rect -2016 187922 -1786 187930
rect -2674 187722 -2006 187922
rect -1806 187722 -1786 187922
rect -2016 187708 -1786 187722
rect -5202 187052 -1206 187076
rect -5202 186780 -1502 187052
rect -1230 186780 -1206 187052
rect -5202 186760 -1206 186780
rect -5202 186756 -1526 186760
rect 303888 186356 304300 189038
rect 303888 186038 303926 186356
rect 304244 186038 304300 186356
rect -5974 184800 -3762 185120
rect -2016 184922 -1786 184930
rect -2674 184722 -2006 184922
rect -1806 184722 -1786 184922
rect -2016 184708 -1786 184722
rect -5202 184052 -1206 184076
rect -5202 183780 -1502 184052
rect -1230 183780 -1206 184052
rect -5202 183760 -1206 183780
rect -5202 183756 -1526 183760
rect 303888 183356 304300 186038
rect 303888 183038 303926 183356
rect 304244 183038 304300 183356
rect -5974 181800 -3762 182120
rect -2016 181922 -1786 181930
rect -2674 181722 -2006 181922
rect -1806 181722 -1786 181922
rect -2016 181708 -1786 181722
rect -5202 181052 -1206 181076
rect -5202 180780 -1502 181052
rect -1230 180780 -1206 181052
rect -5202 180760 -1206 180780
rect -5202 180756 -1526 180760
rect 303888 180356 304300 183038
rect 303888 180038 303926 180356
rect 304244 180038 304300 180356
rect -5974 178800 -3762 179120
rect -2016 178922 -1786 178930
rect -2674 178722 -2006 178922
rect -1806 178722 -1786 178922
rect -2016 178708 -1786 178722
rect -5202 178052 -1206 178076
rect -5202 177780 -1502 178052
rect -1230 177780 -1206 178052
rect -5202 177760 -1206 177780
rect -5202 177756 -1526 177760
rect 303888 177356 304300 180038
rect 303888 177038 303926 177356
rect 304244 177038 304300 177356
rect -5974 175800 -3762 176120
rect -2016 175922 -1786 175930
rect -2674 175722 -2006 175922
rect -1806 175722 -1786 175922
rect -2016 175708 -1786 175722
rect -5202 175052 -1206 175076
rect -5202 174780 -1502 175052
rect -1230 174780 -1206 175052
rect -5202 174760 -1206 174780
rect -5202 174756 -1526 174760
rect 303888 174356 304300 177038
rect 303888 174038 303926 174356
rect 304244 174038 304300 174356
rect -5974 172800 -3762 173120
rect -2016 172922 -1786 172930
rect -2674 172722 -2006 172922
rect -1806 172722 -1786 172922
rect -2016 172708 -1786 172722
rect -5202 172052 -1206 172076
rect -5202 171780 -1502 172052
rect -1230 171780 -1206 172052
rect -5202 171760 -1206 171780
rect -5202 171756 -1526 171760
rect 303888 171356 304300 174038
rect 303888 171038 303926 171356
rect 304244 171038 304300 171356
rect -5974 169800 -3762 170120
rect -2016 169922 -1786 169930
rect -2674 169722 -2006 169922
rect -1806 169722 -1786 169922
rect -2016 169708 -1786 169722
rect -5202 169052 -1206 169076
rect -5202 168780 -1502 169052
rect -1230 168780 -1206 169052
rect -5202 168760 -1206 168780
rect -5202 168756 -1526 168760
rect 303888 168356 304300 171038
rect 303888 168038 303926 168356
rect 304244 168038 304300 168356
rect -5974 166800 -3762 167120
rect -2016 166922 -1786 166930
rect -2674 166722 -2006 166922
rect -1806 166722 -1786 166922
rect -2016 166708 -1786 166722
rect -5202 166052 -1206 166076
rect -5202 165780 -1502 166052
rect -1230 165780 -1206 166052
rect -5202 165760 -1206 165780
rect -5202 165756 -1526 165760
rect 303888 165356 304300 168038
rect 303888 165038 303926 165356
rect 304244 165038 304300 165356
rect -5974 163800 -3762 164120
rect -2016 163922 -1786 163930
rect -2674 163722 -2006 163922
rect -1806 163722 -1786 163922
rect -2016 163708 -1786 163722
rect -5202 163052 -1206 163076
rect -5202 162780 -1502 163052
rect -1230 162780 -1206 163052
rect -5202 162760 -1206 162780
rect -5202 162756 -1526 162760
rect 303888 162356 304300 165038
rect 303888 162038 303926 162356
rect 304244 162038 304300 162356
rect -5974 160800 -3762 161120
rect -2016 160922 -1786 160930
rect -2674 160722 -2006 160922
rect -1806 160722 -1786 160922
rect -2016 160708 -1786 160722
rect -5202 160052 -1206 160076
rect -5202 159780 -1502 160052
rect -1230 159780 -1206 160052
rect -5202 159760 -1206 159780
rect -5202 159756 -1526 159760
rect 303888 159356 304300 162038
rect 303888 159038 303926 159356
rect 304244 159038 304300 159356
rect -5974 157800 -3762 158120
rect -2016 157922 -1786 157930
rect -2674 157722 -2006 157922
rect -1806 157722 -1786 157922
rect -2016 157708 -1786 157722
rect -5202 157052 -1206 157076
rect -5202 156780 -1502 157052
rect -1230 156780 -1206 157052
rect -5202 156760 -1206 156780
rect -5202 156756 -1526 156760
rect 303888 156356 304300 159038
rect 303888 156038 303926 156356
rect 304244 156038 304300 156356
rect -5974 154800 -3762 155120
rect -2016 154922 -1786 154930
rect -2674 154722 -2006 154922
rect -1806 154722 -1786 154922
rect -2016 154708 -1786 154722
rect -5202 154052 -1206 154076
rect -5202 153780 -1502 154052
rect -1230 153780 -1206 154052
rect -5202 153760 -1206 153780
rect -5202 153756 -1526 153760
rect 303888 153356 304300 156038
rect 303888 153038 303926 153356
rect 304244 153038 304300 153356
rect -5974 151800 -3762 152120
rect -2016 151922 -1786 151930
rect -2674 151722 -2006 151922
rect -1806 151722 -1786 151922
rect -2016 151708 -1786 151722
rect -5202 151052 -1206 151076
rect -5202 150780 -1502 151052
rect -1230 150780 -1206 151052
rect -5202 150760 -1206 150780
rect -5202 150756 -1526 150760
rect 303888 150356 304300 153038
rect 303888 150038 303926 150356
rect 304244 150038 304300 150356
rect -5974 148800 -3762 149120
rect -2016 148922 -1786 148930
rect -2674 148722 -2006 148922
rect -1806 148722 -1786 148922
rect -2016 148708 -1786 148722
rect -5202 148052 -1206 148076
rect -5202 147780 -1502 148052
rect -1230 147780 -1206 148052
rect -5202 147760 -1206 147780
rect -5202 147756 -1526 147760
rect 303888 147356 304300 150038
rect 303888 147038 303926 147356
rect 304244 147038 304300 147356
rect -5974 145800 -3762 146120
rect -2016 145922 -1786 145930
rect -2674 145722 -2006 145922
rect -1806 145722 -1786 145922
rect -2016 145708 -1786 145722
rect -5202 145052 -1206 145076
rect -5202 144780 -1502 145052
rect -1230 144780 -1206 145052
rect -5202 144760 -1206 144780
rect -5202 144756 -1526 144760
rect 303888 144356 304300 147038
rect 303888 144038 303926 144356
rect 304244 144038 304300 144356
rect -5974 142800 -3762 143120
rect -2016 142922 -1786 142930
rect -2674 142722 -2006 142922
rect -1806 142722 -1786 142922
rect -2016 142708 -1786 142722
rect -5202 142052 -1206 142076
rect -5202 141780 -1502 142052
rect -1230 141780 -1206 142052
rect -5202 141760 -1206 141780
rect -5202 141756 -1526 141760
rect 303888 141356 304300 144038
rect 303888 141038 303926 141356
rect 304244 141038 304300 141356
rect -5974 139800 -3762 140120
rect -2016 139922 -1786 139930
rect -2674 139722 -2006 139922
rect -1806 139722 -1786 139922
rect -2016 139708 -1786 139722
rect -5202 139052 -1206 139076
rect -5202 138780 -1502 139052
rect -1230 138780 -1206 139052
rect -5202 138760 -1206 138780
rect -5202 138756 -1526 138760
rect 303888 138356 304300 141038
rect 303888 138038 303926 138356
rect 304244 138038 304300 138356
rect -5974 136800 -3762 137120
rect -2016 136922 -1786 136930
rect -2674 136722 -2006 136922
rect -1806 136722 -1786 136922
rect -2016 136708 -1786 136722
rect -5202 136052 -1206 136076
rect -5202 135780 -1502 136052
rect -1230 135780 -1206 136052
rect -5202 135760 -1206 135780
rect -5202 135756 -1526 135760
rect 303888 135356 304300 138038
rect 303888 135038 303926 135356
rect 304244 135038 304300 135356
rect -5974 133800 -3762 134120
rect -2016 133922 -1786 133930
rect -2674 133722 -2006 133922
rect -1806 133722 -1786 133922
rect -2016 133708 -1786 133722
rect -5202 133052 -1206 133076
rect -5202 132780 -1502 133052
rect -1230 132780 -1206 133052
rect -5202 132760 -1206 132780
rect -5202 132756 -1526 132760
rect 303888 132356 304300 135038
rect 303888 132038 303926 132356
rect 304244 132038 304300 132356
rect -5974 130800 -3762 131120
rect -2016 130922 -1786 130930
rect -2674 130722 -2006 130922
rect -1806 130722 -1786 130922
rect -2016 130708 -1786 130722
rect -5202 130052 -1206 130076
rect -5202 129780 -1502 130052
rect -1230 129780 -1206 130052
rect -5202 129760 -1206 129780
rect -5202 129756 -1526 129760
rect 303888 129356 304300 132038
rect 303888 129038 303926 129356
rect 304244 129038 304300 129356
rect -5974 127800 -3762 128120
rect -2016 127922 -1786 127930
rect -2674 127722 -2006 127922
rect -1806 127722 -1786 127922
rect -2016 127708 -1786 127722
rect -5202 127052 -1206 127076
rect -5202 126780 -1502 127052
rect -1230 126780 -1206 127052
rect -5202 126760 -1206 126780
rect -5202 126756 -1526 126760
rect 303888 126356 304300 129038
rect 303888 126038 303926 126356
rect 304244 126038 304300 126356
rect -5974 124800 -3762 125120
rect -2016 124922 -1786 124930
rect -2674 124722 -2006 124922
rect -1806 124722 -1786 124922
rect -2016 124708 -1786 124722
rect -5202 124052 -1206 124076
rect -5202 123780 -1502 124052
rect -1230 123780 -1206 124052
rect -5202 123760 -1206 123780
rect -5202 123756 -1526 123760
rect 303888 123356 304300 126038
rect 303888 123038 303926 123356
rect 304244 123038 304300 123356
rect -5974 121800 -3762 122120
rect -2016 121922 -1786 121930
rect -2674 121722 -2006 121922
rect -1806 121722 -1786 121922
rect -2016 121708 -1786 121722
rect -5202 121052 -1206 121076
rect -5202 120780 -1502 121052
rect -1230 120780 -1206 121052
rect -5202 120760 -1206 120780
rect -5202 120756 -1526 120760
rect 303888 120356 304300 123038
rect 303888 120038 303926 120356
rect 304244 120038 304300 120356
rect -5974 118800 -3762 119120
rect -2016 118922 -1786 118930
rect -2674 118722 -2006 118922
rect -1806 118722 -1786 118922
rect -2016 118708 -1786 118722
rect -5202 118052 -1206 118076
rect -5202 117780 -1502 118052
rect -1230 117780 -1206 118052
rect -5202 117760 -1206 117780
rect -5202 117756 -1526 117760
rect 303888 117356 304300 120038
rect 303888 117038 303926 117356
rect 304244 117038 304300 117356
rect -5974 115800 -3762 116120
rect -2016 115922 -1786 115930
rect -2674 115722 -2006 115922
rect -1806 115722 -1786 115922
rect -2016 115708 -1786 115722
rect -5202 115052 -1206 115076
rect -5202 114780 -1502 115052
rect -1230 114780 -1206 115052
rect -5202 114760 -1206 114780
rect -5202 114756 -1526 114760
rect 303888 114356 304300 117038
rect 303888 114038 303926 114356
rect 304244 114038 304300 114356
rect -5974 112800 -3762 113120
rect -2016 112922 -1786 112930
rect -2674 112722 -2006 112922
rect -1806 112722 -1786 112922
rect -2016 112708 -1786 112722
rect -5202 112052 -1206 112076
rect -5202 111780 -1502 112052
rect -1230 111780 -1206 112052
rect -5202 111760 -1206 111780
rect -5202 111756 -1526 111760
rect 303888 111356 304300 114038
rect 303888 111038 303926 111356
rect 304244 111038 304300 111356
rect -5974 109800 -3762 110120
rect -2016 109922 -1786 109930
rect -2674 109722 -2006 109922
rect -1806 109722 -1786 109922
rect -2016 109708 -1786 109722
rect -5202 109052 -1206 109076
rect -5202 108780 -1502 109052
rect -1230 108780 -1206 109052
rect -5202 108760 -1206 108780
rect -5202 108756 -1526 108760
rect 303888 108356 304300 111038
rect 303888 108038 303926 108356
rect 304244 108038 304300 108356
rect -5974 106800 -3762 107120
rect -2016 106922 -1786 106930
rect -2674 106722 -2006 106922
rect -1806 106722 -1786 106922
rect -2016 106708 -1786 106722
rect -5202 106052 -1206 106076
rect -5202 105780 -1502 106052
rect -1230 105780 -1206 106052
rect -5202 105760 -1206 105780
rect -5202 105756 -1526 105760
rect 303888 105356 304300 108038
rect 303888 105038 303926 105356
rect 304244 105038 304300 105356
rect -5974 103800 -3762 104120
rect -2016 103922 -1786 103930
rect -2674 103722 -2006 103922
rect -1806 103722 -1786 103922
rect -2016 103708 -1786 103722
rect -5202 103052 -1206 103076
rect -5202 102780 -1502 103052
rect -1230 102780 -1206 103052
rect -5202 102760 -1206 102780
rect -5202 102756 -1526 102760
rect 303888 102356 304300 105038
rect 303888 102038 303926 102356
rect 304244 102038 304300 102356
rect -5974 100800 -3762 101120
rect -2016 100922 -1786 100930
rect -2674 100722 -2006 100922
rect -1806 100722 -1786 100922
rect -2016 100708 -1786 100722
rect -5202 100052 -1206 100076
rect -5202 99780 -1502 100052
rect -1230 99780 -1206 100052
rect -5202 99760 -1206 99780
rect -5202 99756 -1526 99760
rect 303888 99356 304300 102038
rect 303888 99038 303926 99356
rect 304244 99038 304300 99356
rect -5974 97800 -3762 98120
rect -2016 97922 -1786 97930
rect -2674 97722 -2006 97922
rect -1806 97722 -1786 97922
rect -2016 97708 -1786 97722
rect -5202 97052 -1206 97076
rect -5202 96780 -1502 97052
rect -1230 96780 -1206 97052
rect -5202 96760 -1206 96780
rect -5202 96756 -1526 96760
rect 303888 96356 304300 99038
rect 303888 96038 303926 96356
rect 304244 96038 304300 96356
rect -5974 94800 -3762 95120
rect -2016 94922 -1786 94930
rect -2674 94722 -2006 94922
rect -1806 94722 -1786 94922
rect -2016 94708 -1786 94722
rect 303888 93356 304300 96038
rect 303888 93038 303926 93356
rect 304244 93038 304300 93356
rect -5974 91800 -3762 92120
rect -2016 91922 -1786 91930
rect -2674 91722 -2006 91922
rect -1806 91722 -1786 91922
rect -2016 91708 -1786 91722
rect -5202 91052 -1206 91076
rect -5202 90780 -1502 91052
rect -1230 90780 -1206 91052
rect -5202 90760 -1206 90780
rect -5202 90756 -1526 90760
rect 303888 90356 304300 93038
rect 303888 90038 303926 90356
rect 304244 90038 304300 90356
rect -5974 88800 -3762 89120
rect -2016 88922 -1786 88930
rect -2674 88722 -2006 88922
rect -1806 88722 -1786 88922
rect -2016 88708 -1786 88722
rect -5202 88052 -1206 88076
rect -5202 87780 -1502 88052
rect -1230 87780 -1206 88052
rect -5202 87760 -1206 87780
rect -5202 87756 -1526 87760
rect 303888 87356 304300 90038
rect 303888 87038 303926 87356
rect 304244 87038 304300 87356
rect -5974 85800 -3762 86120
rect -2016 85922 -1786 85930
rect -2674 85722 -2006 85922
rect -1806 85722 -1786 85922
rect -2016 85708 -1786 85722
rect -5202 85052 -1206 85076
rect -5202 84780 -1502 85052
rect -1230 84780 -1206 85052
rect -5202 84760 -1206 84780
rect -5202 84756 -1526 84760
rect 303888 84356 304300 87038
rect 303888 84038 303926 84356
rect 304244 84038 304300 84356
rect -5974 82800 -3762 83120
rect -2016 82922 -1786 82930
rect -2674 82722 -2006 82922
rect -1806 82722 -1786 82922
rect -2016 82708 -1786 82722
rect -5202 82052 -1206 82076
rect -5202 81780 -1502 82052
rect -1230 81780 -1206 82052
rect -5202 81760 -1206 81780
rect -5202 81756 -1526 81760
rect 303888 81356 304300 84038
rect 303888 81038 303926 81356
rect 304244 81038 304300 81356
rect -5974 79800 -3762 80120
rect -2016 79922 -1786 79930
rect -2674 79722 -2006 79922
rect -1806 79722 -1786 79922
rect -2016 79708 -1786 79722
rect -5202 79052 -1206 79076
rect -5202 78780 -1502 79052
rect -1230 78780 -1206 79052
rect -5202 78760 -1206 78780
rect -5202 78756 -1526 78760
rect 303888 78356 304300 81038
rect 303888 78038 303926 78356
rect 304244 78038 304300 78356
rect -5974 76800 -3762 77120
rect -2016 76922 -1786 76930
rect -2674 76722 -2006 76922
rect -1806 76722 -1786 76922
rect -2016 76708 -1786 76722
rect -5202 76052 -1206 76076
rect -5202 75780 -1502 76052
rect -1230 75780 -1206 76052
rect -5202 75760 -1206 75780
rect -5202 75756 -1526 75760
rect 303888 75356 304300 78038
rect 303888 75038 303926 75356
rect 304244 75038 304300 75356
rect -5974 73800 -3762 74120
rect -2016 73922 -1786 73930
rect -2674 73722 -2006 73922
rect -1806 73722 -1786 73922
rect -2016 73708 -1786 73722
rect -5202 73052 -1206 73076
rect -5202 72780 -1502 73052
rect -1230 72780 -1206 73052
rect -5202 72760 -1206 72780
rect -5202 72756 -1526 72760
rect 303888 72356 304300 75038
rect 303888 72038 303926 72356
rect 304244 72038 304300 72356
rect -5974 70800 -3762 71120
rect -2016 70922 -1786 70930
rect -2674 70722 -2006 70922
rect -1806 70722 -1786 70922
rect -2016 70708 -1786 70722
rect -5202 70052 -1206 70076
rect -5202 69780 -1502 70052
rect -1230 69780 -1206 70052
rect -5202 69760 -1206 69780
rect -5202 69756 -1526 69760
rect 303888 69356 304300 72038
rect 303888 69038 303926 69356
rect 304244 69038 304300 69356
rect -5974 67800 -3762 68120
rect -2016 67922 -1786 67930
rect -2674 67722 -2006 67922
rect -1806 67722 -1786 67922
rect -2016 67708 -1786 67722
rect -5202 67052 -1206 67076
rect -5202 66780 -1502 67052
rect -1230 66780 -1206 67052
rect -5202 66760 -1206 66780
rect -5202 66756 -1526 66760
rect 303888 66356 304300 69038
rect 303888 66038 303926 66356
rect 304244 66038 304300 66356
rect -5974 64800 -3762 65120
rect -2016 64922 -1786 64930
rect -2674 64722 -2006 64922
rect -1806 64722 -1786 64922
rect -2016 64708 -1786 64722
rect -5202 64052 -1206 64076
rect -5202 63780 -1502 64052
rect -1230 63780 -1206 64052
rect -5202 63760 -1206 63780
rect -5202 63756 -1526 63760
rect 303888 63356 304300 66038
rect 303888 63038 303926 63356
rect 304244 63038 304300 63356
rect -5974 61800 -3762 62120
rect -2016 61922 -1786 61930
rect -2674 61722 -2006 61922
rect -1806 61722 -1786 61922
rect -2016 61708 -1786 61722
rect -5202 61052 -1206 61076
rect -5202 60780 -1502 61052
rect -1230 60780 -1206 61052
rect -5202 60760 -1206 60780
rect -5202 60756 -1526 60760
rect 303888 60356 304300 63038
rect 303888 60038 303926 60356
rect 304244 60038 304300 60356
rect -5974 58800 -3762 59120
rect -2016 58922 -1786 58930
rect -2674 58722 -2006 58922
rect -1806 58722 -1786 58922
rect -2016 58708 -1786 58722
rect -5202 58052 -1206 58076
rect -5202 57780 -1502 58052
rect -1230 57780 -1206 58052
rect -5202 57760 -1206 57780
rect -5202 57756 -1526 57760
rect 303888 57356 304300 60038
rect 303888 57038 303926 57356
rect 304244 57038 304300 57356
rect -2016 55922 -1786 55930
rect -2674 55722 -2006 55922
rect -1806 55722 -1786 55922
rect -2016 55708 -1786 55722
rect -5202 55052 -1206 55076
rect -5202 54780 -1502 55052
rect -1230 54780 -1206 55052
rect -5202 54760 -1206 54780
rect -5202 54756 -1526 54760
rect 303888 54356 304300 57038
rect 303888 54038 303926 54356
rect 304244 54038 304300 54356
rect -5974 52800 -3762 53120
rect -2016 52922 -1786 52930
rect -2674 52722 -2006 52922
rect -1806 52722 -1786 52922
rect -2016 52708 -1786 52722
rect -5202 52052 -1206 52076
rect -5202 51780 -1502 52052
rect -1230 51780 -1206 52052
rect -5202 51760 -1206 51780
rect -5202 51756 -1526 51760
rect 303888 51356 304300 54038
rect 303888 51038 303926 51356
rect 304244 51038 304300 51356
rect -5974 49800 -3762 50120
rect -2016 49922 -1786 49930
rect -2674 49722 -2006 49922
rect -1806 49722 -1786 49922
rect -2016 49708 -1786 49722
rect -5202 49052 -1206 49076
rect -5202 48780 -1502 49052
rect -1230 48780 -1206 49052
rect -5202 48760 -1206 48780
rect -5202 48756 -1526 48760
rect 303888 48356 304300 51038
rect 303888 48038 303926 48356
rect 304244 48038 304300 48356
rect -5974 46800 -3762 47120
rect -2016 46922 -1786 46930
rect -2674 46722 -2006 46922
rect -1806 46722 -1786 46922
rect -2016 46708 -1786 46722
rect -5202 46052 -1206 46076
rect -5202 45780 -1502 46052
rect -1230 45780 -1206 46052
rect -5202 45760 -1206 45780
rect -5202 45756 -1526 45760
rect 303888 45356 304300 48038
rect 303888 45038 303926 45356
rect 304244 45038 304300 45356
rect -5974 43800 -3762 44120
rect -2016 43922 -1786 43930
rect -2674 43722 -2006 43922
rect -1806 43722 -1786 43922
rect -2016 43708 -1786 43722
rect -5202 43052 -1206 43076
rect -5202 42780 -1502 43052
rect -1230 42780 -1206 43052
rect -5202 42760 -1206 42780
rect -5202 42756 -1526 42760
rect 303888 42356 304300 45038
rect 303888 42038 303926 42356
rect 304244 42038 304300 42356
rect -5974 40800 -3762 41120
rect -2016 40922 -1786 40930
rect -2674 40722 -2006 40922
rect -1806 40722 -1786 40922
rect -2016 40708 -1786 40722
rect -5202 40052 -1206 40076
rect -5202 39780 -1502 40052
rect -1230 39780 -1206 40052
rect -5202 39760 -1206 39780
rect -5202 39756 -1526 39760
rect 303888 39356 304300 42038
rect 303888 39038 303926 39356
rect 304244 39038 304300 39356
rect -5974 37800 -3762 38120
rect -2044 37922 -1762 37940
rect -2674 37722 -2006 37922
rect -1806 37722 -1762 37922
rect -2044 37700 -1762 37722
rect -5202 37052 -1206 37076
rect -5202 36780 -1502 37052
rect -1230 36780 -1206 37052
rect -5202 36760 -1206 36780
rect -5202 36756 -1526 36760
rect 303888 36356 304300 39038
rect 303888 36038 303926 36356
rect 304244 36038 304300 36356
rect -5974 34800 -3762 35120
rect -2030 34930 -1788 34970
rect -2030 34922 -1786 34930
rect -2674 34722 -2006 34922
rect -1806 34722 -1786 34922
rect -2030 34708 -1786 34722
rect -2030 34702 -1788 34708
rect -2004 34690 -1788 34702
rect -5202 34052 -1206 34076
rect -5202 33780 -1502 34052
rect -1230 33780 -1206 34052
rect -5202 33760 -1206 33780
rect -5202 33756 -1526 33760
rect 303888 33356 304300 36038
rect 303888 33038 303926 33356
rect 304244 33038 304300 33356
rect -5974 31800 -3762 32120
rect -2046 31922 -1772 31996
rect -2674 31722 -2006 31922
rect -1806 31722 -1772 31922
rect -2046 31696 -1772 31722
rect -5202 31052 -1206 31076
rect -5202 30780 -1502 31052
rect -1230 30780 -1206 31052
rect -5202 30760 -1206 30780
rect -5202 30756 -1526 30760
rect 303888 30356 304300 33038
rect 303888 30038 303926 30356
rect 304244 30038 304300 30356
rect -5974 28800 -3762 29120
rect -2016 28922 -1778 28946
rect -2674 28722 -2006 28922
rect -1806 28722 -1778 28922
rect -2016 28696 -1778 28722
rect -5202 28052 -1206 28076
rect -5202 27780 -1502 28052
rect -1230 27780 -1206 28052
rect -5202 27760 -1206 27780
rect -5202 27756 -1526 27760
rect 303888 27356 304300 30038
rect 303888 27038 303926 27356
rect 304244 27038 304300 27356
rect -5974 25800 -3762 26120
rect -2050 25932 -1806 25934
rect -2050 25922 -1780 25932
rect -2674 25722 -2006 25922
rect -1806 25722 -1780 25922
rect -2050 25704 -1780 25722
rect -2050 25692 -1806 25704
rect -5202 25052 -1206 25076
rect -5202 24780 -1502 25052
rect -1230 24780 -1206 25052
rect -5202 24760 -1206 24780
rect -5202 24756 -1526 24760
rect 303888 24356 304300 27038
rect 303888 24038 303926 24356
rect 304244 24038 304300 24356
rect -5974 22800 -3762 23120
rect -2026 22930 -1792 22942
rect -2026 22922 -1786 22930
rect -2674 22722 -2006 22922
rect -1806 22722 -1786 22922
rect -2026 22708 -1786 22722
rect -2026 22706 -1792 22708
rect -5202 22052 -1206 22076
rect -5202 21780 -1502 22052
rect -1230 21780 -1206 22052
rect -5202 21760 -1206 21780
rect -5202 21756 -1526 21760
rect 303888 21356 304300 24038
rect 303888 21038 303926 21356
rect 304244 21038 304300 21356
rect 303888 20952 304300 21038
rect -5974 19800 -3762 20120
rect -5202 19052 -1206 19076
rect -5202 18780 -1502 19052
rect -1230 18780 -1206 19052
rect -5202 18760 -1206 18780
rect -780 18794 1738 18904
rect -5202 18756 -1526 18760
rect -6094 17942 -5984 17960
rect -5994 17742 -5984 17942
rect -6094 17734 -5984 17742
rect -780 16796 -670 18794
rect 2328 18466 2548 19498
rect 5328 18810 5548 19606
rect 7470 18892 7720 18910
rect 8328 18892 8548 19654
rect 7470 18890 8548 18892
rect 5316 18784 5566 18810
rect 5316 18566 5328 18784
rect 5546 18566 5566 18784
rect 7470 18672 7482 18890
rect 7700 18672 8548 18890
rect 10692 18836 10942 18858
rect 11328 18836 11548 19678
rect 10692 18834 11548 18836
rect 7470 18652 7720 18672
rect 10692 18616 10712 18834
rect 10930 18616 11548 18834
rect 13790 18930 14040 18950
rect 14328 18930 14548 19678
rect 13790 18928 14548 18930
rect 13790 18710 13802 18928
rect 14020 18710 14548 18928
rect 16900 18816 17150 18824
rect 17328 18816 17548 19672
rect 19850 19194 20100 19202
rect 20328 19194 20548 19678
rect 19850 19192 20548 19194
rect 19850 18974 19870 19192
rect 20088 18974 20548 19192
rect 19850 18944 20100 18974
rect 13790 18692 14040 18710
rect 10692 18600 10942 18616
rect 16900 18598 16912 18816
rect 17130 18598 17548 18816
rect 22880 18672 23142 18674
rect 16900 18596 17548 18598
rect 22872 18658 23188 18672
rect 23328 18658 23548 19678
rect 25908 19012 26226 19028
rect 26328 19012 26548 19678
rect 29328 19158 29548 19678
rect 25908 19010 26548 19012
rect 25908 18792 25944 19010
rect 26162 18792 26548 19010
rect 29074 19060 29548 19158
rect 29074 18842 29084 19060
rect 29302 18842 29548 19060
rect 32328 18996 32548 19678
rect 35328 19066 35548 19596
rect 38328 19226 38548 19634
rect 38312 19218 38562 19226
rect 35298 19054 35584 19066
rect 32302 18986 32578 18996
rect 29074 18828 29428 18842
rect 25908 18762 26226 18792
rect 32302 18768 32328 18986
rect 32546 18768 32578 18986
rect 35298 18836 35328 19054
rect 35546 18836 35584 19054
rect 38312 19000 38328 19218
rect 38546 19000 38562 19218
rect 38312 18968 38562 19000
rect 41328 18898 41548 19678
rect 44328 18936 44548 19672
rect 47328 19154 47548 19678
rect 47292 19130 47590 19154
rect 44320 18922 44570 18936
rect 35298 18828 35584 18836
rect 41310 18872 41582 18898
rect 32302 18742 32578 18768
rect 35328 18758 35548 18828
rect 16900 18566 17150 18596
rect 5316 18552 5566 18566
rect 2316 18438 2566 18466
rect 2316 18220 2328 18438
rect 2546 18220 2566 18438
rect 22872 18440 22898 18658
rect 23116 18440 23548 18658
rect 41310 18654 41328 18872
rect 41546 18654 41582 18872
rect 44320 18704 44328 18922
rect 44546 18704 44570 18922
rect 47292 18912 47328 19130
rect 47546 18912 47590 19130
rect 47292 18900 47590 18912
rect 50328 19022 50548 19654
rect 53328 19064 53548 19678
rect 56328 19240 56548 19666
rect 56328 19162 56968 19240
rect 53328 19042 53770 19064
rect 50328 19010 50750 19022
rect 47318 18886 47568 18900
rect 50328 18792 50516 19010
rect 50734 18792 50750 19010
rect 53328 18824 53538 19042
rect 53756 18824 53770 19042
rect 56328 18944 56616 19162
rect 56834 18944 56968 19162
rect 56328 18942 56858 18944
rect 56590 18922 56858 18942
rect 53328 18822 53770 18824
rect 53520 18806 53770 18822
rect 59328 18866 59548 19678
rect 59618 18866 59882 18890
rect 50500 18764 50750 18792
rect 44320 18678 44570 18704
rect 41310 18618 41582 18654
rect 59328 18648 59630 18866
rect 59848 18648 59882 18866
rect 59328 18646 59882 18648
rect 59618 18638 59882 18646
rect 62328 18866 62548 19678
rect 65328 18882 65548 19644
rect 68328 18992 68548 19638
rect 71328 19060 71548 19630
rect 71914 19060 72174 19076
rect 68290 18952 68580 18992
rect 65740 18882 65978 18896
rect 65328 18880 65978 18882
rect 62328 18834 62946 18866
rect 62328 18790 62974 18834
rect 62328 18572 62632 18790
rect 62850 18572 62974 18790
rect 65328 18662 65742 18880
rect 65960 18662 65978 18880
rect 68290 18734 68328 18952
rect 68546 18734 68580 18952
rect 71328 18842 71928 19060
rect 72146 18842 72174 19060
rect 71328 18840 72174 18842
rect 71914 18828 72174 18840
rect 74328 19030 74548 19676
rect 75054 19030 75306 19042
rect 74328 18812 75078 19030
rect 75296 18812 75306 19030
rect 74328 18810 75306 18812
rect 75054 18798 75306 18810
rect 68290 18726 68580 18734
rect 65740 18648 65978 18662
rect 62328 18570 62974 18572
rect 62572 18542 62974 18570
rect 62604 18530 62876 18542
rect 22872 18438 23548 18440
rect 22872 18406 23188 18438
rect 71910 18292 72162 18536
rect 77328 18306 77548 19678
rect 80328 18906 80548 19676
rect 80328 18904 81410 18906
rect 80328 18686 81190 18904
rect 81408 18720 81410 18904
rect 81408 18686 81430 18720
rect 81172 18482 81430 18686
rect 83328 18404 83548 19662
rect 84252 18404 84516 18424
rect 83328 18402 84516 18404
rect 78078 18306 78330 18312
rect 2316 18208 2566 18220
rect 77328 18088 78098 18306
rect 78316 18088 78330 18306
rect 83328 18184 84274 18402
rect 84492 18184 84516 18402
rect 84252 18164 84516 18184
rect 86328 18314 86548 19678
rect 89328 18838 89548 19632
rect 90400 18838 90652 18856
rect 89328 18836 90652 18838
rect 89328 18618 90412 18836
rect 90630 18618 90652 18836
rect 90400 18608 90652 18618
rect 92328 18794 92548 19624
rect 95328 18876 95548 19632
rect 96442 18876 96684 18884
rect 95328 18874 96684 18876
rect 93536 18794 93788 18810
rect 92328 18792 93788 18794
rect 92328 18574 93556 18792
rect 93774 18574 93788 18792
rect 95328 18656 96454 18874
rect 96672 18656 96684 18874
rect 96442 18650 96684 18656
rect 93536 18562 93788 18574
rect 98328 18502 98548 19638
rect 101328 18740 101548 19610
rect 102658 18740 102952 18774
rect 99574 18502 99854 18534
rect 101328 18522 102712 18740
rect 102930 18522 102952 18740
rect 104328 18756 104548 19632
rect 107328 19032 107548 19624
rect 108892 19032 109134 19040
rect 107328 18814 108902 19032
rect 109120 18814 109134 19032
rect 107328 18812 109134 18814
rect 108892 18808 109134 18812
rect 110328 18936 110548 19646
rect 113328 18984 113548 19658
rect 114930 18984 115200 19008
rect 111936 18936 112184 18948
rect 110328 18934 112184 18936
rect 105620 18756 105914 18790
rect 104328 18754 105914 18756
rect 104328 18536 105676 18754
rect 105894 18536 105914 18754
rect 110328 18716 111948 18934
rect 112166 18716 112184 18934
rect 113328 18766 114954 18984
rect 115172 18766 115200 18984
rect 113328 18764 115200 18766
rect 114930 18744 115200 18764
rect 116328 18978 116548 19612
rect 117942 18978 118250 18998
rect 116328 18976 118250 18978
rect 116328 18758 117968 18976
rect 118186 18758 118250 18976
rect 111936 18712 112184 18716
rect 117942 18686 118250 18758
rect 119328 18864 119548 19678
rect 121114 18864 121400 18884
rect 119328 18646 121150 18864
rect 121368 18646 121400 18864
rect 119328 18644 121400 18646
rect 121114 18598 121400 18644
rect 122328 18852 122548 19658
rect 125328 18942 125548 19678
rect 127190 18942 127500 18970
rect 124096 18852 124354 18864
rect 122328 18850 124354 18852
rect 122328 18632 124118 18850
rect 124336 18632 124354 18850
rect 125328 18724 127242 18942
rect 127460 18724 127500 18942
rect 125328 18722 127500 18724
rect 127190 18678 127500 18722
rect 128328 18814 128548 19644
rect 131328 18866 131548 19674
rect 133376 18866 133686 18894
rect 130210 18814 130520 18858
rect 128328 18812 130520 18814
rect 124096 18624 124354 18632
rect 128328 18594 130250 18812
rect 130468 18594 130520 18812
rect 131328 18648 133412 18866
rect 133630 18648 133686 18866
rect 131328 18646 133686 18648
rect 133376 18602 133686 18646
rect 130210 18566 130520 18594
rect 101328 18520 102952 18522
rect 98328 18500 99854 18502
rect 87330 18314 87580 18326
rect 86328 18096 87336 18314
rect 87554 18096 87580 18314
rect 98328 18282 99598 18500
rect 99816 18282 99854 18500
rect 102658 18468 102952 18520
rect 105620 18484 105914 18536
rect 99574 18244 99854 18282
rect 86328 18094 87580 18096
rect 77328 18086 78330 18088
rect 87330 18086 87580 18094
rect 134328 18242 134548 19658
rect 137328 18600 137548 19614
rect 140328 18668 140548 19678
rect 143328 18844 143548 19674
rect 145538 18844 145832 18860
rect 143328 18842 145832 18844
rect 142542 18668 142852 18692
rect 139492 18600 139802 18606
rect 137328 18382 139552 18600
rect 139770 18382 139802 18600
rect 140328 18450 142600 18668
rect 142818 18450 142852 18668
rect 143328 18624 145578 18842
rect 145796 18624 145832 18842
rect 146328 18844 146548 19666
rect 148714 18844 149008 18874
rect 146328 18842 149008 18844
rect 146328 18624 148754 18842
rect 148972 18624 149008 18842
rect 145538 18580 145832 18624
rect 148714 18594 149008 18624
rect 149328 18774 149548 19658
rect 152328 18858 152548 19658
rect 155328 18998 155548 19658
rect 157794 18998 158088 19008
rect 155328 18996 158088 18998
rect 154754 18858 155048 18876
rect 151732 18774 152026 18802
rect 149328 18556 151772 18774
rect 151990 18556 152026 18774
rect 152328 18640 154792 18858
rect 155010 18640 155048 18858
rect 155328 18778 157844 18996
rect 158062 18778 158088 18996
rect 157794 18728 158088 18778
rect 158328 18758 158548 19678
rect 161328 18890 161548 19666
rect 164328 19028 164548 19666
rect 167328 19136 167548 19658
rect 160862 18758 161156 18778
rect 152328 18638 155048 18640
rect 154754 18596 155048 18638
rect 149328 18554 152026 18556
rect 151732 18522 152026 18554
rect 158328 18540 160886 18758
rect 161104 18540 161156 18758
rect 161328 18670 163556 18890
rect 164328 18808 166148 19028
rect 167328 18916 169082 19136
rect 158328 18538 161156 18540
rect 160862 18498 161156 18538
rect 163238 18486 163458 18670
rect 140328 18448 142852 18450
rect 142542 18400 142852 18448
rect 163202 18458 163496 18486
rect 137328 18380 139802 18382
rect 139492 18314 139802 18380
rect 136442 18242 136752 18286
rect 134328 18240 136752 18242
rect 78078 18068 78330 18086
rect 84246 17732 84526 18028
rect 134328 18022 136468 18240
rect 136686 18022 136752 18240
rect 163202 18240 163238 18458
rect 163456 18240 163496 18458
rect 163202 18206 163496 18240
rect 165928 18202 166148 18808
rect 136442 17994 136752 18022
rect 165896 18174 166190 18202
rect 165896 17956 165928 18174
rect 166146 17956 166190 18174
rect 165896 17922 166190 17956
rect 168862 17446 169082 18916
rect 170328 18490 170548 19642
rect 173328 19136 173548 19678
rect 174332 19136 174626 19162
rect 173328 19134 174626 19136
rect 173328 18916 174366 19134
rect 174584 18916 174626 19134
rect 174332 18882 174626 18916
rect 176328 18846 176548 19628
rect 176292 18812 176586 18846
rect 176292 18594 176328 18812
rect 176546 18594 176586 18812
rect 176292 18566 176586 18594
rect 173060 18490 173354 18508
rect 170328 18488 173354 18490
rect 170328 18270 173082 18488
rect 173300 18270 173354 18488
rect 173060 18228 173354 18270
rect 179328 17860 179548 19678
rect 182328 18782 182548 19658
rect 182328 18562 184230 18782
rect 182444 17860 182738 17894
rect 179328 17858 182738 17860
rect 179328 17640 182474 17858
rect 182692 17640 182738 17858
rect 182444 17614 182738 17640
rect 168824 17420 169118 17446
rect 168824 17202 168864 17420
rect 169082 17202 169118 17420
rect 168824 17166 169118 17202
rect 184010 17190 184230 18562
rect 185328 18060 185548 19678
rect 185290 18036 185584 18060
rect 185290 17818 185328 18036
rect 185546 17818 185584 18036
rect 185290 17780 185584 17818
rect 188328 17686 188548 19658
rect 191328 18626 191548 19634
rect 191328 18406 193684 18626
rect 188280 17658 188574 17686
rect 188280 17440 188328 17658
rect 188546 17440 188574 17658
rect 188280 17406 188574 17440
rect 183972 17152 184266 17190
rect 183972 16934 184010 17152
rect 184228 16934 184266 17152
rect 193464 17048 193684 18406
rect 194328 17930 194548 19624
rect 197328 17956 197548 19660
rect 200328 18804 200548 19624
rect 200328 18584 202222 18804
rect 200892 17956 201204 18006
rect 196770 17930 197064 17956
rect 194328 17928 197064 17930
rect 194328 17710 196794 17928
rect 197012 17710 197064 17928
rect 197328 17738 200916 17956
rect 201134 17738 201204 17956
rect 197328 17736 201204 17738
rect 196770 17676 197064 17710
rect 200892 17700 201204 17736
rect 183972 16910 184266 16934
rect 193426 17018 193720 17048
rect -4334 16686 -670 16796
rect 193426 16800 193466 17018
rect 193684 16800 193720 17018
rect 202002 16902 202222 18584
rect 203328 17752 203548 19670
rect 206328 18470 206548 19678
rect 206300 18454 206560 18470
rect 206300 18236 206328 18454
rect 206546 18236 206560 18454
rect 206300 18216 206560 18236
rect 209328 18098 209548 19652
rect 212328 18884 212548 19634
rect 212328 18664 214124 18884
rect 213128 18098 213386 18108
rect 209328 17880 213156 18098
rect 213374 17880 213386 18098
rect 209328 17878 213386 17880
rect 213128 17848 213386 17878
rect 206974 17752 207242 17790
rect 203328 17750 207242 17752
rect 203328 17532 207000 17750
rect 207218 17532 207242 17750
rect 206974 17516 207242 17532
rect 213904 17278 214124 18664
rect 215328 18576 215548 19666
rect 218328 18894 218548 19678
rect 218328 18674 220908 18894
rect 215300 18562 215570 18576
rect 215300 18344 215328 18562
rect 215546 18344 215570 18562
rect 215300 18338 215570 18344
rect 213898 17268 214144 17278
rect 213898 17050 213904 17268
rect 214122 17050 214144 17268
rect 220688 17238 220908 18674
rect 221328 17730 221548 19666
rect 224328 18428 224548 19656
rect 227328 18940 227548 19674
rect 229636 18940 229916 18952
rect 227328 18938 229916 18940
rect 227328 18720 229658 18938
rect 229876 18720 229916 18938
rect 229636 18700 229916 18720
rect 227174 18428 227460 18436
rect 224328 18210 227194 18428
rect 227412 18210 227460 18428
rect 224328 18208 227460 18210
rect 227174 18192 227460 18208
rect 230328 18304 230548 19648
rect 233328 18702 233548 19678
rect 233310 18688 233574 18702
rect 233310 18470 233328 18688
rect 233546 18470 233574 18688
rect 233310 18442 233574 18470
rect 234638 18304 234884 18322
rect 230328 18302 234884 18304
rect 230328 18084 234650 18302
rect 234868 18084 234884 18302
rect 234638 18062 234884 18084
rect 236328 18016 236548 19498
rect 239328 18534 239548 19610
rect 242328 18578 242548 19678
rect 245328 18598 245548 19678
rect 248328 19090 248548 19654
rect 248328 18870 249886 19090
rect 242314 18570 242552 18578
rect 241664 18534 241902 18544
rect 239328 18316 241672 18534
rect 241890 18316 241902 18534
rect 242314 18352 242328 18570
rect 242546 18352 242552 18570
rect 245328 18378 248930 18598
rect 242314 18346 242552 18352
rect 239328 18314 241902 18316
rect 241664 18312 241902 18314
rect 240890 18016 241174 18054
rect 236328 18014 241174 18016
rect 236328 17796 240916 18014
rect 241134 17796 241174 18014
rect 240890 17770 241174 17796
rect 221292 17710 221614 17730
rect 221292 17492 221328 17710
rect 221546 17492 221614 17710
rect 221292 17460 221614 17492
rect 213898 17032 214144 17050
rect 220666 17228 220962 17238
rect 220666 17010 220688 17228
rect 220906 17010 220962 17228
rect 248710 17090 248930 18378
rect 249666 17866 249886 18870
rect 251328 18510 251548 19678
rect 254328 18736 254548 19678
rect 254314 18700 254612 18736
rect 253898 18510 254148 18520
rect 251328 18508 254148 18510
rect 251328 18290 253926 18508
rect 254144 18290 254148 18508
rect 254314 18482 254328 18700
rect 254546 18482 254612 18700
rect 254314 18462 254612 18482
rect 257328 18576 257548 19670
rect 260328 19116 260548 19678
rect 260328 18896 261264 19116
rect 257328 18356 260272 18576
rect 253898 18276 254148 18290
rect 249648 17860 249898 17866
rect 249648 17642 249668 17860
rect 249886 17642 249898 17860
rect 249648 17622 249898 17642
rect 260052 17258 260272 18356
rect 261044 18136 261264 18896
rect 261022 18124 261294 18136
rect 261022 17906 261044 18124
rect 261262 17906 261294 18124
rect 261022 17878 261294 17906
rect 263328 17964 263548 19678
rect 266328 18560 266548 19620
rect 268990 18560 269262 18570
rect 266328 18342 269032 18560
rect 269250 18342 269262 18560
rect 266328 18340 269262 18342
rect 268990 18312 269262 18340
rect 269328 18292 269548 19594
rect 269322 18268 269594 18292
rect 269322 18050 269328 18268
rect 269546 18050 269594 18268
rect 269322 18034 269594 18050
rect 265852 17964 266124 17980
rect 263328 17962 266146 17964
rect 263328 17744 265870 17962
rect 266088 17744 266146 17962
rect 265852 17722 266124 17744
rect 272328 17582 272548 19648
rect 275328 18206 275548 19648
rect 278328 18698 278548 19670
rect 279642 18698 279942 18730
rect 278328 18480 279676 18698
rect 279894 18480 279942 18698
rect 278328 18478 279942 18480
rect 279642 18444 279942 18478
rect 278800 18206 279208 18308
rect 275328 17988 278878 18206
rect 279096 17988 279208 18206
rect 275328 17986 279208 17988
rect 278800 17946 279208 17986
rect 277670 17582 277952 17624
rect 272328 17364 277694 17582
rect 277912 17364 277952 17582
rect 272328 17362 277952 17364
rect 277670 17336 277952 17362
rect 281328 17512 281548 19678
rect 284328 18176 284548 19678
rect 287328 18228 287548 19670
rect 290328 18982 290548 19678
rect 290286 18954 290586 18982
rect 290286 18736 290328 18954
rect 290546 18736 290586 18954
rect 290286 18696 290586 18736
rect 292376 18228 292676 18260
rect 287328 18226 292676 18228
rect 284308 18136 284608 18176
rect 284308 17918 284328 18136
rect 284546 17918 284608 18136
rect 287328 18008 292408 18226
rect 292626 18008 292676 18226
rect 292376 17974 292676 18008
rect 284308 17890 284608 17918
rect 293328 17724 293548 19642
rect 296328 18328 296548 19654
rect 299328 19100 299548 19678
rect 305362 19100 305616 19106
rect 299328 19098 305616 19100
rect 299328 18880 305386 19098
rect 305604 18880 305616 19098
rect 305362 18850 305616 18880
rect 303267 18717 303269 18718
rect 303268 18395 303269 18717
rect 303267 18394 303269 18395
rect 296328 18108 300470 18328
rect 299228 17724 299528 17758
rect 293328 17722 299528 17724
rect 286910 17512 287210 17550
rect 281328 17294 286930 17512
rect 287148 17294 287210 17512
rect 293328 17504 299258 17722
rect 299476 17504 299528 17722
rect 299228 17472 299528 17504
rect 281328 17292 287210 17294
rect 286910 17264 287210 17292
rect 260030 17246 260302 17258
rect 220666 17000 220962 17010
rect 248702 17076 248952 17090
rect 193426 16768 193720 16800
rect 201984 16894 202244 16902
rect -4334 13976 -4224 16686
rect 201984 16676 202004 16894
rect 202222 16676 202244 16894
rect 248702 16858 248712 17076
rect 248930 16858 248952 17076
rect 260030 17028 260054 17246
rect 260272 17028 260302 17246
rect 300250 17140 300470 18108
rect 303866 17264 304186 17288
rect 260030 17000 260302 17028
rect 300208 17104 300508 17140
rect 248702 16846 248952 16858
rect 300208 16886 300252 17104
rect 300470 16886 300508 17104
rect 300208 16854 300508 16886
rect 303866 16992 303890 17264
rect 304162 16992 304186 17264
rect 201984 16656 202244 16676
rect 302888 16410 303316 16448
rect 302888 16088 302940 16410
rect 303274 16088 303316 16410
rect 302888 16036 303316 16088
rect 303866 15692 304186 16992
rect 26 15642 390 15664
rect 26 15322 48 15642
rect 368 15322 390 15642
rect 303682 15396 303866 15668
rect 26 15298 390 15322
<< via4 >>
rect -5522 321756 -5202 322076
rect -1502 321780 -1230 322052
rect 302448 324538 302768 324598
rect 302448 324338 302502 324538
rect 302502 324338 302712 324538
rect 302712 324338 302768 324538
rect 302448 324278 302768 324338
rect 303950 321062 304222 321334
rect -6294 319800 -5974 320120
rect -3762 319800 -3442 320120
rect -2994 319662 -2674 319982
rect -5522 318756 -5202 319076
rect -1502 318780 -1230 319052
rect 303950 318062 304222 318334
rect -6294 316800 -5974 317120
rect -3762 316800 -3442 317120
rect -2994 316662 -2674 316982
rect -5522 315756 -5202 316076
rect -1502 315780 -1230 316052
rect 303950 315062 304222 315334
rect -6294 313800 -5974 314120
rect -3762 313800 -3442 314120
rect -2994 313662 -2674 313982
rect -5522 312756 -5202 313076
rect -1502 312780 -1230 313052
rect 303950 312062 304222 312334
rect -6294 310800 -5974 311120
rect -3762 310800 -3442 311120
rect -2994 310662 -2674 310982
rect -5522 309756 -5202 310076
rect -1502 309780 -1230 310052
rect 303950 309062 304222 309334
rect -6294 307800 -5974 308120
rect -3762 307800 -3442 308120
rect -2994 307662 -2674 307982
rect -5522 306756 -5202 307076
rect -1502 306780 -1230 307052
rect 303950 306062 304222 306334
rect -6294 304800 -5974 305120
rect -3762 304800 -3442 305120
rect -2994 304662 -2674 304982
rect -5522 303756 -5202 304076
rect -1502 303780 -1230 304052
rect 303950 303062 304222 303334
rect -6294 301800 -5974 302120
rect -3762 301800 -3442 302120
rect -2994 301662 -2674 301982
rect -5522 300756 -5202 301076
rect -1502 300780 -1230 301052
rect 303950 300062 304222 300334
rect -6294 298800 -5974 299120
rect -3762 298800 -3442 299120
rect -2994 298662 -2674 298982
rect -5522 297756 -5202 298076
rect -1502 297780 -1230 298052
rect 303950 297062 304222 297334
rect -6294 295800 -5974 296120
rect -3762 295800 -3442 296120
rect -2994 295662 -2674 295982
rect -5522 294756 -5202 295076
rect -1502 294780 -1230 295052
rect 303950 294062 304222 294334
rect -6294 292800 -5974 293120
rect -3762 292800 -3442 293120
rect -2994 292662 -2674 292982
rect -5522 291756 -5202 292076
rect -1502 291780 -1230 292052
rect 303950 291062 304222 291334
rect -6294 289800 -5974 290120
rect -3762 289800 -3442 290120
rect -2994 289662 -2674 289982
rect -5522 288756 -5202 289076
rect -1502 288780 -1230 289052
rect 303950 288062 304222 288334
rect -6294 286800 -5974 287120
rect -3762 286800 -3442 287120
rect -2994 286662 -2674 286982
rect -5522 285756 -5202 286076
rect -1502 285780 -1230 286052
rect 303950 285062 304222 285334
rect -6294 283800 -5974 284120
rect -3762 283800 -3442 284120
rect -2994 283662 -2674 283982
rect -5522 282756 -5202 283076
rect -1502 282780 -1230 283052
rect 303950 282062 304222 282334
rect -6294 280800 -5974 281120
rect -3762 280800 -3442 281120
rect -2994 280662 -2674 280982
rect -5522 279756 -5202 280076
rect -1502 279780 -1230 280052
rect 303950 279062 304222 279334
rect -6294 277800 -5974 278120
rect -3762 277800 -3442 278120
rect -2994 277662 -2674 277982
rect -5522 276756 -5202 277076
rect -1502 276780 -1230 277052
rect 303950 276062 304222 276334
rect -6294 274800 -5974 275120
rect -3762 274800 -3442 275120
rect -2994 274662 -2674 274982
rect -5522 273756 -5202 274076
rect -1502 273780 -1230 274052
rect 303950 273062 304222 273334
rect -6294 271800 -5974 272120
rect -3762 271800 -3442 272120
rect -2994 271662 -2674 271982
rect -5522 270756 -5202 271076
rect -1502 270780 -1230 271052
rect 303950 270062 304222 270334
rect -6294 268800 -5974 269120
rect -3762 268800 -3442 269120
rect -2994 268662 -2674 268982
rect -5522 267756 -5202 268076
rect -1502 267780 -1230 268052
rect 303950 267062 304222 267334
rect -6294 265800 -5974 266120
rect -3762 265800 -3442 266120
rect -2994 265662 -2674 265982
rect -5522 264756 -5202 265076
rect -1502 264780 -1230 265052
rect 303950 264062 304222 264334
rect -6294 262800 -5974 263120
rect -3762 262800 -3442 263120
rect -2994 262662 -2674 262982
rect -5522 261756 -5202 262076
rect -1502 261780 -1230 262052
rect 303950 261062 304222 261334
rect -6294 259800 -5974 260120
rect -3762 259800 -3442 260120
rect -2994 259662 -2674 259982
rect -5522 258756 -5202 259076
rect -1502 258780 -1230 259052
rect 303950 258062 304222 258334
rect -6294 256800 -5974 257120
rect -3762 256800 -3442 257120
rect -2994 256662 -2674 256982
rect -5522 255756 -5202 256076
rect -1502 255780 -1230 256052
rect 303950 255062 304222 255334
rect -6294 253800 -5974 254120
rect -3762 253800 -3442 254120
rect -2994 253662 -2674 253982
rect -5522 252756 -5202 253076
rect -1502 252780 -1230 253052
rect 303950 252062 304222 252334
rect -6294 250800 -5974 251120
rect -3762 250800 -3442 251120
rect -2994 250662 -2674 250982
rect -5522 249756 -5202 250076
rect -1502 249780 -1230 250052
rect 303950 249062 304222 249334
rect -6294 247800 -5974 248120
rect -3762 247800 -3442 248120
rect -2994 247662 -2674 247982
rect 303950 246062 304222 246334
rect -6294 244800 -5974 245120
rect -3762 244800 -3442 245120
rect -2994 244662 -2674 244982
rect -5522 243756 -5202 244076
rect -1502 243780 -1230 244052
rect 303950 243062 304222 243334
rect -6294 241800 -5974 242120
rect -3762 241800 -3442 242120
rect -2994 241662 -2674 241982
rect -5522 240756 -5202 241076
rect -1502 240780 -1230 241052
rect 303950 240062 304222 240334
rect -6294 238800 -5974 239120
rect -3762 238800 -3442 239120
rect -2994 238662 -2674 238982
rect -5522 237756 -5202 238076
rect -1502 237780 -1230 238052
rect 303950 237062 304222 237334
rect -6294 235800 -5974 236120
rect -3762 235800 -3442 236120
rect -2994 235662 -2674 235982
rect -5522 234756 -5202 235076
rect -1502 234780 -1230 235052
rect 303950 234062 304222 234334
rect -6294 232800 -5974 233120
rect -3762 232800 -3442 233120
rect -2994 232662 -2674 232982
rect -5522 231756 -5202 232076
rect -1502 231780 -1230 232052
rect 303950 231062 304222 231334
rect -6294 229800 -5974 230120
rect -3762 229800 -3442 230120
rect -2994 229662 -2674 229982
rect -5522 228756 -5202 229076
rect -1502 228780 -1230 229052
rect 303950 228062 304222 228334
rect -6294 226800 -5974 227120
rect -3762 226800 -3442 227120
rect -2994 226662 -2674 226982
rect -5522 225756 -5202 226076
rect -1502 225780 -1230 226052
rect 303950 225062 304222 225334
rect -6294 223800 -5974 224120
rect -3762 223800 -3442 224120
rect -2994 223662 -2674 223982
rect -5522 222756 -5202 223076
rect -1502 222780 -1230 223052
rect 303950 222062 304222 222334
rect -6294 220800 -5974 221120
rect -3762 220800 -3442 221120
rect -2994 220662 -2674 220982
rect -5522 219756 -5202 220076
rect -1502 219780 -1230 220052
rect 303950 219062 304222 219334
rect -6294 217800 -5974 218120
rect -3762 217800 -3442 218120
rect -2994 217662 -2674 217982
rect -5522 216756 -5202 217076
rect -1502 216780 -1230 217052
rect 303950 216062 304222 216334
rect -6294 214800 -5974 215120
rect -3762 214800 -3442 215120
rect -2994 214662 -2674 214982
rect -5522 213756 -5202 214076
rect -1502 213780 -1230 214052
rect 303950 213062 304222 213334
rect -6294 211800 -5974 212120
rect -3762 211800 -3442 212120
rect -2994 211662 -2674 211982
rect -5522 210756 -5202 211076
rect -1502 210780 -1230 211052
rect 303950 210062 304222 210334
rect -2994 208662 -2674 208982
rect -5522 207756 -5202 208076
rect -1502 207780 -1230 208052
rect 303950 207062 304222 207334
rect -6294 205800 -5974 206120
rect -3762 205800 -3442 206120
rect -2994 205662 -2674 205982
rect -5522 204756 -5202 205076
rect -1502 204780 -1230 205052
rect 303950 204062 304222 204334
rect -6294 202800 -5974 203120
rect -3762 202800 -3442 203120
rect -2994 202662 -2674 202982
rect -5522 201756 -5202 202076
rect -1502 201780 -1230 202052
rect 303950 201062 304222 201334
rect -6294 199800 -5974 200120
rect -3762 199800 -3442 200120
rect -2994 199662 -2674 199982
rect -5522 198756 -5202 199076
rect -1502 198780 -1230 199052
rect 303950 198062 304222 198334
rect -6294 196800 -5974 197120
rect -3762 196800 -3442 197120
rect -2994 196662 -2674 196982
rect -5522 195756 -5202 196076
rect -1502 195780 -1230 196052
rect 303950 195062 304222 195334
rect -6294 193800 -5974 194120
rect -3762 193800 -3442 194120
rect -2994 193662 -2674 193982
rect -5522 192756 -5202 193076
rect -1502 192780 -1230 193052
rect 303950 192062 304222 192334
rect -6294 190800 -5974 191120
rect -3762 190800 -3442 191120
rect -2994 190662 -2674 190982
rect -5522 189756 -5202 190076
rect -1502 189780 -1230 190052
rect 303950 189062 304222 189334
rect -6294 187800 -5974 188120
rect -3762 187800 -3442 188120
rect -2994 187662 -2674 187982
rect -5522 186756 -5202 187076
rect -1502 186780 -1230 187052
rect 303950 186062 304222 186334
rect -6294 184800 -5974 185120
rect -3762 184800 -3442 185120
rect -2994 184662 -2674 184982
rect -5522 183756 -5202 184076
rect -1502 183780 -1230 184052
rect 303950 183062 304222 183334
rect -6294 181800 -5974 182120
rect -3762 181800 -3442 182120
rect -2994 181662 -2674 181982
rect -5522 180756 -5202 181076
rect -1502 180780 -1230 181052
rect 303950 180062 304222 180334
rect -6294 178800 -5974 179120
rect -3762 178800 -3442 179120
rect -2994 178662 -2674 178982
rect -5522 177756 -5202 178076
rect -1502 177780 -1230 178052
rect 303950 177062 304222 177334
rect -6294 175800 -5974 176120
rect -3762 175800 -3442 176120
rect -2994 175662 -2674 175982
rect -5522 174756 -5202 175076
rect -1502 174780 -1230 175052
rect 303950 174062 304222 174334
rect -6294 172800 -5974 173120
rect -3762 172800 -3442 173120
rect -2994 172662 -2674 172982
rect -5522 171756 -5202 172076
rect -1502 171780 -1230 172052
rect 303950 171062 304222 171334
rect -6294 169800 -5974 170120
rect -3762 169800 -3442 170120
rect -2994 169662 -2674 169982
rect -5522 168756 -5202 169076
rect -1502 168780 -1230 169052
rect 303950 168062 304222 168334
rect -6294 166800 -5974 167120
rect -3762 166800 -3442 167120
rect -2994 166662 -2674 166982
rect -5522 165756 -5202 166076
rect -1502 165780 -1230 166052
rect 303950 165062 304222 165334
rect -6294 163800 -5974 164120
rect -3762 163800 -3442 164120
rect -2994 163662 -2674 163982
rect -5522 162756 -5202 163076
rect -1502 162780 -1230 163052
rect 303950 162062 304222 162334
rect -6294 160800 -5974 161120
rect -3762 160800 -3442 161120
rect -2994 160662 -2674 160982
rect -5522 159756 -5202 160076
rect -1502 159780 -1230 160052
rect 303950 159062 304222 159334
rect -6294 157800 -5974 158120
rect -3762 157800 -3442 158120
rect -2994 157662 -2674 157982
rect -5522 156756 -5202 157076
rect -1502 156780 -1230 157052
rect 303950 156062 304222 156334
rect -6294 154800 -5974 155120
rect -3762 154800 -3442 155120
rect -2994 154662 -2674 154982
rect -5522 153756 -5202 154076
rect -1502 153780 -1230 154052
rect 303950 153062 304222 153334
rect -6294 151800 -5974 152120
rect -3762 151800 -3442 152120
rect -2994 151662 -2674 151982
rect -5522 150756 -5202 151076
rect -1502 150780 -1230 151052
rect 303950 150062 304222 150334
rect -6294 148800 -5974 149120
rect -3762 148800 -3442 149120
rect -2994 148662 -2674 148982
rect -5522 147756 -5202 148076
rect -1502 147780 -1230 148052
rect 303950 147062 304222 147334
rect -6294 145800 -5974 146120
rect -3762 145800 -3442 146120
rect -2994 145662 -2674 145982
rect -5522 144756 -5202 145076
rect -1502 144780 -1230 145052
rect 303950 144062 304222 144334
rect -6294 142800 -5974 143120
rect -3762 142800 -3442 143120
rect -2994 142662 -2674 142982
rect -5522 141756 -5202 142076
rect -1502 141780 -1230 142052
rect 303950 141062 304222 141334
rect -6294 139800 -5974 140120
rect -3762 139800 -3442 140120
rect -2994 139662 -2674 139982
rect -5522 138756 -5202 139076
rect -1502 138780 -1230 139052
rect 303950 138062 304222 138334
rect -6294 136800 -5974 137120
rect -3762 136800 -3442 137120
rect -2994 136662 -2674 136982
rect -5522 135756 -5202 136076
rect -1502 135780 -1230 136052
rect 303950 135062 304222 135334
rect -6294 133800 -5974 134120
rect -3762 133800 -3442 134120
rect -2994 133662 -2674 133982
rect -5522 132756 -5202 133076
rect -1502 132780 -1230 133052
rect 303950 132062 304222 132334
rect -6294 130800 -5974 131120
rect -3762 130800 -3442 131120
rect -2994 130662 -2674 130982
rect -5522 129756 -5202 130076
rect -1502 129780 -1230 130052
rect 303950 129062 304222 129334
rect -6294 127800 -5974 128120
rect -3762 127800 -3442 128120
rect -2994 127662 -2674 127982
rect -5522 126756 -5202 127076
rect -1502 126780 -1230 127052
rect 303950 126062 304222 126334
rect -6294 124800 -5974 125120
rect -3762 124800 -3442 125120
rect -2994 124662 -2674 124982
rect -5522 123756 -5202 124076
rect -1502 123780 -1230 124052
rect 303950 123062 304222 123334
rect -6294 121800 -5974 122120
rect -3762 121800 -3442 122120
rect -2994 121662 -2674 121982
rect -5522 120756 -5202 121076
rect -1502 120780 -1230 121052
rect 303950 120062 304222 120334
rect -6294 118800 -5974 119120
rect -3762 118800 -3442 119120
rect -2994 118662 -2674 118982
rect -5522 117756 -5202 118076
rect -1502 117780 -1230 118052
rect 303950 117062 304222 117334
rect -6294 115800 -5974 116120
rect -3762 115800 -3442 116120
rect -2994 115662 -2674 115982
rect -5522 114756 -5202 115076
rect -1502 114780 -1230 115052
rect 303950 114062 304222 114334
rect -6294 112800 -5974 113120
rect -3762 112800 -3442 113120
rect -2994 112662 -2674 112982
rect -5522 111756 -5202 112076
rect -1502 111780 -1230 112052
rect 303950 111062 304222 111334
rect -6294 109800 -5974 110120
rect -3762 109800 -3442 110120
rect -2994 109662 -2674 109982
rect -5522 108756 -5202 109076
rect -1502 108780 -1230 109052
rect 303950 108062 304222 108334
rect -6294 106800 -5974 107120
rect -3762 106800 -3442 107120
rect -2994 106662 -2674 106982
rect -5522 105756 -5202 106076
rect -1502 105780 -1230 106052
rect 303950 105062 304222 105334
rect -6294 103800 -5974 104120
rect -3762 103800 -3442 104120
rect -2994 103662 -2674 103982
rect -5522 102756 -5202 103076
rect -1502 102780 -1230 103052
rect 303950 102062 304222 102334
rect -6294 100800 -5974 101120
rect -3762 100800 -3442 101120
rect -2994 100662 -2674 100982
rect -5522 99756 -5202 100076
rect -1502 99780 -1230 100052
rect 303950 99062 304222 99334
rect -6294 97800 -5974 98120
rect -3762 97800 -3442 98120
rect -2994 97662 -2674 97982
rect -5522 96756 -5202 97076
rect -1502 96780 -1230 97052
rect 303950 96062 304222 96334
rect -6294 94800 -5974 95120
rect -3762 94800 -3442 95120
rect -2994 94662 -2674 94982
rect 303950 93062 304222 93334
rect -6294 91800 -5974 92120
rect -3762 91800 -3442 92120
rect -2994 91662 -2674 91982
rect -5522 90756 -5202 91076
rect -1502 90780 -1230 91052
rect 303950 90062 304222 90334
rect -6294 88800 -5974 89120
rect -3762 88800 -3442 89120
rect -2994 88662 -2674 88982
rect -5522 87756 -5202 88076
rect -1502 87780 -1230 88052
rect 303950 87062 304222 87334
rect -6294 85800 -5974 86120
rect -3762 85800 -3442 86120
rect -2994 85662 -2674 85982
rect -5522 84756 -5202 85076
rect -1502 84780 -1230 85052
rect 303950 84062 304222 84334
rect -6294 82800 -5974 83120
rect -3762 82800 -3442 83120
rect -2994 82662 -2674 82982
rect -5522 81756 -5202 82076
rect -1502 81780 -1230 82052
rect 303950 81062 304222 81334
rect -6294 79800 -5974 80120
rect -3762 79800 -3442 80120
rect -2994 79662 -2674 79982
rect -5522 78756 -5202 79076
rect -1502 78780 -1230 79052
rect 303950 78062 304222 78334
rect -6294 76800 -5974 77120
rect -3762 76800 -3442 77120
rect -2994 76662 -2674 76982
rect -5522 75756 -5202 76076
rect -1502 75780 -1230 76052
rect 303950 75062 304222 75334
rect -6294 73800 -5974 74120
rect -3762 73800 -3442 74120
rect -2994 73662 -2674 73982
rect -5522 72756 -5202 73076
rect -1502 72780 -1230 73052
rect 303950 72062 304222 72334
rect -6294 70800 -5974 71120
rect -3762 70800 -3442 71120
rect -2994 70662 -2674 70982
rect -5522 69756 -5202 70076
rect -1502 69780 -1230 70052
rect 303950 69062 304222 69334
rect -6294 67800 -5974 68120
rect -3762 67800 -3442 68120
rect -2994 67662 -2674 67982
rect -5522 66756 -5202 67076
rect -1502 66780 -1230 67052
rect 303950 66062 304222 66334
rect -6294 64800 -5974 65120
rect -3762 64800 -3442 65120
rect -2994 64662 -2674 64982
rect -5522 63756 -5202 64076
rect -1502 63780 -1230 64052
rect 303950 63062 304222 63334
rect -6294 61800 -5974 62120
rect -3762 61800 -3442 62120
rect -2994 61662 -2674 61982
rect -5522 60756 -5202 61076
rect -1502 60780 -1230 61052
rect 303950 60062 304222 60334
rect -6294 58800 -5974 59120
rect -3762 58800 -3442 59120
rect -2994 58662 -2674 58982
rect -5522 57756 -5202 58076
rect -1502 57780 -1230 58052
rect 303950 57062 304222 57334
rect -2994 55662 -2674 55982
rect -5522 54756 -5202 55076
rect -1502 54780 -1230 55052
rect 303950 54062 304222 54334
rect -6294 52800 -5974 53120
rect -3762 52800 -3442 53120
rect -2994 52662 -2674 52982
rect -5522 51756 -5202 52076
rect -1502 51780 -1230 52052
rect 303950 51062 304222 51334
rect -6294 49800 -5974 50120
rect -3762 49800 -3442 50120
rect -2994 49662 -2674 49982
rect -5522 48756 -5202 49076
rect -1502 48780 -1230 49052
rect 303950 48062 304222 48334
rect -6294 46800 -5974 47120
rect -3762 46800 -3442 47120
rect -2994 46662 -2674 46982
rect -5522 45756 -5202 46076
rect -1502 45780 -1230 46052
rect 303950 45062 304222 45334
rect -6294 43800 -5974 44120
rect -3762 43800 -3442 44120
rect -2994 43662 -2674 43982
rect -5522 42756 -5202 43076
rect -1502 42780 -1230 43052
rect 303950 42062 304222 42334
rect -6294 40800 -5974 41120
rect -3762 40800 -3442 41120
rect -2994 40662 -2674 40982
rect -5522 39756 -5202 40076
rect -1502 39780 -1230 40052
rect 303950 39062 304222 39334
rect -6294 37800 -5974 38120
rect -3762 37800 -3442 38120
rect -2994 37662 -2674 37982
rect -5522 36756 -5202 37076
rect -1502 36780 -1230 37052
rect 303950 36062 304222 36334
rect -6294 34800 -5974 35120
rect -3762 34800 -3442 35120
rect -2994 34662 -2674 34982
rect -5522 33756 -5202 34076
rect -1502 33780 -1230 34052
rect 303950 33062 304222 33334
rect -6294 31800 -5974 32120
rect -3762 31800 -3442 32120
rect -2994 31662 -2674 31982
rect -5522 30756 -5202 31076
rect -1502 30780 -1230 31052
rect 303950 30062 304222 30334
rect -6294 28800 -5974 29120
rect -3762 28800 -3442 29120
rect -2994 28662 -2674 28982
rect -5522 27756 -5202 28076
rect -1502 27780 -1230 28052
rect 303950 27062 304222 27334
rect -6294 25800 -5974 26120
rect -3762 25800 -3442 26120
rect -2994 25662 -2674 25982
rect -5522 24756 -5202 25076
rect -1502 24780 -1230 25052
rect 303950 24062 304222 24334
rect -6294 22800 -5974 23120
rect -3762 22800 -3442 23120
rect -2994 22662 -2674 22982
rect -5522 21756 -5202 22076
rect -1502 21780 -1230 22052
rect 303950 21062 304222 21334
rect -6294 19800 -5974 20120
rect -3762 19800 -3442 20120
rect -5522 18756 -5202 19076
rect -1502 18780 -1230 19052
rect -6414 17942 -6094 18002
rect -6414 17742 -6204 17942
rect -6204 17742 -6094 17942
rect -6414 17682 -6094 17742
rect 302945 18717 303267 18718
rect 302945 18395 302946 18717
rect 302946 18395 303267 18717
rect 302945 18394 303267 18395
rect 303890 16992 304162 17264
rect 302940 16088 302942 16410
rect 302942 16088 303274 16410
rect 48 15582 368 15642
rect 48 15382 102 15582
rect 102 15382 312 15582
rect 312 15382 368 15582
rect 48 15322 368 15382
rect 303866 15372 304186 15692
<< metal5 >>
rect -2946 326542 -2626 326564
rect -1526 326542 -1206 326564
rect -2946 326222 305854 326542
rect -5546 322076 -5178 322100
rect -5546 321756 -5522 322076
rect -5202 321756 -5178 322076
rect -5546 321732 -5178 321756
rect -6318 320120 -5950 320144
rect -6318 319800 -6294 320120
rect -5974 319800 -5950 320120
rect -6318 319776 -5950 319800
rect -3786 320120 -3418 320144
rect -2946 320120 -2626 326222
rect -1526 326068 -1206 326222
rect -1526 324636 -1206 324684
rect 302448 324636 302768 324994
rect -1928 324598 304434 324636
rect -1928 324316 302448 324598
rect -3786 319800 -3762 320120
rect -3442 319982 -2626 320120
rect -3442 319800 -2994 319982
rect -3786 319776 -3418 319800
rect -3018 319662 -2994 319800
rect -2674 319662 -2626 319982
rect -3018 319638 -2626 319662
rect -5546 319076 -5178 319100
rect -5546 318756 -5522 319076
rect -5202 318756 -5178 319076
rect -5546 318732 -5178 318756
rect -6318 317120 -5950 317144
rect -6318 316800 -6294 317120
rect -5974 316800 -5950 317120
rect -6318 316776 -5950 316800
rect -3786 317120 -3418 317144
rect -2946 317120 -2626 319638
rect -3786 316800 -3762 317120
rect -3442 316982 -2626 317120
rect -3442 316800 -2994 316982
rect -3786 316776 -3418 316800
rect -3018 316662 -2994 316800
rect -2674 316662 -2626 316982
rect -1526 322052 -1206 324316
rect 302424 324278 302448 324316
rect 302768 324316 304434 324598
rect 302768 324278 302792 324316
rect 302424 324254 302792 324278
rect 303926 322140 304246 324316
rect -1526 321780 -1502 322052
rect -1230 321780 -1206 322052
rect -1526 319052 -1206 321780
rect 303888 321334 304300 322140
rect 303888 321062 303950 321334
rect 304222 321062 304300 321334
rect 288 320218 854 320538
rect -1526 318780 -1502 319052
rect -1230 318780 -1206 319052
rect -1526 316960 -1206 318780
rect -3018 316638 -2626 316662
rect -1528 316640 -1206 316960
rect -5546 316076 -5178 316100
rect -5546 315756 -5522 316076
rect -5202 315756 -5178 316076
rect -5546 315732 -5178 315756
rect -6318 314120 -5950 314144
rect -6318 313800 -6294 314120
rect -5974 313800 -5950 314120
rect -6318 313776 -5950 313800
rect -3786 314120 -3418 314144
rect -2946 314120 -2626 316638
rect -3786 313800 -3762 314120
rect -3442 313982 -2626 314120
rect -3442 313800 -2994 313982
rect -3786 313776 -3418 313800
rect -3018 313662 -2994 313800
rect -2674 313662 -2626 313982
rect -1526 316052 -1206 316640
rect -1526 315780 -1502 316052
rect -1230 315780 -1206 316052
rect -1526 313960 -1206 315780
rect -3018 313638 -2626 313662
rect -1528 313640 -1206 313960
rect -5546 313076 -5178 313100
rect -5546 312756 -5522 313076
rect -5202 312756 -5178 313076
rect -5546 312732 -5178 312756
rect -6318 311120 -5950 311144
rect -6318 310800 -6294 311120
rect -5974 310800 -5950 311120
rect -6318 310776 -5950 310800
rect -3786 311120 -3418 311144
rect -2946 311120 -2626 313638
rect -3786 310800 -3762 311120
rect -3442 310982 -2626 311120
rect -3442 310800 -2994 310982
rect -3786 310776 -3418 310800
rect -3018 310662 -2994 310800
rect -2674 310662 -2626 310982
rect -1526 313052 -1206 313640
rect -1526 312780 -1502 313052
rect -1230 312780 -1206 313052
rect -1526 310960 -1206 312780
rect -3018 310638 -2626 310662
rect -1528 310640 -1206 310960
rect -5546 310076 -5178 310100
rect -5546 309756 -5522 310076
rect -5202 309756 -5178 310076
rect -5546 309732 -5178 309756
rect -6318 308120 -5950 308144
rect -6318 307800 -6294 308120
rect -5974 307800 -5950 308120
rect -6318 307776 -5950 307800
rect -3786 308120 -3418 308144
rect -2946 308120 -2626 310638
rect -3786 307800 -3762 308120
rect -3442 307982 -2626 308120
rect -3442 307800 -2994 307982
rect -3786 307776 -3418 307800
rect -3018 307662 -2994 307800
rect -2674 307662 -2626 307982
rect -1526 310052 -1206 310640
rect -1526 309780 -1502 310052
rect -1230 309780 -1206 310052
rect -1526 307960 -1206 309780
rect -3018 307638 -2626 307662
rect -1528 307640 -1206 307960
rect -5546 307076 -5178 307100
rect -5546 306756 -5522 307076
rect -5202 306756 -5178 307076
rect -5546 306732 -5178 306756
rect -6318 305120 -5950 305144
rect -6318 304800 -6294 305120
rect -5974 304800 -5950 305120
rect -6318 304776 -5950 304800
rect -3786 305120 -3418 305144
rect -2946 305120 -2626 307638
rect -3786 304800 -3762 305120
rect -3442 304982 -2626 305120
rect -3442 304800 -2994 304982
rect -3786 304776 -3418 304800
rect -3018 304662 -2994 304800
rect -2674 304662 -2626 304982
rect -1526 307052 -1206 307640
rect -1526 306780 -1502 307052
rect -1230 306780 -1206 307052
rect -1526 304960 -1206 306780
rect -3018 304638 -2626 304662
rect -1528 304640 -1206 304960
rect -5546 304076 -5178 304100
rect -5546 303756 -5522 304076
rect -5202 303756 -5178 304076
rect -5546 303732 -5178 303756
rect -6318 302120 -5950 302144
rect -6318 301800 -6294 302120
rect -5974 301800 -5950 302120
rect -6318 301776 -5950 301800
rect -3786 302120 -3418 302144
rect -2946 302120 -2626 304638
rect -3786 301800 -3762 302120
rect -3442 301982 -2626 302120
rect -3442 301800 -2994 301982
rect -3786 301776 -3418 301800
rect -3018 301662 -2994 301800
rect -2674 301662 -2626 301982
rect -1526 304052 -1206 304640
rect -1526 303780 -1502 304052
rect -1230 303780 -1206 304052
rect -1526 301960 -1206 303780
rect -3018 301638 -2626 301662
rect -1528 301640 -1206 301960
rect -5546 301076 -5178 301100
rect -5546 300756 -5522 301076
rect -5202 300756 -5178 301076
rect -5546 300732 -5178 300756
rect -6318 299120 -5950 299144
rect -6318 298800 -6294 299120
rect -5974 298800 -5950 299120
rect -6318 298776 -5950 298800
rect -3786 299120 -3418 299144
rect -2946 299120 -2626 301638
rect -3786 298800 -3762 299120
rect -3442 298982 -2626 299120
rect -3442 298800 -2994 298982
rect -3786 298776 -3418 298800
rect -3018 298662 -2994 298800
rect -2674 298662 -2626 298982
rect -1526 301052 -1206 301640
rect -1526 300780 -1502 301052
rect -1230 300780 -1206 301052
rect -1526 298960 -1206 300780
rect -3018 298638 -2626 298662
rect -1528 298640 -1206 298960
rect -5546 298076 -5178 298100
rect -5546 297756 -5522 298076
rect -5202 297756 -5178 298076
rect -5546 297732 -5178 297756
rect -6318 296120 -5950 296144
rect -6318 295800 -6294 296120
rect -5974 295800 -5950 296120
rect -6318 295776 -5950 295800
rect -3786 296120 -3418 296144
rect -2946 296120 -2626 298638
rect -3786 295800 -3762 296120
rect -3442 295982 -2626 296120
rect -3442 295800 -2994 295982
rect -3786 295776 -3418 295800
rect -3018 295662 -2994 295800
rect -2674 295662 -2626 295982
rect -1526 298052 -1206 298640
rect -1526 297780 -1502 298052
rect -1230 297780 -1206 298052
rect -1526 295960 -1206 297780
rect -3018 295638 -2626 295662
rect -1528 295640 -1206 295960
rect -5546 295076 -5178 295100
rect -5546 294756 -5522 295076
rect -5202 294756 -5178 295076
rect -5546 294732 -5178 294756
rect -6318 293120 -5950 293144
rect -6318 292800 -6294 293120
rect -5974 292800 -5950 293120
rect -6318 292776 -5950 292800
rect -3786 293120 -3418 293144
rect -2946 293120 -2626 295638
rect -3786 292800 -3762 293120
rect -3442 292982 -2626 293120
rect -3442 292800 -2994 292982
rect -3786 292776 -3418 292800
rect -3018 292662 -2994 292800
rect -2674 292662 -2626 292982
rect -1526 295052 -1206 295640
rect -1526 294780 -1502 295052
rect -1230 294780 -1206 295052
rect -1526 292960 -1206 294780
rect -3018 292638 -2626 292662
rect -1528 292640 -1206 292960
rect -5546 292076 -5178 292100
rect -5546 291756 -5522 292076
rect -5202 291756 -5178 292076
rect -5546 291732 -5178 291756
rect -6318 290120 -5950 290144
rect -6318 289800 -6294 290120
rect -5974 289800 -5950 290120
rect -6318 289776 -5950 289800
rect -3786 290120 -3418 290144
rect -2946 290120 -2626 292638
rect -3786 289800 -3762 290120
rect -3442 289982 -2626 290120
rect -3442 289800 -2994 289982
rect -3786 289776 -3418 289800
rect -3018 289662 -2994 289800
rect -2674 289662 -2626 289982
rect -1526 292052 -1206 292640
rect -1526 291780 -1502 292052
rect -1230 291780 -1206 292052
rect -1526 289960 -1206 291780
rect -3018 289638 -2626 289662
rect -1528 289640 -1206 289960
rect -5546 289076 -5178 289100
rect -5546 288756 -5522 289076
rect -5202 288756 -5178 289076
rect -5546 288732 -5178 288756
rect -6318 287120 -5950 287144
rect -6318 286800 -6294 287120
rect -5974 286800 -5950 287120
rect -6318 286776 -5950 286800
rect -3786 287120 -3418 287144
rect -2946 287120 -2626 289638
rect -3786 286800 -3762 287120
rect -3442 286982 -2626 287120
rect -3442 286800 -2994 286982
rect -3786 286776 -3418 286800
rect -3018 286662 -2994 286800
rect -2674 286662 -2626 286982
rect -1526 289052 -1206 289640
rect -1526 288780 -1502 289052
rect -1230 288780 -1206 289052
rect -1526 286960 -1206 288780
rect -3018 286638 -2626 286662
rect -1528 286640 -1206 286960
rect -5546 286076 -5178 286100
rect -5546 285756 -5522 286076
rect -5202 285756 -5178 286076
rect -5546 285732 -5178 285756
rect -6318 284120 -5950 284144
rect -6318 283800 -6294 284120
rect -5974 283800 -5950 284120
rect -6318 283776 -5950 283800
rect -3786 284120 -3418 284144
rect -2946 284120 -2626 286638
rect -3786 283800 -3762 284120
rect -3442 283982 -2626 284120
rect -3442 283800 -2994 283982
rect -3786 283776 -3418 283800
rect -3018 283662 -2994 283800
rect -2674 283662 -2626 283982
rect -1526 286052 -1206 286640
rect -1526 285780 -1502 286052
rect -1230 285780 -1206 286052
rect -1526 283960 -1206 285780
rect -3018 283638 -2626 283662
rect -1528 283640 -1206 283960
rect -5546 283076 -5178 283100
rect -5546 282756 -5522 283076
rect -5202 282756 -5178 283076
rect -5546 282732 -5178 282756
rect -6318 281120 -5950 281144
rect -6318 280800 -6294 281120
rect -5974 280800 -5950 281120
rect -6318 280776 -5950 280800
rect -3786 281120 -3418 281144
rect -2946 281120 -2626 283638
rect -3786 280800 -3762 281120
rect -3442 280982 -2626 281120
rect -3442 280800 -2994 280982
rect -3786 280776 -3418 280800
rect -3018 280662 -2994 280800
rect -2674 280662 -2626 280982
rect -1526 283052 -1206 283640
rect -1526 282780 -1502 283052
rect -1230 282780 -1206 283052
rect -1526 280960 -1206 282780
rect -3018 280638 -2626 280662
rect -1528 280640 -1206 280960
rect -5546 280076 -5178 280100
rect -5546 279756 -5522 280076
rect -5202 279756 -5178 280076
rect -5546 279732 -5178 279756
rect -6318 278120 -5950 278144
rect -6318 277800 -6294 278120
rect -5974 277800 -5950 278120
rect -6318 277776 -5950 277800
rect -3786 278120 -3418 278144
rect -2946 278120 -2626 280638
rect -3786 277800 -3762 278120
rect -3442 277982 -2626 278120
rect -3442 277800 -2994 277982
rect -3786 277776 -3418 277800
rect -3018 277662 -2994 277800
rect -2674 277662 -2626 277982
rect -1526 280052 -1206 280640
rect -1526 279780 -1502 280052
rect -1230 279780 -1206 280052
rect -1526 277960 -1206 279780
rect -3018 277638 -2626 277662
rect -1528 277640 -1206 277960
rect -5546 277076 -5178 277100
rect -5546 276756 -5522 277076
rect -5202 276756 -5178 277076
rect -5546 276732 -5178 276756
rect -6318 275120 -5950 275144
rect -6318 274800 -6294 275120
rect -5974 274800 -5950 275120
rect -6318 274776 -5950 274800
rect -3786 275120 -3418 275144
rect -2946 275120 -2626 277638
rect -3786 274800 -3762 275120
rect -3442 274982 -2626 275120
rect -3442 274800 -2994 274982
rect -3786 274776 -3418 274800
rect -3018 274662 -2994 274800
rect -2674 274662 -2626 274982
rect -1526 277052 -1206 277640
rect -1526 276780 -1502 277052
rect -1230 276780 -1206 277052
rect -1526 274960 -1206 276780
rect -3018 274638 -2626 274662
rect -1528 274640 -1206 274960
rect -5546 274076 -5178 274100
rect -5546 273756 -5522 274076
rect -5202 273756 -5178 274076
rect -5546 273732 -5178 273756
rect -6318 272120 -5950 272144
rect -6318 271800 -6294 272120
rect -5974 271800 -5950 272120
rect -6318 271776 -5950 271800
rect -3786 272120 -3418 272144
rect -2946 272120 -2626 274638
rect -3786 271800 -3762 272120
rect -3442 271982 -2626 272120
rect -3442 271800 -2994 271982
rect -3786 271776 -3418 271800
rect -3018 271662 -2994 271800
rect -2674 271662 -2626 271982
rect -1526 274052 -1206 274640
rect -1526 273780 -1502 274052
rect -1230 273780 -1206 274052
rect -1526 271960 -1206 273780
rect -3018 271638 -2626 271662
rect -1528 271640 -1206 271960
rect -5546 271076 -5178 271100
rect -5546 270756 -5522 271076
rect -5202 270756 -5178 271076
rect -5546 270732 -5178 270756
rect -6318 269120 -5950 269144
rect -6318 268800 -6294 269120
rect -5974 268800 -5950 269120
rect -6318 268776 -5950 268800
rect -3786 269120 -3418 269144
rect -2946 269120 -2626 271638
rect -3786 268800 -3762 269120
rect -3442 268982 -2626 269120
rect -3442 268800 -2994 268982
rect -3786 268776 -3418 268800
rect -3018 268662 -2994 268800
rect -2674 268662 -2626 268982
rect -1526 271052 -1206 271640
rect -1526 270780 -1502 271052
rect -1230 270780 -1206 271052
rect -1526 268960 -1206 270780
rect -3018 268638 -2626 268662
rect -1528 268640 -1206 268960
rect -5546 268076 -5178 268100
rect -5546 267756 -5522 268076
rect -5202 267756 -5178 268076
rect -5546 267732 -5178 267756
rect -6318 266120 -5950 266144
rect -6318 265800 -6294 266120
rect -5974 265800 -5950 266120
rect -6318 265776 -5950 265800
rect -3786 266120 -3418 266144
rect -2946 266120 -2626 268638
rect -3786 265800 -3762 266120
rect -3442 265982 -2626 266120
rect -3442 265800 -2994 265982
rect -3786 265776 -3418 265800
rect -3018 265662 -2994 265800
rect -2674 265662 -2626 265982
rect -1526 268052 -1206 268640
rect -1526 267780 -1502 268052
rect -1230 267780 -1206 268052
rect -1526 265960 -1206 267780
rect -3018 265638 -2626 265662
rect -1528 265640 -1206 265960
rect -5546 265076 -5178 265100
rect -5546 264756 -5522 265076
rect -5202 264756 -5178 265076
rect -5546 264732 -5178 264756
rect -6318 263120 -5950 263144
rect -6318 262800 -6294 263120
rect -5974 262800 -5950 263120
rect -6318 262776 -5950 262800
rect -3786 263120 -3418 263144
rect -2946 263120 -2626 265638
rect -3786 262800 -3762 263120
rect -3442 262982 -2626 263120
rect -3442 262800 -2994 262982
rect -3786 262776 -3418 262800
rect -3018 262662 -2994 262800
rect -2674 262662 -2626 262982
rect -1526 265052 -1206 265640
rect -1526 264780 -1502 265052
rect -1230 264780 -1206 265052
rect -1526 262960 -1206 264780
rect -3018 262638 -2626 262662
rect -1528 262640 -1206 262960
rect -5546 262076 -5178 262100
rect -5546 261756 -5522 262076
rect -5202 261756 -5178 262076
rect -5546 261732 -5178 261756
rect -6318 260120 -5950 260144
rect -6318 259800 -6294 260120
rect -5974 259800 -5950 260120
rect -6318 259776 -5950 259800
rect -3786 260120 -3418 260144
rect -2946 260120 -2626 262638
rect -3786 259800 -3762 260120
rect -3442 259982 -2626 260120
rect -3442 259800 -2994 259982
rect -3786 259776 -3418 259800
rect -3018 259662 -2994 259800
rect -2674 259662 -2626 259982
rect -1526 262052 -1206 262640
rect -1526 261780 -1502 262052
rect -1230 261780 -1206 262052
rect -1526 259960 -1206 261780
rect -3018 259638 -2626 259662
rect -1528 259640 -1206 259960
rect -5546 259076 -5178 259100
rect -5546 258756 -5522 259076
rect -5202 258756 -5178 259076
rect -5546 258732 -5178 258756
rect -6318 257120 -5950 257144
rect -6318 256800 -6294 257120
rect -5974 256800 -5950 257120
rect -6318 256776 -5950 256800
rect -3786 257120 -3418 257144
rect -2946 257120 -2626 259638
rect -3786 256800 -3762 257120
rect -3442 256982 -2626 257120
rect -3442 256800 -2994 256982
rect -3786 256776 -3418 256800
rect -3018 256662 -2994 256800
rect -2674 256662 -2626 256982
rect -1526 259052 -1206 259640
rect -1526 258780 -1502 259052
rect -1230 258780 -1206 259052
rect -1526 256960 -1206 258780
rect -3018 256638 -2626 256662
rect -1528 256640 -1206 256960
rect -5546 256076 -5178 256100
rect -5546 255756 -5522 256076
rect -5202 255756 -5178 256076
rect -5546 255732 -5178 255756
rect -6318 254120 -5950 254144
rect -6318 253800 -6294 254120
rect -5974 253800 -5950 254120
rect -6318 253776 -5950 253800
rect -3786 254120 -3418 254144
rect -2946 254120 -2626 256638
rect -3786 253800 -3762 254120
rect -3442 253982 -2626 254120
rect -3442 253800 -2994 253982
rect -3786 253776 -3418 253800
rect -3018 253662 -2994 253800
rect -2674 253662 -2626 253982
rect -1526 256052 -1206 256640
rect -1526 255780 -1502 256052
rect -1230 255780 -1206 256052
rect -1526 253960 -1206 255780
rect -3018 253638 -2626 253662
rect -1528 253640 -1206 253960
rect -5546 253076 -5178 253100
rect -5546 252756 -5522 253076
rect -5202 252756 -5178 253076
rect -5546 252732 -5178 252756
rect -6318 251120 -5950 251144
rect -6318 250800 -6294 251120
rect -5974 250800 -5950 251120
rect -6318 250776 -5950 250800
rect -3786 251120 -3418 251144
rect -2946 251120 -2626 253638
rect -3786 250800 -3762 251120
rect -3442 250982 -2626 251120
rect -3442 250800 -2994 250982
rect -3786 250776 -3418 250800
rect -3018 250662 -2994 250800
rect -2674 250662 -2626 250982
rect -1526 253052 -1206 253640
rect -1526 252780 -1502 253052
rect -1230 252780 -1206 253052
rect -1526 250960 -1206 252780
rect -3018 250638 -2626 250662
rect -1528 250640 -1206 250960
rect -5546 250076 -5178 250100
rect -5546 249756 -5522 250076
rect -5202 249756 -5178 250076
rect -5546 249732 -5178 249756
rect -6318 248120 -5950 248144
rect -6318 247800 -6294 248120
rect -5974 247800 -5950 248120
rect -6318 247776 -5950 247800
rect -3786 248120 -3418 248144
rect -2946 248120 -2626 250638
rect -3786 247800 -3762 248120
rect -3442 247982 -2626 248120
rect -3442 247800 -2994 247982
rect -3786 247776 -3418 247800
rect -3018 247662 -2994 247800
rect -2674 247662 -2626 247982
rect -1526 250052 -1206 250640
rect -1526 249780 -1502 250052
rect -1230 249780 -1206 250052
rect -1526 247960 -1206 249780
rect -3018 247638 -2626 247662
rect -1528 247640 -1206 247960
rect -6318 245120 -5950 245144
rect -6318 244800 -6294 245120
rect -5974 244800 -5950 245120
rect -6318 244776 -5950 244800
rect -3786 245120 -3418 245144
rect -2946 245120 -2626 247638
rect -3786 244800 -3762 245120
rect -3442 244982 -2626 245120
rect -3442 244800 -2994 244982
rect -3786 244776 -3418 244800
rect -3018 244662 -2994 244800
rect -2674 244662 -2626 244982
rect -1526 244960 -1206 247640
rect -3018 244638 -2626 244662
rect -1528 244640 -1206 244960
rect -5546 244076 -5178 244100
rect -5546 243756 -5522 244076
rect -5202 243756 -5178 244076
rect -5546 243732 -5178 243756
rect -6318 242120 -5950 242144
rect -6318 241800 -6294 242120
rect -5974 241800 -5950 242120
rect -6318 241776 -5950 241800
rect -3786 242120 -3418 242144
rect -2946 242120 -2626 244638
rect -3786 241800 -3762 242120
rect -3442 241982 -2626 242120
rect -3442 241800 -2994 241982
rect -3786 241776 -3418 241800
rect -3018 241662 -2994 241800
rect -2674 241662 -2626 241982
rect -1526 244052 -1206 244640
rect -1526 243780 -1502 244052
rect -1230 243780 -1206 244052
rect -1526 241960 -1206 243780
rect -3018 241638 -2626 241662
rect -1528 241640 -1206 241960
rect -5546 241076 -5178 241100
rect -5546 240756 -5522 241076
rect -5202 240756 -5178 241076
rect -5546 240732 -5178 240756
rect -6318 239120 -5950 239144
rect -6318 238800 -6294 239120
rect -5974 238800 -5950 239120
rect -6318 238776 -5950 238800
rect -3786 239120 -3418 239144
rect -2946 239120 -2626 241638
rect -3786 238800 -3762 239120
rect -3442 238982 -2626 239120
rect -3442 238800 -2994 238982
rect -3786 238776 -3418 238800
rect -3018 238662 -2994 238800
rect -2674 238662 -2626 238982
rect -1526 241052 -1206 241640
rect -1526 240780 -1502 241052
rect -1230 240780 -1206 241052
rect -1526 238960 -1206 240780
rect -3018 238638 -2626 238662
rect -1528 238640 -1206 238960
rect -5546 238076 -5178 238100
rect -5546 237756 -5522 238076
rect -5202 237756 -5178 238076
rect -5546 237732 -5178 237756
rect -6318 236120 -5950 236144
rect -6318 235800 -6294 236120
rect -5974 235800 -5950 236120
rect -6318 235776 -5950 235800
rect -3786 236120 -3418 236144
rect -2946 236120 -2626 238638
rect -3786 235800 -3762 236120
rect -3442 235982 -2626 236120
rect -3442 235800 -2994 235982
rect -3786 235776 -3418 235800
rect -3018 235662 -2994 235800
rect -2674 235662 -2626 235982
rect -1526 238052 -1206 238640
rect -1526 237780 -1502 238052
rect -1230 237780 -1206 238052
rect -1526 235960 -1206 237780
rect -3018 235638 -2626 235662
rect -1528 235640 -1206 235960
rect -5546 235076 -5178 235100
rect -5546 234756 -5522 235076
rect -5202 234756 -5178 235076
rect -5546 234732 -5178 234756
rect -6318 233120 -5950 233144
rect -6318 232800 -6294 233120
rect -5974 232800 -5950 233120
rect -6318 232776 -5950 232800
rect -3786 233120 -3418 233144
rect -2946 233120 -2626 235638
rect -3786 232800 -3762 233120
rect -3442 232982 -2626 233120
rect -3442 232800 -2994 232982
rect -3786 232776 -3418 232800
rect -3018 232662 -2994 232800
rect -2674 232662 -2626 232982
rect -1526 235052 -1206 235640
rect -1526 234780 -1502 235052
rect -1230 234780 -1206 235052
rect -1526 232960 -1206 234780
rect -3018 232638 -2626 232662
rect -1528 232640 -1206 232960
rect -5546 232076 -5178 232100
rect -5546 231756 -5522 232076
rect -5202 231756 -5178 232076
rect -5546 231732 -5178 231756
rect -6318 230120 -5950 230144
rect -6318 229800 -6294 230120
rect -5974 229800 -5950 230120
rect -6318 229776 -5950 229800
rect -3786 230120 -3418 230144
rect -2946 230120 -2626 232638
rect -3786 229800 -3762 230120
rect -3442 229982 -2626 230120
rect -3442 229800 -2994 229982
rect -3786 229776 -3418 229800
rect -3018 229662 -2994 229800
rect -2674 229662 -2626 229982
rect -1526 232052 -1206 232640
rect -1526 231780 -1502 232052
rect -1230 231780 -1206 232052
rect -1526 229960 -1206 231780
rect -3018 229638 -2626 229662
rect -1528 229640 -1206 229960
rect -5546 229076 -5178 229100
rect -5546 228756 -5522 229076
rect -5202 228756 -5178 229076
rect -5546 228732 -5178 228756
rect -6318 227120 -5950 227144
rect -6318 226800 -6294 227120
rect -5974 226800 -5950 227120
rect -6318 226776 -5950 226800
rect -3786 227120 -3418 227144
rect -2946 227120 -2626 229638
rect -3786 226800 -3762 227120
rect -3442 226982 -2626 227120
rect -3442 226800 -2994 226982
rect -3786 226776 -3418 226800
rect -3018 226662 -2994 226800
rect -2674 226662 -2626 226982
rect -1526 229052 -1206 229640
rect -1526 228780 -1502 229052
rect -1230 228780 -1206 229052
rect -1526 226960 -1206 228780
rect -3018 226638 -2626 226662
rect -1528 226640 -1206 226960
rect -5546 226076 -5178 226100
rect -5546 225756 -5522 226076
rect -5202 225756 -5178 226076
rect -5546 225732 -5178 225756
rect -6318 224120 -5950 224144
rect -6318 223800 -6294 224120
rect -5974 223800 -5950 224120
rect -6318 223776 -5950 223800
rect -3786 224120 -3418 224144
rect -2946 224120 -2626 226638
rect -3786 223800 -3762 224120
rect -3442 223982 -2626 224120
rect -3442 223800 -2994 223982
rect -3786 223776 -3418 223800
rect -3018 223662 -2994 223800
rect -2674 223662 -2626 223982
rect -1526 226052 -1206 226640
rect -1526 225780 -1502 226052
rect -1230 225780 -1206 226052
rect -1526 223960 -1206 225780
rect -3018 223638 -2626 223662
rect -1528 223640 -1206 223960
rect -5546 223076 -5178 223100
rect -5546 222756 -5522 223076
rect -5202 222756 -5178 223076
rect -5546 222732 -5178 222756
rect -6318 221120 -5950 221144
rect -6318 220800 -6294 221120
rect -5974 220800 -5950 221120
rect -6318 220776 -5950 220800
rect -3786 221120 -3418 221144
rect -2946 221120 -2626 223638
rect -3786 220800 -3762 221120
rect -3442 220982 -2626 221120
rect -3442 220800 -2994 220982
rect -3786 220776 -3418 220800
rect -3018 220662 -2994 220800
rect -2674 220662 -2626 220982
rect -1526 223052 -1206 223640
rect -1526 222780 -1502 223052
rect -1230 222780 -1206 223052
rect -1526 220960 -1206 222780
rect -3018 220638 -2626 220662
rect -1528 220640 -1206 220960
rect -5546 220076 -5178 220100
rect -5546 219756 -5522 220076
rect -5202 219756 -5178 220076
rect -5546 219732 -5178 219756
rect -6318 218120 -5950 218144
rect -6318 217800 -6294 218120
rect -5974 217800 -5950 218120
rect -6318 217776 -5950 217800
rect -3786 218120 -3418 218144
rect -2946 218120 -2626 220638
rect -3786 217800 -3762 218120
rect -3442 217982 -2626 218120
rect -3442 217800 -2994 217982
rect -3786 217776 -3418 217800
rect -3018 217662 -2994 217800
rect -2674 217662 -2626 217982
rect -1526 220052 -1206 220640
rect -1526 219780 -1502 220052
rect -1230 219780 -1206 220052
rect -1526 217960 -1206 219780
rect -3018 217638 -2626 217662
rect -1528 217640 -1206 217960
rect -5546 217076 -5178 217100
rect -5546 216756 -5522 217076
rect -5202 216756 -5178 217076
rect -5546 216732 -5178 216756
rect -6318 215120 -5950 215144
rect -6318 214800 -6294 215120
rect -5974 214800 -5950 215120
rect -6318 214776 -5950 214800
rect -3786 215120 -3418 215144
rect -2946 215120 -2626 217638
rect -3786 214800 -3762 215120
rect -3442 214982 -2626 215120
rect -3442 214800 -2994 214982
rect -3786 214776 -3418 214800
rect -3018 214662 -2994 214800
rect -2674 214662 -2626 214982
rect -1526 217052 -1206 217640
rect -1526 216780 -1502 217052
rect -1230 216780 -1206 217052
rect -1526 214960 -1206 216780
rect -3018 214638 -2626 214662
rect -1528 214640 -1206 214960
rect -5546 214076 -5178 214100
rect -5546 213756 -5522 214076
rect -5202 213756 -5178 214076
rect -5546 213732 -5178 213756
rect -6318 212120 -5950 212144
rect -6318 211800 -6294 212120
rect -5974 211800 -5950 212120
rect -6318 211776 -5950 211800
rect -3786 212120 -3418 212144
rect -2946 212120 -2626 214638
rect -3786 211800 -3762 212120
rect -3442 211982 -2626 212120
rect -3442 211800 -2994 211982
rect -3786 211776 -3418 211800
rect -3018 211662 -2994 211800
rect -2674 211662 -2626 211982
rect -1526 214052 -1206 214640
rect -1526 213780 -1502 214052
rect -1230 213780 -1206 214052
rect -1526 211960 -1206 213780
rect -3018 211638 -2626 211662
rect -1528 211640 -1206 211960
rect -5546 211076 -5178 211100
rect -5546 210756 -5522 211076
rect -5202 210756 -5178 211076
rect -5546 210732 -5178 210756
rect -2946 209120 -2626 211638
rect -3120 208982 -2626 209120
rect -3120 208800 -2994 208982
rect -3018 208662 -2994 208800
rect -2674 208662 -2626 208982
rect -1526 211052 -1206 211640
rect -1526 210780 -1502 211052
rect -1230 210780 -1206 211052
rect -1526 208960 -1206 210780
rect -3018 208638 -2626 208662
rect -1528 208640 -1206 208960
rect -5546 208076 -5178 208100
rect -5546 207756 -5522 208076
rect -5202 207756 -5178 208076
rect -5546 207732 -5178 207756
rect -6318 206120 -5950 206144
rect -6318 205800 -6294 206120
rect -5974 205800 -5950 206120
rect -6318 205776 -5950 205800
rect -3786 206120 -3418 206144
rect -2946 206120 -2626 208638
rect -3786 205800 -3762 206120
rect -3442 205982 -2626 206120
rect -3442 205800 -2994 205982
rect -3786 205776 -3418 205800
rect -3018 205662 -2994 205800
rect -2674 205662 -2626 205982
rect -1526 208052 -1206 208640
rect -1526 207780 -1502 208052
rect -1230 207780 -1206 208052
rect -1526 205960 -1206 207780
rect -3018 205638 -2626 205662
rect -1528 205640 -1206 205960
rect -5546 205076 -5178 205100
rect -5546 204756 -5522 205076
rect -5202 204756 -5178 205076
rect -5546 204732 -5178 204756
rect -6318 203120 -5950 203144
rect -6318 202800 -6294 203120
rect -5974 202800 -5950 203120
rect -6318 202776 -5950 202800
rect -3786 203120 -3418 203144
rect -2946 203120 -2626 205638
rect -3786 202800 -3762 203120
rect -3442 202982 -2626 203120
rect -3442 202800 -2994 202982
rect -3786 202776 -3418 202800
rect -3018 202662 -2994 202800
rect -2674 202662 -2626 202982
rect -1526 205052 -1206 205640
rect -1526 204780 -1502 205052
rect -1230 204780 -1206 205052
rect -1526 202960 -1206 204780
rect -3018 202638 -2626 202662
rect -1528 202640 -1206 202960
rect -5546 202076 -5178 202100
rect -5546 201756 -5522 202076
rect -5202 201756 -5178 202076
rect -5546 201732 -5178 201756
rect -6318 200120 -5950 200144
rect -6318 199800 -6294 200120
rect -5974 199800 -5950 200120
rect -6318 199776 -5950 199800
rect -3786 200120 -3418 200144
rect -2946 200120 -2626 202638
rect -3786 199800 -3762 200120
rect -3442 199982 -2626 200120
rect -3442 199800 -2994 199982
rect -3786 199776 -3418 199800
rect -3018 199662 -2994 199800
rect -2674 199662 -2626 199982
rect -1526 202052 -1206 202640
rect -1526 201780 -1502 202052
rect -1230 201780 -1206 202052
rect -1526 199960 -1206 201780
rect -3018 199638 -2626 199662
rect -1528 199640 -1206 199960
rect -5546 199076 -5178 199100
rect -5546 198756 -5522 199076
rect -5202 198756 -5178 199076
rect -5546 198732 -5178 198756
rect -6318 197120 -5950 197144
rect -6318 196800 -6294 197120
rect -5974 196800 -5950 197120
rect -6318 196776 -5950 196800
rect -3786 197120 -3418 197144
rect -2946 197120 -2626 199638
rect -3786 196800 -3762 197120
rect -3442 196982 -2626 197120
rect -3442 196800 -2994 196982
rect -3786 196776 -3418 196800
rect -3018 196662 -2994 196800
rect -2674 196662 -2626 196982
rect -1526 199052 -1206 199640
rect -1526 198780 -1502 199052
rect -1230 198780 -1206 199052
rect -1526 196960 -1206 198780
rect -3018 196638 -2626 196662
rect -1528 196640 -1206 196960
rect -5546 196076 -5178 196100
rect -5546 195756 -5522 196076
rect -5202 195756 -5178 196076
rect -5546 195732 -5178 195756
rect -6318 194120 -5950 194144
rect -6318 193800 -6294 194120
rect -5974 193800 -5950 194120
rect -6318 193776 -5950 193800
rect -3786 194120 -3418 194144
rect -2946 194120 -2626 196638
rect -3786 193800 -3762 194120
rect -3442 193982 -2626 194120
rect -3442 193800 -2994 193982
rect -3786 193776 -3418 193800
rect -3018 193662 -2994 193800
rect -2674 193662 -2626 193982
rect -1526 196052 -1206 196640
rect -1526 195780 -1502 196052
rect -1230 195780 -1206 196052
rect -1526 193960 -1206 195780
rect -3018 193638 -2626 193662
rect -1528 193640 -1206 193960
rect -5546 193076 -5178 193100
rect -5546 192756 -5522 193076
rect -5202 192756 -5178 193076
rect -5546 192732 -5178 192756
rect -6318 191120 -5950 191144
rect -6318 190800 -6294 191120
rect -5974 190800 -5950 191120
rect -6318 190776 -5950 190800
rect -3786 191120 -3418 191144
rect -2946 191120 -2626 193638
rect -3786 190800 -3762 191120
rect -3442 190982 -2626 191120
rect -3442 190800 -2994 190982
rect -3786 190776 -3418 190800
rect -3018 190662 -2994 190800
rect -2674 190662 -2626 190982
rect -1526 193052 -1206 193640
rect -1526 192780 -1502 193052
rect -1230 192780 -1206 193052
rect -1526 190960 -1206 192780
rect -3018 190638 -2626 190662
rect -1528 190640 -1206 190960
rect -5546 190076 -5178 190100
rect -5546 189756 -5522 190076
rect -5202 189756 -5178 190076
rect -5546 189732 -5178 189756
rect -6318 188120 -5950 188144
rect -6318 187800 -6294 188120
rect -5974 187800 -5950 188120
rect -6318 187776 -5950 187800
rect -3786 188120 -3418 188144
rect -2946 188120 -2626 190638
rect -3786 187800 -3762 188120
rect -3442 187982 -2626 188120
rect -3442 187800 -2994 187982
rect -3786 187776 -3418 187800
rect -3018 187662 -2994 187800
rect -2674 187662 -2626 187982
rect -1526 190052 -1206 190640
rect -1526 189780 -1502 190052
rect -1230 189780 -1206 190052
rect -1526 187960 -1206 189780
rect -3018 187638 -2626 187662
rect -1528 187640 -1206 187960
rect -5546 187076 -5178 187100
rect -5546 186756 -5522 187076
rect -5202 186756 -5178 187076
rect -5546 186732 -5178 186756
rect -6318 185120 -5950 185144
rect -6318 184800 -6294 185120
rect -5974 184800 -5950 185120
rect -6318 184776 -5950 184800
rect -3786 185120 -3418 185144
rect -2946 185120 -2626 187638
rect -3786 184800 -3762 185120
rect -3442 184982 -2626 185120
rect -3442 184800 -2994 184982
rect -3786 184776 -3418 184800
rect -3018 184662 -2994 184800
rect -2674 184662 -2626 184982
rect -1526 187052 -1206 187640
rect -1526 186780 -1502 187052
rect -1230 186780 -1206 187052
rect -1526 184960 -1206 186780
rect -3018 184638 -2626 184662
rect -1528 184640 -1206 184960
rect -5546 184076 -5178 184100
rect -5546 183756 -5522 184076
rect -5202 183756 -5178 184076
rect -5546 183732 -5178 183756
rect -6318 182120 -5950 182144
rect -6318 181800 -6294 182120
rect -5974 181800 -5950 182120
rect -6318 181776 -5950 181800
rect -3786 182120 -3418 182144
rect -2946 182120 -2626 184638
rect -3786 181800 -3762 182120
rect -3442 181982 -2626 182120
rect -3442 181800 -2994 181982
rect -3786 181776 -3418 181800
rect -3018 181662 -2994 181800
rect -2674 181662 -2626 181982
rect -1526 184052 -1206 184640
rect -1526 183780 -1502 184052
rect -1230 183780 -1206 184052
rect -1526 181960 -1206 183780
rect -3018 181638 -2626 181662
rect -1528 181640 -1206 181960
rect -5546 181076 -5178 181100
rect -5546 180756 -5522 181076
rect -5202 180756 -5178 181076
rect -5546 180732 -5178 180756
rect -6318 179120 -5950 179144
rect -6318 178800 -6294 179120
rect -5974 178800 -5950 179120
rect -6318 178776 -5950 178800
rect -3786 179120 -3418 179144
rect -2946 179120 -2626 181638
rect -3786 178800 -3762 179120
rect -3442 178982 -2626 179120
rect -3442 178800 -2994 178982
rect -3786 178776 -3418 178800
rect -3018 178662 -2994 178800
rect -2674 178662 -2626 178982
rect -1526 181052 -1206 181640
rect -1526 180780 -1502 181052
rect -1230 180780 -1206 181052
rect -1526 178960 -1206 180780
rect -3018 178638 -2626 178662
rect -1528 178640 -1206 178960
rect -5546 178076 -5178 178100
rect -5546 177756 -5522 178076
rect -5202 177756 -5178 178076
rect -5546 177732 -5178 177756
rect -6318 176120 -5950 176144
rect -6318 175800 -6294 176120
rect -5974 175800 -5950 176120
rect -6318 175776 -5950 175800
rect -3786 176120 -3418 176144
rect -2946 176120 -2626 178638
rect -3786 175800 -3762 176120
rect -3442 175982 -2626 176120
rect -3442 175800 -2994 175982
rect -3786 175776 -3418 175800
rect -3018 175662 -2994 175800
rect -2674 175662 -2626 175982
rect -1526 178052 -1206 178640
rect -1526 177780 -1502 178052
rect -1230 177780 -1206 178052
rect -1526 175960 -1206 177780
rect -3018 175638 -2626 175662
rect -1528 175640 -1206 175960
rect -5546 175076 -5178 175100
rect -5546 174756 -5522 175076
rect -5202 174756 -5178 175076
rect -5546 174732 -5178 174756
rect -6318 173120 -5950 173144
rect -6318 172800 -6294 173120
rect -5974 172800 -5950 173120
rect -6318 172776 -5950 172800
rect -3786 173120 -3418 173144
rect -2946 173120 -2626 175638
rect -3786 172800 -3762 173120
rect -3442 172982 -2626 173120
rect -3442 172800 -2994 172982
rect -3786 172776 -3418 172800
rect -3018 172662 -2994 172800
rect -2674 172662 -2626 172982
rect -1526 175052 -1206 175640
rect -1526 174780 -1502 175052
rect -1230 174780 -1206 175052
rect -1526 172960 -1206 174780
rect -3018 172638 -2626 172662
rect -1528 172640 -1206 172960
rect -5546 172076 -5178 172100
rect -5546 171756 -5522 172076
rect -5202 171756 -5178 172076
rect -5546 171732 -5178 171756
rect -6318 170120 -5950 170144
rect -6318 169800 -6294 170120
rect -5974 169800 -5950 170120
rect -6318 169776 -5950 169800
rect -3786 170120 -3418 170144
rect -2946 170120 -2626 172638
rect -3786 169800 -3762 170120
rect -3442 169982 -2626 170120
rect -3442 169800 -2994 169982
rect -3786 169776 -3418 169800
rect -3018 169662 -2994 169800
rect -2674 169662 -2626 169982
rect -1526 172052 -1206 172640
rect -1526 171780 -1502 172052
rect -1230 171780 -1206 172052
rect -1526 169960 -1206 171780
rect -3018 169638 -2626 169662
rect -1528 169640 -1206 169960
rect -5546 169076 -5178 169100
rect -5546 168756 -5522 169076
rect -5202 168756 -5178 169076
rect -5546 168732 -5178 168756
rect -6318 167120 -5950 167144
rect -6318 166800 -6294 167120
rect -5974 166800 -5950 167120
rect -6318 166776 -5950 166800
rect -3786 167120 -3418 167144
rect -2946 167120 -2626 169638
rect -3786 166800 -3762 167120
rect -3442 166982 -2626 167120
rect -3442 166800 -2994 166982
rect -3786 166776 -3418 166800
rect -3018 166662 -2994 166800
rect -2674 166662 -2626 166982
rect -1526 169052 -1206 169640
rect -1526 168780 -1502 169052
rect -1230 168780 -1206 169052
rect -1526 166960 -1206 168780
rect -3018 166638 -2626 166662
rect -1528 166640 -1206 166960
rect -5546 166076 -5178 166100
rect -5546 165756 -5522 166076
rect -5202 165756 -5178 166076
rect -5546 165732 -5178 165756
rect -6318 164120 -5950 164144
rect -6318 163800 -6294 164120
rect -5974 163800 -5950 164120
rect -6318 163776 -5950 163800
rect -3786 164120 -3418 164144
rect -2946 164120 -2626 166638
rect -3786 163800 -3762 164120
rect -3442 163982 -2626 164120
rect -3442 163800 -2994 163982
rect -3786 163776 -3418 163800
rect -3018 163662 -2994 163800
rect -2674 163662 -2626 163982
rect -1526 166052 -1206 166640
rect -1526 165780 -1502 166052
rect -1230 165780 -1206 166052
rect -1526 163960 -1206 165780
rect -3018 163638 -2626 163662
rect -1528 163640 -1206 163960
rect -5546 163076 -5178 163100
rect -5546 162756 -5522 163076
rect -5202 162756 -5178 163076
rect -5546 162732 -5178 162756
rect -6318 161120 -5950 161144
rect -6318 160800 -6294 161120
rect -5974 160800 -5950 161120
rect -6318 160776 -5950 160800
rect -3786 161120 -3418 161144
rect -2946 161120 -2626 163638
rect -3786 160800 -3762 161120
rect -3442 160982 -2626 161120
rect -3442 160800 -2994 160982
rect -3786 160776 -3418 160800
rect -3018 160662 -2994 160800
rect -2674 160662 -2626 160982
rect -1526 163052 -1206 163640
rect -1526 162780 -1502 163052
rect -1230 162780 -1206 163052
rect -1526 160960 -1206 162780
rect -3018 160638 -2626 160662
rect -1528 160640 -1206 160960
rect -5546 160076 -5178 160100
rect -5546 159756 -5522 160076
rect -5202 159756 -5178 160076
rect -5546 159732 -5178 159756
rect -6318 158120 -5950 158144
rect -6318 157800 -6294 158120
rect -5974 157800 -5950 158120
rect -6318 157776 -5950 157800
rect -3786 158120 -3418 158144
rect -2946 158120 -2626 160638
rect -3786 157800 -3762 158120
rect -3442 157982 -2626 158120
rect -3442 157800 -2994 157982
rect -3786 157776 -3418 157800
rect -3018 157662 -2994 157800
rect -2674 157662 -2626 157982
rect -1526 160052 -1206 160640
rect -1526 159780 -1502 160052
rect -1230 159780 -1206 160052
rect -1526 157960 -1206 159780
rect -3018 157638 -2626 157662
rect -1528 157640 -1206 157960
rect -5546 157076 -5178 157100
rect -5546 156756 -5522 157076
rect -5202 156756 -5178 157076
rect -5546 156732 -5178 156756
rect -6318 155120 -5950 155144
rect -6318 154800 -6294 155120
rect -5974 154800 -5950 155120
rect -6318 154776 -5950 154800
rect -3786 155120 -3418 155144
rect -2946 155120 -2626 157638
rect -3786 154800 -3762 155120
rect -3442 154982 -2626 155120
rect -3442 154800 -2994 154982
rect -3786 154776 -3418 154800
rect -3018 154662 -2994 154800
rect -2674 154662 -2626 154982
rect -1526 157052 -1206 157640
rect -1526 156780 -1502 157052
rect -1230 156780 -1206 157052
rect -1526 154960 -1206 156780
rect -3018 154638 -2626 154662
rect -1528 154640 -1206 154960
rect -5546 154076 -5178 154100
rect -5546 153756 -5522 154076
rect -5202 153756 -5178 154076
rect -5546 153732 -5178 153756
rect -6318 152120 -5950 152144
rect -6318 151800 -6294 152120
rect -5974 151800 -5950 152120
rect -6318 151776 -5950 151800
rect -3786 152120 -3418 152144
rect -2946 152120 -2626 154638
rect -3786 151800 -3762 152120
rect -3442 151982 -2626 152120
rect -3442 151800 -2994 151982
rect -3786 151776 -3418 151800
rect -3018 151662 -2994 151800
rect -2674 151662 -2626 151982
rect -1526 154052 -1206 154640
rect -1526 153780 -1502 154052
rect -1230 153780 -1206 154052
rect -1526 151960 -1206 153780
rect -3018 151638 -2626 151662
rect -1528 151640 -1206 151960
rect -5546 151076 -5178 151100
rect -5546 150756 -5522 151076
rect -5202 150756 -5178 151076
rect -5546 150732 -5178 150756
rect -6318 149120 -5950 149144
rect -6318 148800 -6294 149120
rect -5974 148800 -5950 149120
rect -6318 148776 -5950 148800
rect -3786 149120 -3418 149144
rect -2946 149120 -2626 151638
rect -3786 148800 -3762 149120
rect -3442 148982 -2626 149120
rect -3442 148800 -2994 148982
rect -3786 148776 -3418 148800
rect -3018 148662 -2994 148800
rect -2674 148662 -2626 148982
rect -1526 151052 -1206 151640
rect -1526 150780 -1502 151052
rect -1230 150780 -1206 151052
rect -1526 148960 -1206 150780
rect -3018 148638 -2626 148662
rect -1528 148640 -1206 148960
rect -5546 148076 -5178 148100
rect -5546 147756 -5522 148076
rect -5202 147756 -5178 148076
rect -5546 147732 -5178 147756
rect -6318 146120 -5950 146144
rect -6318 145800 -6294 146120
rect -5974 145800 -5950 146120
rect -6318 145776 -5950 145800
rect -3786 146120 -3418 146144
rect -2946 146120 -2626 148638
rect -3786 145800 -3762 146120
rect -3442 145982 -2626 146120
rect -3442 145800 -2994 145982
rect -3786 145776 -3418 145800
rect -3018 145662 -2994 145800
rect -2674 145662 -2626 145982
rect -1526 148052 -1206 148640
rect -1526 147780 -1502 148052
rect -1230 147780 -1206 148052
rect -1526 145960 -1206 147780
rect -3018 145638 -2626 145662
rect -1528 145640 -1206 145960
rect -5546 145076 -5178 145100
rect -5546 144756 -5522 145076
rect -5202 144756 -5178 145076
rect -5546 144732 -5178 144756
rect -6318 143120 -5950 143144
rect -6318 142800 -6294 143120
rect -5974 142800 -5950 143120
rect -6318 142776 -5950 142800
rect -3786 143120 -3418 143144
rect -2946 143120 -2626 145638
rect -3786 142800 -3762 143120
rect -3442 142982 -2626 143120
rect -3442 142800 -2994 142982
rect -3786 142776 -3418 142800
rect -3018 142662 -2994 142800
rect -2674 142662 -2626 142982
rect -1526 145052 -1206 145640
rect -1526 144780 -1502 145052
rect -1230 144780 -1206 145052
rect -1526 142960 -1206 144780
rect -3018 142638 -2626 142662
rect -1528 142640 -1206 142960
rect -5546 142076 -5178 142100
rect -5546 141756 -5522 142076
rect -5202 141756 -5178 142076
rect -5546 141732 -5178 141756
rect -6318 140120 -5950 140144
rect -6318 139800 -6294 140120
rect -5974 139800 -5950 140120
rect -6318 139776 -5950 139800
rect -3786 140120 -3418 140144
rect -2946 140120 -2626 142638
rect -3786 139800 -3762 140120
rect -3442 139982 -2626 140120
rect -3442 139800 -2994 139982
rect -3786 139776 -3418 139800
rect -3018 139662 -2994 139800
rect -2674 139662 -2626 139982
rect -1526 142052 -1206 142640
rect -1526 141780 -1502 142052
rect -1230 141780 -1206 142052
rect -1526 139960 -1206 141780
rect -3018 139638 -2626 139662
rect -1528 139640 -1206 139960
rect -5546 139076 -5178 139100
rect -5546 138756 -5522 139076
rect -5202 138756 -5178 139076
rect -5546 138732 -5178 138756
rect -6318 137120 -5950 137144
rect -6318 136800 -6294 137120
rect -5974 136800 -5950 137120
rect -6318 136776 -5950 136800
rect -3786 137120 -3418 137144
rect -2946 137120 -2626 139638
rect -3786 136800 -3762 137120
rect -3442 136982 -2626 137120
rect -3442 136800 -2994 136982
rect -3786 136776 -3418 136800
rect -3018 136662 -2994 136800
rect -2674 136662 -2626 136982
rect -1526 139052 -1206 139640
rect -1526 138780 -1502 139052
rect -1230 138780 -1206 139052
rect -1526 136960 -1206 138780
rect -3018 136638 -2626 136662
rect -1528 136640 -1206 136960
rect -5546 136076 -5178 136100
rect -5546 135756 -5522 136076
rect -5202 135756 -5178 136076
rect -5546 135732 -5178 135756
rect -6318 134120 -5950 134144
rect -6318 133800 -6294 134120
rect -5974 133800 -5950 134120
rect -6318 133776 -5950 133800
rect -3786 134120 -3418 134144
rect -2946 134120 -2626 136638
rect -3786 133800 -3762 134120
rect -3442 133982 -2626 134120
rect -3442 133800 -2994 133982
rect -3786 133776 -3418 133800
rect -3018 133662 -2994 133800
rect -2674 133662 -2626 133982
rect -1526 136052 -1206 136640
rect -1526 135780 -1502 136052
rect -1230 135780 -1206 136052
rect -1526 133960 -1206 135780
rect -3018 133638 -2626 133662
rect -1528 133640 -1206 133960
rect -5546 133076 -5178 133100
rect -5546 132756 -5522 133076
rect -5202 132756 -5178 133076
rect -5546 132732 -5178 132756
rect -6318 131120 -5950 131144
rect -6318 130800 -6294 131120
rect -5974 130800 -5950 131120
rect -6318 130776 -5950 130800
rect -3786 131120 -3418 131144
rect -2946 131120 -2626 133638
rect -3786 130800 -3762 131120
rect -3442 130982 -2626 131120
rect -3442 130800 -2994 130982
rect -3786 130776 -3418 130800
rect -3018 130662 -2994 130800
rect -2674 130662 -2626 130982
rect -1526 133052 -1206 133640
rect -1526 132780 -1502 133052
rect -1230 132780 -1206 133052
rect -1526 130960 -1206 132780
rect -3018 130638 -2626 130662
rect -1528 130640 -1206 130960
rect -5546 130076 -5178 130100
rect -5546 129756 -5522 130076
rect -5202 129756 -5178 130076
rect -5546 129732 -5178 129756
rect -6318 128120 -5950 128144
rect -6318 127800 -6294 128120
rect -5974 127800 -5950 128120
rect -6318 127776 -5950 127800
rect -3786 128120 -3418 128144
rect -2946 128120 -2626 130638
rect -3786 127800 -3762 128120
rect -3442 127982 -2626 128120
rect -3442 127800 -2994 127982
rect -3786 127776 -3418 127800
rect -3018 127662 -2994 127800
rect -2674 127662 -2626 127982
rect -1526 130052 -1206 130640
rect -1526 129780 -1502 130052
rect -1230 129780 -1206 130052
rect -1526 127960 -1206 129780
rect -3018 127638 -2626 127662
rect -1528 127640 -1206 127960
rect -5546 127076 -5178 127100
rect -5546 126756 -5522 127076
rect -5202 126756 -5178 127076
rect -5546 126732 -5178 126756
rect -6318 125120 -5950 125144
rect -6318 124800 -6294 125120
rect -5974 124800 -5950 125120
rect -6318 124776 -5950 124800
rect -3786 125120 -3418 125144
rect -2946 125120 -2626 127638
rect -3786 124800 -3762 125120
rect -3442 124982 -2626 125120
rect -3442 124800 -2994 124982
rect -3786 124776 -3418 124800
rect -3018 124662 -2994 124800
rect -2674 124662 -2626 124982
rect -1526 127052 -1206 127640
rect -1526 126780 -1502 127052
rect -1230 126780 -1206 127052
rect -1526 124960 -1206 126780
rect -3018 124638 -2626 124662
rect -1528 124640 -1206 124960
rect -5546 124076 -5178 124100
rect -5546 123756 -5522 124076
rect -5202 123756 -5178 124076
rect -5546 123732 -5178 123756
rect -6318 122120 -5950 122144
rect -6318 121800 -6294 122120
rect -5974 121800 -5950 122120
rect -6318 121776 -5950 121800
rect -3786 122120 -3418 122144
rect -2946 122120 -2626 124638
rect -3786 121800 -3762 122120
rect -3442 121982 -2626 122120
rect -3442 121800 -2994 121982
rect -3786 121776 -3418 121800
rect -3018 121662 -2994 121800
rect -2674 121662 -2626 121982
rect -1526 124052 -1206 124640
rect -1526 123780 -1502 124052
rect -1230 123780 -1206 124052
rect -1526 121960 -1206 123780
rect -3018 121638 -2626 121662
rect -1528 121640 -1206 121960
rect -5546 121076 -5178 121100
rect -5546 120756 -5522 121076
rect -5202 120756 -5178 121076
rect -5546 120732 -5178 120756
rect -6318 119120 -5950 119144
rect -6318 118800 -6294 119120
rect -5974 118800 -5950 119120
rect -6318 118776 -5950 118800
rect -3786 119120 -3418 119144
rect -2946 119120 -2626 121638
rect -3786 118800 -3762 119120
rect -3442 118982 -2626 119120
rect -3442 118800 -2994 118982
rect -3786 118776 -3418 118800
rect -3018 118662 -2994 118800
rect -2674 118662 -2626 118982
rect -1526 121052 -1206 121640
rect -1526 120780 -1502 121052
rect -1230 120780 -1206 121052
rect -1526 118960 -1206 120780
rect -3018 118638 -2626 118662
rect -1528 118640 -1206 118960
rect -5546 118076 -5178 118100
rect -5546 117756 -5522 118076
rect -5202 117756 -5178 118076
rect -5546 117732 -5178 117756
rect -6318 116120 -5950 116144
rect -6318 115800 -6294 116120
rect -5974 115800 -5950 116120
rect -6318 115776 -5950 115800
rect -3786 116120 -3418 116144
rect -2946 116120 -2626 118638
rect -3786 115800 -3762 116120
rect -3442 115982 -2626 116120
rect -3442 115800 -2994 115982
rect -3786 115776 -3418 115800
rect -3018 115662 -2994 115800
rect -2674 115662 -2626 115982
rect -1526 118052 -1206 118640
rect -1526 117780 -1502 118052
rect -1230 117780 -1206 118052
rect -1526 115960 -1206 117780
rect -3018 115638 -2626 115662
rect -1528 115640 -1206 115960
rect -5546 115076 -5178 115100
rect -5546 114756 -5522 115076
rect -5202 114756 -5178 115076
rect -5546 114732 -5178 114756
rect -6318 113120 -5950 113144
rect -6318 112800 -6294 113120
rect -5974 112800 -5950 113120
rect -6318 112776 -5950 112800
rect -3786 113120 -3418 113144
rect -2946 113120 -2626 115638
rect -3786 112800 -3762 113120
rect -3442 112982 -2626 113120
rect -3442 112800 -2994 112982
rect -3786 112776 -3418 112800
rect -3018 112662 -2994 112800
rect -2674 112662 -2626 112982
rect -1526 115052 -1206 115640
rect -1526 114780 -1502 115052
rect -1230 114780 -1206 115052
rect -1526 112960 -1206 114780
rect -3018 112638 -2626 112662
rect -1528 112640 -1206 112960
rect -5546 112076 -5178 112100
rect -5546 111756 -5522 112076
rect -5202 111756 -5178 112076
rect -5546 111732 -5178 111756
rect -6318 110120 -5950 110144
rect -6318 109800 -6294 110120
rect -5974 109800 -5950 110120
rect -6318 109776 -5950 109800
rect -3786 110120 -3418 110144
rect -2946 110120 -2626 112638
rect -3786 109800 -3762 110120
rect -3442 109982 -2626 110120
rect -3442 109800 -2994 109982
rect -3786 109776 -3418 109800
rect -3018 109662 -2994 109800
rect -2674 109662 -2626 109982
rect -1526 112052 -1206 112640
rect -1526 111780 -1502 112052
rect -1230 111780 -1206 112052
rect -1526 109960 -1206 111780
rect -3018 109638 -2626 109662
rect -1528 109640 -1206 109960
rect -5546 109076 -5178 109100
rect -5546 108756 -5522 109076
rect -5202 108756 -5178 109076
rect -5546 108732 -5178 108756
rect -6318 107120 -5950 107144
rect -6318 106800 -6294 107120
rect -5974 106800 -5950 107120
rect -6318 106776 -5950 106800
rect -3786 107120 -3418 107144
rect -2946 107120 -2626 109638
rect -3786 106800 -3762 107120
rect -3442 106982 -2626 107120
rect -3442 106800 -2994 106982
rect -3786 106776 -3418 106800
rect -3018 106662 -2994 106800
rect -2674 106662 -2626 106982
rect -1526 109052 -1206 109640
rect -1526 108780 -1502 109052
rect -1230 108780 -1206 109052
rect -1526 106960 -1206 108780
rect -3018 106638 -2626 106662
rect -1528 106640 -1206 106960
rect -5546 106076 -5178 106100
rect -5546 105756 -5522 106076
rect -5202 105756 -5178 106076
rect -5546 105732 -5178 105756
rect -6318 104120 -5950 104144
rect -6318 103800 -6294 104120
rect -5974 103800 -5950 104120
rect -6318 103776 -5950 103800
rect -3786 104120 -3418 104144
rect -2946 104120 -2626 106638
rect -3786 103800 -3762 104120
rect -3442 103982 -2626 104120
rect -3442 103800 -2994 103982
rect -3786 103776 -3418 103800
rect -3018 103662 -2994 103800
rect -2674 103662 -2626 103982
rect -1526 106052 -1206 106640
rect -1526 105780 -1502 106052
rect -1230 105780 -1206 106052
rect -1526 103960 -1206 105780
rect -3018 103638 -2626 103662
rect -1528 103640 -1206 103960
rect -5546 103076 -5178 103100
rect -5546 102756 -5522 103076
rect -5202 102756 -5178 103076
rect -5546 102732 -5178 102756
rect -6318 101120 -5950 101144
rect -6318 100800 -6294 101120
rect -5974 100800 -5950 101120
rect -6318 100776 -5950 100800
rect -3786 101120 -3418 101144
rect -2946 101120 -2626 103638
rect -3786 100800 -3762 101120
rect -3442 100982 -2626 101120
rect -3442 100800 -2994 100982
rect -3786 100776 -3418 100800
rect -3018 100662 -2994 100800
rect -2674 100662 -2626 100982
rect -1526 103052 -1206 103640
rect -1526 102780 -1502 103052
rect -1230 102780 -1206 103052
rect -1526 100960 -1206 102780
rect -3018 100638 -2626 100662
rect -1528 100640 -1206 100960
rect -5546 100076 -5178 100100
rect -5546 99756 -5522 100076
rect -5202 99756 -5178 100076
rect -5546 99732 -5178 99756
rect -6318 98120 -5950 98144
rect -6318 97800 -6294 98120
rect -5974 97800 -5950 98120
rect -6318 97776 -5950 97800
rect -3786 98120 -3418 98144
rect -2946 98120 -2626 100638
rect -3786 97800 -3762 98120
rect -3442 97982 -2626 98120
rect -3442 97800 -2994 97982
rect -3786 97776 -3418 97800
rect -3018 97662 -2994 97800
rect -2674 97662 -2626 97982
rect -1526 100052 -1206 100640
rect -1526 99780 -1502 100052
rect -1230 99780 -1206 100052
rect -1526 97960 -1206 99780
rect -3018 97638 -2626 97662
rect -1528 97640 -1206 97960
rect -5546 97076 -5178 97100
rect -5546 96756 -5522 97076
rect -5202 96756 -5178 97076
rect -5546 96732 -5178 96756
rect -6318 95120 -5950 95144
rect -6318 94800 -6294 95120
rect -5974 94800 -5950 95120
rect -6318 94776 -5950 94800
rect -3786 95120 -3418 95144
rect -2946 95120 -2626 97638
rect -3786 94800 -3762 95120
rect -3442 94982 -2626 95120
rect -3442 94800 -2994 94982
rect -3786 94776 -3418 94800
rect -3018 94662 -2994 94800
rect -2674 94662 -2626 94982
rect -1526 97052 -1206 97640
rect -1526 96780 -1502 97052
rect -1230 96780 -1206 97052
rect -1526 94960 -1206 96780
rect -3018 94638 -2626 94662
rect -1528 94640 -1206 94960
rect -6318 92120 -5950 92144
rect -6318 91800 -6294 92120
rect -5974 91800 -5950 92120
rect -6318 91776 -5950 91800
rect -3786 92120 -3418 92144
rect -2946 92120 -2626 94638
rect -3786 91800 -3762 92120
rect -3442 91982 -2626 92120
rect -3442 91800 -2994 91982
rect -3786 91776 -3418 91800
rect -3018 91662 -2994 91800
rect -2674 91662 -2626 91982
rect -1526 91960 -1206 94640
rect -3018 91638 -2626 91662
rect -1528 91640 -1206 91960
rect -5546 91076 -5178 91100
rect -5546 90756 -5522 91076
rect -5202 90756 -5178 91076
rect -5546 90732 -5178 90756
rect -6318 89120 -5950 89144
rect -6318 88800 -6294 89120
rect -5974 88800 -5950 89120
rect -6318 88776 -5950 88800
rect -3786 89120 -3418 89144
rect -2946 89120 -2626 91638
rect -3786 88800 -3762 89120
rect -3442 88982 -2626 89120
rect -3442 88800 -2994 88982
rect -3786 88776 -3418 88800
rect -3018 88662 -2994 88800
rect -2674 88662 -2626 88982
rect -1526 91052 -1206 91640
rect -1526 90780 -1502 91052
rect -1230 90780 -1206 91052
rect -1526 88960 -1206 90780
rect -3018 88638 -2626 88662
rect -1528 88640 -1206 88960
rect -5546 88076 -5178 88100
rect -5546 87756 -5522 88076
rect -5202 87756 -5178 88076
rect -5546 87732 -5178 87756
rect -6318 86120 -5950 86144
rect -6318 85800 -6294 86120
rect -5974 85800 -5950 86120
rect -6318 85776 -5950 85800
rect -3786 86120 -3418 86144
rect -2946 86120 -2626 88638
rect -3786 85800 -3762 86120
rect -3442 85982 -2626 86120
rect -3442 85800 -2994 85982
rect -3786 85776 -3418 85800
rect -3018 85662 -2994 85800
rect -2674 85662 -2626 85982
rect -1526 88052 -1206 88640
rect -1526 87780 -1502 88052
rect -1230 87780 -1206 88052
rect -1526 85960 -1206 87780
rect -3018 85638 -2626 85662
rect -1528 85640 -1206 85960
rect -5546 85076 -5178 85100
rect -5546 84756 -5522 85076
rect -5202 84756 -5178 85076
rect -5546 84732 -5178 84756
rect -6318 83120 -5950 83144
rect -6318 82800 -6294 83120
rect -5974 82800 -5950 83120
rect -6318 82776 -5950 82800
rect -3786 83120 -3418 83144
rect -2946 83120 -2626 85638
rect -3786 82800 -3762 83120
rect -3442 82982 -2626 83120
rect -3442 82800 -2994 82982
rect -3786 82776 -3418 82800
rect -3018 82662 -2994 82800
rect -2674 82662 -2626 82982
rect -1526 85052 -1206 85640
rect -1526 84780 -1502 85052
rect -1230 84780 -1206 85052
rect -1526 82960 -1206 84780
rect -3018 82638 -2626 82662
rect -1528 82640 -1206 82960
rect -5546 82076 -5178 82100
rect -5546 81756 -5522 82076
rect -5202 81756 -5178 82076
rect -5546 81732 -5178 81756
rect -6318 80120 -5950 80144
rect -6318 79800 -6294 80120
rect -5974 79800 -5950 80120
rect -6318 79776 -5950 79800
rect -3786 80120 -3418 80144
rect -2946 80120 -2626 82638
rect -3786 79800 -3762 80120
rect -3442 79982 -2626 80120
rect -3442 79800 -2994 79982
rect -3786 79776 -3418 79800
rect -3018 79662 -2994 79800
rect -2674 79662 -2626 79982
rect -1526 82052 -1206 82640
rect -1526 81780 -1502 82052
rect -1230 81780 -1206 82052
rect -1526 79960 -1206 81780
rect -3018 79638 -2626 79662
rect -1528 79640 -1206 79960
rect -5546 79076 -5178 79100
rect -5546 78756 -5522 79076
rect -5202 78756 -5178 79076
rect -5546 78732 -5178 78756
rect -6318 77120 -5950 77144
rect -6318 76800 -6294 77120
rect -5974 76800 -5950 77120
rect -6318 76776 -5950 76800
rect -3786 77120 -3418 77144
rect -2946 77120 -2626 79638
rect -3786 76800 -3762 77120
rect -3442 76982 -2626 77120
rect -3442 76800 -2994 76982
rect -3786 76776 -3418 76800
rect -3018 76662 -2994 76800
rect -2674 76662 -2626 76982
rect -1526 79052 -1206 79640
rect -1526 78780 -1502 79052
rect -1230 78780 -1206 79052
rect -1526 76960 -1206 78780
rect -3018 76638 -2626 76662
rect -1528 76640 -1206 76960
rect -5546 76076 -5178 76100
rect -5546 75756 -5522 76076
rect -5202 75756 -5178 76076
rect -5546 75732 -5178 75756
rect -6318 74120 -5950 74144
rect -6318 73800 -6294 74120
rect -5974 73800 -5950 74120
rect -6318 73776 -5950 73800
rect -3786 74120 -3418 74144
rect -2946 74120 -2626 76638
rect -3786 73800 -3762 74120
rect -3442 73982 -2626 74120
rect -3442 73800 -2994 73982
rect -3786 73776 -3418 73800
rect -3018 73662 -2994 73800
rect -2674 73662 -2626 73982
rect -1526 76052 -1206 76640
rect -1526 75780 -1502 76052
rect -1230 75780 -1206 76052
rect -1526 73960 -1206 75780
rect -3018 73638 -2626 73662
rect -1528 73640 -1206 73960
rect -5546 73076 -5178 73100
rect -5546 72756 -5522 73076
rect -5202 72756 -5178 73076
rect -5546 72732 -5178 72756
rect -6318 71120 -5950 71144
rect -6318 70800 -6294 71120
rect -5974 70800 -5950 71120
rect -6318 70776 -5950 70800
rect -3786 71120 -3418 71144
rect -2946 71120 -2626 73638
rect -3786 70800 -3762 71120
rect -3442 70982 -2626 71120
rect -3442 70800 -2994 70982
rect -3786 70776 -3418 70800
rect -3018 70662 -2994 70800
rect -2674 70662 -2626 70982
rect -1526 73052 -1206 73640
rect -1526 72780 -1502 73052
rect -1230 72780 -1206 73052
rect -1526 70960 -1206 72780
rect -3018 70638 -2626 70662
rect -1528 70640 -1206 70960
rect -5546 70076 -5178 70100
rect -5546 69756 -5522 70076
rect -5202 69756 -5178 70076
rect -5546 69732 -5178 69756
rect -6318 68120 -5950 68144
rect -6318 67800 -6294 68120
rect -5974 67800 -5950 68120
rect -6318 67776 -5950 67800
rect -3786 68120 -3418 68144
rect -2946 68120 -2626 70638
rect -3786 67800 -3762 68120
rect -3442 67982 -2626 68120
rect -3442 67800 -2994 67982
rect -3786 67776 -3418 67800
rect -3018 67662 -2994 67800
rect -2674 67662 -2626 67982
rect -1526 70052 -1206 70640
rect -1526 69780 -1502 70052
rect -1230 69780 -1206 70052
rect -1526 67960 -1206 69780
rect -3018 67638 -2626 67662
rect -1528 67640 -1206 67960
rect -5546 67076 -5178 67100
rect -5546 66756 -5522 67076
rect -5202 66756 -5178 67076
rect -5546 66732 -5178 66756
rect -6318 65120 -5950 65144
rect -6318 64800 -6294 65120
rect -5974 64800 -5950 65120
rect -6318 64776 -5950 64800
rect -3786 65120 -3418 65144
rect -2946 65120 -2626 67638
rect -3786 64800 -3762 65120
rect -3442 64982 -2626 65120
rect -3442 64800 -2994 64982
rect -3786 64776 -3418 64800
rect -3018 64662 -2994 64800
rect -2674 64662 -2626 64982
rect -1526 67052 -1206 67640
rect -1526 66780 -1502 67052
rect -1230 66780 -1206 67052
rect -1526 64960 -1206 66780
rect -3018 64638 -2626 64662
rect -1528 64640 -1206 64960
rect -5546 64076 -5178 64100
rect -5546 63756 -5522 64076
rect -5202 63756 -5178 64076
rect -5546 63732 -5178 63756
rect -6318 62120 -5950 62144
rect -6318 61800 -6294 62120
rect -5974 61800 -5950 62120
rect -6318 61776 -5950 61800
rect -3786 62120 -3418 62144
rect -2946 62120 -2626 64638
rect -3786 61800 -3762 62120
rect -3442 61982 -2626 62120
rect -3442 61800 -2994 61982
rect -3786 61776 -3418 61800
rect -3018 61662 -2994 61800
rect -2674 61662 -2626 61982
rect -1526 64052 -1206 64640
rect -1526 63780 -1502 64052
rect -1230 63780 -1206 64052
rect -1526 61960 -1206 63780
rect -3018 61638 -2626 61662
rect -1528 61640 -1206 61960
rect -5546 61076 -5178 61100
rect -5546 60756 -5522 61076
rect -5202 60756 -5178 61076
rect -5546 60732 -5178 60756
rect -6318 59120 -5950 59144
rect -6318 58800 -6294 59120
rect -5974 58800 -5950 59120
rect -6318 58776 -5950 58800
rect -3786 59120 -3418 59144
rect -2946 59120 -2626 61638
rect -3786 58800 -3762 59120
rect -3442 58982 -2626 59120
rect -3442 58800 -2994 58982
rect -3786 58776 -3418 58800
rect -3018 58662 -2994 58800
rect -2674 58662 -2626 58982
rect -1526 61052 -1206 61640
rect -1526 60780 -1502 61052
rect -1230 60780 -1206 61052
rect -1526 58960 -1206 60780
rect -3018 58638 -2626 58662
rect -1528 58640 -1206 58960
rect -5546 58076 -5178 58100
rect -5546 57756 -5522 58076
rect -5202 57756 -5178 58076
rect -5546 57732 -5178 57756
rect -2946 56120 -2626 58638
rect -3120 55982 -2626 56120
rect -3120 55800 -2994 55982
rect -3018 55662 -2994 55800
rect -2674 55662 -2626 55982
rect -1526 58052 -1206 58640
rect -1526 57780 -1502 58052
rect -1230 57780 -1206 58052
rect -1526 55960 -1206 57780
rect -3018 55638 -2626 55662
rect -1528 55640 -1206 55960
rect -5546 55076 -5178 55100
rect -5546 54756 -5522 55076
rect -5202 54756 -5178 55076
rect -5546 54732 -5178 54756
rect -6318 53120 -5950 53144
rect -6318 52800 -6294 53120
rect -5974 52800 -5950 53120
rect -6318 52776 -5950 52800
rect -3786 53120 -3418 53144
rect -2946 53120 -2626 55638
rect -3786 52800 -3762 53120
rect -3442 52982 -2626 53120
rect -3442 52800 -2994 52982
rect -3786 52776 -3418 52800
rect -3018 52662 -2994 52800
rect -2674 52662 -2626 52982
rect -1526 55052 -1206 55640
rect -1526 54780 -1502 55052
rect -1230 54780 -1206 55052
rect -1526 52960 -1206 54780
rect -3018 52638 -2626 52662
rect -1528 52640 -1206 52960
rect -5546 52076 -5178 52100
rect -5546 51756 -5522 52076
rect -5202 51756 -5178 52076
rect -5546 51732 -5178 51756
rect -6318 50120 -5950 50144
rect -6318 49800 -6294 50120
rect -5974 49800 -5950 50120
rect -6318 49776 -5950 49800
rect -3786 50120 -3418 50144
rect -2946 50120 -2626 52638
rect -3786 49800 -3762 50120
rect -3442 49982 -2626 50120
rect -3442 49800 -2994 49982
rect -3786 49776 -3418 49800
rect -3018 49662 -2994 49800
rect -2674 49662 -2626 49982
rect -1526 52052 -1206 52640
rect -1526 51780 -1502 52052
rect -1230 51780 -1206 52052
rect -1526 49960 -1206 51780
rect -3018 49638 -2626 49662
rect -1528 49640 -1206 49960
rect -5546 49076 -5178 49100
rect -5546 48756 -5522 49076
rect -5202 48756 -5178 49076
rect -5546 48732 -5178 48756
rect -6318 47120 -5950 47144
rect -6318 46800 -6294 47120
rect -5974 46800 -5950 47120
rect -6318 46776 -5950 46800
rect -3786 47120 -3418 47144
rect -2946 47120 -2626 49638
rect -3786 46800 -3762 47120
rect -3442 46982 -2626 47120
rect -3442 46800 -2994 46982
rect -3786 46776 -3418 46800
rect -3018 46662 -2994 46800
rect -2674 46662 -2626 46982
rect -1526 49052 -1206 49640
rect -1526 48780 -1502 49052
rect -1230 48780 -1206 49052
rect -1526 46960 -1206 48780
rect -3018 46638 -2626 46662
rect -1528 46640 -1206 46960
rect -5546 46076 -5178 46100
rect -5546 45756 -5522 46076
rect -5202 45756 -5178 46076
rect -5546 45732 -5178 45756
rect -6318 44120 -5950 44144
rect -6318 43800 -6294 44120
rect -5974 43800 -5950 44120
rect -6318 43776 -5950 43800
rect -3786 44120 -3418 44144
rect -2946 44120 -2626 46638
rect -3786 43800 -3762 44120
rect -3442 43982 -2626 44120
rect -3442 43800 -2994 43982
rect -3786 43776 -3418 43800
rect -3018 43662 -2994 43800
rect -2674 43662 -2626 43982
rect -1526 46052 -1206 46640
rect -1526 45780 -1502 46052
rect -1230 45780 -1206 46052
rect -1526 43960 -1206 45780
rect -3018 43638 -2626 43662
rect -1528 43640 -1206 43960
rect -5546 43076 -5178 43100
rect -5546 42756 -5522 43076
rect -5202 42756 -5178 43076
rect -5546 42732 -5178 42756
rect -6318 41120 -5950 41144
rect -6318 40800 -6294 41120
rect -5974 40800 -5950 41120
rect -6318 40776 -5950 40800
rect -3786 41120 -3418 41144
rect -2946 41120 -2626 43638
rect -3786 40800 -3762 41120
rect -3442 40982 -2626 41120
rect -3442 40800 -2994 40982
rect -3786 40776 -3418 40800
rect -3018 40662 -2994 40800
rect -2674 40662 -2626 40982
rect -1526 43052 -1206 43640
rect -1526 42780 -1502 43052
rect -1230 42780 -1206 43052
rect -1526 40960 -1206 42780
rect -3018 40638 -2626 40662
rect -1528 40640 -1206 40960
rect -5546 40076 -5178 40100
rect -5546 39756 -5522 40076
rect -5202 39756 -5178 40076
rect -5546 39732 -5178 39756
rect -6318 38120 -5950 38144
rect -6318 37800 -6294 38120
rect -5974 37800 -5950 38120
rect -6318 37776 -5950 37800
rect -3786 38120 -3418 38144
rect -2946 38120 -2626 40638
rect -3786 37800 -3762 38120
rect -3442 37982 -2626 38120
rect -3442 37800 -2994 37982
rect -3786 37776 -3418 37800
rect -3018 37662 -2994 37800
rect -2674 37662 -2626 37982
rect -1526 40052 -1206 40640
rect -1526 39780 -1502 40052
rect -1230 39780 -1206 40052
rect -1526 37960 -1206 39780
rect -3018 37638 -2626 37662
rect -1528 37640 -1206 37960
rect -5546 37076 -5178 37100
rect -5546 36756 -5522 37076
rect -5202 36756 -5178 37076
rect -5546 36732 -5178 36756
rect -6318 35120 -5950 35144
rect -6318 34800 -6294 35120
rect -5974 34800 -5950 35120
rect -6318 34776 -5950 34800
rect -3786 35120 -3418 35144
rect -2946 35120 -2626 37638
rect -3786 34800 -3762 35120
rect -3442 34982 -2626 35120
rect -3442 34800 -2994 34982
rect -3786 34776 -3418 34800
rect -3018 34662 -2994 34800
rect -2674 34662 -2626 34982
rect -1526 37052 -1206 37640
rect -1526 36780 -1502 37052
rect -1230 36780 -1206 37052
rect -1526 34960 -1206 36780
rect -3018 34638 -2626 34662
rect -1528 34640 -1206 34960
rect -5546 34076 -5178 34100
rect -5546 33756 -5522 34076
rect -5202 33756 -5178 34076
rect -5546 33732 -5178 33756
rect -6318 32120 -5950 32144
rect -6318 31800 -6294 32120
rect -5974 31800 -5950 32120
rect -6318 31776 -5950 31800
rect -3786 32120 -3418 32144
rect -2946 32120 -2626 34638
rect -3786 31800 -3762 32120
rect -3442 31982 -2626 32120
rect -3442 31800 -2994 31982
rect -3786 31776 -3418 31800
rect -3018 31662 -2994 31800
rect -2674 31662 -2626 31982
rect -1526 34052 -1206 34640
rect -1526 33780 -1502 34052
rect -1230 33780 -1206 34052
rect -1526 31960 -1206 33780
rect -3018 31638 -2626 31662
rect -1528 31640 -1206 31960
rect -5546 31076 -5178 31100
rect -5546 30756 -5522 31076
rect -5202 30756 -5178 31076
rect -5546 30732 -5178 30756
rect -6318 29120 -5950 29144
rect -6318 28800 -6294 29120
rect -5974 28800 -5950 29120
rect -6318 28776 -5950 28800
rect -3786 29120 -3418 29144
rect -2946 29120 -2626 31638
rect -3786 28800 -3762 29120
rect -3442 28982 -2626 29120
rect -3442 28800 -2994 28982
rect -3786 28776 -3418 28800
rect -3018 28662 -2994 28800
rect -2674 28662 -2626 28982
rect -1526 31052 -1206 31640
rect -1526 30780 -1502 31052
rect -1230 30780 -1206 31052
rect -1526 28960 -1206 30780
rect -3018 28638 -2626 28662
rect -1528 28640 -1206 28960
rect -5546 28076 -5178 28100
rect -5546 27756 -5522 28076
rect -5202 27756 -5178 28076
rect -5546 27732 -5178 27756
rect -6318 26120 -5950 26144
rect -6318 25800 -6294 26120
rect -5974 25800 -5950 26120
rect -6318 25776 -5950 25800
rect -3786 26120 -3418 26144
rect -2946 26120 -2626 28638
rect -3786 25800 -3762 26120
rect -3442 25982 -2626 26120
rect -3442 25800 -2994 25982
rect -3786 25776 -3418 25800
rect -3018 25662 -2994 25800
rect -2674 25662 -2626 25982
rect -1526 28052 -1206 28640
rect -1526 27780 -1502 28052
rect -1230 27780 -1206 28052
rect -1526 25960 -1206 27780
rect -3018 25638 -2626 25662
rect -1528 25640 -1206 25960
rect -5546 25076 -5178 25100
rect -5546 24756 -5522 25076
rect -5202 24756 -5178 25076
rect -5546 24732 -5178 24756
rect -6318 23120 -5950 23144
rect -6318 22800 -6294 23120
rect -5974 22800 -5950 23120
rect -6318 22776 -5950 22800
rect -3786 23120 -3418 23144
rect -2946 23120 -2626 25638
rect -3786 22800 -3762 23120
rect -3442 22982 -2626 23120
rect -3442 22800 -2994 22982
rect -3786 22776 -3418 22800
rect -3018 22662 -2994 22800
rect -2674 22662 -2626 22982
rect -1526 25052 -1206 25640
rect -1526 24780 -1502 25052
rect -1230 24780 -1206 25052
rect -1526 22960 -1206 24780
rect -3018 22638 -2626 22662
rect -1528 22640 -1206 22960
rect -5546 22076 -5178 22100
rect -5546 21756 -5522 22076
rect -5202 21756 -5178 22076
rect -5546 21732 -5178 21756
rect -6318 20120 -5950 20144
rect -6318 19800 -6294 20120
rect -5974 19800 -5950 20120
rect -6318 19776 -5950 19800
rect -3786 20120 -3418 20144
rect -2946 20120 -2626 22638
rect -3786 19800 -3762 20120
rect -3442 19800 -2626 20120
rect -1526 22052 -1206 22640
rect -1526 21780 -1502 22052
rect -1230 21780 -1206 22052
rect -1526 19960 -1206 21780
rect 303888 318334 304300 321062
rect 303888 318062 303950 318334
rect 304222 318062 304300 318334
rect 303888 315334 304300 318062
rect 303888 315062 303950 315334
rect 304222 315062 304300 315334
rect 303888 312334 304300 315062
rect 303888 312062 303950 312334
rect 304222 312062 304300 312334
rect 303888 309334 304300 312062
rect 303888 309062 303950 309334
rect 304222 309062 304300 309334
rect 303888 306334 304300 309062
rect 303888 306062 303950 306334
rect 304222 306062 304300 306334
rect 303888 303334 304300 306062
rect 303888 303062 303950 303334
rect 304222 303062 304300 303334
rect 303888 300334 304300 303062
rect 303888 300062 303950 300334
rect 304222 300062 304300 300334
rect 303888 297334 304300 300062
rect 303888 297062 303950 297334
rect 304222 297062 304300 297334
rect 303888 294334 304300 297062
rect 303888 294062 303950 294334
rect 304222 294062 304300 294334
rect 303888 291334 304300 294062
rect 303888 291062 303950 291334
rect 304222 291062 304300 291334
rect 303888 288334 304300 291062
rect 303888 288062 303950 288334
rect 304222 288062 304300 288334
rect 303888 285334 304300 288062
rect 303888 285062 303950 285334
rect 304222 285062 304300 285334
rect 303888 282334 304300 285062
rect 303888 282062 303950 282334
rect 304222 282062 304300 282334
rect 303888 279334 304300 282062
rect 303888 279062 303950 279334
rect 304222 279062 304300 279334
rect 303888 276334 304300 279062
rect 303888 276062 303950 276334
rect 304222 276062 304300 276334
rect 303888 273334 304300 276062
rect 303888 273062 303950 273334
rect 304222 273062 304300 273334
rect 303888 270334 304300 273062
rect 303888 270062 303950 270334
rect 304222 270062 304300 270334
rect 303888 267334 304300 270062
rect 303888 267062 303950 267334
rect 304222 267062 304300 267334
rect 303888 264334 304300 267062
rect 303888 264062 303950 264334
rect 304222 264062 304300 264334
rect 303888 261334 304300 264062
rect 303888 261062 303950 261334
rect 304222 261062 304300 261334
rect 303888 258334 304300 261062
rect 303888 258062 303950 258334
rect 304222 258062 304300 258334
rect 303888 255334 304300 258062
rect 303888 255062 303950 255334
rect 304222 255062 304300 255334
rect 303888 252334 304300 255062
rect 303888 252062 303950 252334
rect 304222 252062 304300 252334
rect 303888 249334 304300 252062
rect 303888 249062 303950 249334
rect 304222 249062 304300 249334
rect 303888 246334 304300 249062
rect 303888 246062 303950 246334
rect 304222 246062 304300 246334
rect 303888 243334 304300 246062
rect 303888 243062 303950 243334
rect 304222 243062 304300 243334
rect 303888 240334 304300 243062
rect 303888 240062 303950 240334
rect 304222 240062 304300 240334
rect 303888 237334 304300 240062
rect 303888 237062 303950 237334
rect 304222 237062 304300 237334
rect 303888 234334 304300 237062
rect 303888 234062 303950 234334
rect 304222 234062 304300 234334
rect 303888 231334 304300 234062
rect 303888 231062 303950 231334
rect 304222 231062 304300 231334
rect 303888 228334 304300 231062
rect 303888 228062 303950 228334
rect 304222 228062 304300 228334
rect 303888 225334 304300 228062
rect 303888 225062 303950 225334
rect 304222 225062 304300 225334
rect 303888 222334 304300 225062
rect 303888 222062 303950 222334
rect 304222 222062 304300 222334
rect 303888 219334 304300 222062
rect 303888 219062 303950 219334
rect 304222 219062 304300 219334
rect 303888 216334 304300 219062
rect 303888 216062 303950 216334
rect 304222 216062 304300 216334
rect 303888 213334 304300 216062
rect 303888 213062 303950 213334
rect 304222 213062 304300 213334
rect 303888 210334 304300 213062
rect 303888 210062 303950 210334
rect 304222 210062 304300 210334
rect 303888 207334 304300 210062
rect 303888 207062 303950 207334
rect 304222 207062 304300 207334
rect 303888 204334 304300 207062
rect 303888 204062 303950 204334
rect 304222 204062 304300 204334
rect 303888 201334 304300 204062
rect 303888 201062 303950 201334
rect 304222 201062 304300 201334
rect 303888 198334 304300 201062
rect 303888 198062 303950 198334
rect 304222 198062 304300 198334
rect 303888 195334 304300 198062
rect 303888 195062 303950 195334
rect 304222 195062 304300 195334
rect 303888 192334 304300 195062
rect 303888 192062 303950 192334
rect 304222 192062 304300 192334
rect 303888 189334 304300 192062
rect 303888 189062 303950 189334
rect 304222 189062 304300 189334
rect 303888 186334 304300 189062
rect 303888 186062 303950 186334
rect 304222 186062 304300 186334
rect 303888 183334 304300 186062
rect 303888 183062 303950 183334
rect 304222 183062 304300 183334
rect 303888 180334 304300 183062
rect 303888 180062 303950 180334
rect 304222 180062 304300 180334
rect 303888 177334 304300 180062
rect 303888 177062 303950 177334
rect 304222 177062 304300 177334
rect 303888 174334 304300 177062
rect 303888 174062 303950 174334
rect 304222 174062 304300 174334
rect 303888 171334 304300 174062
rect 303888 171062 303950 171334
rect 304222 171062 304300 171334
rect 303888 168334 304300 171062
rect 303888 168062 303950 168334
rect 304222 168062 304300 168334
rect 303888 165334 304300 168062
rect 303888 165062 303950 165334
rect 304222 165062 304300 165334
rect 303888 162334 304300 165062
rect 303888 162062 303950 162334
rect 304222 162062 304300 162334
rect 303888 159334 304300 162062
rect 303888 159062 303950 159334
rect 304222 159062 304300 159334
rect 303888 156334 304300 159062
rect 303888 156062 303950 156334
rect 304222 156062 304300 156334
rect 303888 153334 304300 156062
rect 303888 153062 303950 153334
rect 304222 153062 304300 153334
rect 303888 150334 304300 153062
rect 303888 150062 303950 150334
rect 304222 150062 304300 150334
rect 303888 147334 304300 150062
rect 303888 147062 303950 147334
rect 304222 147062 304300 147334
rect 303888 144334 304300 147062
rect 303888 144062 303950 144334
rect 304222 144062 304300 144334
rect 303888 141334 304300 144062
rect 303888 141062 303950 141334
rect 304222 141062 304300 141334
rect 303888 138334 304300 141062
rect 303888 138062 303950 138334
rect 304222 138062 304300 138334
rect 303888 135334 304300 138062
rect 303888 135062 303950 135334
rect 304222 135062 304300 135334
rect 303888 132334 304300 135062
rect 303888 132062 303950 132334
rect 304222 132062 304300 132334
rect 303888 129334 304300 132062
rect 303888 129062 303950 129334
rect 304222 129062 304300 129334
rect 303888 126334 304300 129062
rect 303888 126062 303950 126334
rect 304222 126062 304300 126334
rect 303888 123334 304300 126062
rect 303888 123062 303950 123334
rect 304222 123062 304300 123334
rect 303888 120334 304300 123062
rect 303888 120062 303950 120334
rect 304222 120062 304300 120334
rect 303888 117334 304300 120062
rect 303888 117062 303950 117334
rect 304222 117062 304300 117334
rect 303888 114334 304300 117062
rect 303888 114062 303950 114334
rect 304222 114062 304300 114334
rect 303888 111334 304300 114062
rect 303888 111062 303950 111334
rect 304222 111062 304300 111334
rect 303888 108334 304300 111062
rect 303888 108062 303950 108334
rect 304222 108062 304300 108334
rect 303888 105334 304300 108062
rect 303888 105062 303950 105334
rect 304222 105062 304300 105334
rect 303888 102334 304300 105062
rect 303888 102062 303950 102334
rect 304222 102062 304300 102334
rect 303888 99334 304300 102062
rect 303888 99062 303950 99334
rect 304222 99062 304300 99334
rect 303888 96334 304300 99062
rect 303888 96062 303950 96334
rect 304222 96062 304300 96334
rect 303888 93334 304300 96062
rect 303888 93062 303950 93334
rect 304222 93062 304300 93334
rect 303888 90334 304300 93062
rect 303888 90062 303950 90334
rect 304222 90062 304300 90334
rect 303888 87334 304300 90062
rect 303888 87062 303950 87334
rect 304222 87062 304300 87334
rect 303888 84334 304300 87062
rect 303888 84062 303950 84334
rect 304222 84062 304300 84334
rect 303888 81334 304300 84062
rect 303888 81062 303950 81334
rect 304222 81062 304300 81334
rect 303888 78334 304300 81062
rect 303888 78062 303950 78334
rect 304222 78062 304300 78334
rect 303888 75334 304300 78062
rect 303888 75062 303950 75334
rect 304222 75062 304300 75334
rect 303888 72334 304300 75062
rect 303888 72062 303950 72334
rect 304222 72062 304300 72334
rect 303888 69334 304300 72062
rect 303888 69062 303950 69334
rect 304222 69062 304300 69334
rect 303888 66334 304300 69062
rect 303888 66062 303950 66334
rect 304222 66062 304300 66334
rect 303888 63334 304300 66062
rect 303888 63062 303950 63334
rect 304222 63062 304300 63334
rect 303888 60334 304300 63062
rect 303888 60062 303950 60334
rect 304222 60062 304300 60334
rect 303888 57334 304300 60062
rect 303888 57062 303950 57334
rect 304222 57062 304300 57334
rect 303888 54334 304300 57062
rect 303888 54062 303950 54334
rect 304222 54062 304300 54334
rect 303888 51334 304300 54062
rect 303888 51062 303950 51334
rect 304222 51062 304300 51334
rect 303888 48334 304300 51062
rect 303888 48062 303950 48334
rect 304222 48062 304300 48334
rect 303888 45334 304300 48062
rect 303888 45062 303950 45334
rect 304222 45062 304300 45334
rect 303888 42334 304300 45062
rect 303888 42062 303950 42334
rect 304222 42062 304300 42334
rect 303888 39334 304300 42062
rect 303888 39062 303950 39334
rect 304222 39062 304300 39334
rect 303888 36334 304300 39062
rect 303888 36062 303950 36334
rect 304222 36062 304300 36334
rect 303888 33334 304300 36062
rect 303888 33062 303950 33334
rect 304222 33062 304300 33334
rect 303888 30334 304300 33062
rect 303888 30062 303950 30334
rect 304222 30062 304300 30334
rect 303888 27334 304300 30062
rect 303888 27062 303950 27334
rect 304222 27062 304300 27334
rect 303888 24334 304300 27062
rect 303888 24062 303950 24334
rect 304222 24062 304300 24334
rect 303888 21372 304300 24062
rect 303888 21334 304304 21372
rect 303888 21062 303950 21334
rect 304222 21062 304304 21334
rect 303888 21004 304304 21062
rect 303888 20952 304300 21004
rect -3786 19776 -3418 19800
rect -5546 19076 -5178 19100
rect -5546 18756 -5522 19076
rect -5202 18756 -5178 19076
rect -5546 18732 -5178 18756
rect -6414 18026 -6094 18186
rect -6438 18002 -6070 18026
rect -6438 17682 -6414 18002
rect -6094 17960 -6070 18002
rect -6094 17734 -5984 17960
rect -6094 17682 -6070 17734
rect -6438 17658 -6070 17682
rect -6414 17374 -6094 17658
rect -2946 17288 -2626 19800
rect -1528 19640 -1206 19960
rect -1526 19052 -1206 19640
rect -1526 18780 -1502 19052
rect -1230 18780 -1206 19052
rect 303926 19273 304246 20952
rect -1526 18760 -1206 18780
rect 289572 18760 289952 18790
rect 303926 18768 304262 19273
rect 302310 18760 304262 18768
rect -1578 18718 304262 18760
rect -1578 18440 302945 18718
rect 289572 18422 289952 18440
rect 301985 18395 302945 18440
rect 302921 18394 302945 18395
rect 303267 18446 304262 18718
rect 303267 18395 303850 18446
rect 303267 18394 303291 18395
rect 302921 18370 303291 18394
rect 305436 17288 305756 326222
rect -2982 17264 305756 17288
rect -2982 16992 303890 17264
rect 304162 16992 305756 17264
rect -2982 16968 305756 16992
rect -2946 16904 -2626 16968
rect 644 16874 964 16968
rect 3644 16874 3964 16968
rect 6644 16874 6964 16968
rect 9644 16874 9964 16968
rect 12644 16874 12964 16968
rect 15644 16874 15964 16968
rect 18644 16874 18964 16968
rect 21644 16874 21964 16968
rect 24644 16874 24964 16968
rect 27644 16874 27964 16968
rect 30644 16874 30964 16968
rect 33644 16874 33964 16968
rect 36644 16874 36964 16968
rect 39644 16874 39964 16968
rect 42644 16874 42964 16968
rect 45644 16874 45964 16968
rect 48644 16874 48964 16968
rect 51644 16874 51964 16968
rect 54644 16874 54964 16968
rect 57644 16874 57964 16968
rect 60644 16874 60964 16968
rect 63644 16874 63964 16968
rect 66644 16874 66964 16968
rect 69644 16874 69964 16968
rect 72644 16874 72964 16968
rect 75644 16874 75964 16968
rect 78644 16874 78964 16968
rect 81644 16874 81964 16968
rect 84644 16874 84964 16968
rect 87644 16874 87964 16968
rect 90644 16874 90964 16968
rect 93644 16874 93964 16968
rect 96644 16874 96964 16968
rect 99644 16874 99964 16968
rect 102644 16874 102964 16968
rect 105644 16874 105964 16968
rect 108644 16874 108964 16968
rect 111644 16874 111964 16968
rect 114644 16874 114964 16968
rect 117644 16874 117964 16968
rect 120644 16874 120964 16968
rect 123644 16874 123964 16968
rect 126644 16874 126964 16968
rect 129644 16874 129964 16968
rect 132644 16874 132964 16968
rect 135644 16874 135964 16968
rect 138644 16874 138964 16968
rect 141644 16874 141964 16968
rect 144644 16874 144964 16968
rect 147644 16874 147964 16968
rect 150644 16874 150964 16968
rect 153644 16874 153964 16968
rect 156644 16874 156964 16968
rect 159644 16874 159964 16968
rect 162644 16874 162964 16968
rect 165644 16874 165964 16968
rect 168644 16874 168964 16968
rect 171644 16874 171964 16968
rect 174644 16874 174964 16968
rect 177644 16874 177964 16968
rect 180644 16874 180964 16968
rect 183644 16874 183964 16968
rect 186644 16874 186964 16968
rect 189644 16874 189964 16968
rect 192644 16874 192964 16968
rect 195644 16874 195964 16968
rect 198644 16874 198964 16968
rect 201644 16874 201964 16968
rect 204644 16874 204964 16968
rect 207644 16874 207964 16968
rect 210644 16874 210964 16968
rect 213644 16874 213964 16968
rect 216644 16874 216964 16968
rect 219644 16874 219964 16968
rect 222644 16874 222964 16968
rect 225644 16874 225964 16968
rect 228644 16874 228964 16968
rect 231644 16874 231964 16968
rect 234644 16874 234964 16968
rect 237644 16874 237964 16968
rect 240644 16874 240964 16968
rect 243644 16874 243964 16968
rect 246644 16874 246964 16968
rect 249644 16874 249964 16968
rect 252644 16874 252964 16968
rect 255644 16874 255964 16968
rect 258644 16874 258964 16968
rect 261644 16874 261964 16968
rect 264644 16874 264964 16968
rect 270644 16874 270964 16968
rect 273644 16874 273964 16968
rect 276644 16874 276964 16968
rect 279644 16874 279964 16968
rect 282644 16874 282964 16968
rect 285644 16874 285964 16968
rect 288644 16874 288964 16968
rect 291644 16874 291964 16968
rect 294644 16874 294964 16968
rect 297644 16874 297964 16968
rect 300644 16874 300964 16968
rect 302888 16410 303316 16448
rect 302888 16088 302940 16410
rect 303274 16088 303316 16410
rect 302888 16064 303316 16088
rect 306874 16048 307194 16842
rect 303842 15692 304210 15716
rect 24 15642 392 15666
rect 24 15322 48 15642
rect 368 15322 836 15642
rect 303842 15372 303866 15692
rect 304186 15372 304210 15692
rect 303842 15348 304210 15372
rect 24 15298 392 15322
use pixel_array100x100_fill  pixel_array100x100_fill_0
timestamp 1758314889
transform 1 0 2108 0 1 317378
box -3000 -298600 300740 5000
use shift_registerC  shift_registerC_0
timestamp 1758314889
transform 1 0 58 0 1 590
box -1076 -4 307988 16000
use shift_registerC  shift_registerC_1
timestamp 1758314889
transform 0 1 -21068 -1 0 323980
box -1076 -4 307988 16000
<< labels >>
rlabel metal5 -2842 18750 -2834 18760 1 VDD
port 1 n
rlabel metal5 -1354 19538 -1354 19538 1 GND
port 2 n
rlabel space 306642 6498 306642 6498 1 COL_ENA
port 3 n
rlabel metal3 306826 6496 306826 6496 1 COL_ENA
port 3 n
rlabel metal3 306748 10568 306748 10568 1 COL_RST
port 4 n
rlabel metal3 306704 14532 306704 14532 1 COL_DIN
port 5 n
rlabel metal3 306718 2558 306718 2558 1 COL_CLK
port 6 n
rlabel metal4 -4276 14472 -4276 14472 1 CSA_VREF
port 8 n
rlabel metal2 304782 19400 304782 19400 1 ARRAY_OUT
port 9 n
rlabel metal2 1414 325058 1414 325058 1 NB1
port 10 n
rlabel metal2 2166 325646 2166 325646 1 NB2
port 11 n
rlabel metal4 -7482 325904 -7482 325904 1 VBIAS
port 12 n
rlabel metal2 -7646 325424 -7614 325458 1 VREF
port 13 n
rlabel metal3 942 325236 942 325236 1 SF_IB
port 14 n
rlabel metal3 -7150 17524 -7150 17524 1 ROW_DIN
port 16 n
rlabel metal3 -11058 17572 -11058 17572 1 ROW_RST
port 17 n
rlabel metal3 -15162 17518 -15162 17518 1 ROW_ENA
port 18 n
rlabel metal3 -19086 17484 -19086 17484 1 ROW_CLK
port 19 n
rlabel metal5 666 320402 666 320402 1 gring
port 20 n
<< end >>
