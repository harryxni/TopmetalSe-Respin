* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt pixel gring VDD GND VREF ROW_SEL NB1 VBIAS NB2 AMP_IN SF_IB PIX_OUT CSA_VREF
X0 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5 pd=7.5 as=25.284374 ps=56.25 w=2 l=2
X1 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.2925 pd=2.2 as=1.57 ps=12.3 w=0.65 l=0.65
X2 a_4120_n520# VBIAS a_4120_n750# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.995 ps=8.8 w=1 l=0.8
X3 a_5720_n730# a_4600_n810# GND VDD sky130_fd_pr__pfet_01v8_lvt ad=0.25 pd=1.5 as=0.35 ps=2.7 w=1 l=1
X4 VDD SF_IB a_5720_n730# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.25 ps=1.5 w=1 l=1
X5 a_5460_10# a_4350_10# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X6 a_3860_n520# VBIAS a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.76 ps=8.8 w=1 l=0.8
X7 VDD a_4120_n520# a_4600_n810# GND sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=1
X8 a_4350_10# a_3860_n520# a_3860_n520# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X9 a_4120_n750# AMP_IN a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=1.995 pd=8.8 as=1.4 ps=7.4 w=7 l=0.15
X10 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.119375 pd=7.15 as=0 ps=0 w=2 l=3.35
X11 a_4120_n520# a_3860_n520# a_5460_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X12 GND NB1 a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0.42 pd=3.1 as=0.42 ps=3.1 w=1.2 l=1
X13 a_5750_n920# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=0.6 pd=2.95 as=5.4 ps=9.4 w=2 l=1
X14 a_4050_n2590# VREF a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=1.4 pd=7.4 as=1.76 ps=8.8 w=7 l=0.15
X15 a_4600_n810# NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1.15
X16 AMP_IN a_4600_n810# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VDD a_4350_10# a_4350_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X18 VDD a_5720_n730# a_5750_n920# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.6 ps=2.95 w=1 l=0.15
X19 AMP_IN CSA_VREF a_4600_n810# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.294 pd=2.24 as=0.273 ps=2.14 w=0.42 l=8
X20 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=10.715 pd=15.9 as=0 ps=0 w=2.6 l=0.35
.ends

.subckt pixel_array VBIAS VREF NB2 SF_IB CSA_VREF NB1 ROW_SEL0 ROW_SEL1 ROW_SEL2 PIX0_IN
+ GRING PIX1_IN PIX2_IN PIX3_IN PIX4_IN PIX5_IN PIX6_IN PIX_OUT0 PIX7_IN PIX_OUT1
+ PIX8_IN PIX_OUT2 ARRAY_OUT COL_SEL0 COL_SEl1 COL_SEL2 VDD GND
Xpixel_0 GRING VDD GND VREF ROW_SEL0 NB1 VBIAS NB2 PIX0_IN SF_IB PIX_OUT0 CSA_VREF
+ pixel
Xpixel_1 GRING VDD GND VREF ROW_SEL0 NB1 VBIAS NB2 PIX1_IN SF_IB PIX_OUT1 CSA_VREF
+ pixel
Xpixel_2 GRING VDD GND VREF ROW_SEL0 NB1 VBIAS NB2 PIX2_IN SF_IB PIX_OUT2 CSA_VREF
+ pixel
Xpixel_3 GRING VDD GND VREF ROW_SEL1 NB1 VBIAS NB2 PIX3_IN SF_IB PIX_OUT0 CSA_VREF
+ pixel
Xpixel_5 GRING VDD GND VREF ROW_SEL1 NB1 VBIAS NB2 PIX5_IN SF_IB PIX_OUT2 CSA_VREF
+ pixel
Xpixel_4 GRING VDD GND VREF ROW_SEL1 NB1 VBIAS NB2 PIX4_IN SF_IB PIX_OUT1 CSA_VREF
+ pixel
Xpixel_6 GRING VDD GND VREF ROW_SEL2 NB1 VBIAS NB2 PIX6_IN SF_IB PIX_OUT0 CSA_VREF
+ pixel
Xpixel_7 GRING VDD GND VREF ROW_SEL2 NB1 VBIAS NB2 PIX7_IN SF_IB PIX_OUT1 CSA_VREF
+ pixel
Xpixel_8 GRING VDD GND VREF ROW_SEL2 NB1 VBIAS NB2 PIX8_IN SF_IB PIX_OUT2 CSA_VREF
+ pixel
X0 PIX_OUT2 COL_SEL2 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X1 PIX_OUT1 COL_SEl1 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X2 PIX_OUT0 COL_SEL0 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
.ends

.subckt marker_pixel gring VDD GND VREF ROW_SEL NB1 VBIAS NB2 AMP_IN SF_IB PIX_OUT
+ CSA_VREF
X0 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5 pd=7.5 as=25.284374 ps=56.25 w=2 l=2
X1 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.2925 pd=2.2 as=1.57 ps=12.3 w=0.65 l=0.65
X2 a_4120_n520# VBIAS a_4120_n750# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.995 ps=8.8 w=1 l=0.8
X3 a_5720_n730# a_4600_n810# GND VDD sky130_fd_pr__pfet_01v8_lvt ad=0.25 pd=1.5 as=0.35 ps=2.7 w=1 l=1
X4 VDD SF_IB a_5720_n730# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.25 ps=1.5 w=1 l=1
X5 a_5460_10# a_4350_10# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X6 a_3860_n520# VBIAS a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.76 ps=8.8 w=1 l=0.8
X7 VDD a_4120_n520# a_4600_n810# GND sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=1
X8 a_4350_10# a_3860_n520# a_3860_n520# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X9 a_4120_n750# AMP_IN a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=1.995 pd=8.8 as=1.4 ps=7.4 w=7 l=0.15
X10 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.119375 pd=7.15 as=0 ps=0 w=2 l=3.35
X11 a_4120_n520# a_3860_n520# a_5460_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X12 GND NB1 a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0.42 pd=3.1 as=0.42 ps=3.1 w=1.2 l=1
X13 a_5750_n920# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=0.6 pd=2.95 as=5.4 ps=9.4 w=2 l=1
X14 a_4050_n2590# a_4020_n2258# a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=1.4 pd=7.4 as=1.76 ps=8.8 w=7 l=0.15
X15 a_4600_n810# NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1.15
X16 AMP_IN a_4600_n810# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VDD a_4350_10# a_4350_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X18 VDD a_5720_n730# a_5750_n920# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.6 ps=2.95 w=1 l=0.15
X19 AMP_IN CSA_VREF a_4600_n810# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.294 pd=2.24 as=0.273 ps=2.14 w=0.42 l=8
X20 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=10.715 pd=15.9 as=0 ps=0 w=2.6 l=0.35
.ends

.subckt pixel_array100x100 VBIAS VREF NB2 NB1 ROW_SEL[0] GRING ROW_SEL[1] ROW_SEL[2]
+ ROW_SEL[3] ROW_SEL[4] ROW_SEL[5] ROW_SEL[6] ROW_SEL[7] ROW_SEL[8] ROW_SEL[9] ROW_SEL[10]
+ ROW_SEL[11] ROW_SEL[12] ROW_SEL[13] ROW_SEL[14] ROW_SEL[15] ROW_SEL[16] ROW_SEL[17]
+ ROW_SEL[18] ROW_SEL[19] ROW_SEL[20] ROW_SEL[21] ROW_SEL[22] ROW_SEL[23] ROW_SEL[24]
+ ROW_SEL[25] ROW_SEL[26] ROW_SEL[27] ROW_SEL[28] ROW_SEL[29] ROW_SEL[30] ROW_SEL[31]
+ ROW_SEL[32] ROW_SEL[33] ROW_SEL[34] ROW_SEL[35] ROW_SEL[36] ROW_SEL[37] ROW_SEL[38]
+ ROW_SEL[39] ROW_SEL[40] ROW_SEL[41] ROW_SEL[42] ROW_SEL[43] ROW_SEL[44] ROW_SEL[45]
+ ROW_SEL[46] ROW_SEL[47] ROW_SEL[48] ROW_SEL[49] ROW_SEL[50] ROW_SEL[51] ROW_SEL[52]
+ ROW_SEL[53] ROW_SEL[54] ROW_SEL[55] ROW_SEL[56] ROW_SEL[57] ROW_SEL[58] ROW_SEL[59]
+ ROW_SEL[60] ROW_SEL[61] ROW_SEL[62] ROW_SEL[63] ROW_SEL[64] ROW_SEL[65] ROW_SEL[66]
+ ROW_SEL[67] ROW_SEL[68] ROW_SEL[69] ROW_SEL[70] ROW_SEL[71] ROW_SEL[72] ROW_SEL[73]
+ ROW_SEL[74] ROW_SEL[75] ROW_SEL[76] ROW_SEL[77] ROW_SEL[78] ROW_SEL[79] ROW_SEL[80]
+ ROW_SEL[81] ROW_SEL[82] ROW_SEL[83] ROW_SEL[84] ROW_SEL[85] ROW_SEL[86] ROW_SEL[87]
+ ROW_SEL[88] ROW_SEL[89] ROW_SEL[90] ROW_SEL[91] ROW_SEL[92] ROW_SEL[93] ROW_SEL[94]
+ ROW_SEL[95] ROW_SEL[96] ROW_SEL[97] ROW_SEL[98] COL_SEL[0] CSA_VREF ROW_SEL[99]
+ COL_SEL[1] COL_SEL[2] COL_SEL[3] COL_SEL[4] COL_SEL[5] COL_SEL[6] COL_SEL[7] COL_SEL[8]
+ COL_SEL[9] COL_SEL[10] COL_SEL[11] COL_SEL[12] COL_SEL[13] COL_SEL[14] COL_SEL[15]
+ COL_SEL[16] COL_SEL[17] COL_SEL[18] COL_SEL[19] COL_SEL[20] COL_SEL[21] COL_SEL[22]
+ COL_SEL[23] COL_SEL[24] COL_SEL[25] COL_SEL[26] COL_SEL[27] COL_SEL[28] COL_SEL[29]
+ COL_SEL[30] COL_SEL[31] COL_SEL[32] COL_SEL[33] COL_SEL[34] COL_SEL[35] COL_SEL[36]
+ COL_SEL[37] COL_SEL[38] COL_SEL[39] COL_SEL[40] COL_SEL[41] COL_SEL[42] COL_SEL[43]
+ COL_SEL[44] COL_SEL[45] COL_SEL[46] COL_SEL[47] COL_SEL[48] COL_SEL[49] COL_SEL[50]
+ COL_SEL[51] COL_SEL[52] COL_SEL[53] COL_SEL[54] COL_SEL[55] COL_SEL[56] COL_SEL[57]
+ COL_SEL[58] COL_SEL[59] COL_SEL[60] COL_SEL[61] COL_SEL[62] COL_SEL[63] COL_SEL[64]
+ COL_SEL[65] COL_SEL[66] COL_SEL[67] COL_SEL[68] COL_SEL[69] COL_SEL[70] COL_SEL[71]
+ COL_SEL[72] COL_SEL[73] COL_SEL[74] COL_SEL[75] COL_SEL[76] COL_SEL[77] COL_SEL[78]
+ COL_SEL[79] COL_SEL[80] COL_SEL[81] COL_SEL[82] COL_SEL[83] COL_SEL[84] COL_SEL[85]
+ COL_SEL[86] COL_SEL[87] COL_SEL[88] COL_SEL[89] COL_SEL[90] COL_SEL[91] COL_SEL[92]
+ COL_SEL[93] COL_SEL[94] COL_SEL[95] COL_SEL[96] COL_SEL[97] COL_SEL[98] ARRAY_OUT
+ COL_SEL[99] SF_IB VDD GND
Xpixel_9273 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9262 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9251 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8572 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8561 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8550 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9295 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9284 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8594 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8583 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7860 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7871 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7882 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7893 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5209 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_514 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_503 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4508 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_4519 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_547 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_536 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_525 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_3807 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_569 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_558 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3818 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_3829 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_7101 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7112 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7123 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_7134 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_7145 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7156 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6400 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6411 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7167 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7178 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7189 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_6422 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6433 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6444 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_6455 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6466 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6477 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5710 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5721 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5732 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_5743 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6488 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_6499 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_5754 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5765 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_5776 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_5787 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5798 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9081 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9081/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9070 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9070/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9092 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9092/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_8380 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8391 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_7690 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_81 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_81/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_70 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_70/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_92 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_92/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5006 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5006/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_5017 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5017/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5028 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5028/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_322 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_311 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_300 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5039 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5039/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_4305 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4316 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_4327 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_355 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_344 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_333 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3615 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_3604 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4338 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_4349 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_399 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_388 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_377 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_366 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_2914 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_2903 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_3648 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3637 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3626 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2947 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_2936 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2925 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_3659 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2969 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2958 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6230 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_6241 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6252 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6263 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_6274 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6285 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6296 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_5540 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5551 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_5562 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5573 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5584 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5595 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4850 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4861 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4872 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_4883 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4894 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1509 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9806 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_9839 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_9828 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9817 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_4102 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_130 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4113 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_4124 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4135 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_163 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_152 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_141 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3423 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3412 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_3401 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4146 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_4157 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4168 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_196 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_185 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_174 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_2722 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_2711 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2700 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_3467 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3456 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3445 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3434 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4179 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2755 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_2744 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2733 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3489 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3478 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2788 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_2777 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2766 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_2799 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_6060 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6060/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6071 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6071/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6082 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6082/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6093 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6093/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5370 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5381 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5392 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_4680 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4691 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3990 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_2018 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2018/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2007 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2007/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1306 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2029 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2029/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1339 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1328 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1317 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9603 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9614 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8902 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9625 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_9636 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9647 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_8946 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_8935 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8924 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8913 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9658 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_9669 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_8979 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_8968 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_8957 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3242 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3231 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3220 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2530 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3275 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3264 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3253 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2563 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2552 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2541 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3297 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_3286 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_1862 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_1851 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1840 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_2596 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2585 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_2574 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1895 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1884 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1873 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8209 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7508 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7519 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_6807 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6818 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6829 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1114 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1103 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_1147 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1136 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_1125 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1169 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_1158 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_9422 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9411 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9400 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8721 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_8710 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9455 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9444 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9433 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8754 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8743 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8732 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_9499 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_9488 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9477 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9466 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8787 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8776 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8765 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8798 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3050 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3050/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3083 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3083/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3072 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3072/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3061 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3061/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2382 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_2371 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2360 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3094 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3094/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1670 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2393 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1692 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1681 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_729 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_718 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_707 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8006 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8006/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8017 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8017/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8028 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8028/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_8039 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8039/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_7305 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7316 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7327 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7338 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7349 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6604 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_6615 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6626 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6637 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6648 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6659 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_5903 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5914 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5925 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5936 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5947 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_5958 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5969 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9230 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9274 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_9263 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9252 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_9241 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8562 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8551 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8540 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9296 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9285 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8595 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8584 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8573 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7850 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7861 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7872 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7883 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7894 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2190 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_504 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4509 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_548 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_537 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_526 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_515 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_559 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_3808 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_3819 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_7102 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7113 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_7124 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_7135 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7146 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6401 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7157 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_7168 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7179 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_6412 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_6423 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6434 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6445 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5700 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6456 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6467 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6478 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5711 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5722 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_5733 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6489 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_5744 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5755 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_5766 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_5777 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5788 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5799 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_9082 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9082/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9071 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9071/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9060 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9060/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9093 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9093/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_8370 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8381 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8392 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7680 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7691 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_6990 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_82 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_82/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_71 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_71/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_60 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_60/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_93 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_93/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5007 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5007/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5018 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5018/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5029 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5029/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_312 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_301 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4306 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4317 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_356 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_345 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_334 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_323 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3616 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_3605 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4328 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_4339 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_389 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_378 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_367 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_2904 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_3649 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3638 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3627 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2937 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_2926 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2915 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2959 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2948 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6220 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_6231 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6242 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6253 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6264 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6275 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6286 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5530 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5541 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6297 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5552 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_5563 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5574 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_5585 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4840 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5596 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4851 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4862 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_4873 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_890 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_4884 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4895 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9829 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_9818 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9807 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_131 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_120 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4103 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4114 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4125 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_164 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_153 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_142 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3424 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3413 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3402 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4136 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_4147 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4158 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4169 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_197 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_186 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_175 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_2712 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2701 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_3457 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3446 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3435 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2756 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_2745 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2734 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2723 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3479 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_3468 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2789 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2778 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2767 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6050 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6050/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6061 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6061/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6072 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6072/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_6083 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6083/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6094 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6094/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_5360 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5371 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5382 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5393 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_4670 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4681 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_4692 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3980 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_3991 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2008 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2008/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_2019 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2019/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1329 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1318 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_1307 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_9604 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_8903 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9615 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_9626 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9637 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9648 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8936 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8925 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8914 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_9659 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8969 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_8958 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8947 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3232 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3221 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_3210 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2531 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_2520 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_3265 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3254 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_3243 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2564 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_2553 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2542 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3298 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3287 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_3276 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1852 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_1841 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1830 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_2597 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2586 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2575 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1896 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_1885 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1874 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1863 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5190 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_7509 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6808 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6819 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1115 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1104 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_1148 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1137 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1126 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_1159 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9423 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_9412 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9401 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_8711 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8700 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9456 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_9445 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9434 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8744 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8733 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8722 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9489 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9478 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9467 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8788 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_8777 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8766 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8755 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_8799 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3040 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3040/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3084 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3084/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3073 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3073/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3062 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3062/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_3051 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3051/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_2372 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2361 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2350 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3095 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3095/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1660 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2394 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2383 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1693 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1682 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1671 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9990 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_719 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_708 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8007 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8007/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8018 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8018/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_8029 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8029/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_7306 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7317 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7328 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7339 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6605 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6616 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6627 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_6638 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6649 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_5904 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5915 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5926 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5937 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5948 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_5959 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9231 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9220 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9264 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9253 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9242 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8563 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8552 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8541 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8530 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9297 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9286 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9275 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8596 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8585 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8574 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7840 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_7851 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_7862 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7873 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7884 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_7895 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2180 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2191 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1490 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_505 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_538 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_527 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_516 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_549 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3809 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7103 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7114 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7125 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7136 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7147 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6402 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7158 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7169 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_6413 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6424 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6435 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_6446 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6457 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6468 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5701 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5712 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5723 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_5734 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6479 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5745 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5756 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_5767 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5778 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5789 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9072 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9072/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9061 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9061/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_9050 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9050/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9094 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9094/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_9083 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9083/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_8360 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_8371 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8382 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_8393 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_7670 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7681 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7692 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6980 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6991 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_72 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_72/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_61 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_61/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_50 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_50/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_94 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_94/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_83 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_83/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5008 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5008/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5019 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5019/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_313 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_302 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4307 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4318 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_346 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_335 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_324 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3606 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4329 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_379 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_368 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_357 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_2905 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_3639 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3628 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3617 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2938 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_2927 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2916 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2949 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6210 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_6221 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_6232 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6243 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6254 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_6265 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6276 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6287 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5520 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5531 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5542 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6298 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_5553 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5564 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_5575 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4830 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5586 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5597 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4841 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4852 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4863 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_4874 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_891 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_880 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4885 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4896 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8190 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9819 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9808 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_121 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_110 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4104 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4115 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4126 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_154 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_143 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_132 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3414 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3403 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4137 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_4148 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4159 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_198 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_187 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_176 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_165 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_2713 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_2702 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_3458 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3447 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3436 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_3425 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2746 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_2735 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2724 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3469 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2779 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2768 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2757 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6040 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6040/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_6051 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6051/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6062 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6062/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6073 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6073/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_6084 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6084/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6095 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6095/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_5350 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5361 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5372 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5383 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5394 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4660 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4671 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4682 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_4693 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3970 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_3981 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_3992 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_2 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_2/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2009 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2009/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1319 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1308 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_9605 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9616 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9627 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9638 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_8937 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_8926 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8915 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8904 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9649 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8959 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8948 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3233 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3222 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3211 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_3200 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2521 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2510 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_3266 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3255 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3244 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2554 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2543 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2532 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3299 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3288 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3277 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_1853 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_1842 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1831 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1820 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2598 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2587 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2576 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_2565 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1886 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_1875 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1864 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1897 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5180 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5191 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_4490 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_6809 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1105 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1138 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1127 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_1116 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_1149 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_9413 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9402 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_8712 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_8701 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9446 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9435 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9424 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8745 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8734 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8723 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_9479 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9468 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9457 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8778 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8767 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8756 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8789 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3041 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3041/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3030 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3030/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3074 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3074/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3063 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3063/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_3052 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3052/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2373 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_2362 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2351 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_2340 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3096 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3096/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_3085 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3085/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1661 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_1650 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_2395 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2384 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1694 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1683 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1672 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9980 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_9991 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_709 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8008 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8008/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8019 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8019/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_7307 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7318 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7329 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_6606 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6617 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6628 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6639 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_5905 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5916 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5927 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5938 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_5949 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_9221 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9210 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_8520 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9265 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_9254 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9243 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9232 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8553 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8542 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8531 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9298 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9287 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9276 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8586 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8575 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8564 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7830 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7841 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_7852 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8597 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_7863 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7874 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7885 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7896 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2181 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2170 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2192 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1491 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1480 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_539 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_528 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_517 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_506 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7104 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7115 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7126 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7137 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7148 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_7159 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_6403 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_6414 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6425 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6436 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_6447 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6458 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6469 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_5702 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5713 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_5724 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_5735 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5746 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_5757 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_5768 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5779 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9040 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9040/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9073 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9073/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9062 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9062/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9051 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9051/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_9095 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9095/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9084 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9084/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8350 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_8361 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8372 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8383 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_8394 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_7660 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7671 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7682 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7693 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_6970 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6981 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_73 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_73/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_62 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_62/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_51 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_51/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_40 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_40/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_6992 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_95 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_95/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_84 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_84/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5009 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5009/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_303 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4308 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_347 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_336 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_325 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_314 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3607 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4319 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_369 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_358 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3629 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3618 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2928 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_2917 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2906 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2939 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6200 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6211 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_6222 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6233 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6244 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_6255 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6266 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6277 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5510 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5521 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5532 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6288 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_6299 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_5543 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_5554 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5565 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_5576 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4820 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4831 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5587 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5598 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4842 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4853 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4864 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_892 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_881 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_870 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4875 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4886 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_4897 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_8180 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8191 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_7490 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9809 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_122 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_111 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_100 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4105 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4116 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_155 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_144 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_133 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3415 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_3404 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4127 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_4138 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_4149 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_188 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_177 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_166 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_2703 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_3448 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3437 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3426 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_199 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2747 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_2736 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2725 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2714 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3459 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2769 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2758 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6030 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6030/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_6041 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6041/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6052 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6052/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6063 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6063/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_6074 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6074/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6085 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6085/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_5340 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5351 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6096 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6096/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_5362 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5373 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5384 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5395 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4650 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4661 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4672 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_4683 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4694 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3960 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3971 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_3982 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3993 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_3/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_1309 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9606 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_9617 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9628 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9639 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_8927 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8916 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8905 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_8949 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8938 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3223 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3212 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_3201 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2522 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_2511 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2500 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_3256 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3245 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3234 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1810 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2555 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_2544 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2533 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3289 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3278 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_3267 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1843 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_1832 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1821 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2588 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_2577 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2566 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1887 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_1876 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1865 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1854 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2599 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1898 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_5170 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5181 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5192 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_4480 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4491 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3790 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_1106 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_1139 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1128 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1117 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9414 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_9403 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_8702 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9447 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_9436 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9425 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8735 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8724 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8713 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9469 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9458 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8779 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_8768 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_8757 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8746 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3031 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3031/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3020 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3020/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2330 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3075 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3075/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3064 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3064/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3053 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3053/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_3042 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3042/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_2363 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2352 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2341 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3097 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3097/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_3086 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3086/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_1651 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1640 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_2396 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2385 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_2374 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1695 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1684 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1673 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1662 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9970 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9981 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9992 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_8009 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8009/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7308 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7319 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_6607 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6618 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6629 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_5906 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_5917 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5928 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5939 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_9222 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9211 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9200 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8510 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9255 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9244 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9233 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8554 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8543 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8532 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8521 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9288 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9277 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9266 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8587 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8576 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8565 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_9299 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_7820 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7831 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_7842 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8598 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_7853 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7864 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7875 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_7886 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7897 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2171 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2160 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_1470 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2193 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_2182 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1492 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1481 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_529 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_518 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_507 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7105 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7116 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7127 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7138 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7149 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6404 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_6415 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6426 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6437 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6448 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6459 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_5703 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5714 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5725 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5736 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5747 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_5758 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5769 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9030 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9030/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9063 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9063/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9052 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9052/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_9041 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9041/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9096 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9096/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9085 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9085/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_9074 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9074/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_8340 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_8351 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8362 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8373 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8384 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8395 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_7650 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7661 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7672 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7683 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7694 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_30 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_30/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_6960 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6971 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6982 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_63 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_63/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_52 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_52/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_41 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_41/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6993 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_96 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_96/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_85 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_85/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_74 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_74/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_304 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4309 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_337 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_326 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_315 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_359 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_348 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3619 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3608 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_2929 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_2918 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2907 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6201 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_6212 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_6223 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6234 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6245 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_6256 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6267 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6278 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5500 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5511 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5522 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_5533 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6289 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_5544 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5555 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_5566 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4810 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4821 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_860 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5577 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5588 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5599 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4832 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4843 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4854 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_4865 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_893 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_882 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_871 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4876 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4887 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_4898 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_8170 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8181 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8192 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7480 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7491 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_6790 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_112 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_101 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4106 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4117 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_145 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_134 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_123 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3405 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4128 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_4139 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_189 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_178 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_167 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_156 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_2704 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_3449 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3438 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3427 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_3416 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2737 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_2726 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2715 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2759 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2748 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6020 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6020/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_6031 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6031/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6042 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6042/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6053 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6053/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6064 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6064/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6075 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6075/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6086 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6086/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5330 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5341 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6097 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6097/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5352 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_5363 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5374 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_5385 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_5396 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4640 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4651 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4662 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_4673 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_690 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_4684 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4695 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3950 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3961 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_3972 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3983 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3994 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_4/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9607 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_9618 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9629 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_8928 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_8917 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8906 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8939 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3224 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3213 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3202 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2512 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2501 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_3257 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3246 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3235 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1800 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2545 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2534 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2523 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3279 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_3268 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_1844 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_1833 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1822 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1811 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2589 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2578 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2567 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_2556 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1877 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_1866 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1855 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1899 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1888 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5160 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5171 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5182 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5193 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_4470 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4481 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_4492 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3791 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3780 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_1129 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1118 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_1107 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_9404 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_8703 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9437 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9426 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9415 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8736 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8725 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8714 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_9459 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9448 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8769 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_8758 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8747 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3032 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3032/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3021 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3021/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_3010 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3010/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2320 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_3065 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3065/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3054 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3054/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_3043 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3043/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2364 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_2353 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2342 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_2331 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3098 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3098/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3087 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3087/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_3076 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3076/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1652 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_1641 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1630 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_2397 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2386 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2375 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1685 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1674 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1663 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_1696 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9960 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9971 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9982 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9993 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_7309 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6608 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6619 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5907 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5918 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5929 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_9212 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9201 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_8511 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8500 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9256 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_9245 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9234 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_9223 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8544 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8533 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8522 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9289 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9278 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9267 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8577 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8566 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8555 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_7810 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7821 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7832 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_7843 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8599 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_8588 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7854 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7865 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_7876 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7887 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7898 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2172 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2161 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2150 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_1460 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2194 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2183 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1493 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1482 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1471 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9790 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_519 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_508 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7106 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7117 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7128 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7139 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6405 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6416 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6427 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_6438 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6449 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_5704 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5715 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5726 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5737 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5748 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_5759 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9031 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9031/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9020 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9020/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9064 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9064/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9053 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9053/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9042 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9042/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_9097 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9097/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9086 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9086/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9075 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9075/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8330 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_8341 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8352 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8363 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8374 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_8385 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8396 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_7640 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_7651 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_7662 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7673 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7684 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_20 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_20/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7695 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_6950 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6961 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6972 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_64 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_64/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_53 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_53/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_42 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_42/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_31 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_31/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6983 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6994 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_97 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_97/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_86 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_86/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_75 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_75/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1290 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_338 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_327 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_316 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_305 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_349 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3609 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2919 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_2908 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6202 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_6213 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6224 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6235 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_6246 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6257 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6268 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5501 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5512 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5523 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6279 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5534 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_5545 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5556 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_5567 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4800 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4811 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4822 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_850 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5578 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5589 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4833 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4844 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4855 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_894 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_883 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_872 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_861 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4866 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4877 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_4888 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_4899 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_8160 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_8171 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8182 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_8193 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_7470 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7481 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7492 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6780 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6791 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_113 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_102 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4107 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_146 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_135 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_124 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3406 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4118 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_4129 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_179 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_168 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_157 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3439 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3428 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3417 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2738 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_2727 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2716 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2705 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_2749 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6010 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6010/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_6021 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6021/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_6032 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6032/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6043 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6043/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6054 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6054/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_6065 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6065/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6076 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6076/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_5320 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5331 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6087 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6087/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_6098 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6098/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_5342 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_5353 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5364 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_5375 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4630 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5386 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5397 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4641 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4652 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4663 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_691 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_680 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4674 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_4685 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4696 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_3940 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3951 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3962 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_3973 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3984 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3995 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_5 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_5/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9608 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_9619 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_8918 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_8907 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8929 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3214 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3203 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2513 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_2502 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_3247 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3236 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_3225 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1801 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2546 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_2535 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2524 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3269 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_3258 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1834 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1823 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1812 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2579 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2568 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2557 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1878 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_1867 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1856 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1845 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_1889 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_5150 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5161 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5172 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5183 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5194 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4460 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4471 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_3770 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4482 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_4493 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3792 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3781 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_1119 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1108 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_9405 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9438 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_9427 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9416 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8726 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8715 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8704 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9449 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8759 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8748 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8737 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3022 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3022/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3011 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3011/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_3000 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3000/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2321 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2310 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_3066 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3066/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3055 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3055/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3044 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3044/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_3033 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3033/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_2354 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2343 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2332 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3099 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3099/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3088 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3088/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3077 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3077/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_1642 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1631 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1620 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2387 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2376 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_2365 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1686 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_1675 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1664 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1653 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2398 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1697 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9950 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9961 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_9972 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9983 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_9994 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4290 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_6609 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5908 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5919 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9213 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9202 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_8501 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9246 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9235 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9224 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8545 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8534 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8523 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8512 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9279 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9268 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9257 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_7800 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8578 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8567 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8556 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_7811 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7822 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_7833 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8589 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_7844 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7855 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_7866 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_7877 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7888 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7899 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2162 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2151 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_2140 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_1461 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_1450 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_2195 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2184 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_2173 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1494 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1483 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1472 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9780 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_9791 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_509 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7107 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7118 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7129 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_6406 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6417 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6428 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6439 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_5705 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5716 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5727 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5738 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_5749 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_9021 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9021/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9010 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9010/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9054 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9054/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9043 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9043/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9032 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9032/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_9098 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9098/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9087 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9087/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9076 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9076/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_9065 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9065/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8320 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_8331 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_8342 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8353 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8364 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_8375 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8386 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7630 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7641 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8397 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_7652 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_7663 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7674 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7685 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6940 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_21 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_21/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_10 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_10/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7696 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_6951 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6962 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6973 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_54 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_54/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_43 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_43/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_32 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_32/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6984 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6995 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_87 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_87/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_76 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_76/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_65 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_65/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_98 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_98/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1291 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1280 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_328 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_317 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_306 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_339 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2909 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6203 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_6214 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6225 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6236 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_6247 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6258 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6269 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_5502 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5513 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_5524 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_5535 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5546 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_5557 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4801 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4812 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_851 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_840 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5568 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5579 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4823 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4834 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4845 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_4856 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_884 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_873 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_862 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_4867 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4878 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_4889 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_895 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8150 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_8161 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8172 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8183 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_8194 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_7460 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7471 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7482 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7493 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_6770 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6781 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_6792 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_103 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4108 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_136 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_125 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_114 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4119 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_169 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_158 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_147 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3429 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3418 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_3407 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_2728 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_2717 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2706 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2739 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6000 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6000/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6011 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6011/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_6022 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6022/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6033 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6033/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6044 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6044/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_6055 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6055/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6066 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6066/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6077 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6077/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5310 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5321 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5332 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6088 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6088/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_6099 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6099/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_5343 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_5354 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5365 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4620 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5376 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_5387 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5398 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4631 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_4642 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4653 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4664 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_692 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_681 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_670 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4675 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4686 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_4697 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_3930 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3941 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3952 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_3963 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_3974 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3985 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3996 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_6 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_6/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7290 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9609 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8919 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_8908 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_3215 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_3204 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2503 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_3248 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3237 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3226 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2536 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2525 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2514 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3259 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1835 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1824 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1813 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1802 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2569 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2558 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_2547 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1868 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_1857 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1846 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1879 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5140 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5151 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_5162 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5173 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5184 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5195 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4450 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4461 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4472 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3760 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4483 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4494 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3793 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3782 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3771 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_1109 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9428 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9417 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9406 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8727 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8716 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8705 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9439 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_8749 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8738 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3023 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3023/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3012 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3012/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_3001 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3001/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2311 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2300 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_3056 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3056/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3045 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3045/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3034 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3034/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1610 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2355 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_2344 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2333 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_2322 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3089 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3089/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3078 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3078/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_3067 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3067/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1643 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_1632 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1621 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2388 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_2377 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2366 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1676 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1665 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1654 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2399 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1698 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1687 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9940 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9951 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_9962 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9973 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9984 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_9995 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4280 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4291 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3590 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5909 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9203 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_8502 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9247 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_9236 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9225 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_9214 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8535 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8524 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8513 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9269 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9258 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8568 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_8557 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8546 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_7801 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7812 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7823 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_7834 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8579 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_7845 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7856 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_7867 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7878 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7889 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2163 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2152 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2141 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_2130 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_1451 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1440 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_2196 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2185 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_2174 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1484 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1473 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1462 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_1495 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9770 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9781 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9792 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7108 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7119 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_6407 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6418 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6429 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_5706 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_5717 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5728 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5739 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_9022 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9022/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9011 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9011/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9000 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9000/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9055 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9055/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9044 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9044/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9033 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9033/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8310 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9088 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9088/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9077 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9077/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9066 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9066/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8321 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_8332 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8343 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9099 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9099/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_8354 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8365 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8376 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8387 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7620 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7631 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_7642 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8398 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_7653 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7664 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7675 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6930 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_11 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_11/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7686 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7697 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_6941 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6952 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6963 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_55 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_55/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_44 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_44/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_33 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_33/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_22 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_22/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6974 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6985 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6996 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_88 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_88/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_77 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_77/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_66 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_66/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_99 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_99/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1292 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1281 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_1270 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_329 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_318 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_307 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6204 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_6215 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6226 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6237 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6248 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6259 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_5503 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5514 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5525 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5536 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5547 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_5558 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4802 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4813 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_841 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_830 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5569 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4824 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4835 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_4846 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_885 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_874 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_863 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_852 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4857 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4868 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_4879 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_896 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8140 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_8151 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8162 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8173 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8184 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8195 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_7450 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7461 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7472 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7483 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7494 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_6760 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6771 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6782 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6793 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_104 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_137 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_126 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_115 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4109 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_159 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_148 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3419 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3408 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_2729 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_2718 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2707 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6001 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6001/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_6012 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6012/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_6023 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6023/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6034 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6034/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6045 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6045/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_6056 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6056/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6067 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6067/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5300 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5311 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5322 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6078 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6078/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_6089 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6089/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_5333 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_5344 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5355 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_5366 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4610 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4621 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5377 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5388 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5399 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4632 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4643 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4654 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_693 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_682 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_671 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_660 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4665 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4676 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4687 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_4698 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3920 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_3931 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3942 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3953 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_3964 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3975 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3986 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_3997 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_7 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_7/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7280 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7291 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_6590 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_8909 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_3205 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_3238 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3227 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_3216 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2537 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_2526 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2515 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2504 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_3249 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1825 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1814 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1803 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2559 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2548 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1869 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_1858 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1847 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1836 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5130 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5141 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_5152 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_5163 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5174 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_5185 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_5196 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4440 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4451 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4462 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_490 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_3761 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_3750 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4473 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_4484 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4495 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3794 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3783 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3772 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xmarker_pixel_0 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 marker_pixel_0/AMP_IN
+ SF_IB pixel_900/PIX_OUT CSA_VREF marker_pixel
Xpixel_9429 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_9418 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9407 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8717 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8706 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8739 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_8728 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3013 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3013/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3002 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3002/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2312 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2301 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_3057 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3057/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3046 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3046/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3035 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3035/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_3024 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3024/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1600 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2345 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2334 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2323 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3079 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3079/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_3068 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3068/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_1633 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1622 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1611 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2378 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2367 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_2356 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1677 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_1666 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1655 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1644 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2389 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1699 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1688 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9941 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9930 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9952 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_9963 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9974 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_9985 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_9996 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4270 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4281 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_4292 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3591 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3580 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2890 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9204 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9237 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9226 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9215 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8536 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8525 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8514 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8503 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9259 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9248 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8569 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_8558 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8547 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_7802 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7813 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_7824 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_7835 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7846 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_7857 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_7868 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7879 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2120 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2153 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2142 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_2131 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1452 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_1441 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1430 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_2197 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2186 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2175 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_2164 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1485 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1474 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1463 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_1496 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9760 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9771 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9782 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9793 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_7109 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6408 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6419 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5707 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5718 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5729 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_9012 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9012/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9001 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9001/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9045 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9045/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9034 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9034/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_9023 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9023/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8300 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9089 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9089/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9078 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9078/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9067 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9067/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_9056 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9056/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8311 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8322 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_8333 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8344 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8355 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_8366 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8377 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7610 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7621 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7632 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8388 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_8399 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_7643 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_7654 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7665 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_7676 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6920 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_6931 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_12 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_12/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7687 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7698 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_6942 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6953 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6964 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_45 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_45/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_34 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_34/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_23 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_23/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6975 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6986 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_6997 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_78 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_78/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_67 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_67/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_56 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_56/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_89 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_89/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1260 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_1293 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1282 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1271 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9590 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_319 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_308 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6205 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6216 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6227 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_6238 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6249 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_5504 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5515 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5526 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5537 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5548 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4803 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_842 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_831 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_820 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5559 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4814 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4825 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_4836 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_4847 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_875 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_864 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_853 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4858 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4869 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_897 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_886 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8130 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_8141 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8152 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8163 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8174 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_8185 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7440 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_8196 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_7451 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_7462 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7473 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7484 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_7495 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_6750 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6761 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6772 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_6783 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6794 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1090 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1090/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_127 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_116 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_105 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_149 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_138 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3409 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2719 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_2708 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6002 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6002/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_6013 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6013/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6024 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6024/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6035 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6035/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_6046 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6046/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6057 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6057/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6068 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6068/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5301 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5312 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5323 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6079 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6079/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5334 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_5345 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5356 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4600 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4611 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_650 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5367 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5378 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5389 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4622 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_4633 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4644 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4655 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3910 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_683 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_672 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_661 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4666 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4677 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_4688 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3921 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_3932 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3943 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_694 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4699 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3954 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_3965 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3976 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3987 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_3998 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_8 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_8/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7270 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7281 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7292 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6580 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6591 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_5890 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_3206 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_3239 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3228 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3217 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2527 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2516 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2505 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1826 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_1815 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1804 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2549 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2538 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1859 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1848 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1837 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5120 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5131 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5142 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_5153 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5164 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_4430 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5175 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_5186 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5197 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4441 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4452 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4463 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_491 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_480 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_3751 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3740 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4474 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_4485 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4496 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_3795 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3784 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3773 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3762 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xmarker_pixel_1 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 marker_pixel_1/AMP_IN
+ SF_IB pixel_901/PIX_OUT CSA_VREF marker_pixel
Xpixel_9419 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9408 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8718 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_8707 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8729 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3014 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3014/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3003 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3003/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2302 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_3047 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3047/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3036 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3036/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_3025 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3025/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1601 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2335 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2324 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_2313 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3069 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3069/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_3058 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3058/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1634 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1623 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1612 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2379 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2368 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2357 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_2346 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1667 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1656 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1645 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_1689 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1678 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9942 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_9931 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9920 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9953 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9964 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9975 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_9986 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9997 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4260 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4271 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_3570 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4282 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_4293 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3592 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3581 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2891 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2880 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_9238 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_9227 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9216 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9205 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_8526 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8515 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8504 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9249 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8559 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8548 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8537 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7803 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7814 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7825 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7836 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7847 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_7858 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7869 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2110 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2154 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2143 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2132 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_2121 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_1442 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1431 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1420 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2187 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2176 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_2165 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1475 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1464 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1453 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2198 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1497 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_1486 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9750 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9761 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_9772 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9783 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_9794 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4090 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4090/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_6409 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5708 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5719 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9013 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9013/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9002 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9002/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9046 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9046/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9035 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9035/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9024 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9024/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8301 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9079 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9079/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9068 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9068/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9057 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9057/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8312 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_8323 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8334 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8345 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8356 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8367 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8378 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7600 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_7611 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7622 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_7633 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8389 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_7644 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7655 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_7666 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6910 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_6921 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7677 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7688 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7699 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_6932 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6943 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6954 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_46 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_46/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_35 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_35/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_24 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_24/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_13 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_13/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6965 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6976 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6987 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_6998 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_79 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_79/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_68 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_68/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_57 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_57/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1250 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_1294 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1283 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1272 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_1261 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_9591 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_9580 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8890 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_309 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6206 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6217 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6228 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6239 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_5505 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5516 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5527 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5538 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_5549 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4804 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_832 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_821 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_810 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4815 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4826 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_4837 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_876 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_865 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_854 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_843 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4848 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4859 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_898 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_887 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8120 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_8131 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_8142 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8153 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8164 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_8175 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8186 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7430 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7441 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8197 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_7452 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_7463 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7474 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7485 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7496 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_6740 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_6751 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6762 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6773 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_6784 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6795 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1091 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1091/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1080 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1080/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_128 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_117 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_106 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_139 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2709 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6003 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6003/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_6014 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6014/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6025 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6025/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6036 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6036/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_6047 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6047/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6058 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6058/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5302 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5313 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6069 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6069/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_5324 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_5335 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5346 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_5357 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4601 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4612 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_640 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5368 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5379 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4623 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4634 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4645 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3900 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_684 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_673 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_662 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_651 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4656 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4667 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4678 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_4689 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3911 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_3922 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3933 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3944 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_695 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3955 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3966 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3977 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_3988 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3999 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_9 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_9/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7260 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7271 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7282 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7293 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_6570 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6581 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_6592 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5880 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5891 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3229 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3218 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_3207 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_2528 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_2517 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2506 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_1816 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_1805 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_2539 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1849 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1838 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1827 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5110 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5121 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5132 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_5143 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_5154 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5165 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4420 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5176 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_5187 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5198 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4431 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_4442 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4453 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_492 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_481 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_470 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_3752 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_3741 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3730 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4464 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_4475 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4486 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_4497 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_3785 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3774 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3763 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_3796 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_7090 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7090/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9409 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8708 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8719 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3004 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3004/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2303 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_3048 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3048/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3037 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3037/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3026 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3026/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_3015 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3015/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2336 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2325 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2314 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3059 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3059/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1624 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1613 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1602 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2369 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2358 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_2347 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1668 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_1657 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1646 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1635 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1679 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9932 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_9921 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9910 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9943 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9954 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9965 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_9976 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_9987 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9998 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4250 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4261 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4272 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3560 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4283 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4294 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3593 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3582 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3571 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2892 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_2881 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2870 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9228 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9217 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9206 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8527 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8516 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8505 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9239 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_8549 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8538 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7804 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7815 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7826 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7837 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7848 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_7859 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2111 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2100 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2144 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2133 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_2122 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1443 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_1432 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1421 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_1410 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2177 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2166 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_2155 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1476 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1465 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1454 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2199 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2188 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_1498 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1487 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9740 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9751 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_9762 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9773 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9784 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_9795 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4080 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4080/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4091 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4091/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3390 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5709 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9003 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9003/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9036 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9036/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9025 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9025/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_9014 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9014/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_9069 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9069/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9058 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9058/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_9047 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9047/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_8302 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_8313 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_8324 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8335 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8346 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_8357 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8368 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7601 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7612 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7623 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8379 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_7634 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_7645 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7656 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6900 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6911 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_6922 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_7667 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7678 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7689 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_6933 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6944 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_6955 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_36 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_36/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_25 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_25/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_14 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_14/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6966 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6977 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_6988 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_69 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_69/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_58 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_58/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_47 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_47/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6999 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1251 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1240 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_1284 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1273 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1262 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_1295 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9592 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_9581 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9570 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8891 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_8880 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6207 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6218 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6229 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_5506 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_5517 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5528 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5539 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_833 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_822 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_811 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_800 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4805 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4816 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_4827 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_4838 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_866 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_855 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_844 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4849 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_899 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_888 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_877 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8110 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_8121 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_8132 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8143 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8154 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8165 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8176 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7420 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7431 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_8187 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8198 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_7442 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_7453 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7464 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7475 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6730 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7486 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7497 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_6741 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6752 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6763 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_6774 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6785 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6796 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_1092 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1092/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1081 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1081/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_1070 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1070/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_118 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_107 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_129 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_6004 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6004/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_6015 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6015/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6026 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6026/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6037 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6037/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6048 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6048/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6059 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6059/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_5303 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5314 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5325 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5336 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5347 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4602 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_641 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_630 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5358 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5369 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4613 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_4624 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4635 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_4646 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3901 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_674 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_663 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_652 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4657 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4668 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_4679 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_3912 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_3923 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3934 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_696 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_685 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3945 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3956 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3967 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3978 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_3989 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_7250 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7261 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7272 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7283 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7294 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_6560 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6571 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6582 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6593 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5870 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5881 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5892 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3219 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3208 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_2518 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2507 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1817 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_1806 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2529 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1839 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1828 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5100 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5111 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5122 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_5133 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_5144 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5155 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_4410 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4421 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5166 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_5177 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5188 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5199 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4432 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4443 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4454 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_482 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_471 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_460 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3742 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3731 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3720 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4465 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4476 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4487 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_493 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3786 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_3775 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3764 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3753 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4498 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3797 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_7080 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7080/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7091 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7091/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_6390 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_8709 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_3005 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3005/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_3038 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3038/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3027 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3027/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_3016 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3016/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2326 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2315 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2304 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_3049 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3049/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1625 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1614 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1603 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2359 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2348 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_2337 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1658 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1647 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1636 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_1669 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9900 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9933 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_9922 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9911 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9944 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9955 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9966 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_9977 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9988 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9999 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4240 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4251 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4262 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_290 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_3561 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_3550 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4273 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_4284 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4295 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3594 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3583 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3572 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2882 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_2871 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2860 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2893 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_9229 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_9218 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9207 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8517 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8506 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8539 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_8528 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7805 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7816 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7827 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7838 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7849 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2101 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_1400 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2145 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2134 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2123 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_2112 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_1433 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1422 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1411 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2178 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2167 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_2156 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1466 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1455 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1444 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2189 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1499 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1488 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_1477 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9730 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9741 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9752 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_9763 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9774 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_9785 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_9796 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4070 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4070/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4081 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4081/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_4092 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4092/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3391 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3380 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2690 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9004 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9004/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9037 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9037/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9026 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9026/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9015 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9015/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_9059 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9059/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9048 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9048/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8303 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_8314 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8325 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8336 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8347 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_8358 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8369 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_7602 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7613 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_7624 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_7635 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7646 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_7657 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6901 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_6912 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7668 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7679 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_6923 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6934 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6945 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_37 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_37/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_26 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_26/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_15 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_15/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6956 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6967 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6978 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_6989 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_59 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_59/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_48 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_48/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1241 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1230 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_1285 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1274 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1263 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_1252 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_1296 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9593 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_9582 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9571 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9560 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_8881 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8870 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8892 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6208 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6219 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5507 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5518 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5529 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_823 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_812 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_801 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4806 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4817 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_4828 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_856 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_845 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_834 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4839 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_889 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_878 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_867 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8100 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8111 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8122 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_8133 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8144 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8155 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_8166 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8177 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7410 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7421 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7432 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8188 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_8199 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_7443 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_7454 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7465 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6720 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7476 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7487 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7498 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_6731 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6742 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6753 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6764 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6775 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6786 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_6797 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_1060 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1060/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_1093 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1093/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1082 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1082/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1071 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1071/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9390 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_119 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_108 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6005 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6005/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6016 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6016/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6027 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6027/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_6038 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6038/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6049 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6049/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_5304 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5315 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5326 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5337 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5348 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4603 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_631 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_620 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5359 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4614 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4625 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_4636 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_675 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_664 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_653 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_642 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4647 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4658 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4669 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_3902 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_3913 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3924 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3935 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_697 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_686 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_3946 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3957 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3968 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_3979 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_7240 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_7251 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_7262 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7273 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7284 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_7295 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_6550 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6561 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6572 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_6583 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6594 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_5860 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5871 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5882 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5893 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3209 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2519 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_2508 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_1807 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1829 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1818 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5101 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5112 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5123 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_5134 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_5145 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5156 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4400 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4411 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_450 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3710 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5167 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5178 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5189 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4422 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_4433 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4444 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_483 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_472 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_461 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_3743 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_3732 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3721 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_4455 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_4466 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4477 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_4488 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_494 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3776 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3765 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3754 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_4499 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3798 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3787 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7070 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7070/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7081 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7081/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7092 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7092/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6380 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6391 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_5690 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_3039 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3039/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3028 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3028/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3017 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3017/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_3006 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3006/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2327 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2316 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2305 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1615 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1604 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2349 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2338 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1659 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1648 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1637 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1626 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9923 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_9912 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9901 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9945 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9934 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_9956 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_9967 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_9978 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9989 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4230 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4241 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4252 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4263 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_291 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_280 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_3551 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3540 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4274 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_4285 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4296 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2850 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3584 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3573 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3562 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2883 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_2872 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2861 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_3595 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2894 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_9219 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9208 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8518 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_8507 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8529 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_7806 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7817 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7828 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7839 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2102 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2135 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2124 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_2113 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1434 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1423 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1412 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_1401 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2168 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2157 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_2146 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1467 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1456 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1445 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2179 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1489 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1478 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9720 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9731 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9742 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_9753 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9764 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9775 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_9786 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9797 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4060 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4060/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4071 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4071/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4082 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4082/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_4093 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4093/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3392 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3381 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_3370 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2691 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2680 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_1990 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9027 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9027/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9016 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9016/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9005 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9005/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9049 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9049/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_9038 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9038/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_8304 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_8315 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8326 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8337 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_8348 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8359 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_7603 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7614 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7625 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7636 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7647 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6902 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_6913 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_7658 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7669 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_6924 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6935 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_6946 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_27 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_27/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_16 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_16/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6957 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6968 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_6979 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_49 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_49/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_38 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_38/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1242 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1231 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1220 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_1275 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1264 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1253 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_1297 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_1286 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9550 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9583 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_9572 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9561 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8882 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_8871 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8860 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9594 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8893 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_6209 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5508 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5519 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_824 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_813 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_802 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4807 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4818 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_857 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_846 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_835 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_4829 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_879 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_868 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_8101 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_8112 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_8123 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8134 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8145 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8156 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8167 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7400 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_7411 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7422 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_8178 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8189 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_7433 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_7444 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7455 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_7466 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6710 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_6721 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7477 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7488 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7499 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_6732 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6743 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6754 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_6765 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6776 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6787 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_6798 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1050 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1050/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_1083 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1083/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1072 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1072/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_1061 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1061/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_1094 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1094/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_9391 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_9380 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8690 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_109 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6006 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6006/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6017 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6017/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6028 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6028/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6039 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6039/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_5305 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5316 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5327 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5338 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_632 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_621 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_610 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5349 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4604 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4615 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4626 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_4637 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_665 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_654 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_643 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4648 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4659 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_3903 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_3914 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3925 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_698 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_687 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_676 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3936 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_3947 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3958 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3969 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_7230 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7241 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_7252 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_7263 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7274 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7285 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7296 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_6540 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_6551 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6562 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6573 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_6584 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6595 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_5850 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5861 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5872 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5883 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5894 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2509 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1808 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_1819 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5102 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5113 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_5124 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_5135 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5146 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_4401 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4412 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_440 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3700 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5157 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_5168 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5179 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4423 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4434 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4445 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_473 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_462 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_451 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3733 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3722 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3711 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4456 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4467 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4478 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_495 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_484 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3777 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_3766 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3755 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3744 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4489 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3799 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3788 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7060 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7060/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7071 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7071/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7082 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7082/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7093 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7093/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_6370 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6381 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_6392 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5680 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5691 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_4990 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_3029 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3029/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3018 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3018/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_3007 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3007/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_2317 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2306 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_1616 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_1605 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_2339 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2328 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1649 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1638 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1627 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9924 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_9913 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9902 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9946 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9935 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9957 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_9968 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9979 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4220 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4231 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_4242 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4253 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_292 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_281 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_270 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_3552 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_3541 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3530 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4264 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_4275 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4286 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2840 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3585 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3574 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3563 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_4297 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2873 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_2862 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2851 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3596 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2895 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2884 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_9209 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8508 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8519 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_7807 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7818 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7829 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_2136 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2125 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2114 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_2103 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_1424 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1413 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1402 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2169 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2158 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_2147 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1457 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1446 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1435 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1479 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1468 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9710 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9721 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9732 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_9743 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9754 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9765 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_9776 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_9787 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9798 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4050 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4050/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4061 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4061/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_3360 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4072 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4072/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_4083 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4083/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4094 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4094/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3393 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3382 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3371 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2692 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_2681 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2670 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_1980 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_1991 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_9028 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9028/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9017 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9017/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9006 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9006/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_9039 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9039/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_8305 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_8316 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8327 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8338 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_8349 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_7604 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7615 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7626 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7637 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7648 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6903 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7659 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_6914 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6925 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6936 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_28 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_28/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_17 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_17/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6947 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6958 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6969 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_39 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_39/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1232 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1221 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_1210 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_1276 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1265 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1254 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_1243 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_1298 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1287 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9540 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9584 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_9573 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9562 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9551 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8872 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8861 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8850 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9595 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8894 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8883 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3190 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5509 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_814 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_803 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4808 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_4819 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_847 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_836 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_825 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_869 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_858 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8102 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_8113 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_8124 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8135 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8146 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_8157 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8168 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7401 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7412 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7423 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8179 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_7434 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_7445 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7456 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6700 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6711 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7467 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7478 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7489 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_6722 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6733 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6744 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_6755 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6766 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6777 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_6788 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_6799 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1051 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1051/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1040 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1040/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_1084 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1084/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1073 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1073/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1062 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1062/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_1095 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1095/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9392 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_9381 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9370 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8680 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8691 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_7990 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_6007 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6007/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6018 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6018/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6029 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6029/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_5306 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_5317 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5328 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5339 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_622 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_611 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_600 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4605 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4616 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_4627 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_666 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_655 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_644 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_633 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4638 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_4649 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3904 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_3915 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_3926 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_699 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_688 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_677 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_3937 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3948 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3959 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_7220 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7231 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_7242 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_7253 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7264 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6530 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7275 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_7286 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7297 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_6541 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6552 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6563 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_6574 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6585 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6596 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_5840 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5851 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_5862 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5873 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5884 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5895 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1809 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5103 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5114 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5125 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5136 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5147 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4402 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_441 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_430 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3701 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5158 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5169 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4413 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_4424 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4435 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_474 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_463 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_452 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_3734 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_3723 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3712 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_4446 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_4457 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4468 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_4479 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_496 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_485 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3767 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3756 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3745 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3789 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3778 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7050 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7050/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7061 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7061/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7072 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7072/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7083 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7083/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7094 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7094/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_6360 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6371 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6382 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6393 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5670 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5681 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5692 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_4980 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4991 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3019 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3019/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3008 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3008/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_2318 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2307 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1606 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2329 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1639 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1628 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1617 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9914 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_9903 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9947 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_9936 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9925 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_9958 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_9969 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4210 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4221 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_4232 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4243 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4254 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_282 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_271 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_260 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3542 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3531 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3520 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4265 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4276 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4287 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_293 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_2841 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_2830 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3575 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3564 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3553 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4298 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2874 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_2863 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2852 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_3597 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_3586 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2896 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2885 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6190 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_8509 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7808 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7819 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_2126 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2115 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2104 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_1425 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1414 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1403 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2159 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2148 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_2137 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1458 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1447 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1436 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_1469 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9700 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9711 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9722 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9733 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_9744 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9755 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9766 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_9777 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9788 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9799 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4040 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4040/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4051 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4051/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4062 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4062/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_3350 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4073 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4073/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_4084 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4084/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4095 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4095/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3394 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3383 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3372 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3361 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2682 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_2671 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2660 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_1970 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2693 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1992 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1981 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9018 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9018/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9007 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9007/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_9029 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9029/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_8306 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8317 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8328 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_8339 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_7605 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7616 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7627 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7638 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6904 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7649 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6915 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6926 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6937 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_18 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_18/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6948 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6959 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_29 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_29/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1200 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_1233 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1222 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1211 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_1266 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1255 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1244 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_1299 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1288 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_1277 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9541 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9530 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9574 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_9563 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9552 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8873 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8862 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8851 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8840 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9596 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9585 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8895 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8884 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3191 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3180 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2490 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_815 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_804 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4809 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_848 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_837 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_826 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_859 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8103 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_8114 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8125 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8136 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8147 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_8158 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7402 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7413 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_8169 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_7424 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_7435 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7446 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_7457 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6701 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_6712 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7468 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7479 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_6723 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6734 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6745 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_6756 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6767 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6778 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_6789 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1041 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1041/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1030 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1030/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_1074 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1074/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1063 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1063/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_1052 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1052/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_1096 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1096/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_1085 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1085/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_9382 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9371 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9360 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_8681 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8670 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9393 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_8692 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7980 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7991 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_6008 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6008/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6019 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6019/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5307 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5318 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5329 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_623 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_612 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_601 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4606 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4617 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_4628 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_656 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_645 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_634 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4639 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3905 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_3916 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_689 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_678 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_667 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3927 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_3938 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3949 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_7210 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7221 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7232 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_7243 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_7254 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7265 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6520 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7276 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7287 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7298 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_6531 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6542 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6553 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6564 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6575 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6586 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_6597 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5830 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5841 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_5852 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_5863 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5874 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_5885 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_5896 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9190 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5104 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5115 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5126 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5137 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_4403 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_431 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_420 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5148 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_5159 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4414 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4425 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_4436 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_464 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_453 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_442 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3724 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3713 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3702 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4447 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4458 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4469 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_497 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_486 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_475 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3768 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_3757 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3746 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3735 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_3779 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_7040 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7040/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_7051 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7051/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_7062 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7062/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7073 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7073/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7084 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7084/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_7095 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7095/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_6350 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6361 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6372 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_6383 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6394 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_5660 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5671 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5682 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5693 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_4970 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4981 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_4992 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3009 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3009/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2308 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_1607 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_2319 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1629 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1618 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9915 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_9904 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9937 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9926 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9948 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_9959 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4200 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4211 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4222 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_4233 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4244 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_283 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_272 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_261 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_250 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3543 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_3532 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3521 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_3510 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4255 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_4266 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4277 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_294 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2831 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_2820 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_3576 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3565 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3554 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_4288 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_4299 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2864 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_2853 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2842 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3598 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3587 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2897 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2886 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2875 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6180 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6191 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_5490 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_7809 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2127 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2116 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2105 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1415 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1404 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2149 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2138 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1448 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1437 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1426 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_1459 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9701 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9712 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9723 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_9734 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_9745 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9756 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_9767 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_9778 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9789 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4030 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4030/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4041 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4041/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4052 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4052/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_3351 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3340 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4063 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4063/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_4074 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4074/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_4085 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4085/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4096 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4096/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_3384 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3373 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3362 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2672 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2661 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2650 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3395 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1971 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_1960 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2694 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2683 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1993 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1982 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9019 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9019/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9008 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9008/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8307 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8318 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_8329 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_7606 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7617 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7628 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7639 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6905 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6916 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6927 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_19 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_19/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_6938 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6949 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1223 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1212 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_1201 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_1267 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1256 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1245 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_1234 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1289 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1278 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9531 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9520 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_8830 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9575 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_9564 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9553 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9542 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8863 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8852 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8841 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9597 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9586 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8896 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8885 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8874 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3192 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3181 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_3170 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2491 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2480 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_1790 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_805 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_838 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_827 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_816 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_849 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8104 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_8115 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8126 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8137 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_8148 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8159 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_7403 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7414 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7425 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7436 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7447 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6702 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7458 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7469 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_6713 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6724 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6735 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_6746 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6757 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6768 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_6779 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1042 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1042/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1031 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1031/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1020 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1020/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_1075 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1075/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1064 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1064/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1053 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1053/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_1097 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1097/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_1086 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1086/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9350 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9383 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_9372 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9361 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8671 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8660 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9394 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8693 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_8682 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7970 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7981 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7992 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6009 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6009/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5308 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5319 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_613 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_602 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4607 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4618 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_657 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_646 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_635 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_624 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4629 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3906 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_3917 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_679 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_668 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_3928 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3939 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_7200 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_7211 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7222 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_7233 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_7244 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7255 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6510 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_6521 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7266 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_7277 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7288 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7299 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_6532 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6543 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6554 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_6565 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6576 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6587 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5820 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5831 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5842 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6598 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_5853 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5864 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_5875 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_5886 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5897 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9191 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_9180 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8490 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5105 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5116 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5127 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5138 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_432 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_421 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_410 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5149 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4404 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4415 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4426 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_465 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_454 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_443 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_3725 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_3714 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3703 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4437 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_4448 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4459 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_498 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_487 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_476 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3758 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3747 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3736 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_3769 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_7030 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7030/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7041 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7041/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_7052 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7052/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_7063 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7063/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7074 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7074/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7085 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7085/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7096 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7096/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_6340 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_6351 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6362 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6373 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_6384 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6395 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_5650 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5661 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5672 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5683 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5694 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4960 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4971 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4982 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_4993 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_2309 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1619 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1608 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_9905 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9938 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_9927 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9916 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9949 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4201 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_240 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3500 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4212 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_4223 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4234 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4245 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_273 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_262 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_251 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3533 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3522 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3511 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4256 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4267 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4278 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_295 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_284 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_2821 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2810 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_3566 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3555 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3544 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4289 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2865 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_2854 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2843 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2832 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3599 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3588 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3577 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2898 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2887 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2876 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6170 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6181 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_6192 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5480 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5491 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_4790 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_2117 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2106 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_1416 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_1405 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_2139 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2128 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1449 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1438 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1427 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9702 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9713 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9724 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_9735 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9746 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9757 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_9768 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9779 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4020 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4020/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4031 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4031/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_4042 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4042/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4053 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4053/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_3341 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3330 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4064 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4064/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_4075 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4075/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4086 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4086/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2640 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3385 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3374 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3363 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_3352 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4097 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4097/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2673 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_2662 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2651 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3396 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_1961 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_1950 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_2695 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2684 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1994 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1983 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1972 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9009 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9009/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8308 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8319 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_7607 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7618 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7629 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_6906 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6917 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6928 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6939 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1224 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1213 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1202 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_1257 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1246 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1235 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1279 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1268 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9532 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_9521 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9510 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_8820 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9565 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_9554 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9543 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8864 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_8853 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8842 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8831 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9598 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9587 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9576 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8897 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_8886 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8875 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3193 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3182 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3171 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_3160 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2481 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2470 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_1780 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2492 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1791 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_806 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_839 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_828 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_817 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8105 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_8116 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8127 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8138 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_8149 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_7404 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7415 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7426 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7437 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7448 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6703 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7459 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_6714 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6725 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6736 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_6747 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6758 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6769 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_1032 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1032/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1021 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1021/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_1010 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1010/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_1065 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1065/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1054 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1054/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_1043 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1043/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_1098 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1098/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1087 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1087/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_1076 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1076/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_9340 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9373 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9362 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9351 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8672 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8661 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8650 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9395 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9384 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8694 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8683 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7960 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7971 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7982 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7993 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5309 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_614 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_603 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4608 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_4619 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_647 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_636 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_625 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_3907 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_669 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_658 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3918 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_3929 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_7201 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7212 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7223 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_7234 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_7245 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7256 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6500 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6511 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7267 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7278 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7289 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_6522 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6533 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6544 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_6555 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6566 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6577 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_6588 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5810 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5821 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5832 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_5843 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6599 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_5854 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5865 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_5876 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_5887 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5898 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9192 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_9181 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9170 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8480 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8491 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_7790 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5106 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_5117 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5128 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_422 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_411 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_400 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5139 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_4405 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4416 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_4427 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_455 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_444 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_433 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3715 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_3704 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4438 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_4449 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_499 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_488 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_477 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_466 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3759 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_3748 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3737 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3726 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7020 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7020/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7031 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7031/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_7042 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7042/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_7053 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7053/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7064 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7064/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7075 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7075/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_7086 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7086/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7097 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7097/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_6330 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_6341 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6352 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6363 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_6374 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6385 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6396 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_5640 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5651 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_5662 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5673 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5684 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5695 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4950 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4961 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4972 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_4983 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4994 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1609 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9906 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_9939 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_9928 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9917 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_4202 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_230 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4213 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_4224 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4235 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_274 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_263 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_252 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_241 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3534 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_3523 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3512 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_3501 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4246 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_4257 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4268 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_296 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_285 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_2822 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_2811 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2800 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_3567 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3556 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3545 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_4279 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2855 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_2844 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2833 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3589 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3578 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2899 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2888 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_2877 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2866 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6160 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6171 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6182 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6193 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5470 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5481 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5492 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_4780 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4791 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2118 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2107 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1406 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2129 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1439 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1428 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1417 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9703 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9714 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_9725 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_9736 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9747 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_9758 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_9769 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4010 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4010/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4021 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4021/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_4032 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4032/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4043 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4043/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_3342 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3331 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3320 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4054 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4054/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_4065 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4065/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4076 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4076/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4087 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4087/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2630 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3375 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3364 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3353 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4098 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4098/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2663 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2652 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2641 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3397 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_3386 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_1962 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_1951 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1940 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_2696 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2685 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_2674 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1995 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1984 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1973 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8309 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7608 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7619 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_6907 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6918 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6929 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1214 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1203 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_1258 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1247 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1236 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_1225 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1269 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9522 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9511 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9500 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8821 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_8810 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9566 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_9555 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9544 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9533 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8854 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8843 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8832 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_9599 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_9588 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9577 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8887 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8876 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8865 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8898 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3150 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3183 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3172 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3161 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2482 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_2471 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2460 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3194 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1770 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2493 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1792 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1781 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_829 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_818 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_807 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8106 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8117 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8128 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_8139 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_7405 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7416 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7427 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7438 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7449 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6704 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_6715 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6726 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6737 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6748 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6759 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1033 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1033/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1022 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1022/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1011 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1011/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_1000 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1000/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_1066 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1066/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1055 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1055/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1044 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1044/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_1099 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1099/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1088 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1088/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_1077 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1077/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9341 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9330 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9374 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_9363 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9352 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8662 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8651 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8640 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9396 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9385 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8695 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8684 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8673 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7950 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7961 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7972 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7983 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7994 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2290 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_604 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4609 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_648 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_637 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_626 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_615 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_3908 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_659 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_3919 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_7202 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7213 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_7224 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_7235 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7246 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6501 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_6512 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7257 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_7268 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7279 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_6523 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6534 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6545 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5800 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6556 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6567 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6578 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5811 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5822 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_5833 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6589 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_5844 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5855 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_5866 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_5877 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5888 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5899 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_9182 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9171 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9160 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9193 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_8470 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8481 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8492 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7780 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7791 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_5107 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5118 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5129 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_423 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_412 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_401 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4406 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4417 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_456 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_445 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_434 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_3716 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_3705 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4428 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_4439 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_489 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_478 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_467 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3749 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3738 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3727 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7010 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7010/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7021 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7021/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7032 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7032/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_7043 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7043/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_7054 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7054/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7065 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7065/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6320 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7076 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7076/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7087 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7087/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7098 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7098/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_6331 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6342 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6353 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6364 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6375 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6386 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5630 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5641 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6397 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5652 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_5663 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5674 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_5685 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4940 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5696 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4951 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4962 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_4973 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_990 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_4984 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4995 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9929 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_9918 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9907 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_231 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_220 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4203 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4214 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4225 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_4236 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_264 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_253 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_242 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3524 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3513 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3502 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4247 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4258 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4269 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_297 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_286 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_275 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_2812 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2801 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_3557 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3546 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3535 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2856 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_2845 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2834 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2823 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3579 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_3568 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2889 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2878 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2867 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6150 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6161 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6172 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_6183 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6194 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_5460 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5471 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5482 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5493 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_4770 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4781 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_4792 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_2108 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_1407 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_2119 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1429 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1418 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9704 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9715 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_9726 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9737 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9748 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_9759 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4000 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4000/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4011 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4011/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4022 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4022/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_4033 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4033/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4044 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4044/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_3332 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3321 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_3310 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4055 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4055/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_4066 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4066/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4077 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4077/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2631 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_2620 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_3376 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3365 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3354 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_3343 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4088 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4088/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_4099 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4099/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2664 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_2653 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2642 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3398 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3387 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_1952 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_1941 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1930 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_2697 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2686 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2675 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1996 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_1985 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1974 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1963 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5290 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_7609 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_7609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6908 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6919 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1215 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1204 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_1248 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1237 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1226 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_1259 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9523 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_9512 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9501 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_8811 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8800 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9556 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_9545 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9534 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8855 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_8844 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8833 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8822 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9589 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9578 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9567 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8888 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_8877 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8866 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8899 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3140 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3184 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3173 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3162 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_3151 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_2472 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2461 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2450 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3195 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1771 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_1760 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2494 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2483 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1793 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1782 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_819 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_808 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8107 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8118 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_8129 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_7406 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7417 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7428 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7439 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6705 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6716 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6727 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_6738 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6749 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1023 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1023/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1012 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1012/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_1001 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1001/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_1056 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1056/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1045 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1045/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_1034 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1034/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1089 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1089/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1078 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1078/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_1067 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1067/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_9331 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9320 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9364 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9353 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9342 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8663 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8652 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8641 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8630 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9397 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9386 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9375 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8696 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8685 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8674 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7940 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_7951 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_7962 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7973 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7984 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_7995 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2280 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2291 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1590 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_605 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_638 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_627 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_616 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_649 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3909 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_3909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7203 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7214 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7225 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7236 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7247 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6502 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7258 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7269 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_6513 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6524 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6535 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_6546 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6557 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6568 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_6579 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5801 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5812 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5823 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_5834 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_5845 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5856 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_5867 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5878 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5889 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9183 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_9172 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9161 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_9150 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9194 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8460 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_8471 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8482 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_8493 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_7770 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7781 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7792 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5108 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5119 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_413 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_402 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4407 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4418 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_446 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_435 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_424 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3706 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4429 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_479 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_468 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_457 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3739 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3728 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3717 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7000 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7000/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_7011 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7011/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7022 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7022/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_7033 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7033/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_7044 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7044/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7055 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7055/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6310 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7066 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7066/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_7077 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7077/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7088 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7088/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_6321 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_6332 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6343 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6354 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7099 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7099/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_6365 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6376 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6387 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5620 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5631 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5642 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6398 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_5653 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5664 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_5675 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4930 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5686 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5697 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4941 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4952 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4963 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_4974 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_991 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_980 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4985 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4996 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8290 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9919 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9908 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_221 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_210 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4204 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4215 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4226 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_265 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_254 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_243 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_232 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3525 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_3514 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3503 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4237 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_4248 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4259 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_298 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_287 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_276 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_2813 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_2802 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_3558 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3547 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3536 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2846 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_2835 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2824 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3569 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2879 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2868 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2857 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6140 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_6151 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6162 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6173 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_6184 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6195 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_5450 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5461 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5472 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5483 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5494 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4760 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4771 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4782 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_4793 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_2109 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_2109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1419 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1408 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_9705 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9716 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9727 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9738 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_9749 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4001 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4001/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4012 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4012/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_4023 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4023/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4034 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4034/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_3333 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3322 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3311 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_3300 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4045 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4045/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_4056 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4056/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4067 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4067/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4078 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4078/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2621 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2610 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_3366 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3355 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3344 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4089 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4089/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1920 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2654 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2643 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2632 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3399 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3388 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3377 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_1953 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_1942 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1931 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_2698 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2687 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2676 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_2665 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1986 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_1975 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1964 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1997 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5280 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5291 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_4590 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_6909 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_6909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1205 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1249 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1238 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1227 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_1216 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9513 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9502 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_8812 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_8801 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9557 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_9546 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9535 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9524 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8845 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8834 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8823 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_9579 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9568 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_8878 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8867 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8856 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8889 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3141 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3130 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3174 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3163 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_3152 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2473 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_2462 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2451 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_2440 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3196 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_3185 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1761 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_1750 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_2495 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2484 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1794 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1783 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1772 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_809 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8108 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8119 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_7407 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7418 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7429 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_6706 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6717 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6728 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6739 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1024 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1024/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1013 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1013/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1002 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1002/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_1057 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1057/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1046 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1046/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1035 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1035/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1079 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1079/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1068 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1068/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9321 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9310 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_8620 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9365 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_9354 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9343 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9332 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8653 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8642 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8631 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9398 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9387 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9376 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8697 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_8686 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8675 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8664 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7930 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7941 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_7952 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_7963 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7974 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7985 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7996 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2281 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2270 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2292 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1591 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1580 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_639 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_628 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_617 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_606 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7204 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7215 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7226 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7237 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6503 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7248 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_7259 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_6514 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6525 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6536 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_6547 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6558 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6569 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_5802 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5813 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_5824 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_5835 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5846 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_5857 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_5868 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5879 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9140 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9173 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9162 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9151 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_9195 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9184 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8450 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_8461 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8472 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8483 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_8494 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_7760 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7771 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7782 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7793 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5109 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_5109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_414 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_403 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4408 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_447 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_436 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_425 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_3707 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4419 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_469 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_458 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3729 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3718 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7001 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7001/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7012 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7012/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7023 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7023/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_7034 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7034/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_7045 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7045/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7056 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7056/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6300 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6311 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7067 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7067/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7078 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7078/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7089 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7089/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_6322 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6333 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6344 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_6355 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6366 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6377 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5610 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5621 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5632 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6388 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_6399 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_5643 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_5654 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5665 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_5676 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4920 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4931 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5687 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5698 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4942 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4953 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4964 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_992 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_981 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_970 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4975 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4986 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_4997 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_8280 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8291 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_7590 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9909 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_9909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_222 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_211 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_200 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4205 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4216 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_4227 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_255 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_244 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_233 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3515 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_3504 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4238 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_4249 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_288 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_277 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_266 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_2803 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_3548 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3537 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3526 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_299 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2847 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_2836 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2825 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2814 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3559 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2869 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2858 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6130 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_6141 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6152 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6163 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_6174 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6185 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6196 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_5440 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5451 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_5462 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5473 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5484 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5495 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4750 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4761 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4772 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_4783 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4794 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1409 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_1409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9706 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_9717 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9728 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9739 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_4002 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4002/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4013 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4013/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_4024 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4024/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4035 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4035/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_3323 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3312 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_3301 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4046 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4046/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_4057 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4057/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4068 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4068/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2622 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_2611 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2600 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_3367 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3356 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3345 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3334 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4079 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4079/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1910 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2655 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_2644 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2633 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3389 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3378 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_1943 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_1932 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1921 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2688 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_2677 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2666 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1987 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_1976 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1965 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1954 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2699 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1998 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_5270 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5281 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5292 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_4580 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4591 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3890 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_1206 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_1239 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1228 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1217 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9514 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_9503 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_8802 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9547 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_9536 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9525 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8846 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_8835 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8824 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8813 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9569 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9558 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8879 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_8868 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_8857 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3131 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3120 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2430 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3175 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3164 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3153 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_3142 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_2463 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2452 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2441 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3197 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_3186 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_1762 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_1751 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1740 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_2496 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2485 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_2474 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1795 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1784 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1773 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8109 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_8109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7408 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7419 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_6707 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6718 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6729 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1014 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1014/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1003 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1003/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_1047 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1047/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1036 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1036/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_1025 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1025/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1069 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1069/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_1058 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1058/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_9322 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9311 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9300 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8610 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9355 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9344 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9333 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8654 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8643 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8632 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8621 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9399 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_9388 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9377 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9366 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8687 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8676 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8665 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_7920 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7931 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_7942 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8698 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_7953 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7964 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7975 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_7986 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7997 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2271 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2260 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_1570 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2293 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_2282 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1592 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1581 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_629 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_618 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_607 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7205 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7216 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7227 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7238 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7249 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6504 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_6515 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6526 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6537 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6548 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6559 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_5803 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5814 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5825 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5836 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5847 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_5858 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5869 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9130 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9163 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9152 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_9141 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9196 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9185 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_9174 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_8440 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_8451 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8462 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8473 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8484 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8495 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_7750 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7761 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7772 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7783 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7794 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2090 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2090/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_404 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4409 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_4409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_437 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_426 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_415 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_459 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_448 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3719 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3708 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7002 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7002/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7013 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7013/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_7024 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7024/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_7035 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7035/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7046 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7046/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6301 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7057 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7057/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_7068 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7068/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7079 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7079/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_6312 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_6323 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6334 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6345 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5600 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6356 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6367 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6378 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5611 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5622 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_5633 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6389 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_5644 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5655 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_5666 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4910 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4921 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_960 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5677 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5688 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5699 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4932 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4943 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4954 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_4965 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_993 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_982 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_971 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4976 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4987 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_4998 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_8270 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8281 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8292 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7580 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7591 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_6890 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_212 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_201 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4206 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4217 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_256 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_245 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_234 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_223 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3516 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_3505 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4228 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_4239 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_289 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_278 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_267 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_2804 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_3549 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3538 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3527 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2837 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_2826 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2815 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2859 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2848 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6120 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_6131 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6142 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6153 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6164 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6175 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6186 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5430 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5441 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6197 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5452 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_5463 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5474 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_4740 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5485 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_5496 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4751 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4762 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_4773 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_790 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_4784 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4795 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9707 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_9718 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9729 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_4003 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4003/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4014 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4014/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4025 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4025/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_3324 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3313 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3302 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4036 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4036/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_4047 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4047/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4058 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4058/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4069 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4069/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2612 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2601 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_3357 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3346 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3335 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1911 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_1900 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2645 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2634 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2623 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3379 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_3368 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_1944 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_1933 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1922 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_2689 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2678 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2667 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_2656 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1977 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_1966 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1955 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1999 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1988 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5260 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5271 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5282 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5293 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_4570 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4581 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_3880 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4592 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3891 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1229 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1218 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_1207 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_9504 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_8803 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9548 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_9537 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9526 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9515 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8836 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8825 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8814 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_9559 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8869 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_8858 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8847 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3132 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3121 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_3110 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2420 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_3165 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3154 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_3143 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2464 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_2453 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2442 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_2431 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3198 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3187 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_3176 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1752 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_1741 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1730 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_2497 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2486 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2475 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1785 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1774 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1763 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_1796 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_5090 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5090/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_7409 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_7409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6708 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6719 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1004 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1004/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_1048 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1048/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1037 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1037/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1026 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1026/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_1015 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1015/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1059 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1059/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9312 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9301 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_8611 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8600 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9356 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_9345 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9334 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_9323 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8644 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8633 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8622 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9389 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9378 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9367 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8688 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_8677 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8666 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8655 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_7910 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7921 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7932 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_7943 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8699 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_7954 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7965 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_7976 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7987 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7998 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2272 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2261 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2250 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_1560 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2294 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2283 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1593 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1582 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1571 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9890 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_619 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_608 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7206 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7217 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7228 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7239 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6505 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6516 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6527 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_6538 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6549 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_5804 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5815 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5826 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5837 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5848 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_5859 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9131 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9120 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9164 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9153 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9142 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8430 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9197 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9186 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9175 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8441 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8452 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8463 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8474 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_8485 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8496 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_7740 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_7751 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_7762 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7773 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7784 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_7795 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2080 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2080/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2091 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2091/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1390 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_405 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_438 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_427 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_416 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_449 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3709 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_3709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7003 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7003/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7014 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7014/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7025 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7025/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7036 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7036/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7047 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7047/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6302 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7058 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7058/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7069 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7069/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_6313 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6324 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6335 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_6346 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6357 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6368 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5601 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5612 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5623 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6379 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5634 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_5645 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5656 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_5667 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4900 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4911 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4922 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_950 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5678 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5689 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4933 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4944 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4955 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_994 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_983 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_972 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_961 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4966 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4977 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_4988 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_4999 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_8260 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_8271 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8282 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_8293 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_7570 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7581 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7592 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6880 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6891 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_213 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_202 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4207 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4218 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_246 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_235 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_224 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3506 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4229 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_279 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_268 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_257 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3539 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3528 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3517 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2838 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_2827 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2816 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2805 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_2849 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6110 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_6121 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_6132 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6143 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6154 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_6165 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6176 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6187 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5420 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5431 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5442 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6198 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_5453 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5464 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_5475 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4730 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5486 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5497 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4741 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4752 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4763 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_791 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_780 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4774 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_4785 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4796 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8090 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8090/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9708 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_9719 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_4004 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4004/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4015 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4015/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4026 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4026/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_3314 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3303 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4037 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4037/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_4048 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4048/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4059 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4059/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2613 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_2602 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_3358 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3347 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3336 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_3325 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1901 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2646 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_2635 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2624 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3369 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_1934 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1923 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1912 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2679 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2668 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2657 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1978 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_1967 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1956 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1945 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_1989 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_5250 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5261 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5272 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5283 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5294 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4560 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4571 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4582 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3870 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4593 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3892 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3881 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_1219 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1208 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_9505 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9538 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_9527 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9516 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8837 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_8826 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8815 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8804 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9549 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8859 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8848 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3122 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3111 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_3100 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2421 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2410 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_3166 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3155 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3144 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_3133 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_2454 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2443 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2432 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3199 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3188 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3177 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_1753 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_1742 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1731 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1720 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2487 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2476 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_2465 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1786 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_1775 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1764 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_2498 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1797 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5080 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5080/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5091 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5091/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_4390 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_6709 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_6709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1005 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1005/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1038 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1038/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1027 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1027/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_1016 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1016/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_1049 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1049/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_9313 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9302 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_8601 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9346 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9335 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9324 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8645 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8634 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8623 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8612 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9379 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9368 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9357 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_7900 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8678 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8667 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8656 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_7911 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7922 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_7933 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8689 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_7944 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7955 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_7966 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_7977 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7988 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7999 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2262 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2251 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_2240 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_1561 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_1550 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_2295 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2284 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_2273 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1594 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1583 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1572 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9880 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_9891 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_609 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7207 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7218 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7229 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_6506 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6517 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6528 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6539 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_5805 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5816 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5827 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5838 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_5849 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_9121 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9110 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_8420 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9154 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9143 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9132 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8431 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9198 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9187 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9176 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_9165 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8442 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8453 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8464 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_8475 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8486 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7730 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7741 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8497 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_7752 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_7763 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7774 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7785 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7796 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2081 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2081/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2070 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2070/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2092 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2092/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1391 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1380 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_428 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_417 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_406 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_439 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_7004 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7004/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7015 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7015/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7026 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7026/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7037 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7037/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7048 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7048/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_7059 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7059/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_6303 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_6314 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6325 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6336 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_6347 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6358 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6369 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_5602 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5613 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_5624 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_5635 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5646 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_5657 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4901 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4912 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_951 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_940 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5668 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5679 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4923 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4934 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4945 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_4956 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_984 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_973 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_962 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_4967 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4978 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_4989 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_995 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8250 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_8261 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8272 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8283 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_8294 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_7560 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7571 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7582 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7593 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_6870 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6881 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_6892 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_203 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4208 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_247 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_236 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_225 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_214 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3507 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4219 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_269 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_258 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3529 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3518 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2828 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_2817 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2806 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2839 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6100 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6111 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_6122 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6133 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6144 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_6155 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6166 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6177 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5410 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5421 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5432 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6188 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_6199 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_5443 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_5454 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5465 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4720 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4731 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5476 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_5487 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5498 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4742 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4753 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4764 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_792 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_781 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_770 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4775 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4786 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_4797 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_8080 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8080/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8091 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8091/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_7390 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9709 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_9709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_4005 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4005/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4016 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4016/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_3315 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_3304 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4027 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4027/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_4038 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4038/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_4049 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4049/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2603 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_3348 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3337 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3326 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_1902 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2636 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2625 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2614 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3359 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1935 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1924 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1913 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_2669 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2658 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_2647 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1968 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_1957 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1946 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1979 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5240 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5251 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_5262 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5273 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5284 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5295 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4550 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4561 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4572 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3871 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_3860 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4583 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4594 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3893 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3882 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1209 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_1209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9539 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_9528 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9517 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9506 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8827 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8816 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8805 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_8849 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8838 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3123 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3112 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_3101 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2411 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2400 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_3156 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3145 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3134 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1710 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2455 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_2444 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2433 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_2422 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3189 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3178 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_3167 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1743 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_1732 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1721 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2488 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_2477 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2466 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1776 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1765 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1754 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2499 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1798 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1787 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5070 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5070/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5081 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5081/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5092 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5092/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_4380 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4391 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3690 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_1039 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1039/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1028 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1028/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1017 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1017/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_1006 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1006/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_9303 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_8602 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9347 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_9336 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9325 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_9314 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8635 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8624 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8613 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9369 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9358 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8679 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_8668 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_8657 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8646 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_7901 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7912 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7923 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_7934 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_7945 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7956 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_7967 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7978 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7989 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2230 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_2263 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2252 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2241 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1551 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1540 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_2296 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2285 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_2274 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1595 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1584 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1573 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1562 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9870 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9881 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9892 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7208 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7219 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_6507 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6518 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6529 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_5806 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_5817 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5828 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5839 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_9122 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9111 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9100 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8410 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9155 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9144 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9133 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8432 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8421 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9188 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9177 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9166 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8443 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9199 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_8454 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8465 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8476 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8487 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7720 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7731 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_7742 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8498 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_7753 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7764 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7775 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_7786 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7797 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2071 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2071/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2060 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2060/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_1370 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2093 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2093/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_2082 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2082/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1392 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1381 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_429 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_418 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_407 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7005 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7005/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7016 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7016/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7027 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7027/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7038 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7038/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7049 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7049/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6304 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_6315 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6326 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6337 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6348 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6359 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_5603 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5614 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5625 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5636 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5647 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_5658 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4902 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4913 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_941 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_930 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5669 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4924 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4935 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_4946 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_985 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_974 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_963 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_952 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4957 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4968 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_4979 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_996 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8240 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_8251 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8262 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8273 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8284 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8295 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_7550 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7561 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7572 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7583 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7594 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_6860 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6871 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6882 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6893 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_204 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4209 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_4209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_237 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_226 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_215 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_259 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_248 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3519 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3508 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_2829 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_2818 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2807 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6101 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_6112 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_6123 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6134 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6145 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_6156 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6167 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5400 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5411 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5422 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_5433 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6178 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_6189 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_5444 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5455 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_5466 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4710 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4721 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_760 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5477 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5488 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5499 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4732 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4743 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4754 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_793 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_782 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_771 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4765 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4776 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4787 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_4798 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_8070 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8070/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8081 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8081/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8092 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8092/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7380 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7391 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_6690 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_4006 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4006/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4017 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4017/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_3305 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4028 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4028/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_4039 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4039/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2604 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_3349 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3338 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3327 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_3316 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2637 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_2626 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2615 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1925 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1914 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1903 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2659 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2648 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1969 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_1958 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1947 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1936 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5230 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5241 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_5252 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_5263 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5274 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_5285 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_5296 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4540 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4551 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4562 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_4573 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_590 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_3861 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_3850 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4584 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4595 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3894 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3883 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3872 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9529 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_9518 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9507 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8828 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_8817 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8806 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8839 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3113 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3102 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2412 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2401 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_3157 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3146 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3135 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_3124 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1700 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2445 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2434 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2423 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3179 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_3168 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_1744 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_1733 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1722 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1711 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2478 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2467 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_2456 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1777 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_1766 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1755 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_2489 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1799 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1788 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5060 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5060/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5071 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5071/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5082 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5082/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5093 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5093/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_4370 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4381 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_4392 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3691 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3680 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2990 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_1029 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1029/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1018 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1018/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_1007 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1007/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_9304 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9337 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9326 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9315 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8636 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8625 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8614 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8603 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9359 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9348 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8669 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_8658 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8647 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_7902 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7913 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_7924 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_7935 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7946 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_7957 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_7968 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7979 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2220 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2253 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2242 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_2231 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1552 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_1541 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1530 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_2297 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2286 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2275 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_2264 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1585 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1574 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1563 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_1596 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9860 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9871 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9882 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9893 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_7209 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_7209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6508 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6519 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5807 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5818 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5829 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_9112 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9101 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_8411 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8400 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9145 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9134 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_9123 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8433 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8422 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9189 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9178 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9167 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_9156 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8444 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8455 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_8466 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8477 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7710 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7721 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7732 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8488 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_8499 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_7743 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_7754 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7765 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_7776 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7787 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7798 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2072 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2072/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2061 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2061/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2050 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2050/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_1360 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2094 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2094/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2083 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2083/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1393 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1382 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1371 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9690 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_419 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_408 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7006 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7006/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7017 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7017/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7028 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7028/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7039 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7039/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6305 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6316 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6327 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_6338 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6349 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_5604 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5615 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5626 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5637 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5648 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4903 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_942 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_931 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_920 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5659 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4914 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4925 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_4936 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_4947 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_975 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_964 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_953 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4958 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4969 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_997 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_986 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8230 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_8241 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8252 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8263 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8274 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_8285 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7540 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_7551 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8296 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_7562 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7573 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7584 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_7595 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_6850 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6861 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6872 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_6883 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6894 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1190 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_238 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_227 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_216 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_205 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_249 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3509 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_3509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2819 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_2808 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6102 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_6113 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6124 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6135 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_6146 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6157 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6168 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5401 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5412 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5423 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6179 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5434 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_5445 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5456 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4700 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4711 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4722 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_750 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5467 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5478 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5489 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4733 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4744 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4755 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_783 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_772 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_761 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4766 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4777 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_4788 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_794 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4799 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_8060 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8060/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_8071 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8071/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8082 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8082/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_8093 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8093/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_7370 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7381 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7392 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6680 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6691 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_5990 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_4007 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4007/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_3306 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4018 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4018/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_4029 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4029/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3339 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3328 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3317 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2627 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2616 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2605 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1926 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_1915 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1904 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2649 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2638 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1959 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1948 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1937 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5220 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5231 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5242 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_5253 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5264 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_5275 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4530 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5286 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5297 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4541 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4552 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4563 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_591 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_580 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_3862 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_3851 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4574 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_4585 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4596 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_3840 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3895 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3884 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3873 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9519 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9508 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8818 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8818/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_8807 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8807/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8829 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8829/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3114 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3103 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2402 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_3147 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3136 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_3125 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1701 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2446 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_2435 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2424 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_2413 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3169 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_3158 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1734 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1723 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1712 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2479 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2468 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2457 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1767 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1756 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1745 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_1789 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1778 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5050 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5050/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5061 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5061/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5072 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5072/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5083 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5083/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5094 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5094/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4360 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4371 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_3670 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4382 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_4393 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3692 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3681 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2991 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2980 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_1019 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1019/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1008 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1008/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_9338 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_9327 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9316 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9305 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_8626 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8626/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8615 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8615/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8604 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8604/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9349 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8659 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8659/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8648 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8648/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8637 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8637/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7903 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7914 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7925 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7936 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7947 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_7958 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7969 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2221 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2210 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2254 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2243 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2232 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1542 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1531 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1520 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2287 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2276 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_2265 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1586 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_1575 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1564 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1553 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2298 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1597 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9850 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9861 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_9872 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9883 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_9894 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4190 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_6509 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_6509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5808 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5819 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9113 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9102 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_8401 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8401/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9146 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9135 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9124 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8434 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8434/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8423 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8423/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8412 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8412/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9179 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9168 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9157 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_7700 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8445 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8445/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8456 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8456/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8467 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8467/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8478 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8478/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7711 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7722 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_7733 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8489 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8489/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_7744 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7755 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_7766 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_7777 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7788 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7799 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2062 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2062/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2051 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2051/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_2040 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2040/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_1361 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_1350 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_2095 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2095/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2084 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2084/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_2073 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2073/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1394 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1383 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1372 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9691 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_9680 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8990 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8990/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_409 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7007 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7007/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7018 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7018/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7029 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7029/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_6306 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6317 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6328 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6339 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_5605 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5616 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5627 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5638 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_5649 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4904 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_932 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_921 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_910 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4915 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4926 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_4937 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_976 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_965 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_954 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_943 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4948 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4959 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_998 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_987 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8220 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8220/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_8231 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8231/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_8242 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8242/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8253 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8253/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8264 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8264/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_8275 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8275/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8286 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8286/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7530 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7541 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8297 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8297/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_7552 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_7563 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7574 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6840 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_7585 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7596 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_6851 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6862 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6873 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_6884 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6895 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1191 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1180 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_228 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_217 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_206 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_239 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2809 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_2809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6103 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_6114 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6125 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6136 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_6147 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6158 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5402 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5413 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_5424 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6169 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_5435 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5446 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_5457 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4701 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4712 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_751 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_740 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5468 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5479 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4723 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4734 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4745 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_784 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_773 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_762 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_4756 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4767 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4778 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_4789 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_795 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8050 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8050/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_8061 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8061/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8072 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8072/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8083 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8083/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_8094 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8094/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_7360 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7371 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7382 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7393 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_6670 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6681 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_6692 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5980 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5991 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_4008 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4008/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_4019 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4019/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3329 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3318 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_3307 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_2628 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_2617 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2606 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_1916 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_1905 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_2639 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1949 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1938 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1927 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5210 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5221 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5232 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_5243 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_5254 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5265 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4520 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5276 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_5287 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5298 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4531 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_4542 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4553 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4564 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_592 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_581 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_570 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_3852 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4575 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4586 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_4597 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_3830 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3841 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3885 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3874 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3863 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_3896 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_7190 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9509 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_9509/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8808 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8808/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8819 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8819/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3104 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2403 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_3148 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3137 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_3126 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_3115 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2436 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2425 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2414 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3159 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1735 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1724 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1713 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1702 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2469 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2458 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_2447 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1768 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_1757 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1746 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1779 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5040 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5040/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5051 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5051/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_5062 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5062/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5073 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5073/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5084 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5084/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5095 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5095/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4350 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4361 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4372 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3660 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4383 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4394 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3693 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3682 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3671 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2992 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_2981 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2970 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_1009 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_1009/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9328 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9328/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9317 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9317/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9306 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9306/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8627 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8627/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8616 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8616/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8605 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8605/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9339 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9339/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_8649 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8649/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8638 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8638/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7904 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7915 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7926 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7937 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7948 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_7959 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2211 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2200 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_1510 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2244 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2233 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_2222 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1543 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_1532 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1521 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2288 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_2277 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2266 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_2255 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1576 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1565 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1554 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2299 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1598 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1587 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9840 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9840/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9851 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9851/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_9862 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9862/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9873 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9873/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9884 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9884/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_9895 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9895/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_4180 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4191 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3490 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5809 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_5809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_9103 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9103/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_8402 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8402/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9136 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9136/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9125 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9125/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_9114 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9114/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8435 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8435/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8424 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8424/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8413 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8413/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9169 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9169/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9158 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9158/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_9147 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9147/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_8446 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8446/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_8457 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8457/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8468 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8468/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7701 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7712 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7723 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8479 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8479/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_7734 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_7745 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7756 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_7767 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7778 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7789 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2063 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2063/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2052 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2052/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2041 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2041/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_2030 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2030/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_1351 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1340 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_2096 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2096/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2085 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2085/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_2074 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2074/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1384 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1373 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1362 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_1395 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9692 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9692/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_9670 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9670/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9681 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9681/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8991 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8991/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_8980 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8980/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7008 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7008/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7019 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7019/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_6307 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6318 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6329 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_5606 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_900 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5617 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5628 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5639 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_933 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_922 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_911 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4905 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4916 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_4927 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_4938 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_966 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_955 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_944 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4949 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_999 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_988 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_977 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8210 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8210/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_8221 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8221/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_8232 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8232/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8243 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8243/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8254 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8254/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8265 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8265/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8276 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8276/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7520 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7531 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_7542 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8287 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8287/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8298 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8298/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_7553 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7564 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7575 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6830 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7586 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7597 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_6841 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6852 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6863 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_6874 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6885 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6896 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_1192 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1181 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_1170 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_229 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_218 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_207 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6104 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_6115 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6126 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6137 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6148 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6159 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_5403 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5414 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5425 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5436 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5447 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4702 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4713 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_741 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_730 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5458 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5469 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4724 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4735 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_4746 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_774 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_763 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_752 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4757 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4768 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_4779 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_796 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_785 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8040 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8040/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_8051 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8051/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8062 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8062/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8073 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8073/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8084 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8084/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8095 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8095/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_7350 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7361 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7372 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7383 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7394 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_6660 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6671 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6682 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6693 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5970 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5981 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5992 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_4009 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_4009/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_3319 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3308 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_2618 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2607 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1917 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_1906 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2629 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1939 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1928 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5200 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5211 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5222 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_5233 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_5244 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5255 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_5266 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4510 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4521 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5277 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5288 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5299 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4532 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4543 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4554 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_593 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_582 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_571 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_560 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3853 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4565 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4576 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4587 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_3820 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_3831 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3842 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3886 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_3875 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3864 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_4598 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3897 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_7180 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7191 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_6490 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_8809 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_8809/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_3105 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_3138 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_3127 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_3116 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2437 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_2426 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2415 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2404 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_3149 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1725 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1714 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1703 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2459 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2448 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1758 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1747 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1736 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_1769 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_5030 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5030/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5041 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5041/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_5052 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5052/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_5063 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5063/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5074 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5074/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_5085 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5085/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_5096 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5096/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4340 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4351 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4362 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_390 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_3661 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_3650 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4373 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_4384 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4395 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3694 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3683 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3672 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2982 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_2971 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2960 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2993 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_9329 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9329/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_9318 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9318/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9307 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9307/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8617 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8617/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8606 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8606/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8639 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8639/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_8628 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8628/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7905 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7916 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7927 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7938 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7949 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2212 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2201 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_1500 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2245 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2234 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2223 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1533 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1522 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1511 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2278 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2267 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_2256 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1577 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_1566 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1555 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1544 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2289 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1599 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1588 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9841 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9841/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9830 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9830/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9852 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9852/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_9863 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9863/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9874 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9874/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_9885 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9885/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_9896 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9896/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_4170 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4181 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_4192 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3491 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3480 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2790 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_9104 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9104/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9137 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9137/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9126 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9126/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9115 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9115/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8425 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8425/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8414 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8414/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8403 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8403/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9159 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9159/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9148 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9148/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8436 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8436/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8447 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8447/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_8458 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8458/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8469 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8469/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_7702 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7713 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_7724 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_7735 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7746 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_7757 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_7768 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7779 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2020 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2020/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2053 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2053/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2042 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2042/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_2031 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2031/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1341 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1330 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_2086 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2086/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2075 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2075/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_2064 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2064/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1385 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1374 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1363 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_1352 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2097 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2097/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_1396 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9693 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9693/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_9660 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9660/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9671 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9671/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9682 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9682/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_8981 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8981/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8970 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8970/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8992 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8992/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7009 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_7009/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6308 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6319 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5607 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5618 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5629 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_923 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_912 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_901 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4906 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4917 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_4928 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_967 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_956 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_945 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_934 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4939 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_989 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_978 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8200 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8200/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8211 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8211/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8222 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8222/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_8233 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8233/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8244 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8244/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8255 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8255/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_8266 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8266/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8277 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8277/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7510 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7521 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7532 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8288 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8288/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_8299 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8299/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_7543 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_7554 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7565 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6820 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7576 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7587 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7598 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_6831 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6842 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6853 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6864 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6875 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6886 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_6897 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_1160 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_1193 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1182 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_1171 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9490 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9490/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_219 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_208 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6105 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6116 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6127 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_6138 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6149 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_5404 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5415 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5426 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5437 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5448 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4703 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_742 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_731 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_720 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5459 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4714 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4725 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_4736 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_775 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_764 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_753 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4747 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4758 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4769 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_797 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_786 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8030 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8030/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_8041 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8041/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8052 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8052/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8063 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8063/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8074 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8074/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_8085 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8085/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7340 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_8096 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8096/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_7351 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_7362 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7373 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7384 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_7395 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_6650 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6661 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6672 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_6683 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6694 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_5960 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5971 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5982 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5993 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3309 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_3309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2619 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_2608 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_1907 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1929 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1918 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5201 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5212 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5223 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_5234 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_5245 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5256 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4500 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4511 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_550 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5267 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5278 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5289 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4522 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_4533 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4544 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4555 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3810 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_583 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_572 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_561 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_4566 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4577 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_4588 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3821 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_3832 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3843 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_594 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3876 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3865 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3854 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_4599 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3898 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3887 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7170 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7181 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7192 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6480 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6491 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_5790 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_3139 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3128 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3117 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_3106 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2427 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2416 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2405 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1726 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_1715 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1704 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2449 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2438 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1759 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1748 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1737 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5020 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5020/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5031 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5031/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5042 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5042/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_5053 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5053/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5064 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5064/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_5075 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5075/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_5086 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5086/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5097 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5097/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4330 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4341 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4352 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4363 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_391 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_380 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_3651 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3640 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4374 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_4385 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4396 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2950 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3695 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3684 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3673 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3662 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2983 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_2972 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2961 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2994 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_9319 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9319/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9308 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9308/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8618 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8618/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_8607 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8607/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8629 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8629/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_7906 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7917 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7928 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7939 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2202 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2235 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2224 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_2213 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1534 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1523 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1512 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_1501 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2279 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2268 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2257 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_2246 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1567 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1556 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1545 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_1589 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1578 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9842 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9842/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_9831 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9831/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9820 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9820/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9853 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9853/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9864 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9864/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9875 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9875/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_9886 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9886/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9897 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9897/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_4160 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4171 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4182 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_4193 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3492 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3481 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_3470 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2791 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2780 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_9127 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9127/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9116 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9116/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9105 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9105/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_8426 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8426/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8415 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8415/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8404 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8404/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9149 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9149/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_9138 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9138/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_8437 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8437/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_8448 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8448/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8459 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8459/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_7703 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7714 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7725 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7736 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7747 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_7758 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7769 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2010 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2010/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2054 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2054/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2043 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2043/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2032 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2032/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_2021 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2021/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_1342 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1331 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1320 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_2087 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2087/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2076 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2076/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_2065 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2065/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1375 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1364 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1353 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2098 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2098/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1397 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_1386 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9650 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9650/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9661 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9661/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_9672 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9672/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9683 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9683/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_8982 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8982/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_8971 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8971/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8960 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8960/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9694 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9694/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8993 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8993/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_6309 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_6309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5608 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5619 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_924 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_913 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_902 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4907 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4918 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_4929 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_957 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_946 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_935 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_979 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_968 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_8201 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8201/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_8212 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8212/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_8223 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8223/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8234 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8234/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8245 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8245/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8256 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8256/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8267 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8267/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7500 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_7511 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7522 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_7533 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8278 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8278/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8289 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8289/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_7544 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7555 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_7566 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6810 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_6821 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7577 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7588 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7599 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_6832 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6843 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6854 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_6865 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6876 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6887 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_6898 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1150 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_1183 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1172 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_1161 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_1194 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_9491 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9491/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_9480 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9480/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8790 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8790/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_209 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_6106 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6117 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6128 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6139 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_5405 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5416 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5427 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5438 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_4704 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_732 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_721 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_710 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5449 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4715 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4726 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_4737 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_765 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_754 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_743 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4748 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4759 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_798 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_787 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_776 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8020 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8020/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_8031 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8031/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_8042 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8042/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8053 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8053/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8064 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8064/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_8075 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8075/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8086 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8086/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7330 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7341 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_8097 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8097/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_7352 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_7363 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7374 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7385 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7396 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_6640 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_6651 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6662 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6673 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_6684 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6695 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_5950 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5961 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5972 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5983 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5994 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2609 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_2609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1908 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_1919 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5202 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5213 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_5224 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_5235 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5246 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_5257 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4501 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4512 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_540 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5268 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5279 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4523 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4534 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4545 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3800 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_584 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_573 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_562 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_551 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3844 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4556 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4567 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4578 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_3811 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_3822 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3833 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_595 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3877 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_3866 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3855 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_4589 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3899 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3888 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7160 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_7171 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_7182 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7193 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_6470 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6481 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_6492 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5780 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5791 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3129 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3118 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_3107 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_2428 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_2417 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2406 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_1716 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_1705 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_2439 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1749 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1738 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1727 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5010 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5010/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5021 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5021/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5032 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5032/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_5043 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5043/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_5054 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5054/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5065 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5065/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4320 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5076 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5076/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_5087 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5087/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5098 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5098/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4331 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_4342 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4353 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_392 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_381 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_370 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_3652 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_3641 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3630 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4364 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_4375 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4386 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_4397 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2940 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3685 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3674 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3663 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2973 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_2962 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2951 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3696 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2995 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2984 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_9309 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_9309/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8608 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8608/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8619 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8619/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_7907 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7918 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7929 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_2203 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2236 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2225 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2214 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1524 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1513 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1502 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2269 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2258 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_2247 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1568 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_1557 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1546 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1535 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1579 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9832 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9832/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_9821 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9821/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9810 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9810/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9843 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9843/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9854 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9854/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9865 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9865/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_9876 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9876/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_9887 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9887/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9898 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9898/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_4150 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4161 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_3460 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4172 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_4183 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_4194 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3493 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3482 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3471 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2792 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_2781 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2770 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9128 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9128/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_9117 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9117/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9106 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9106/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8416 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8416/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8405 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8405/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9139 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9139/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_8427 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8427/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8438 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8438/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_8449 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8449/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_7704 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7715 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7726 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7737 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7748 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_7759 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2011 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2011/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2000 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2000/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2044 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2044/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2033 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2033/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_2022 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2022/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1332 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1321 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_1310 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_2077 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2077/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2066 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2066/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_2055 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2055/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1376 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_1365 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1354 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_1343 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2099 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2099/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2088 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2088/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_1398 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1387 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9640 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9640/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9684 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9684/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_9651 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9651/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_9662 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9662/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9673 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9673/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8972 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8972/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8961 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8961/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8950 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8950/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9695 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9695/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8994 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8994/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8983 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8983/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3290 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5609 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_5609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_914 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_914/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_903 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_903/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4908 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_4919 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_958 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_958/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_947 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_947/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_936 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_936/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_925 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_925/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_969 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_969/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_8202 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8202/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_8213 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8213/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_8224 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8224/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8235 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8235/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8246 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8246/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_8257 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8257/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8268 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8268/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7501 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7512 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7523 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8279 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8279/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_7534 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_7545 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7556 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6800 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6811 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7567 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7578 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7589 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_6822 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6833 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6844 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_6855 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6866 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6877 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_6888 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_6899 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1151 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_1140 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_1184 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1173 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_1162 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_1195 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9492 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9492/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_9481 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9481/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9470 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9470/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8780 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8780/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8791 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8791/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_6107 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_6118 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_6129 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_5406 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_5417 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5428 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5439 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_733 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_733/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_722 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_722/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_711 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_711/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_700 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_700/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4705 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4716 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_4727 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_766 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_766/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_755 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_755/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_744 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_744/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4738 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_4749 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_799 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_799/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_788 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_788/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_777 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_777/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8010 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8010/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_8021 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8021/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_8032 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8032/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8043 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8043/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8054 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8054/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8065 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8065/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8076 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8076/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7320 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7331 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_8087 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8087/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8098 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8098/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_7342 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_7353 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7364 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7375 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6630 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7386 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7397 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_6641 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6652 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6663 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_6674 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6685 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6696 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_5940 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5951 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_5962 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5973 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5984 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5995 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1909 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_1909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5203 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5214 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5225 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5236 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5247 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4502 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_541 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_541/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_530 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_530/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5258 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5269 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4513 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_4524 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4535 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_4546 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3801 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_574 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_574/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_563 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_563/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_552 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_552/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4557 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4568 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_4579 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_3812 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_3823 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3834 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_596 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_596/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_585 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_585/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3867 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3856 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3845 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_3889 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3878 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7150 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_7161 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_7172 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_7183 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_7194 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_6460 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6471 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6482 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6493 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5770 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5781 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5792 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3119 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_3108 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_2418 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2407 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1717 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_1706 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2429 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1739 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1728 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5000 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5000/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5011 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5011/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5022 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5022/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_5033 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5033/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_5044 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5044/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5055 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5055/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_4310 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5066 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5066/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_5077 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5077/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5088 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5088/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5099 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5099/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4321 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_4332 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4343 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4354 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_382 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_382/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_371 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_371/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_360 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_360/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3642 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3631 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3620 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4365 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4376 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4387 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_393 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_393/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_2941 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_2930 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3686 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_3675 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3664 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3653 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4398 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2974 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_2963 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2952 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_3697 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2996 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2985 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6290 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_8609 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_8609/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7908 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7919 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_2226 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2215 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2204 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_1525 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1514 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1503 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2259 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2248 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_2237 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1558 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1547 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1536 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_1569 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9833 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9833/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_9822 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9822/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9811 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9811/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9800 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9800/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9844 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9844/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9855 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9855/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9866 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9866/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_9877 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9877/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9888 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9888/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9899 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9899/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_4140 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4151 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_4162 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_190 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_190/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_3450 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_4173 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_4184 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_4195 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_3494 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_3483 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3472 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3461 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2782 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_2771 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2760 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2793 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_9118 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9118/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9107 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9107/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8417 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8417/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8406 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8406/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_9129 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9129/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_8428 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8428/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_8439 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8439/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_7705 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7716 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7727 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7738 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7749 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2001 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2001/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_1300 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_2045 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2045/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2034 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2034/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2023 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2023/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_2012 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2012/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_1333 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1322 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1311 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2078 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2078/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2067 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2067/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_2056 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2056/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1366 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1355 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1344 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2089 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2089/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1399 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1388 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_1377 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9630 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9630/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9641 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9641/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9652 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9652/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_9663 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9663/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9674 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9674/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_8973 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8973/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_8962 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8962/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8951 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8951/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8940 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8940/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9696 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9696/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9685 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9685/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8995 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8995/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8984 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8984/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3291 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3280 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2590 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_915 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_915/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_904 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_904/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4909 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_4909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_948 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_948/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_937 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_937/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_926 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_926/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_959 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_959/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8203 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8203/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_8214 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8214/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8225 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8225/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8236 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8236/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8247 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8247/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_8258 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8258/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7502 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7513 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_7524 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8269 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8269/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_7535 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7546 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_7557 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6801 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_6812 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7568 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7579 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_6823 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6834 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6845 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_6856 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6867 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6878 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_6889 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1141 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_1130 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_1174 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_1163 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_1152 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_1196 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_1185 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_9482 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9482/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9471 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9471/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9460 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9460/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_8781 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8781/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8770 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8770/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9493 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9493/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_8792 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8792/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_6108 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_6119 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5407 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5418 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5429 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_723 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_723/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_712 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_712/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_701 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_701/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4706 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4717 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_4728 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_756 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_756/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_745 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_745/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_734 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_734/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4739 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_789 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_789/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_778 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_778/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_767 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_767/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8000 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8000/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_8011 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8011/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8022 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8022/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_8033 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8033/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8044 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8044/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8055 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8055/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_8066 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8066/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8077 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8077/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7310 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7321 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7332 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8088 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8088/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_8099 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8099/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_7343 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_7354 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7365 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6620 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7376 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7387 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7398 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_6631 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6642 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6653 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6664 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6675 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6686 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_6697 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5930 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5941 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_5952 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_5963 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5974 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_5985 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_5996 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9290 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9290/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5204 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5215 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5226 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5237 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_5248 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4503 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_531 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_531/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_520 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_520/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5259 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4514 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4525 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_4536 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_575 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_575/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_564 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_564/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_553 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_553/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_542 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_542/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4547 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4558 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4569 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_3802 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_3813 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3824 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_597 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_597/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_586 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_586/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_3868 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_3857 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3846 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3835 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_3879 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_7140 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_7151 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_7162 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_7173 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_7184 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_7195 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_6450 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6461 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6472 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_6483 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6494 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_5760 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5771 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5782 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5793 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3109 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_3109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2419 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_2408 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_1707 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1729 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1718 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5001 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5001/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_5012 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5012/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5023 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5023/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_5034 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5034/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_5045 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5045/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5056 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5056/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4300 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4311 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5067 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5067/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5078 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5078/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5089 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5089/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4322 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_4333 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4344 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_383 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_383/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_372 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_372/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_361 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_361/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_350 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_350/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3643 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_3632 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3621 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_3610 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4355 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_4366 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4377 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_4388 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_394 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_394/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2931 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_2920 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_3676 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3665 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3654 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_4399 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2964 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_2953 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2942 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3698 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3687 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2997 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2986 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2975 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6280 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6291 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_5590 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_7909 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_7909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2227 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2216 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2205 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1515 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1504 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2249 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2238 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1559 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1548 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1537 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1526 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9823 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9823/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_9812 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9812/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9801 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9801/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9845 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9845/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9834 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9834/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_9856 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9856/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_9867 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9867/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_9878 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9878/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9889 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9889/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_4130 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4141 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_4152 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_191 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_191/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_180 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_180/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_3451 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3440 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_4163 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_4174 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_4185 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_4196 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_3484 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3473 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3462 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2783 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_2772 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2761 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2750 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3495 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2794 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_9119 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9119/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_9108 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9108/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8407 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8407/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8429 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8429/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_8418 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8418/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7706 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7717 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7728 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7739 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2002 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2002/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2035 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2035/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2024 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2024/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_2013 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2013/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1323 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1312 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_1301 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_2068 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2068/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2057 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2057/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_2046 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2046/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1367 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_1356 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1345 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_1334 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_2079 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2079/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1389 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1378 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_9620 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9620/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9631 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9631/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_8930 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8930/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9642 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9642/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_9653 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9653/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9664 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9664/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9675 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9675/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8963 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8963/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8952 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8952/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8941 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8941/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9697 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9697/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9686 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9686/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8996 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8996/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8985 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8985/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8974 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8974/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3292 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3281 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_3270 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2591 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2580 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_1890 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_905 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_905/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_949 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_949/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_938 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_938/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_927 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_927/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_916 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_916/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8204 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8204/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_8215 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8215/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8226 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8226/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8237 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8237/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_8248 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8248/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8259 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8259/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_7503 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7503/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7514 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7514/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7525 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7525/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7536 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7536/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7547 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7547/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6802 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7558 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7558/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7569 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7569/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_6813 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6824 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6835 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_6846 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6857 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6868 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_6879 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1142 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_1131 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_1120 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_1175 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_1164 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_1153 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_1197 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_1186 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9450 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9450/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9483 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9483/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_9472 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9472/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9461 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9461/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8771 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8771/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8760 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8760/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9494 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9494/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8793 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8793/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_8782 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8782/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6109 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_6109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5408 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5419 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_724 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_724/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_713 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_713/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_702 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_702/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4707 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4718 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_757 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_757/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_746 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_746/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_735 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_735/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_4729 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_779 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_779/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_768 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_768/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_8001 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8001/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_8012 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8012/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_8023 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8023/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8034 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8034/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8045 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8045/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8056 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8056/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8067 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8067/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7300 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7300/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_7311 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7311/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7322 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7322/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_8078 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8078/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8089 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8089/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_7333 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7333/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_7344 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7344/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7355 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7355/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_7366 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7366/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6610 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_6621 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7377 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7377/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7388 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7388/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7399 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7399/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_6632 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6643 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6654 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_6665 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6676 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6687 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5920 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5931 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5942 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6698 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_5953 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5964 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_5975 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_5986 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5997 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9291 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9291/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_9280 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9280/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8590 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8590/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5205 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5216 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5227 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5238 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_532 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_532/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_521 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_521/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_510 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_510/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5249 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4504 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4515 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4526 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_4537 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_565 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_565/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_554 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_554/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_543 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_543/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4548 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4559 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_3803 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_3814 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3825 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_598 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_598/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_587 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_587/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_576 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_576/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3858 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3847 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3836 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_3869 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_7130 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7130/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_7141 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7141/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_7152 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7152/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_7163 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7163/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_7174 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7174/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_7185 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7185/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_7196 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7196/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_6440 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_6451 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6462 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6473 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_6484 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6495 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_5750 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5761 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5772 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5783 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5794 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2409 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_2409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1708 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_1719 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_5002 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5002/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5013 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5013/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_5024 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5024/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_5035 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5035/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5046 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5046/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_4301 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_340 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_340/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3600 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_5057 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5057/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_5068 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5068/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5079 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5079/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4312 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_4323 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4334 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4345 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_373 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_373/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_362 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_362/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_351 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_351/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3633 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3622 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3611 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4356 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4367 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4378 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_395 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_395/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_384 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_384/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_2932 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_2921 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2910 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_3666 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3655 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3644 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4389 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2965 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_2954 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2943 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_3699 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3688 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3677 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2998 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2987 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2976 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6270 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6281 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_6292 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5580 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5591 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_4890 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_2217 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2206 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_1516 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_1505 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_2239 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2228 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1549 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1538 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1527 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9824 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9824/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_9813 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9813/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_9802 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9802/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9846 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9846/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9835 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9835/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9857 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9857/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_9868 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9868/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9879 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9879/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_4120 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4131 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_4142 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_4153 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_181 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_181/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_170 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_170/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_3441 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3430 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_4164 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_4175 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_4186 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_192 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_192/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_2740 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3485 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_3474 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3463 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_3452 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_4197 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2773 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_2762 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2751 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3496 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2795 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2784 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_9109 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_9109/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8408 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8408/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8419 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8419/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_7707 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7707/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7718 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7718/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7729 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7729/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_2036 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2036/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2025 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2025/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_2014 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2014/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_2003 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2003/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_1324 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1313 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1302 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_2069 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2069/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2058 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2058/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_2047 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2047/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1357 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1346 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1335 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1379 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1368 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9610 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9610/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9621 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9621/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9632 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9632/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_8920 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8920/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9643 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9643/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_9654 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9654/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9665 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9665/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8964 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8964/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_8953 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8953/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8942 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8942/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8931 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8931/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9698 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9698/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9687 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9687/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9676 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9676/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8997 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8997/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_8986 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8986/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8975 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8975/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3260 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3293 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3282 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3271 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2581 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2570 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_1880 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2592 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1891 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_906 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_906/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_939 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_939/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_928 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_928/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_917 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_917/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8205 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8205/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_8216 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8216/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8227 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8227/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8238 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8238/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_8249 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8249/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_7504 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7504/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7515 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7515/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7526 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7526/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7537 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7537/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7548 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7548/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6803 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7559 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7559/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_6814 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6825 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6836 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_6847 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6858 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6869 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_1132 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_1121 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_1110 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_1165 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_1154 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_1143 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_1198 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_1187 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_1176 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_9440 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9440/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9473 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9473/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_9462 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9462/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_9451 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9451/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8772 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8772/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_8761 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8761/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_8750 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8750/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_9495 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9495/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_9484 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9484/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8794 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8794/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8783 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8783/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3090 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3090/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5409 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_5409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_714 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_714/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_703 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_703/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4708 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_4719 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_747 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_747/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_736 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_736/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_725 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_725/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_769 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_769/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_758 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_758/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_8002 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8002/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_8013 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8013/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_8024 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8024/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_8035 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8035/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_8046 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8046/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_8057 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8057/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8068 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8068/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7301 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7301/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_7312 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7312/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7323 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7323/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8079 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8079/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_7334 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7334/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_7345 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7345/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_7356 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7356/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6600 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6611 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7367 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7367/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_7378 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7378/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_7389 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7389/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_6622 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_6633 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6644 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5910 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_6655 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6666 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6677 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_6688 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5921 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_5932 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_5943 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6699 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_5954 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_5965 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_5976 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_5987 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5998 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9292 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9292/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_9281 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9281/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_9270 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9270/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_8580 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8580/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8591 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8591/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_7890 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7890/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5206 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_5217 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_5228 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_5239 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_522 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_522/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_511 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_511/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_500 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_500/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4505 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_4516 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_4527 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_566 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_566/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_555 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_555/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_544 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_544/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_533 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_533/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4538 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_4549 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3804 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_3815 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_599 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_599/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_588 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_588/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_577 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_577/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_3859 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_3848 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_3826 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_3837 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7120 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7120/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7131 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7131/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_7142 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7142/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_7153 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7153/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_7164 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7164/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_7175 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7175/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_7186 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7186/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_7197 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7197/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_6430 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_6441 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_6452 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6463 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_6474 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_6485 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6496 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_5740 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_5751 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_5762 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_5773 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_5784 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_5795 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1709 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_1709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_5003 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5003/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_5014 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5014/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_5025 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5025/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_5036 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5036/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_5047 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5047/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4302 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_330 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_330/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5058 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5058/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_5069 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5069/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4313 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_4324 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4335 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_374 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_374/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_363 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_363/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_352 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_352/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_341 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_341/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3634 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_3623 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_3612 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_3601 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4346 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_4357 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_4368 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_4379 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_396 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_396/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_385 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_385/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_2922 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_2911 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_2900 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_3667 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3656 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_3645 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2955 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_2944 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_2933 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3689 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3678 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2999 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2988 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_2977 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2966 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_6260 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_6271 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_6282 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_6293 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_5570 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_5581 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_5592 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_4880 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_4891 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2218 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_2207 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_1506 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_2229 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1539 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1528 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1517 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_9814 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9814/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_9803 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9803/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_9847 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9847/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_9836 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9836/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_9825 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9825/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_9858 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9858/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_9869 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9869/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_4110 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4121 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_4132 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_4143 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_182 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_182/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_171 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_171/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_160 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_160/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3442 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3431 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_3420 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_4154 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_4165 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_4176 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_4187 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_193 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_193/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_2730 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_3475 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_3464 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3453 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_4198 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2774 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_2763 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_2752 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2741 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3497 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_3486 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2796 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_2785 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_6090 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6090/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_8409 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_8409/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_7708 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7708/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_7719 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7719/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_2026 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2026/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_2015 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2015/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_2004 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2004/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_1314 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_1303 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_2059 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2059/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_2048 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2048/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_2037 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2037/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1358 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_1347 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_1336 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_1325 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_1369 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_9600 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9600/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9611 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9611/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_9622 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9622/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_8921 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8921/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_8910 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8910/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_9633 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9633/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_9644 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9644/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_9655 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9655/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_9666 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9666/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8954 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8954/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_8943 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8943/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8932 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8932/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_9699 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9699/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_9688 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9688/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_9677 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9677/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8987 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8987/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_8976 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8976/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8965 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8965/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_8998 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8998/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3250 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3283 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_3272 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_3261 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2582 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_2571 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_2560 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_3294 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1870 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2593 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1892 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1881 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_929 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_929/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_918 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_918/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_907 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_907/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8206 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8206/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_8217 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8217/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8228 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8228/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_8239 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8239/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_7505 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7505/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_7516 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7516/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_7527 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7527/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_7538 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7538/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7549 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7549/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_6804 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_6815 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_6826 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_6837 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_6848 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6859 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_1133 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_1122 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_1111 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_1100 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_1166 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_1155 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_1144 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_1199 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_1188 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_1177 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_9441 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9441/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9430 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9430/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9474 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9474/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_9463 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9463/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_9452 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9452/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8762 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8762/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_8751 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8751/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_8740 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8740/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_9496 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9496/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9485 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9485/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8795 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8795/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_8784 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8784/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_8773 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8773/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3091 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3091/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_3080 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3080/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_2390 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_715 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_715/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_704 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_704/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4709 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_4709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_748 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_748/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_737 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_737/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_726 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_726/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_759 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_759/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_8003 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8003/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_8014 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8014/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_8025 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8025/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_8036 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8036/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_8047 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8047/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_8058 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8058/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7302 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7302/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7313 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7313/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_8069 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8069/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_7324 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7324/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_7335 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7335/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_7346 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7346/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_7357 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7357/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6601 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_6612 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_7368 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7368/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_7379 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7379/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_6623 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_6634 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_6645 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5900 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_6656 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_6667 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6678 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5911 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_5922 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_5933 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_6689 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_5944 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_5955 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_5966 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_5977 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_5988 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_5999 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_9282 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9282/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_9271 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9271/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_9260 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9260/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_8581 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8581/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_8570 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8570/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_9293 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9293/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_8592 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8592/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_7880 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7880/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_7891 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7891/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_5207 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_5218 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_5229 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_523 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_523/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_512 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_512/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_501 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_501/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_4506 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_4517 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_4528 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_556 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_556/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_545 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_545/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_534 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_534/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_4539 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_3805 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_3816 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_589 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_589/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_578 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_578/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_567 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_567/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_3849 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_3827 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_3838 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_7110 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7110/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7121 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7121/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_7132 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7132/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_7143 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7143/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_7154 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7154/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_7165 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7165/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6420 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_7176 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7176/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_7187 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7187/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_7198 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7198/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_6431 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_6442 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6453 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_6464 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_6475 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6486 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5730 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_5741 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_5752 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_6497 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_5763 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_5774 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_5785 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_5796 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_9090 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9090/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_90 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_90/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_5004 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5004/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_5015 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5015/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_5026 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5026/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_5037 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5037/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_331 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_331/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_320 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_320/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5048 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5048/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_5059 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5059/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4303 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4314 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_4325 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_4336 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_364 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_364/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_353 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_353/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_342 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_342/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3624 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3613 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_3602 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4347 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_4358 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_4369 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_397 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_397/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_386 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_386/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_375 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_375/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_2923 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_2912 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_2901 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_3657 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_3646 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_3635 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2956 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_2945 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_2934 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_3679 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_3668 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2989 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2978 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_2967 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_6250 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_6261 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_6272 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_6283 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_6294 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_5560 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_5571 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_5582 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_5593 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_4870 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_4881 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_4892 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_2208 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_1507 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_2219 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1529 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_1518 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_9815 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9815/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_9804 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9804/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_9837 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9837/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_9826 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9826/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_9848 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9848/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_9859 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9859/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_4100 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4111 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4122 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_4133 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_4144 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_172 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_172/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_161 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_161/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_150 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_150/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3432 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3421 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_3410 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_4155 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_4166 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_4177 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_194 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_194/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_183 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_183/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_2731 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_2720 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_3476 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_3465 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_3454 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_3443 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_4188 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_4199 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_2764 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_2753 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_2742 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_3498 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_3487 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2797 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_2786 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_2775 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_6080 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6080/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_6091 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6091/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_5390 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_7709 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_7709/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_2027 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2027/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_2016 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2016/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_2005 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2005/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_1315 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_1304 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_2049 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2049/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_2038 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2038/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1348 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_1337 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_1326 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_1359 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_9601 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9601/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9612 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9612/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_9623 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9623/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_8911 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8911/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_8900 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8900/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_9634 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9634/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_9645 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9645/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_9656 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9656/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8955 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8955/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_8944 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8944/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_8933 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8933/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_8922 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8922/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_9689 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9689/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9667 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9667/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_9678 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9678/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8988 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8988/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_8977 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8977/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_8966 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8966/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_8999 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8999/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3251 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3240 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3284 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_3273 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_3262 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2572 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_2561 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_2550 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_3295 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_1871 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_1860 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2594 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_2583 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1893 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_1882 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_919 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_919/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_908 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_908/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8207 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8207/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_8218 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8218/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_8229 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8229/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_7506 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7506/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_7517 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7517/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_7528 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7528/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_7539 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7539/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_6805 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_6816 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_6827 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_6838 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_6849 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1123 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_1112 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_1101 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_1156 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_1145 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_1134 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_1189 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_1178 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_1167 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_9431 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9431/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9420 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9420/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_8730 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8730/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_9464 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9464/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_9453 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9453/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_9442 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9442/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8763 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8763/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_8752 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8752/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_8741 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8741/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_9497 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9497/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9486 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9486/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_9475 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9475/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8796 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8796/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_8785 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8785/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_8774 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8774/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3092 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3092/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_3081 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3081/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_3070 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3070/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2391 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_2380 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_1690 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_705 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_705/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_738 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_738/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_727 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_727/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_716 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_716/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_749 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_749/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_8004 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8004/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_8015 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8015/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_8026 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8026/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_8037 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8037/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_8048 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8048/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_8059 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8059/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_7303 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7303/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7314 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7314/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_7325 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7325/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_7336 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7336/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_7347 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7347/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6602 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_7358 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7358/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_7369 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7369/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_6613 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_6624 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_6635 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5901 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_6646 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_6657 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6668 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_6679 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_5912 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_5923 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_5934 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_5945 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_5956 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_5967 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_5978 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_5989 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_9283 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9283/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_9272 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9272/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_9261 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9261/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_9250 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9250/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_8571 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8571/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_8560 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8560/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_9294 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9294/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_8593 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8593/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_8582 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_8582/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_7870 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7870/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_7881 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7881/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_7892 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_7892/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5208 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_5219 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_5219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_513 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_513/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_502 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_502/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_4507 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_4518 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_557 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_557/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_546 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_546/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_535 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_535/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_524 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_524/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_4529 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_4529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_3806 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_579 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_579/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_568 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_568/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_3817 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_3828 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_3839 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_3839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_7100 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7100/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_7111 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7111/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_7122 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7122/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_7133 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7133/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_7144 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7144/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_7155 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7155/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_6410 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_7166 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7166/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_7177 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7177/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_7188 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7188/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_7199 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_7199/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_6421 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_6432 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_6443 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_6454 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_6465 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_6476 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6487 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_5720 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_5731 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_5742 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_6498 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_6498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_5753 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_5764 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_5775 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_5786 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_5797 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_5797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_9091 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9091/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_9080 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_9080/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_8390 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_8390/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_91 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_91/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_80 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_80/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5005 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5005/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_5016 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5016/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_5027 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5027/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_5038 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5038/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_321 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_321/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_310 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_310/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_5049 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_5049/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4304 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_4315 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_4326 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_365 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_365/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_354 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_354/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_343 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_343/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_332 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_332/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3625 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_3614 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_3603 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_4337 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_4348 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_4359 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_4359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_398 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_398/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_387 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_387/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_376 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_376/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_2913 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_2902 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_3658 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_3647 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_3636 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_2946 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_2935 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_2924 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_3669 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_3669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_2979 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_2968 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_2957 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_2957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_6240 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_6251 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6251/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_6262 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6262/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_6273 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6273/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_6284 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6284/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_6295 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_6295/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_5550 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5550/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_5561 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5561/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_5572 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5572/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_5583 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5583/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_5594 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_5594/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_4860 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4860/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_4871 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4871/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_4882 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4882/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_4893 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_4893/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_2209 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_2209/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_1519 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1519/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_1508 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_1508/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_9805 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9805/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_9838 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9838/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_9827 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9827/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_9816 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9816/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9849 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_9849/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_4101 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4101/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_140 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_140/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3400 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3400/AMP_IN SF_IB pixel_900/PIX_OUT
+ CSA_VREF pixel
Xpixel_4112 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4112/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_4123 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4123/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_4134 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4134/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_173 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_173/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_162 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_162/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_151 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_151/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3433 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3433/AMP_IN SF_IB pixel_33/PIX_OUT
+ CSA_VREF pixel
Xpixel_3422 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3422/AMP_IN SF_IB pixel_22/PIX_OUT
+ CSA_VREF pixel
Xpixel_3411 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3411/AMP_IN SF_IB pixel_11/PIX_OUT
+ CSA_VREF pixel
Xpixel_4145 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4145/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_4156 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4156/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_4167 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4167/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_4178 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4178/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_195 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_195/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_184 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_184/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_2721 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2721/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_2710 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2710/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_3466 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3466/AMP_IN SF_IB pixel_66/PIX_OUT
+ CSA_VREF pixel
Xpixel_3455 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3455/AMP_IN SF_IB pixel_55/PIX_OUT
+ CSA_VREF pixel
Xpixel_3444 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3444/AMP_IN SF_IB pixel_44/PIX_OUT
+ CSA_VREF pixel
Xpixel_4189 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_4189/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_2765 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2765/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_2754 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2754/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_2743 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2743/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_2732 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2732/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_3499 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3499/AMP_IN SF_IB pixel_99/PIX_OUT
+ CSA_VREF pixel
Xpixel_3488 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3488/AMP_IN SF_IB pixel_88/PIX_OUT
+ CSA_VREF pixel
Xpixel_3477 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_3477/AMP_IN SF_IB pixel_77/PIX_OUT
+ CSA_VREF pixel
Xpixel_2798 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2798/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_2787 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2787/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_2776 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_2776/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_6070 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6070/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_6081 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6081/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_6092 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_6092/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_5380 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5380/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_5391 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_5391/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_4690 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_4690/AMP_IN SF_IB pixel_90/PIX_OUT
+ CSA_VREF pixel
Xpixel_2017 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2017/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_2006 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2006/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_1305 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1305/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_2039 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2039/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_2028 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_2028/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_1349 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1349/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_1338 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1338/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_1327 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1327/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_1316 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_1316/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_9602 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9602/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_9613 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9613/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_8912 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8912/AMP_IN SF_IB pixel_12/PIX_OUT
+ CSA_VREF pixel
Xpixel_8901 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8901/AMP_IN SF_IB pixel_901/PIX_OUT
+ CSA_VREF pixel
Xpixel_9624 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9624/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_9635 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9635/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_9646 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9646/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_9657 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9657/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_8945 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8945/AMP_IN SF_IB pixel_45/PIX_OUT
+ CSA_VREF pixel
Xpixel_8934 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8934/AMP_IN SF_IB pixel_34/PIX_OUT
+ CSA_VREF pixel
Xpixel_8923 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8923/AMP_IN SF_IB pixel_23/PIX_OUT
+ CSA_VREF pixel
Xpixel_9668 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9668/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9679 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_9679/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_8978 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8978/AMP_IN SF_IB pixel_78/PIX_OUT
+ CSA_VREF pixel
Xpixel_8967 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8967/AMP_IN SF_IB pixel_67/PIX_OUT
+ CSA_VREF pixel
Xpixel_8956 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8956/AMP_IN SF_IB pixel_56/PIX_OUT
+ CSA_VREF pixel
Xpixel_8989 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_8989/AMP_IN SF_IB pixel_89/PIX_OUT
+ CSA_VREF pixel
Xpixel_3241 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3241/AMP_IN SF_IB pixel_41/PIX_OUT
+ CSA_VREF pixel
Xpixel_3230 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3230/AMP_IN SF_IB pixel_30/PIX_OUT
+ CSA_VREF pixel
Xpixel_2540 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2540/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
Xpixel_3274 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3274/AMP_IN SF_IB pixel_74/PIX_OUT
+ CSA_VREF pixel
Xpixel_3263 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3263/AMP_IN SF_IB pixel_63/PIX_OUT
+ CSA_VREF pixel
Xpixel_3252 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3252/AMP_IN SF_IB pixel_52/PIX_OUT
+ CSA_VREF pixel
Xpixel_2573 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2573/AMP_IN SF_IB pixel_73/PIX_OUT
+ CSA_VREF pixel
Xpixel_2562 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2562/AMP_IN SF_IB pixel_62/PIX_OUT
+ CSA_VREF pixel
Xpixel_2551 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2551/AMP_IN SF_IB pixel_51/PIX_OUT
+ CSA_VREF pixel
Xpixel_3296 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3296/AMP_IN SF_IB pixel_96/PIX_OUT
+ CSA_VREF pixel
Xpixel_3285 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_3285/AMP_IN SF_IB pixel_85/PIX_OUT
+ CSA_VREF pixel
Xpixel_1861 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1861/AMP_IN SF_IB pixel_61/PIX_OUT
+ CSA_VREF pixel
Xpixel_1850 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1850/AMP_IN SF_IB pixel_50/PIX_OUT
+ CSA_VREF pixel
Xpixel_2595 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2595/AMP_IN SF_IB pixel_95/PIX_OUT
+ CSA_VREF pixel
Xpixel_2584 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_2584/AMP_IN SF_IB pixel_84/PIX_OUT
+ CSA_VREF pixel
Xpixel_1894 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1894/AMP_IN SF_IB pixel_94/PIX_OUT
+ CSA_VREF pixel
Xpixel_1883 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1883/AMP_IN SF_IB pixel_83/PIX_OUT
+ CSA_VREF pixel
Xpixel_1872 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_1872/AMP_IN SF_IB pixel_72/PIX_OUT
+ CSA_VREF pixel
Xpixel_909 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_909/AMP_IN SF_IB pixel_9/PIX_OUT
+ CSA_VREF pixel
Xpixel_8208 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8208/AMP_IN SF_IB pixel_8/PIX_OUT
+ CSA_VREF pixel
Xpixel_8219 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_8219/AMP_IN SF_IB pixel_19/PIX_OUT
+ CSA_VREF pixel
Xpixel_7507 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7507/AMP_IN SF_IB pixel_7/PIX_OUT
+ CSA_VREF pixel
Xpixel_7518 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7518/AMP_IN SF_IB pixel_18/PIX_OUT
+ CSA_VREF pixel
Xpixel_7529 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_7529/AMP_IN SF_IB pixel_29/PIX_OUT
+ CSA_VREF pixel
Xpixel_6806 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6806/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_6817 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6817/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_6828 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6828/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_6839 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_6839/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_1124 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1124/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_1113 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1113/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_1102 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1102/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_1157 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1157/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_1146 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1146/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_1135 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1135/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_1179 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1179/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_1168 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_1168/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_9432 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9432/AMP_IN SF_IB pixel_32/PIX_OUT
+ CSA_VREF pixel
Xpixel_9421 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9421/AMP_IN SF_IB pixel_21/PIX_OUT
+ CSA_VREF pixel
Xpixel_9410 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9410/AMP_IN SF_IB pixel_10/PIX_OUT
+ CSA_VREF pixel
Xpixel_8720 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8720/AMP_IN SF_IB pixel_20/PIX_OUT
+ CSA_VREF pixel
Xpixel_9465 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9465/AMP_IN SF_IB pixel_65/PIX_OUT
+ CSA_VREF pixel
Xpixel_9454 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9454/AMP_IN SF_IB pixel_54/PIX_OUT
+ CSA_VREF pixel
Xpixel_9443 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9443/AMP_IN SF_IB pixel_43/PIX_OUT
+ CSA_VREF pixel
Xpixel_8753 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8753/AMP_IN SF_IB pixel_53/PIX_OUT
+ CSA_VREF pixel
Xpixel_8742 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8742/AMP_IN SF_IB pixel_42/PIX_OUT
+ CSA_VREF pixel
Xpixel_8731 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8731/AMP_IN SF_IB pixel_31/PIX_OUT
+ CSA_VREF pixel
Xpixel_9498 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9498/AMP_IN SF_IB pixel_98/PIX_OUT
+ CSA_VREF pixel
Xpixel_9487 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9487/AMP_IN SF_IB pixel_87/PIX_OUT
+ CSA_VREF pixel
Xpixel_9476 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_9476/AMP_IN SF_IB pixel_76/PIX_OUT
+ CSA_VREF pixel
Xpixel_8797 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8797/AMP_IN SF_IB pixel_97/PIX_OUT
+ CSA_VREF pixel
Xpixel_8786 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8786/AMP_IN SF_IB pixel_86/PIX_OUT
+ CSA_VREF pixel
Xpixel_8775 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8775/AMP_IN SF_IB pixel_75/PIX_OUT
+ CSA_VREF pixel
Xpixel_8764 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_8764/AMP_IN SF_IB pixel_64/PIX_OUT
+ CSA_VREF pixel
Xpixel_3093 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3093/AMP_IN SF_IB pixel_93/PIX_OUT
+ CSA_VREF pixel
Xpixel_3082 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3082/AMP_IN SF_IB pixel_82/PIX_OUT
+ CSA_VREF pixel
Xpixel_3071 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3071/AMP_IN SF_IB pixel_71/PIX_OUT
+ CSA_VREF pixel
Xpixel_3060 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_3060/AMP_IN SF_IB pixel_60/PIX_OUT
+ CSA_VREF pixel
Xpixel_2381 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2381/AMP_IN SF_IB pixel_81/PIX_OUT
+ CSA_VREF pixel
Xpixel_2370 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2370/AMP_IN SF_IB pixel_70/PIX_OUT
+ CSA_VREF pixel
Xpixel_2392 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_2392/AMP_IN SF_IB pixel_92/PIX_OUT
+ CSA_VREF pixel
Xpixel_1691 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1691/AMP_IN SF_IB pixel_91/PIX_OUT
+ CSA_VREF pixel
Xpixel_1680 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_1680/AMP_IN SF_IB pixel_80/PIX_OUT
+ CSA_VREF pixel
Xpixel_706 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_706/AMP_IN SF_IB pixel_6/PIX_OUT
+ CSA_VREF pixel
Xpixel_739 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_739/AMP_IN SF_IB pixel_39/PIX_OUT
+ CSA_VREF pixel
Xpixel_728 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_728/AMP_IN SF_IB pixel_28/PIX_OUT
+ CSA_VREF pixel
Xpixel_717 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_717/AMP_IN SF_IB pixel_17/PIX_OUT
+ CSA_VREF pixel
Xpixel_8005 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8005/AMP_IN SF_IB pixel_5/PIX_OUT
+ CSA_VREF pixel
Xpixel_8016 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8016/AMP_IN SF_IB pixel_16/PIX_OUT
+ CSA_VREF pixel
Xpixel_8027 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8027/AMP_IN SF_IB pixel_27/PIX_OUT
+ CSA_VREF pixel
Xpixel_8038 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8038/AMP_IN SF_IB pixel_38/PIX_OUT
+ CSA_VREF pixel
Xpixel_8049 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_8049/AMP_IN SF_IB pixel_49/PIX_OUT
+ CSA_VREF pixel
Xpixel_7304 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7304/AMP_IN SF_IB pixel_4/PIX_OUT
+ CSA_VREF pixel
Xpixel_7315 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7315/AMP_IN SF_IB pixel_15/PIX_OUT
+ CSA_VREF pixel
Xpixel_7326 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7326/AMP_IN SF_IB pixel_26/PIX_OUT
+ CSA_VREF pixel
Xpixel_7337 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7337/AMP_IN SF_IB pixel_37/PIX_OUT
+ CSA_VREF pixel
Xpixel_7348 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7348/AMP_IN SF_IB pixel_48/PIX_OUT
+ CSA_VREF pixel
Xpixel_6603 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6603/AMP_IN SF_IB pixel_3/PIX_OUT
+ CSA_VREF pixel
Xpixel_7359 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_7359/AMP_IN SF_IB pixel_59/PIX_OUT
+ CSA_VREF pixel
Xpixel_6614 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6614/AMP_IN SF_IB pixel_14/PIX_OUT
+ CSA_VREF pixel
Xpixel_6625 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6625/AMP_IN SF_IB pixel_25/PIX_OUT
+ CSA_VREF pixel
Xpixel_6636 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6636/AMP_IN SF_IB pixel_36/PIX_OUT
+ CSA_VREF pixel
Xpixel_6647 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6647/AMP_IN SF_IB pixel_47/PIX_OUT
+ CSA_VREF pixel
Xpixel_6658 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6658/AMP_IN SF_IB pixel_58/PIX_OUT
+ CSA_VREF pixel
Xpixel_6669 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_6669/AMP_IN SF_IB pixel_69/PIX_OUT
+ CSA_VREF pixel
Xpixel_5902 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5902/AMP_IN SF_IB pixel_2/PIX_OUT
+ CSA_VREF pixel
Xpixel_5913 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5913/AMP_IN SF_IB pixel_13/PIX_OUT
+ CSA_VREF pixel
Xpixel_5924 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5924/AMP_IN SF_IB pixel_24/PIX_OUT
+ CSA_VREF pixel
Xpixel_5935 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5935/AMP_IN SF_IB pixel_35/PIX_OUT
+ CSA_VREF pixel
Xpixel_5946 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5946/AMP_IN SF_IB pixel_46/PIX_OUT
+ CSA_VREF pixel
Xpixel_5957 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5957/AMP_IN SF_IB pixel_57/PIX_OUT
+ CSA_VREF pixel
Xpixel_5968 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5968/AMP_IN SF_IB pixel_68/PIX_OUT
+ CSA_VREF pixel
Xpixel_5979 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_5979/AMP_IN SF_IB pixel_79/PIX_OUT
+ CSA_VREF pixel
Xpixel_9240 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_9240/AMP_IN SF_IB pixel_40/PIX_OUT
+ CSA_VREF pixel
X0 pixel_83/PIX_OUT COL_SEL[83] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X1 pixel_79/PIX_OUT COL_SEL[79] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X2 pixel_75/PIX_OUT COL_SEL[75] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X3 pixel_71/PIX_OUT COL_SEL[71] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X4 pixel_67/PIX_OUT COL_SEL[67] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X5 pixel_26/PIX_OUT COL_SEL[26] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X6 pixel_64/PIX_OUT COL_SEL[64] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X7 pixel_22/PIX_OUT COL_SEL[22] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X8 pixel_18/PIX_OUT COL_SEL[18] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X9 pixel_60/PIX_OUT COL_SEL[60] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X10 pixel_14/PIX_OUT COL_SEL[14] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X11 pixel_10/PIX_OUT COL_SEL[10] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X12 pixel_86/PIX_OUT COL_SEL[86] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X13 pixel_82/PIX_OUT COL_SEL[82] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X14 pixel_78/PIX_OUT COL_SEL[78] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X15 pixel_74/PIX_OUT COL_SEL[74] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X16 pixel_70/PIX_OUT COL_SEL[70] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X17 pixel_33/PIX_OUT COL_SEL[33] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X18 pixel_29/PIX_OUT COL_SEL[29] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X19 pixel_25/PIX_OUT COL_SEL[25] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X20 pixel_21/PIX_OUT COL_SEL[21] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X21 pixel_17/PIX_OUT COL_SEL[17] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X22 pixel_93/PIX_OUT COL_SEL[93] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X23 pixel_89/PIX_OUT COL_SEL[89] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X24 pixel_85/PIX_OUT COL_SEL[85] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X25 pixel_81/PIX_OUT COL_SEL[81] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X26 pixel_77/PIX_OUT COL_SEL[77] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X27 pixel_36/PIX_OUT COL_SEL[36] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X28 pixel_32/PIX_OUT COL_SEL[32] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X29 pixel_28/PIX_OUT COL_SEL[28] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X30 pixel_24/PIX_OUT COL_SEL[24] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X31 pixel_20/PIX_OUT COL_SEL[20] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X32 pixel_3/PIX_OUT COL_SEL[3] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X33 pixel_96/PIX_OUT COL_SEL[96] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X34 pixel_92/PIX_OUT COL_SEL[92] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X35 pixel_88/PIX_OUT COL_SEL[88] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X36 pixel_84/PIX_OUT COL_SEL[84] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X37 pixel_80/PIX_OUT COL_SEL[80] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X38 pixel_43/PIX_OUT COL_SEL[43] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X39 pixel_900/PIX_OUT COL_SEL[0] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X40 pixel_39/PIX_OUT COL_SEL[39] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X41 pixel_35/PIX_OUT COL_SEL[35] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X42 pixel_31/PIX_OUT COL_SEL[31] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X43 pixel_27/PIX_OUT COL_SEL[27] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X44 pixel_2/PIX_OUT COL_SEL[2] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X45 pixel_99/PIX_OUT COL_SEL[99] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X46 pixel_95/PIX_OUT COL_SEL[95] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X47 pixel_91/PIX_OUT COL_SEL[91] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X48 pixel_87/PIX_OUT COL_SEL[87] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X49 pixel_46/PIX_OUT COL_SEL[46] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X50 pixel_42/PIX_OUT COL_SEL[42] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X51 pixel_38/PIX_OUT COL_SEL[38] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X52 pixel_34/PIX_OUT COL_SEL[34] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X53 pixel_30/PIX_OUT COL_SEL[30] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X54 pixel_901/PIX_OUT COL_SEL[1] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X55 pixel_98/PIX_OUT COL_SEL[98] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X56 pixel_94/PIX_OUT COL_SEL[94] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X57 pixel_90/PIX_OUT COL_SEL[90] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X58 pixel_53/PIX_OUT COL_SEL[53] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X59 pixel_49/PIX_OUT COL_SEL[49] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X60 pixel_45/PIX_OUT COL_SEL[45] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X61 pixel_41/PIX_OUT COL_SEL[41] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X62 pixel_37/PIX_OUT COL_SEL[37] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X63 pixel_97/PIX_OUT COL_SEL[97] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X64 pixel_56/PIX_OUT COL_SEL[56] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X65 pixel_52/PIX_OUT COL_SEL[52] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X66 pixel_6/PIX_OUT COL_SEL[6] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X67 pixel_48/PIX_OUT COL_SEL[48] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X68 pixel_44/PIX_OUT COL_SEL[44] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X69 pixel_40/PIX_OUT COL_SEL[40] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X70 pixel_63/PIX_OUT COL_SEL[63] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X71 pixel_59/PIX_OUT COL_SEL[59] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X72 pixel_55/PIX_OUT COL_SEL[55] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X73 pixel_13/PIX_OUT COL_SEL[13] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X74 pixel_9/PIX_OUT COL_SEL[9] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X75 pixel_51/PIX_OUT COL_SEL[51] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X76 pixel_5/PIX_OUT COL_SEL[5] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X77 pixel_47/PIX_OUT COL_SEL[47] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X78 pixel_73/PIX_OUT COL_SEL[73] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X79 pixel_69/PIX_OUT COL_SEL[69] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X80 pixel_66/PIX_OUT COL_SEL[66] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X81 pixel_62/PIX_OUT COL_SEL[62] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X82 pixel_16/PIX_OUT COL_SEL[16] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X83 pixel_12/PIX_OUT COL_SEL[12] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X84 pixel_58/PIX_OUT COL_SEL[58] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X85 pixel_54/PIX_OUT COL_SEL[54] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X86 pixel_8/PIX_OUT COL_SEL[8] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X87 pixel_50/PIX_OUT COL_SEL[50] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X88 pixel_4/PIX_OUT COL_SEL[4] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X89 pixel_76/PIX_OUT COL_SEL[76] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X90 pixel_72/PIX_OUT COL_SEL[72] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X91 pixel_68/PIX_OUT COL_SEL[68] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X92 pixel_23/PIX_OUT COL_SEL[23] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X93 pixel_19/PIX_OUT COL_SEL[19] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X94 pixel_65/PIX_OUT COL_SEL[65] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X95 pixel_61/PIX_OUT COL_SEL[61] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X96 pixel_15/PIX_OUT COL_SEL[15] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X97 pixel_11/PIX_OUT COL_SEL[11] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X98 pixel_57/PIX_OUT COL_SEL[57] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X99 pixel_7/PIX_OUT COL_SEL[7] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt shift_registerC COL_SEL[0] COL_SEL[10] COL_SEL[11] COL_SEL[12] COL_SEL[13]
+ COL_SEL[14] COL_SEL[15] COL_SEL[16] COL_SEL[17] COL_SEL[18] COL_SEL[19] COL_SEL[1]
+ COL_SEL[20] COL_SEL[21] COL_SEL[22] COL_SEL[23] COL_SEL[24] COL_SEL[25] COL_SEL[26]
+ COL_SEL[27] COL_SEL[28] COL_SEL[29] COL_SEL[2] COL_SEL[30] COL_SEL[31] COL_SEL[32]
+ COL_SEL[33] COL_SEL[34] COL_SEL[35] COL_SEL[36] COL_SEL[37] COL_SEL[38] COL_SEL[39]
+ COL_SEL[3] COL_SEL[40] COL_SEL[41] COL_SEL[42] COL_SEL[43] COL_SEL[44] COL_SEL[45]
+ COL_SEL[46] COL_SEL[47] COL_SEL[48] COL_SEL[49] COL_SEL[4] COL_SEL[50] COL_SEL[51]
+ COL_SEL[52] COL_SEL[53] COL_SEL[54] COL_SEL[55] COL_SEL[56] COL_SEL[57] COL_SEL[58]
+ COL_SEL[59] COL_SEL[5] COL_SEL[60] COL_SEL[61] COL_SEL[62] COL_SEL[63] COL_SEL[64]
+ COL_SEL[65] COL_SEL[66] COL_SEL[67] COL_SEL[68] COL_SEL[69] COL_SEL[6] COL_SEL[70]
+ COL_SEL[71] COL_SEL[72] COL_SEL[73] COL_SEL[74] COL_SEL[75] COL_SEL[76] COL_SEL[77]
+ COL_SEL[78] COL_SEL[79] COL_SEL[7] COL_SEL[80] COL_SEL[81] COL_SEL[82] COL_SEL[83]
+ COL_SEL[84] COL_SEL[85] COL_SEL[86] COL_SEL[87] COL_SEL[88] COL_SEL[89] COL_SEL[8]
+ COL_SEL[90] COL_SEL[91] COL_SEL[92] COL_SEL[93] COL_SEL[94] COL_SEL[95] COL_SEL[96]
+ COL_SEL[97] COL_SEL[98] COL_SEL[99] COL_SEL[9] clk data_in data_out ena rst VDD
+ GND
XFILLER_3_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_501_ _727_/Q _726_/Q _503_/S GND GND VDD VDD _502_/A sky130_fd_sc_hd__mux2_1
X_432_ _758_/Q _757_/Q _436_/S GND GND VDD VDD _433_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_363_ _789_/Q _788_/Q _369_/S GND GND VDD VDD _364_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2524 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2629 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1730 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_648 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_415_ _415_/A GND GND VDD VDD _766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3011 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3044 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_2310 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3105 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_3077 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_2343 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1620 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1653 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2993 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1368 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1357 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_7_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_556 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2151 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_220 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_669 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_1_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_680_ _683_/A GND GND VDD VDD _680_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1110 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_1154 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_397 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2220 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2097 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1341 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_732_ _773_/CLK _732_/D _618_/Y GND GND VDD VDD _732_/Q sky130_fd_sc_hd__dfrtp_1
X_663_ _664_/A GND GND VDD VDD _663_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_594_ _596_/A GND GND VDD VDD _594_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_868 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_5 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_3_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1625 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2094 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_359 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2871 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput42 _719_/Q GND GND VDD VDD COL_SEL[44] sky130_fd_sc_hd__clkbuf_1
Xoutput31 _709_/Q GND GND VDD VDD COL_SEL[34] sky130_fd_sc_hd__clkbuf_1
Xoutput20 _699_/Q GND GND VDD VDD COL_SEL[24] sky130_fd_sc_hd__clkbuf_1
Xoutput7 _787_/Q GND GND VDD VDD COL_SEL[12] sky130_fd_sc_hd__clkbuf_1
Xoutput64 _739_/Q GND GND VDD VDD COL_SEL[64] sky130_fd_sc_hd__clkbuf_1
Xoutput53 _729_/Q GND GND VDD VDD COL_SEL[54] sky130_fd_sc_hd__clkbuf_1
Xoutput75 _749_/Q GND GND VDD VDD COL_SEL[74] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput97 _769_/Q GND GND VDD VDD COL_SEL[94] sky130_fd_sc_hd__clkbuf_1
Xoutput86 _759_/Q GND GND VDD VDD COL_SEL[84] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_715_ _795_/CLK _715_/D _596_/Y GND GND VDD VDD _715_/Q sky130_fd_sc_hd__dfrtp_1
X_646_ _646_/A GND GND VDD VDD _646_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_577_ _578_/A GND GND VDD VDD _577_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2657 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_808 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1709 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2189 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_500_ _500_/A GND GND VDD VDD _728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_431_ _431_/A GND GND VDD VDD _759_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_6__f_clk clkbuf_0_clk/X GND GND VDD VDD _775_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_362_ _362_/A GND GND VDD VDD _790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1802 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_963 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1929 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_629_ _633_/A GND GND VDD VDD _629_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1786 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2885 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_414_ _766_/Q _765_/Q _414_/S GND GND VDD VDD _415_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2405 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_2377 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1676 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_281 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_579 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2163 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1509 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_276 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1166 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_8_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_332 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2508 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2232 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_15_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1397 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_445 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_731_ _773_/CLK _731_/D _617_/Y GND GND VDD VDD _731_/Q sky130_fd_sc_hd__dfrtp_1
X_662_ _664_/A GND GND VDD VDD _662_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_836 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_593_ _596_/A GND GND VDD VDD _593_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2585 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_8_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_6 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_3_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput43 _720_/Q GND GND VDD VDD COL_SEL[45] sky130_fd_sc_hd__clkbuf_1
Xoutput32 _710_/Q GND GND VDD VDD COL_SEL[35] sky130_fd_sc_hd__clkbuf_1
Xoutput10 _790_/Q GND GND VDD VDD COL_SEL[15] sky130_fd_sc_hd__clkbuf_1
Xoutput21 _700_/Q GND GND VDD VDD COL_SEL[25] sky130_fd_sc_hd__clkbuf_1
Xoutput8 _788_/Q GND GND VDD VDD COL_SEL[13] sky130_fd_sc_hd__clkbuf_1
Xoutput76 _750_/Q GND GND VDD VDD COL_SEL[75] sky130_fd_sc_hd__clkbuf_1
Xoutput65 _740_/Q GND GND VDD VDD COL_SEL[65] sky130_fd_sc_hd__clkbuf_1
Xoutput54 _730_/Q GND GND VDD VDD COL_SEL[55] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput98 _770_/Q GND GND VDD VDD COL_SEL[95] sky130_fd_sc_hd__clkbuf_1
Xoutput87 _760_/Q GND GND VDD VDD COL_SEL[85] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_714_ _786_/CLK _714_/D _595_/Y GND GND VDD VDD _714_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_611 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_645_ _646_/A GND GND VDD VDD _645_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_576_ _578_/A GND GND VDD VDD _576_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2124 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1401 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1423 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_430_ _759_/Q _758_/Q _436_/S GND GND VDD VDD _431_/A sky130_fd_sc_hd__mux2_1
X_361_ _790_/Q _789_/Q _369_/S GND GND VDD VDD _362_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_920 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_628_ _628_/A GND GND VDD VDD _633_/A sky130_fd_sc_hd__buf_2
XFILLER_18_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_559_ _701_/Q _700_/Q _559_/S GND GND VDD VDD _560_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2488 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_413_ _413_/A GND GND VDD VDD _767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2797 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1705 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_293 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2049 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_981 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3273 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2572 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1893 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2082 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2756 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_388 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_377 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_730_ _774_/CLK _730_/D _615_/Y GND GND VDD VDD _730_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_661_ _664_/A GND GND VDD VDD _661_/Y sky130_fd_sc_hd__inv_2
X_592_ _596_/A GND GND VDD VDD _592_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2807 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_7 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_3_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1173 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_13_317 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_2895 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput33 _711_/Q GND GND VDD VDD COL_SEL[36] sky130_fd_sc_hd__clkbuf_1
Xoutput22 _701_/Q GND GND VDD VDD COL_SEL[26] sky130_fd_sc_hd__clkbuf_1
Xoutput11 _791_/Q GND GND VDD VDD COL_SEL[16] sky130_fd_sc_hd__clkbuf_1
Xoutput9 _789_/Q GND GND VDD VDD COL_SEL[14] sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput55 _731_/Q GND GND VDD VDD COL_SEL[56] sky130_fd_sc_hd__clkbuf_1
Xoutput44 _721_/Q GND GND VDD VDD COL_SEL[46] sky130_fd_sc_hd__clkbuf_1
Xoutput66 _741_/Q GND GND VDD VDD COL_SEL[66] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput99 _771_/Q GND GND VDD VDD COL_SEL[96] sky130_fd_sc_hd__clkbuf_1
Xoutput77 _751_/Q GND GND VDD VDD COL_SEL[76] sky130_fd_sc_hd__clkbuf_1
Xoutput88 _761_/Q GND GND VDD VDD COL_SEL[86] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_713_ _786_/CLK _713_/D _594_/Y GND GND VDD VDD _713_/Q sky130_fd_sc_hd__dfrtp_1
X_644_ _646_/A GND GND VDD VDD _644_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_575_ _578_/A GND GND VDD VDD _575_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2615 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1903 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3285 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_409 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2946 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_360_ _393_/A GND GND VDD VDD _369_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_910 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_627_ _627_/A GND GND VDD VDD _627_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_558_ _558_/A GND GND VDD VDD _702_/D sky130_fd_sc_hd__clkbuf_1
X_489_ _489_/A GND GND VDD VDD _733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1243 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1254 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2710 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_412_ _767_/Q _766_/Q _414_/S GND GND VDD VDD _413_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_809 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2880 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2176 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2237 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2735 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2768 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1261 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_660_ _664_/A GND GND VDD VDD _660_/Y sky130_fd_sc_hd__inv_2
X_591_ _597_/A GND GND VDD VDD _596_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_827 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_304 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2819 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2598 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_8 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_10_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_789_ _791_/CLK _789_/D _688_/Y GND GND VDD VDD _789_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2031 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2086 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1116 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput34 _712_/Q GND GND VDD VDD COL_SEL[37] sky130_fd_sc_hd__clkbuf_1
Xoutput23 _702_/Q GND GND VDD VDD COL_SEL[27] sky130_fd_sc_hd__clkbuf_1
Xoutput12 _792_/Q GND GND VDD VDD COL_SEL[17] sky130_fd_sc_hd__clkbuf_1
Xoutput67 _742_/Q GND GND VDD VDD COL_SEL[67] sky130_fd_sc_hd__clkbuf_1
Xoutput45 _722_/Q GND GND VDD VDD COL_SEL[47] sky130_fd_sc_hd__clkbuf_1
Xoutput56 _732_/Q GND GND VDD VDD COL_SEL[57] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput78 _752_/Q GND GND VDD VDD COL_SEL[77] sky130_fd_sc_hd__clkbuf_1
Xoutput89 _762_/Q GND GND VDD VDD COL_SEL[87] sky130_fd_sc_hd__clkbuf_1
XFILLER_20_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_277 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_712_ _791_/CLK _712_/D _593_/Y GND GND VDD VDD _712_/Q sky130_fd_sc_hd__dfrtp_1
X_643_ _646_/A GND GND VDD VDD _643_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_574_ _578_/A GND GND VDD VDD _574_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2638 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_626_ _627_/A GND GND VDD VDD _626_/Y sky130_fd_sc_hd__inv_2
X_557_ _702_/Q _701_/Q _559_/S GND GND VDD VDD _558_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1745 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_488_ _733_/Q _732_/Q _492_/S GND GND VDD VDD _489_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_2181 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_411_ _411_/A GND GND VDD VDD _768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3037 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_609_ _609_/A GND GND VDD VDD _609_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2265 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_416 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1597 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_1586 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2007 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1537 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_1476 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2051 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2040 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2095 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_780 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_357 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2013 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1284 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_590_ _590_/A GND GND VDD VDD _590_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_9 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_10_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_8 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_788_ _792_/CLK _788_/D _687_/Y GND GND VDD VDD _788_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2043 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2076 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2864 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1128 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput24 _703_/Q GND GND VDD VDD COL_SEL[28] sky130_fd_sc_hd__clkbuf_1
Xoutput13 _793_/Q GND GND VDD VDD COL_SEL[18] sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput46 _723_/Q GND GND VDD VDD COL_SEL[48] sky130_fd_sc_hd__clkbuf_1
Xoutput35 _713_/Q GND GND VDD VDD COL_SEL[38] sky130_fd_sc_hd__clkbuf_1
Xoutput57 _733_/Q GND GND VDD VDD COL_SEL[58] sky130_fd_sc_hd__clkbuf_1
Xoutput68 _743_/Q GND GND VDD VDD COL_SEL[68] sky130_fd_sc_hd__clkbuf_1
Xoutput79 _753_/Q GND GND VDD VDD COL_SEL[78] sky130_fd_sc_hd__clkbuf_1
X_711_ _786_/CLK _711_/D _592_/Y GND GND VDD VDD _711_/Q sky130_fd_sc_hd__dfrtp_1
X_642_ _646_/A GND GND VDD VDD _642_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_573_ _597_/A GND GND VDD VDD _578_/A sky130_fd_sc_hd__buf_2
XFILLER_18_1916 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_1__f_clk clkbuf_0_clk/X GND GND VDD VDD _795_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1415 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2904 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_2959 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_13_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_956 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_444 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_625_ _627_/A GND GND VDD VDD _625_/Y sky130_fd_sc_hd__inv_2
X_556_ _556_/A GND GND VDD VDD _703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1702 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_487_ _487_/A GND GND VDD VDD _734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2723 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_410_ _768_/Q _767_/Q _414_/S GND GND VDD VDD _411_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_2778 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_3005 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_1_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2337 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1625 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_608_ _609_/A GND GND VDD VDD _608_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_539_ _561_/A GND GND VDD VDD _548_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1565 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2965 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1885 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1373 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_2940 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1513 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2069 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1313 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_818 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_787_ _795_/CLK _787_/D _686_/Y GND GND VDD VDD _787_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2055 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1093 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput25 _704_/Q GND GND VDD VDD COL_SEL[29] sky130_fd_sc_hd__clkbuf_1
Xoutput14 _794_/Q GND GND VDD VDD COL_SEL[19] sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput58 _734_/Q GND GND VDD VDD COL_SEL[59] sky130_fd_sc_hd__clkbuf_1
Xoutput36 _714_/Q GND GND VDD VDD COL_SEL[39] sky130_fd_sc_hd__clkbuf_1
Xoutput47 _724_/Q GND GND VDD VDD COL_SEL[49] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput69 _744_/Q GND GND VDD VDD COL_SEL[69] sky130_fd_sc_hd__clkbuf_1
X_710_ _792_/CLK _710_/D _590_/Y GND GND VDD VDD _710_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_641_ _659_/A GND GND VDD VDD _646_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_604 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_572_ _665_/A GND GND VDD VDD _597_/A sky130_fd_sc_hd__buf_2
XFILLER_16_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1630 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2117 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XPHY_0 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_624_ _627_/A GND GND VDD VDD _624_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_555_ _703_/Q _702_/Q _559_/S GND GND VDD VDD _556_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_486_ _734_/Q _733_/Q _492_/S GND GND VDD VDD _487_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1758 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1268 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1648 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_607_ _609_/A GND GND VDD VDD _607_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_538_ _538_/A GND GND VDD VDD _711_/D sky130_fd_sc_hd__clkbuf_1
X_469_ _469_/A GND GND VDD VDD _742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2919 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1087 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2565 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2124 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_2157 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_1401 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_584 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2952 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2741 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2749 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1369 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_2760 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_417 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_786_ _786_/CLK _786_/D _685_/Y GND GND VDD VDD _786_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_340 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2170 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput15 _776_/Q GND GND VDD VDD COL_SEL[1] sky130_fd_sc_hd__clkbuf_1
Xoutput48 _779_/Q GND GND VDD VDD COL_SEL[4] sky130_fd_sc_hd__clkbuf_1
Xoutput37 _778_/Q GND GND VDD VDD COL_SEL[3] sky130_fd_sc_hd__clkbuf_1
Xoutput26 _777_/Q GND GND VDD VDD COL_SEL[2] sky130_fd_sc_hd__clkbuf_1
Xoutput59 _780_/Q GND GND VDD VDD COL_SEL[5] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_4_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_640_ _640_/A GND GND VDD VDD _640_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_571_ _571_/A GND GND VDD VDD _696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1642 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_781 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_769_ _771_/CLK _769_/D _663_/Y GND GND VDD VDD _769_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_1 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1940 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_623_ _627_/A GND GND VDD VDD _623_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_936 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_554_ _554_/A GND GND VDD VDD _704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_485_ _485_/A GND GND VDD VDD _735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2195 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_980 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2950 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2736 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_606_ _609_/A GND GND VDD VDD _606_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_537_ _711_/Q _710_/Q _537_/S GND GND VDD VDD _538_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2202 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2257 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_468_ _742_/Q _741_/Q _470_/S GND GND VDD VDD _469_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1578 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_399_ _399_/A GND GND VDD VDD _773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_920 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2577 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1424 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_clk clkbuf_0_clk/X GND GND VDD VDD _773_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_249 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_2964 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2797 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_360 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_1298 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2772 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3273 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_785_ _792_/CLK _785_/D _683_/Y GND GND VDD VDD _785_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2068 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1145 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1109 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput49 _725_/Q GND GND VDD VDD COL_SEL[50] sky130_fd_sc_hd__clkbuf_1
Xoutput38 _715_/Q GND GND VDD VDD COL_SEL[40] sky130_fd_sc_hd__clkbuf_1
Xoutput27 _705_/Q GND GND VDD VDD COL_SEL[30] sky130_fd_sc_hd__clkbuf_1
Xoutput16 _795_/Q GND GND VDD VDD COL_SEL[20] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_570_ _696_/Q _795_/Q _570_/S GND GND VDD VDD _571_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2090 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_10_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_768_ _775_/CLK _768_/D _662_/Y GND GND VDD VDD _768_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_699_ _786_/CLK _699_/D _577_/Y GND GND VDD VDD _699_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk GND GND VDD VDD clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_15_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_622_ _628_/A GND GND VDD VDD _627_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_553_ _704_/Q _703_/Q _559_/S GND GND VDD VDD _554_/A sky130_fd_sc_hd__mux2_1
X_484_ _735_/Q _734_/Q _492_/S GND GND VDD VDD _485_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_992 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2962 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2494 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1782 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_5_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_605_ _609_/A GND GND VDD VDD _605_/Y sky130_fd_sc_hd__inv_2
X_536_ _536_/A GND GND VDD VDD _712_/D sky130_fd_sc_hd__clkbuf_1
X_467_ _467_/A GND GND VDD VDD _743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_398_ _773_/Q _772_/Q _402_/S GND GND VDD VDD _399_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2852 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2100 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2209 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1469 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_519_ _519_/A GND GND VDD VDD _720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1387 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1970 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2729 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1200 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_851 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1233 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_394 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2784 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_29 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_1_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2573 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_784_ _795_/CLK _784_/D _682_/Y GND GND VDD VDD _784_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_865 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2857 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput39 _716_/Q GND GND VDD VDD COL_SEL[41] sky130_fd_sc_hd__clkbuf_1
Xoutput28 _706_/Q GND GND VDD VDD COL_SEL[31] sky130_fd_sc_hd__clkbuf_1
Xoutput17 _696_/Q GND GND VDD VDD COL_SEL[21] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_249 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1677 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_767_ _771_/CLK _767_/D _661_/Y GND GND VDD VDD _767_/Q sky130_fd_sc_hd__dfrtp_1
X_698_ _795_/CLK _698_/D _576_/Y GND GND VDD VDD _698_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_621_ _621_/A GND GND VDD VDD _621_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_949 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_437 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_415 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_552_ _552_/A GND GND VDD VDD _705_/D sky130_fd_sc_hd__clkbuf_1
X_483_ _505_/A GND GND VDD VDD _492_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2153 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_12_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2974 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1761 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_604_ _628_/A GND GND VDD VDD _609_/A sky130_fd_sc_hd__buf_2
XFILLER_18_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_535_ _712_/Q _711_/Q _537_/S GND GND VDD VDD _536_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1503 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_466_ _743_/Q _742_/Q _470_/S GND GND VDD VDD _467_/A sky130_fd_sc_hd__mux2_1
X_397_ _397_/A GND GND VDD VDD _774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2893 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2524 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1801 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2112 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1509 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_518_ _720_/Q _719_/Q _526_/S GND GND VDD VDD _519_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2045 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_449_ _449_/A GND GND VDD VDD _458_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_785 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1620 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1256 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2796 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1873 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1804 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_921 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_10_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_783_ _795_/CLK _783_/D _681_/Y GND GND VDD VDD _783_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_822 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_354 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1042 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput29 _707_/Q GND GND VDD VDD COL_SEL[32] sky130_fd_sc_hd__clkbuf_1
Xoutput18 _697_/Q GND GND VDD VDD COL_SEL[22] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_766_ _773_/CLK _766_/D _660_/Y GND GND VDD VDD _766_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_697_ _792_/CLK _697_/D _575_/Y GND GND VDD VDD _697_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2611 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_620_ _621_/A GND GND VDD VDD _620_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_551_ _705_/Q _704_/Q _559_/S GND GND VDD VDD _552_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_449 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_482_ _482_/A GND GND VDD VDD _736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_2110 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_749_ _774_/CLK _749_/D _639_/Y GND GND VDD VDD _749_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2986 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_1228 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2474 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1740 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_603_ _665_/A GND GND VDD VDD _628_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_534_ _534_/A GND GND VDD VDD _713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1515 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_465_ _465_/A GND GND VDD VDD _744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_396_ _796_/A _773_/Q _402_/S GND GND VDD VDD _397_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2937 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2783 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2536 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2124 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1581 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_10_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_577 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_517_ _561_/A GND GND VDD VDD _526_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2901 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_448_ _448_/A GND GND VDD VDD _751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_208 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_379_ _379_/A GND GND VDD VDD _782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_742 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_720 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_308 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2208 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1676 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_875 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_897 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3193 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1816 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_561 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_10_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_782_ _791_/CLK _782_/D _680_/Y GND GND VDD VDD _782_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_977 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_834 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_366 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2185 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1451 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1065 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput19 _698_/Q GND GND VDD VDD COL_SEL[23] sky130_fd_sc_hd__clkbuf_1
XFILLER_6_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_765_ _775_/CLK _765_/D _658_/Y GND GND VDD VDD _765_/Q sky130_fd_sc_hd__dfrtp_1
X_696_ _786_/CLK _696_/D _574_/Y GND GND VDD VDD _696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_5 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2870 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_550_ _561_/A GND GND VDD VDD _559_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_17_428 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_481_ _736_/Q _735_/Q _481_/S GND GND VDD VDD _482_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2188 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_748_ _771_/CLK _748_/D _638_/Y GND GND VDD VDD _748_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_450 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_679_ _683_/A GND GND VDD VDD _679_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_602_ _602_/A GND GND VDD VDD _602_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_533_ _713_/Q _712_/Q _537_/S GND GND VDD VDD _534_/A sky130_fd_sc_hd__mux2_1
X_464_ _744_/Q _743_/Q _470_/S GND GND VDD VDD _465_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1527 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_395_ _395_/A GND GND VDD VDD _775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2811 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1004 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2795 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_2__f_clk clkbuf_0_clk/X GND GND VDD VDD _786_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2548 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2129 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_516_ _516_/A GND GND VDD VDD _561_/A sky130_fd_sc_hd__buf_2
XFILLER_18_2058 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1313 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_447_ _751_/Q _750_/Q _447_/S GND GND VDD VDD _448_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_378_ _782_/Q _781_/Q _380_/S GND GND VDD VDD _379_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1379 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2713 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_2685 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2592 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1611 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_353 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_887 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_386 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_375 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2460 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_551 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_584 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_781_ _795_/CLK _781_/D _679_/Y GND GND VDD VDD _781_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1430 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_378 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1463 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2017 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1088 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2083 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_753 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_764_ _771_/CLK _764_/D _657_/Y GND GND VDD VDD _764_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_695_ _695_/A GND GND VDD VDD _695_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_6 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_480_ _480_/A GND GND VDD VDD _737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2181 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_747_ _773_/CLK _747_/D _637_/Y GND GND VDD VDD _747_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_678_ _690_/A GND GND VDD VDD _683_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_462 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2487 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1775 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_11_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_601_ _602_/A GND GND VDD VDD _601_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_532_ _532_/A GND GND VDD VDD _714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_463_ _463_/A GND GND VDD VDD _745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_394_ _775_/Q input1/X _402_/S GND GND VDD VDD _395_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1252 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2801 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2823 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_925 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2516 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1815 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_515_ _515_/A GND GND VDD VDD _721_/D sky130_fd_sc_hd__clkbuf_1
X_446_ _446_/A GND GND VDD VDD _752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_377_ _377_/A GND GND VDD VDD _783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1093 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2697 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1985 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2769 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_10_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_844 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2891 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_429_ _429_/A GND GND VDD VDD _760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xinput1 data_in GND GND VDD VDD input1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3245 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_6_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_780_ _795_/CLK _780_/D _677_/Y GND GND VDD VDD _780_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_313 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1475 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1012 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1117 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_360 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_393 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_763_ _771_/CLK _763_/D _656_/Y GND GND VDD VDD _763_/Q sky130_fd_sc_hd__dfrtp_1
X_694_ _695_/A GND GND VDD VDD _694_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_7 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1250 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1681 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_408 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1481 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1423 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_746_ _773_/CLK _746_/D _636_/Y GND GND VDD VDD _746_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_677_ _677_/A GND GND VDD VDD _677_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1754 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_600_ _602_/A GND GND VDD VDD _600_/Y sky130_fd_sc_hd__inv_2
X_531_ _714_/Q _713_/Q _537_/S GND GND VDD VDD _532_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_462_ _745_/Q _744_/Q _470_/S GND GND VDD VDD _463_/A sky130_fd_sc_hd__mux2_1
X_393_ _393_/A GND GND VDD VDD _402_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_16_1264 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2857 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_729_ _773_/CLK _729_/D _614_/Y GND GND VDD VDD _729_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_2720 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2753 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_948 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1827 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1595 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_514_ _721_/Q _720_/Q _514_/S GND GND VDD VDD _515_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_445_ _752_/Q _751_/Q _447_/S GND GND VDD VDD _446_/A sky130_fd_sc_hd__mux2_1
X_376_ _783_/Q _782_/Q _380_/S GND GND VDD VDD _377_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_701 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1205 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1112 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_428_ _760_/Q _759_/Q _436_/S GND GND VDD VDD _429_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1145 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_359_ _359_/A GND GND VDD VDD _791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xinput2 ena GND GND VDD VDD _516_/A sky130_fd_sc_hd__buf_6
XFILLER_0_2545 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_520 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1690 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2122 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_347 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1487 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1024 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3021 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_762_ _773_/CLK _762_/D _655_/Y GND GND VDD VDD _762_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_693_ _695_/A GND GND VDD VDD _693_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_8 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2604 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1947 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_585 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_745_ _771_/CLK _745_/D _633_/Y GND GND VDD VDD _745_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_676_ _677_/A GND GND VDD VDD _676_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_530_ _530_/A GND GND VDD VDD _715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_461_ _505_/A GND GND VDD VDD _470_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_392_ _392_/A GND GND VDD VDD _776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1276 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_728_ _773_/CLK _728_/D _613_/Y GND GND VDD VDD _728_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_659_ _659_/A GND GND VDD VDD _664_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_2710 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2776 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1839 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_513_ _513_/A GND GND VDD VDD _722_/D sky130_fd_sc_hd__clkbuf_1
X_444_ _444_/A GND GND VDD VDD _753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2916 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_375_ _375_/A GND GND VDD VDD _784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2677 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_581 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1625 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2050 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1228 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2860 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_427_ _449_/A GND GND VDD VDD _436_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_358_ _791_/Q _790_/Q _358_/S GND GND VDD VDD _359_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xinput3 rst GND GND VDD VDD _665_/A sky130_fd_sc_hd__buf_6
XFILLER_20_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1845 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_326 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_2145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1444 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1499 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3077 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2321 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1592 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1606 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_30 _771_/Q GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_761_ _775_/CLK _761_/D _654_/Y GND GND VDD VDD _761_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_692_ _695_/A GND GND VDD VDD _692_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_602 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_9 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1274 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2885 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_744_ _773_/CLK _744_/D _632_/Y GND GND VDD VDD _744_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_675_ _677_/A GND GND VDD VDD _675_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_421 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2936 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_443 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1060 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_281 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_460_ _516_/A GND GND VDD VDD _505_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_391_ _776_/Q _775_/Q _391_/S GND GND VDD VDD _392_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1244 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_1288 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_361 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_2837 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2909 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_727_ _775_/CLK _727_/D _612_/Y GND GND VDD VDD _727_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_658_ _658_/A GND GND VDD VDD _658_/Y sky130_fd_sc_hd__inv_2
X_589_ _590_/A GND GND VDD VDD _589_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2766 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2210 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_512_ _722_/Q _721_/Q _514_/S GND GND VDD VDD _513_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_443_ _753_/Q _752_/Q _447_/S GND GND VDD VDD _444_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_374_ _784_/Q _783_/Q _380_/S GND GND VDD VDD _375_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2928 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1900 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2689 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_1977 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1704 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_836 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_368 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_426_ _426_/A GND GND VDD VDD _761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_357_ _357_/A GND GND VDD VDD _792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_3165 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_4_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1534 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_949 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2157 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_10_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_611 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2680 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_409_ _409_/A GND GND VDD VDD _769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2250 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1621 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2377 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_20 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_2076 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_760_ _773_/CLK _760_/D _652_/Y GND GND VDD VDD _760_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_691_ _695_/A GND GND VDD VDD _691_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_614 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1220 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2897 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_452 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1927 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1640 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_743_ _774_/CLK _743_/D _631_/Y GND GND VDD VDD _743_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_674_ _677_/A GND GND VDD VDD _674_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_956 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1960 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1768 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_390_ _390_/A GND GND VDD VDD _777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_726_ _773_/CLK _726_/D _611_/Y GND GND VDD VDD _726_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_657_ _658_/A GND GND VDD VDD _657_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_588_ _590_/A GND GND VDD VDD _588_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1808 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_511_ _511_/A GND GND VDD VDD _723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_442_ _442_/A GND GND VDD VDD _754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_373_ _373_/A GND GND VDD VDD _785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_709_ _792_/CLK _709_/D _589_/Y GND GND VDD VDD _709_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_594 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2041 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_425_ _761_/Q _760_/Q _425_/S GND GND VDD VDD _426_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1126 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_356_ _792_/Q _791_/Q _358_/S GND GND VDD VDD _357_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2748 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3144 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_589 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_10_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_408_ _769_/Q _768_/Q _414_/S GND GND VDD VDD _409_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2262 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1677 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_12_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1619 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XANTENNA_10 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_21 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_725 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_690_ _690_/A GND GND VDD VDD _695_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_626 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_475 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2618 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1652 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2153 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1416 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_742_ _774_/CLK _742_/D _630_/Y GND GND VDD VDD _742_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_673_ _677_/A GND GND VDD VDD _673_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_968 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1972 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_261 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1747 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_725_ _773_/CLK _725_/D _609_/Y GND GND VDD VDD _725_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_656_ _658_/A GND GND VDD VDD _656_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_587_ _590_/A GND GND VDD VDD _587_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1780 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2223 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_510_ _723_/Q _722_/Q _514_/S GND GND VDD VDD _511_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_441_ _754_/Q _753_/Q _447_/S GND GND VDD VDD _442_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_372_ _785_/Q _784_/Q _380_/S GND GND VDD VDD _373_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_193 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_708_ _792_/CLK _708_/D _588_/Y GND GND VDD VDD _708_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_639_ _640_/A GND GND VDD VDD _639_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_12_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1639 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2064 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1396 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_805 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_304 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2852 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_424_ _424_/A GND GND VDD VDD _762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_355_ _355_/A GND GND VDD VDD _793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3112 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3217 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3178 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3156 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_2444 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1732 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_893 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_clk clkbuf_0_clk/X GND GND VDD VDD _792_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_407_ _407_/A GND GND VDD VDD _770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_11 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_20_332 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XANTENNA_22 _796_/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1491 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1480 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_638 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1108 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_410 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_465 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_487 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1664 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1453 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_501 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_741_ _774_/CLK _741_/D _629_/Y GND GND VDD VDD _741_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_672_ _690_/A GND GND VDD VDD _677_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1984 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_295 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2829 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_724_ _775_/CLK _724_/D _608_/Y GND GND VDD VDD _724_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_655_ _658_/A GND GND VDD VDD _655_/Y sky130_fd_sc_hd__inv_2
X_586_ _590_/A GND GND VDD VDD _586_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2482 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_9_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1792 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2235 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_440_ _440_/A GND GND VDD VDD _755_/D sky130_fd_sc_hd__clkbuf_1
X_371_ _393_/A GND GND VDD VDD _380_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2780 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_707_ _792_/CLK _707_/D _587_/Y GND GND VDD VDD _707_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_638_ _640_/A GND GND VDD VDD _638_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_574 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_569_ _569_/A GND GND VDD VDD _697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2599 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_423_ _762_/Q _761_/Q _425_/S GND GND VDD VDD _424_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_354_ _793_/Q _792_/Q _358_/S GND GND VDD VDD _355_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3124 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2412 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2517 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_371 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_603 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_406_ _770_/Q _769_/Q _414_/S GND GND VDD VDD _407_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_341 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1971 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2297 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XANTENNA_12 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_23 _796_/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1201 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2881 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_8_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_444 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_499 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1621 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1676 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_174 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_740_ _771_/CLK _740_/D _627_/Y GND GND VDD VDD _740_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_557 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_671_ _671_/A GND GND VDD VDD _671_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_937 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_915 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_436 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2929 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1086 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_274 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2185 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_15_2196 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2940 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_723_ _792_/CLK _723_/D _607_/Y GND GND VDD VDD _723_/Q sky130_fd_sc_hd__dfrtp_1
X_654_ _658_/A GND GND VDD VDD _654_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_585_ _597_/A GND GND VDD VDD _590_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_370_ _370_/A GND GND VDD VDD _786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2792 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_13_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_706_ _792_/CLK _706_/D _586_/Y GND GND VDD VDD _706_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_637_ _640_/A GND GND VDD VDD _637_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_568_ _697_/Q _696_/Q _570_/S GND GND VDD VDD _569_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_729 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_499_ _728_/Q _727_/Q _503_/S GND GND VDD VDD _500_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_829 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_422_ _422_/A GND GND VDD VDD _763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_353_ _353_/A GND GND VDD VDD _794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_862 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1817 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_383 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2991 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_320 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_405_ _449_/A GND GND VDD VDD _414_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1983 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3049 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1564 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2150 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_13 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_18_2183 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_24 _796_/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_11_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2069 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1213 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1909 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_15_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2492 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1780 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2040 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1394 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_197 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_186 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_5_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_670_ _671_/A GND GND VDD VDD _670_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1920 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1180 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1285 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_13_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2952 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_333 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_722_ _786_/CLK _722_/D _606_/Y GND GND VDD VDD _722_/Q sky130_fd_sc_hd__dfrtp_1
X_653_ _659_/A GND GND VDD VDD _658_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_584_ _584_/A GND GND VDD VDD _584_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2473 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_705_ _792_/CLK _705_/D _584_/Y GND GND VDD VDD _705_/Q sky130_fd_sc_hd__dfrtp_1
X_636_ _640_/A GND GND VDD VDD _636_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_565 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_567_ _567_/A GND GND VDD VDD _698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_708 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2579 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_498_ _498_/A GND GND VDD VDD _729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1889 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_329 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_421_ _763_/Q _762_/Q _425_/S GND GND VDD VDD _422_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_2844 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1119 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_352_ _794_/Q _793_/Q _358_/S GND GND VDD VDD _353_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_6_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3137 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_852 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_619_ _621_/A GND GND VDD VDD _619_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_538 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1406 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2641 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_404_ _516_/A GND GND VDD VDD _449_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1995 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2349 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_14 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_25 _796_/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2460 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2081 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1340 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2096 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1409 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2880 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_928 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2622 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_950 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1420 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1192 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2964 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_389 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_721_ _786_/CLK _721_/D _605_/Y GND GND VDD VDD _721_/Q sky130_fd_sc_hd__dfrtp_1
X_652_ _652_/A GND GND VDD VDD _652_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_583_ _584_/A GND GND VDD VDD _583_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1061 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_13_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2761 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_704_ _792_/CLK _704_/D _583_/Y GND GND VDD VDD _704_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_635_ _659_/A GND GND VDD VDD _640_/A sky130_fd_sc_hd__buf_2
XFILLER_18_2514 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_566_ _698_/Q _697_/Q _570_/S GND GND VDD VDD _567_/A sky130_fd_sc_hd__mux2_1
X_497_ _729_/Q _728_/Q _503_/S GND GND VDD VDD _498_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2057 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2901 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_420_ _420_/A GND GND VDD VDD _764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_2867 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_351_ _351_/A GND GND VDD VDD _795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2437 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_330 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_618_ _621_/A GND GND VDD VDD _618_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1632 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_549_ _549_/A GND GND VDD VDD _706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_617 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_403_ _403_/A GND GND VDD VDD _771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_355 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_15_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1544 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1649 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_15 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_26 _770_/Q GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_11_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput100 _772_/Q GND GND VDD VDD COL_SEL[97] sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1237 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_892 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1793 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2125 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_144 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1270 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2634 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_962 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2280 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1432 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_720_ _786_/CLK _720_/D _602_/Y GND GND VDD VDD _720_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_651_ _652_/A GND GND VDD VDD _651_/Y sky130_fd_sc_hd__inv_2
X_582_ _584_/A GND GND VDD VDD _582_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2729 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1752 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3300 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_165 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_703_ _795_/CLK _703_/D _582_/Y GND GND VDD VDD _703_/Q sky130_fd_sc_hd__dfrtp_1
X_634_ _665_/A GND GND VDD VDD _659_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2526 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_565_ _565_/A GND GND VDD VDD _699_/D sky130_fd_sc_hd__clkbuf_1
X_496_ _496_/A GND GND VDD VDD _730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_350_ _795_/Q _794_/Q _358_/S GND GND VDD VDD _351_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1704 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_364 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_617_ _621_/A GND GND VDD VDD _617_/Y sky130_fd_sc_hd__inv_2
X_548_ _706_/Q _705_/Q _548_/S GND GND VDD VDD _549_/A sky130_fd_sc_hd__mux2_1
X_479_ _737_/Q _736_/Q _481_/S GND GND VDD VDD _480_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1666 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2972 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2109 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1110 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_11_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_402_ _771_/Q _770_/Q _402_/S GND GND VDD VDD _403_/A sky130_fd_sc_hd__mux2_1
XPHY_40 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_334 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1964 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1556 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_304 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XANTENNA_16 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_20_337 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XANTENNA_27 _665_/A GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_11_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput101 _773_/Q GND GND VDD VDD COL_SEL[98] sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_437 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2010 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1425 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_156 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_429 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2646 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_796_ _796_/A GND GND VDD VDD _796_/X sky130_fd_sc_hd__buf_6
XFILLER_1_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_974 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2292 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1444 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_650_ _652_/A GND GND VDD VDD _650_/Y sky130_fd_sc_hd__inv_2
X_581_ _584_/A GND GND VDD VDD _581_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_779_ _791_/CLK _779_/D _676_/Y GND GND VDD VDD _779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_702_ _792_/CLK _702_/D _581_/Y GND GND VDD VDD _702_/Q sky130_fd_sc_hd__dfrtp_1
X_633_ _633_/A GND GND VDD VDD _633_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_564_ _699_/Q _698_/Q _570_/S GND GND VDD VDD _565_/A sky130_fd_sc_hd__mux2_1
X_495_ _730_/Q _729_/Q _503_/S GND GND VDD VDD _496_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2538 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2240 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2825 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2836 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2428 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_4_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_616_ _628_/A GND GND VDD VDD _621_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_547_ _547_/A GND GND VDD VDD _707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_508 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_478_ _478_/A GND GND VDD VDD _738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1678 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1509 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1100 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2880 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2600 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2633 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XPHY_30 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_401_ _401_/A GND GND VDD VDD _772_/D sky130_fd_sc_hd__clkbuf_1
XPHY_41 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2269 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_641 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2176 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XANTENNA_17 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_28 _771_/Q GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_9_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput102 _796_/A GND GND VDD VDD COL_SEL[99] sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2853 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1228 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2073 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2894 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_529 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1913 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_795_ _795_/CLK _795_/D _695_/Y GND GND VDD VDD _795_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_clk clkbuf_0_clk/X GND GND VDD VDD _771_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1401 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1201 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1173 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_1_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_580_ _584_/A GND GND VDD VDD _580_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_893 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_778_ _791_/CLK _778_/D _675_/Y GND GND VDD VDD _778_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_701_ _795_/CLK _701_/D _580_/Y GND GND VDD VDD _701_/Q sky130_fd_sc_hd__dfrtp_1
X_632_ _633_/A GND GND VDD VDD _632_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_563_ _563_/A GND GND VDD VDD _700_/D sky130_fd_sc_hd__clkbuf_1
X_494_ _505_/A GND GND VDD VDD _503_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_13_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2252 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2915 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_615_ _615_/A GND GND VDD VDD _615_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_546_ _707_/Q _706_/Q _548_/S GND GND VDD VDD _547_/A sky130_fd_sc_hd__mux2_1
X_477_ _738_/Q _737_/Q _481_/S GND GND VDD VDD _478_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_400_ _772_/Q _771_/Q _402_/S GND GND VDD VDD _401_/A sky130_fd_sc_hd__mux2_1
XPHY_31 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_20 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_2656 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1900 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1569 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_529_ _715_/Q _714_/Q _537_/S GND GND VDD VDD _530_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1432 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_18 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_29 _771_/Q GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput103 _784_/Q GND GND VDD VDD COL_SEL[9] sky130_fd_sc_hd__clkbuf_1
XFILLER_5_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_22 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2453 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2045 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1355 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1251 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_11_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2615 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1936 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_794_ _795_/CLK _794_/D _694_/Y GND GND VDD VDD _794_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_943 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2125 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1560 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_15_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_291 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1257 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_305 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_777_ _792_/CLK _777_/D _674_/Y GND GND VDD VDD _777_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2754 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_700_ _792_/CLK _700_/D _578_/Y GND GND VDD VDD _700_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_631_ _633_/A GND GND VDD VDD _631_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_562_ _700_/Q _699_/Q _570_/S GND GND VDD VDD _563_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2507 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_493_ _493_/A GND GND VDD VDD _731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1806 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2264 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_592 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2927 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_813 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_614_ _615_/A GND GND VDD VDD _614_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_545_ _545_/A GND GND VDD VDD _708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1603 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_476_ _476_/A GND GND VDD VDD _739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2997 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_3_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2860 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2624 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XPHY_10 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_21 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_2668 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_32 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1956 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_348 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_528_ _561_/A GND GND VDD VDD _537_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1411 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XANTENNA_19 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
X_459_ _459_/A GND GND VDD VDD _746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1444 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput104 _796_/X GND GND VDD VDD data_out sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_885 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_34 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1731 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1628 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2068 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_974 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_137 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2685 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1005 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_660 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1948 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_793_ _795_/CLK _793_/D _693_/Y GND GND VDD VDD _793_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3161 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1745 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_776_ _791_/CLK _776_/D _673_/Y GND GND VDD VDD _776_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1033 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_630_ _633_/A GND GND VDD VDD _630_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_561_ _561_/A GND GND VDD VDD _570_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_17_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_492_ _731_/Q _730_/Q _492_/S GND GND VDD VDD _493_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_759_ _773_/CLK _759_/D _651_/Y GND GND VDD VDD _759_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1096 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2585 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_10_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_613_ _615_/A GND GND VDD VDD _613_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_346 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_544_ _708_/Q _707_/Q _548_/S GND GND VDD VDD _545_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_357 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_475_ _739_/Q _738_/Q _481_/S GND GND VDD VDD _476_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1648 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2095 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_880 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_11 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_22 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_33 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_327 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1516 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_633 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_4_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_527_ _527_/A GND GND VDD VDD _716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_458_ _746_/Q _745_/Q _458_/S GND GND VDD VDD _459_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1456 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_389_ _777_/Q _776_/Q _391_/S GND GND VDD VDD _390_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_371 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_897 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_46 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_11_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1743 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_953 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1368 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1220 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2570 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1985 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1927 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_792_ _792_/CLK _792_/D _692_/Y GND GND VDD VDD _792_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1061 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2461 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1768 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_775_ _775_/CLK _775_/D _671_/Y GND GND VDD VDD _775_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2082 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_81 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1089 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_137 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_560_ _560_/A GND GND VDD VDD _701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_491_ _491_/A GND GND VDD VDD _732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_758_ _771_/CLK _758_/D _650_/Y GND GND VDD VDD _758_/Q sky130_fd_sc_hd__dfrtp_1
X_689_ _689_/A GND GND VDD VDD _689_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1709 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_826 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_612_ _615_/A GND GND VDD VDD _612_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_543_ _543_/A GND GND VDD VDD _709_/D sky130_fd_sc_hd__clkbuf_1
X_474_ _474_/A GND GND VDD VDD _740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_892 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_12 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_34 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_23 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1513 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1528 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_526_ _716_/Q _715_/Q _526_/S GND GND VDD VDD _527_/A sky130_fd_sc_hd__mux2_1
X_457_ _457_/A GND GND VDD VDD _747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_309 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2169 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1424 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1468 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_388_ _388_/A GND GND VDD VDD _778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_383 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_13_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2445 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1788 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2088 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_921 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_509_ _509_/A GND GND VDD VDD _724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2887 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3261 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_791_ _791_/CLK _791_/D _691_/Y GND GND VDD VDD _791_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_935 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1761 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_470 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_774_ _774_/CLK _774_/D _670_/Y GND GND VDD VDD _796_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2768 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_490_ _732_/Q _731_/Q _492_/S GND GND VDD VDD _491_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_757_ _773_/CLK _757_/D _649_/Y GND GND VDD VDD _757_/Q sky130_fd_sc_hd__dfrtp_1
X_688_ _689_/A GND GND VDD VDD _688_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_611_ _615_/A GND GND VDD VDD _611_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_542_ _709_/Q _708_/Q _548_/S GND GND VDD VDD _543_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_473_ _740_/Q _739_/Q _481_/S GND GND VDD VDD _474_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_13 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_2649 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XPHY_35 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_24 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_1650 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_525_ _525_/A GND GND VDD VDD _717_/D sky130_fd_sc_hd__clkbuf_1
X_456_ _747_/Q _746_/Q _458_/S GND GND VDD VDD _457_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_340 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_387_ _778_/Q _777_/Q _391_/S GND GND VDD VDD _388_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2825 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1723 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1767 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2027 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_966 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_421 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_508_ _724_/Q _723_/Q _514_/S GND GND VDD VDD _509_/A sky130_fd_sc_hd__mux2_1
X_439_ _755_/Q _754_/Q _447_/S GND GND VDD VDD _440_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2608 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_790_ _792_/CLK _790_/D _689_/Y GND GND VDD VDD _790_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2210 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1704 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1759 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_865 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_773_ _773_/CLK _773_/D _669_/Y GND GND VDD VDD _773_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1383 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2293 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2202 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1534 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_756_ _775_/CLK _756_/D _648_/Y GND GND VDD VDD _756_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_687_ _689_/A GND GND VDD VDD _687_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_15_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2577 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_610_ _628_/A GND GND VDD VDD _615_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_839 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_541_ _541_/A GND GND VDD VDD _710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_472_ _505_/A GND GND VDD VDD _481_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_16_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1397 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2979 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_739_ _771_/CLK _739_/D _626_/Y GND GND VDD VDD _739_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_36 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_14 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_25 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1949 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1662 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_614 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_524_ _717_/Q _716_/Q _526_/S GND GND VDD VDD _525_/A sky130_fd_sc_hd__mux2_1
X_455_ _455_/A GND GND VDD VDD _748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_2138 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_386_ _386_/A GND GND VDD VDD _779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput90 _763_/Q GND GND VDD VDD COL_SEL[88] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_878 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_466 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_507_ _507_/A GND GND VDD VDD _725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_438_ _449_/A GND GND VDD VDD _447_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_20_108 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_369_ _786_/Q _785_/Q _369_/S GND GND VDD VDD _370_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2601 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_1861 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1872 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2244 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1587 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_775 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_797 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1229 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1075 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1691 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_772_ _773_/CLK _772_/D _668_/Y GND GND VDD VDD _772_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2041 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1593 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_641 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_755_ _774_/CLK _755_/D _646_/Y GND GND VDD VDD _755_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_686_ _689_/A GND GND VDD VDD _686_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1089 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2501 GND GND VDD VDD sky130_fd_sc_hd__decap_4
Xclkbuf_3_5__f_clk clkbuf_0_clk/X GND GND VDD VDD _774_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_540_ _710_/Q _709_/Q _548_/S GND GND VDD VDD _541_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_306 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_471_ _471_/A GND GND VDD VDD _741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_738_ _771_/CLK _738_/D _625_/Y GND GND VDD VDD _738_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_669_ _671_/A GND GND VDD VDD _669_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XPHY_37 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_15 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_26 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_309 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1674 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1509 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_523_ _523_/A GND GND VDD VDD _718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_454_ _748_/Q _747_/Q _458_/S GND GND VDD VDD _455_/A sky130_fd_sc_hd__mux2_1
X_385_ _779_/Q _778_/Q _391_/S GND GND VDD VDD _386_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1140 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput91 _764_/Q GND GND VDD VDD COL_SEL[89] sky130_fd_sc_hd__clkbuf_1
Xoutput80 _754_/Q GND GND VDD VDD COL_SEL[79] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_813 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_434 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_506_ _725_/Q _724_/Q _514_/S GND GND VDD VDD _507_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_437_ _437_/A GND GND VDD VDD _756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_368_ _368_/A GND GND VDD VDD _787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2657 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1901 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2481 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_676 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1677 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2256 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2234 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1408 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3133 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_771_ _771_/CLK _771_/D _667_/Y GND GND VDD VDD _771_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1396 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1005 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2738 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_281 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_697 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_754_ _775_/CLK _754_/D _645_/Y GND GND VDD VDD _754_/Q sky130_fd_sc_hd__dfrtp_1
X_685_ _689_/A GND GND VDD VDD _685_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_370 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_808 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_470_ _741_/Q _740_/Q _470_/S GND GND VDD VDD _471_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2045 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_1300 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_737_ _771_/CLK _737_/D _624_/Y GND GND VDD VDD _737_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_668_ _671_/A GND GND VDD VDD _668_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2844 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_599_ _602_/A GND GND VDD VDD _599_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_0 _690_/A GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_8_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_38 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_27 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_16 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1620 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_522_ _718_/Q _717_/Q _526_/S GND GND VDD VDD _523_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_453_ _453_/A GND GND VDD VDD _749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_384_ _384_/A GND GND VDD VDD _780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput70 _781_/Q GND GND VDD VDD COL_SEL[6] sky130_fd_sc_hd__clkbuf_1
Xoutput92 _783_/Q GND GND VDD VDD COL_SEL[8] sky130_fd_sc_hd__clkbuf_1
Xoutput81 _782_/Q GND GND VDD VDD COL_SEL[7] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2685 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_836 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1962 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1329 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_505_ _505_/A GND GND VDD VDD _514_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_436_ _756_/Q _755_/Q _436_/S GND GND VDD VDD _437_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_367_ _787_/Q _786_/Q _369_/S GND GND VDD VDD _368_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2869 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_13_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2531 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1957 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2493 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_688 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_928 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2268 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1578 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1280 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_10_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_419_ _764_/Q _763_/Q _425_/S GND GND VDD VDD _420_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1088 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1099 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3084 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2433 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3189 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_770_ _775_/CLK _770_/D _664_/Y GND GND VDD VDD _770_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_109 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_6_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2216 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_753_ _774_/CLK _753_/D _644_/Y GND GND VDD VDD _753_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_684_ _690_/A GND GND VDD VDD _689_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1312 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_473 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_736_ _773_/CLK _736_/D _623_/Y GND GND VDD VDD _736_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_667_ _671_/A GND GND VDD VDD _667_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_330 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_598_ _602_/A GND GND VDD VDD _598_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_897 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_1_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2867 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_1 _690_/A GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_6_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_17 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_28 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_39 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1643 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_521_ _521_/A GND GND VDD VDD _719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_452_ _749_/Q _748_/Q _458_/S GND GND VDD VDD _453_/A sky130_fd_sc_hd__mux2_1
X_383_ _780_/Q _779_/Q _391_/S GND GND VDD VDD _384_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput60 _735_/Q GND GND VDD VDD COL_SEL[60] sky130_fd_sc_hd__clkbuf_1
Xoutput93 _765_/Q GND GND VDD VDD COL_SEL[90] sky130_fd_sc_hd__clkbuf_1
Xoutput82 _755_/Q GND GND VDD VDD COL_SEL[80] sky130_fd_sc_hd__clkbuf_1
Xoutput71 _745_/Q GND GND VDD VDD COL_SEL[70] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_719_ _786_/CLK _719_/D _601_/Y GND GND VDD VDD _719_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_2631 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1974 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2196 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_458 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_504_ _504_/A GND GND VDD VDD _726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_435_ _435_/A GND GND VDD VDD _757_/D sky130_fd_sc_hd__clkbuf_1
X_366_ _366_/A GND GND VDD VDD _788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3211 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_9_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_3244 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_3233 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_3277 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_970 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_1886 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_612 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1116 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_277 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_418_ _418_/A GND GND VDD VDD _765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_349_ _393_/A GND GND VDD VDD _358_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3096 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2384 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2489 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1733 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_486 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2033 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2932 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_1376 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2228 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_752_ _775_/CLK _752_/D _643_/Y GND GND VDD VDD _752_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_683_ _683_/A GND GND VDD VDD _683_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2058 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2902 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_11_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_735_ _771_/CLK _735_/D _621_/Y GND GND VDD VDD _735_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_666_ _690_/A GND GND VDD VDD _671_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_597_ _597_/A GND GND VDD VDD _602_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_2 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_12_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_29 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_18 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1633 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_607 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_520_ _719_/Q _718_/Q _526_/S GND GND VDD VDD _521_/A sky130_fd_sc_hd__mux2_1
X_451_ _451_/A GND GND VDD VDD _750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_382_ _393_/A GND GND VDD VDD _391_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput4 _775_/Q GND GND VDD VDD COL_SEL[0] sky130_fd_sc_hd__clkbuf_1
Xoutput61 _736_/Q GND GND VDD VDD COL_SEL[61] sky130_fd_sc_hd__clkbuf_1
Xoutput50 _726_/Q GND GND VDD VDD COL_SEL[51] sky130_fd_sc_hd__clkbuf_1
Xoutput94 _766_/Q GND GND VDD VDD COL_SEL[91] sky130_fd_sc_hd__clkbuf_1
Xoutput83 _756_/Q GND GND VDD VDD COL_SEL[81] sky130_fd_sc_hd__clkbuf_1
Xoutput72 _746_/Q GND GND VDD VDD COL_SEL[71] sky130_fd_sc_hd__clkbuf_1
XFILLER_4_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_718_ _786_/CLK _718_/D _600_/Y GND GND VDD VDD _718_/Q sky130_fd_sc_hd__dfrtp_1
X_649_ _652_/A GND GND VDD VDD _649_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2698 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1430 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_503_ _726_/Q _725_/Q _503_/S GND GND VDD VDD _504_/A sky130_fd_sc_hd__mux2_1
X_434_ _757_/Q _756_/Q _436_/S GND GND VDD VDD _435_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1227 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_365_ _788_/Q _787_/Q _369_/S GND GND VDD VDD _366_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3201 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2544 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1843 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1810 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1794 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_417_ _765_/Q _764_/Q _425_/S GND GND VDD VDD _418_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_348_ _516_/A GND GND VDD VDD _393_/A sky130_fd_sc_hd__buf_4
XFILLER_18_1068 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2396 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1684 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1789 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_421 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_498 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_837 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3280 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_8_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2265 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_clk clkbuf_0_clk/X GND GND VDD VDD _791_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_751_ _775_/CLK _751_/D _642_/Y GND GND VDD VDD _751_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_682_ _683_/A GND GND VDD VDD _682_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1130 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_74 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_1_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_734_ _773_/CLK _734_/D _620_/Y GND GND VDD VDD _734_/Q sky130_fd_sc_hd__dfrtp_1
X_665_ _665_/A GND GND VDD VDD _690_/A sky130_fd_sc_hd__buf_4
XFILLER_17_844 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_596_ _596_/A GND GND VDD VDD _596_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_343 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_1_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_3 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_12_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_19 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_450_ _750_/Q _749_/Q _458_/S GND GND VDD VDD _451_/A sky130_fd_sc_hd__mux2_1
X_381_ _381_/A GND GND VDD VDD _781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput5 _785_/Q GND GND VDD VDD COL_SEL[10] sky130_fd_sc_hd__clkbuf_1
Xoutput51 _727_/Q GND GND VDD VDD COL_SEL[52] sky130_fd_sc_hd__clkbuf_1
Xoutput40 _717_/Q GND GND VDD VDD COL_SEL[42] sky130_fd_sc_hd__clkbuf_1
Xoutput73 _747_/Q GND GND VDD VDD COL_SEL[72] sky130_fd_sc_hd__clkbuf_1
Xoutput84 _757_/Q GND GND VDD VDD COL_SEL[82] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput62 _737_/Q GND GND VDD VDD COL_SEL[62] sky130_fd_sc_hd__clkbuf_1
Xoutput95 _767_/Q GND GND VDD VDD COL_SEL[92] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_717_ _791_/CLK _717_/D _599_/Y GND GND VDD VDD _717_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_648_ _652_/A GND GND VDD VDD _648_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_579_ _597_/A GND GND VDD VDD _584_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1442 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_416 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_502_ _502_/A GND GND VDD VDD _727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_433_ _433_/A GND GND VDD VDD _758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_364_ _364_/A GND GND VDD VDD _789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1537 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1548 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1261 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2894 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_416_ _449_/A GND GND VDD VDD _425_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1681 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_444 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1592 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2068 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1080 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_566 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3292 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1565 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_13_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_241 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_613 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_750_ _775_/CLK _750_/D _640_/Y GND GND VDD VDD _750_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_681_ _683_/A GND GND VDD VDD _681_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1142 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2742 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2041 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_20 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_97 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_733_ _775_/CLK _733_/D _619_/Y GND GND VDD VDD _733_/Q sky130_fd_sc_hd__dfrtp_1
X_664_ _664_/A GND GND VDD VDD _664_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_856 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_595_ _596_/A GND GND VDD VDD _595_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_355 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_4 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_6_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_380_ _781_/Q _780_/Q _380_/S GND GND VDD VDD _381_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1101 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_347 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput6 _786_/Q GND GND VDD VDD COL_SEL[11] sky130_fd_sc_hd__clkbuf_1
Xoutput52 _728_/Q GND GND VDD VDD COL_SEL[53] sky130_fd_sc_hd__clkbuf_1
Xoutput41 _718_/Q GND GND VDD VDD COL_SEL[43] sky130_fd_sc_hd__clkbuf_1
Xoutput30 _708_/Q GND GND VDD VDD COL_SEL[33] sky130_fd_sc_hd__clkbuf_1
Xoutput74 _748_/Q GND GND VDD VDD COL_SEL[73] sky130_fd_sc_hd__clkbuf_1
Xoutput85 _758_/Q GND GND VDD VDD COL_SEL[83] sky130_fd_sc_hd__clkbuf_1
Xoutput63 _738_/Q GND GND VDD VDD COL_SEL[63] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput96 _768_/Q GND GND VDD VDD COL_SEL[93] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_716_ _786_/CLK _716_/D _598_/Y GND GND VDD VDD _716_/Q sky130_fd_sc_hd__dfrtp_1
X_647_ _659_/A GND GND VDD VDD _652_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_578_ _578_/A GND GND VDD VDD _578_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1955 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
.ends

.subckt array_SR COL_ENA COL_RST COL_DIN COL_CLK COL_DOUT CSA_VREF ARRAY_OUT NB1 NB2
+ VBIAS VREF SF_IB ROW_DIN ROW_CLK ROW_RST gring ROW_ENA VDD GND
Xpixel_array100x100_0 VBIAS VREF NB2 NB1 shift_registerC_1/COL_SEL[0] gring shift_registerC_1/COL_SEL[1]
+ shift_registerC_1/COL_SEL[2] shift_registerC_1/COL_SEL[3] shift_registerC_1/COL_SEL[4]
+ shift_registerC_1/COL_SEL[5] shift_registerC_1/COL_SEL[6] shift_registerC_1/COL_SEL[7]
+ shift_registerC_1/COL_SEL[8] shift_registerC_1/COL_SEL[9] shift_registerC_1/COL_SEL[10]
+ shift_registerC_1/COL_SEL[11] shift_registerC_1/COL_SEL[12] shift_registerC_1/COL_SEL[13]
+ shift_registerC_1/COL_SEL[14] shift_registerC_1/COL_SEL[15] shift_registerC_1/COL_SEL[16]
+ shift_registerC_1/COL_SEL[17] shift_registerC_1/COL_SEL[18] shift_registerC_1/COL_SEL[19]
+ shift_registerC_1/COL_SEL[20] shift_registerC_1/COL_SEL[21] shift_registerC_1/COL_SEL[22]
+ shift_registerC_1/COL_SEL[23] shift_registerC_1/COL_SEL[24] shift_registerC_1/COL_SEL[25]
+ shift_registerC_1/COL_SEL[26] shift_registerC_1/COL_SEL[27] shift_registerC_1/COL_SEL[28]
+ shift_registerC_1/COL_SEL[29] shift_registerC_1/COL_SEL[30] shift_registerC_1/COL_SEL[31]
+ shift_registerC_1/COL_SEL[32] shift_registerC_1/COL_SEL[33] shift_registerC_1/COL_SEL[34]
+ shift_registerC_1/COL_SEL[35] shift_registerC_1/COL_SEL[36] shift_registerC_1/COL_SEL[37]
+ shift_registerC_1/COL_SEL[38] shift_registerC_1/COL_SEL[39] shift_registerC_1/COL_SEL[40]
+ shift_registerC_1/COL_SEL[41] shift_registerC_1/COL_SEL[42] shift_registerC_1/COL_SEL[43]
+ shift_registerC_1/COL_SEL[44] shift_registerC_1/COL_SEL[45] shift_registerC_1/COL_SEL[46]
+ shift_registerC_1/COL_SEL[47] shift_registerC_1/COL_SEL[48] shift_registerC_1/COL_SEL[49]
+ shift_registerC_1/COL_SEL[50] shift_registerC_1/COL_SEL[51] shift_registerC_1/COL_SEL[52]
+ shift_registerC_1/COL_SEL[53] shift_registerC_1/COL_SEL[54] shift_registerC_1/COL_SEL[55]
+ shift_registerC_1/COL_SEL[56] shift_registerC_1/COL_SEL[57] shift_registerC_1/COL_SEL[58]
+ shift_registerC_1/COL_SEL[59] shift_registerC_1/COL_SEL[60] shift_registerC_1/COL_SEL[61]
+ shift_registerC_1/COL_SEL[62] shift_registerC_1/COL_SEL[63] shift_registerC_1/COL_SEL[64]
+ shift_registerC_1/COL_SEL[65] shift_registerC_1/COL_SEL[66] shift_registerC_1/COL_SEL[67]
+ shift_registerC_1/COL_SEL[68] shift_registerC_1/COL_SEL[69] shift_registerC_1/COL_SEL[70]
+ shift_registerC_1/COL_SEL[71] shift_registerC_1/COL_SEL[72] shift_registerC_1/COL_SEL[73]
+ shift_registerC_1/COL_SEL[74] shift_registerC_1/COL_SEL[75] shift_registerC_1/COL_SEL[76]
+ shift_registerC_1/COL_SEL[77] shift_registerC_1/COL_SEL[78] shift_registerC_1/COL_SEL[79]
+ shift_registerC_1/COL_SEL[80] shift_registerC_1/COL_SEL[81] shift_registerC_1/COL_SEL[82]
+ shift_registerC_1/COL_SEL[83] shift_registerC_1/COL_SEL[84] shift_registerC_1/COL_SEL[85]
+ shift_registerC_1/COL_SEL[86] shift_registerC_1/COL_SEL[87] shift_registerC_1/COL_SEL[88]
+ shift_registerC_1/COL_SEL[89] shift_registerC_1/COL_SEL[90] shift_registerC_1/COL_SEL[91]
+ shift_registerC_1/COL_SEL[92] shift_registerC_1/COL_SEL[93] shift_registerC_1/COL_SEL[94]
+ shift_registerC_1/COL_SEL[95] shift_registerC_1/COL_SEL[96] shift_registerC_1/COL_SEL[97]
+ shift_registerC_1/COL_SEL[98] shift_registerC_0/COL_SEL[0] CSA_VREF shift_registerC_1/COL_SEL[99]
+ shift_registerC_0/COL_SEL[1] shift_registerC_0/COL_SEL[2] shift_registerC_0/COL_SEL[3]
+ shift_registerC_0/COL_SEL[4] shift_registerC_0/COL_SEL[5] shift_registerC_0/COL_SEL[6]
+ shift_registerC_0/COL_SEL[7] shift_registerC_0/COL_SEL[8] shift_registerC_0/COL_SEL[9]
+ shift_registerC_0/COL_SEL[10] shift_registerC_0/COL_SEL[11] shift_registerC_0/COL_SEL[12]
+ shift_registerC_0/COL_SEL[13] shift_registerC_0/COL_SEL[14] shift_registerC_0/COL_SEL[15]
+ shift_registerC_0/COL_SEL[16] shift_registerC_0/COL_SEL[17] shift_registerC_0/COL_SEL[18]
+ shift_registerC_0/COL_SEL[19] shift_registerC_0/COL_SEL[20] shift_registerC_0/COL_SEL[21]
+ shift_registerC_0/COL_SEL[22] shift_registerC_0/COL_SEL[23] shift_registerC_0/COL_SEL[24]
+ shift_registerC_0/COL_SEL[25] shift_registerC_0/COL_SEL[26] shift_registerC_0/COL_SEL[27]
+ shift_registerC_0/COL_SEL[28] shift_registerC_0/COL_SEL[29] shift_registerC_0/COL_SEL[30]
+ shift_registerC_0/COL_SEL[31] shift_registerC_0/COL_SEL[32] shift_registerC_0/COL_SEL[33]
+ shift_registerC_0/COL_SEL[34] shift_registerC_0/COL_SEL[35] shift_registerC_0/COL_SEL[36]
+ shift_registerC_0/COL_SEL[37] shift_registerC_0/COL_SEL[38] shift_registerC_0/COL_SEL[39]
+ shift_registerC_0/COL_SEL[40] shift_registerC_0/COL_SEL[41] shift_registerC_0/COL_SEL[42]
+ shift_registerC_0/COL_SEL[43] shift_registerC_0/COL_SEL[44] shift_registerC_0/COL_SEL[45]
+ shift_registerC_0/COL_SEL[46] shift_registerC_0/COL_SEL[47] shift_registerC_0/COL_SEL[48]
+ shift_registerC_0/COL_SEL[49] shift_registerC_0/COL_SEL[50] shift_registerC_0/COL_SEL[51]
+ shift_registerC_0/COL_SEL[52] shift_registerC_0/COL_SEL[53] shift_registerC_0/COL_SEL[54]
+ shift_registerC_0/COL_SEL[55] shift_registerC_0/COL_SEL[56] shift_registerC_0/COL_SEL[57]
+ shift_registerC_0/COL_SEL[58] shift_registerC_0/COL_SEL[59] shift_registerC_0/COL_SEL[60]
+ shift_registerC_0/COL_SEL[61] shift_registerC_0/COL_SEL[62] shift_registerC_0/COL_SEL[63]
+ shift_registerC_0/COL_SEL[64] shift_registerC_0/COL_SEL[65] shift_registerC_0/COL_SEL[66]
+ shift_registerC_0/COL_SEL[67] shift_registerC_0/COL_SEL[68] shift_registerC_0/COL_SEL[69]
+ shift_registerC_0/COL_SEL[70] shift_registerC_0/COL_SEL[71] shift_registerC_0/COL_SEL[72]
+ shift_registerC_0/COL_SEL[73] shift_registerC_0/COL_SEL[74] shift_registerC_0/COL_SEL[75]
+ shift_registerC_0/COL_SEL[76] shift_registerC_0/COL_SEL[77] shift_registerC_0/COL_SEL[78]
+ shift_registerC_0/COL_SEL[79] shift_registerC_0/COL_SEL[80] shift_registerC_0/COL_SEL[81]
+ shift_registerC_0/COL_SEL[82] shift_registerC_0/COL_SEL[83] shift_registerC_0/COL_SEL[84]
+ shift_registerC_0/COL_SEL[85] shift_registerC_0/COL_SEL[86] shift_registerC_0/COL_SEL[87]
+ shift_registerC_0/COL_SEL[88] shift_registerC_0/COL_SEL[89] shift_registerC_0/COL_SEL[90]
+ shift_registerC_0/COL_SEL[91] shift_registerC_0/COL_SEL[92] shift_registerC_0/COL_SEL[93]
+ shift_registerC_0/COL_SEL[94] shift_registerC_0/COL_SEL[95] shift_registerC_0/COL_SEL[96]
+ shift_registerC_0/COL_SEL[97] shift_registerC_0/COL_SEL[98] ARRAY_OUT shift_registerC_0/COL_SEL[99]
+ SF_IB VDD GND pixel_array100x100
Xshift_registerC_0 shift_registerC_0/COL_SEL[0] shift_registerC_0/COL_SEL[10] shift_registerC_0/COL_SEL[11]
+ shift_registerC_0/COL_SEL[12] shift_registerC_0/COL_SEL[13] shift_registerC_0/COL_SEL[14]
+ shift_registerC_0/COL_SEL[15] shift_registerC_0/COL_SEL[16] shift_registerC_0/COL_SEL[17]
+ shift_registerC_0/COL_SEL[18] shift_registerC_0/COL_SEL[19] shift_registerC_0/COL_SEL[1]
+ shift_registerC_0/COL_SEL[20] shift_registerC_0/COL_SEL[21] shift_registerC_0/COL_SEL[22]
+ shift_registerC_0/COL_SEL[23] shift_registerC_0/COL_SEL[24] shift_registerC_0/COL_SEL[25]
+ shift_registerC_0/COL_SEL[26] shift_registerC_0/COL_SEL[27] shift_registerC_0/COL_SEL[28]
+ shift_registerC_0/COL_SEL[29] shift_registerC_0/COL_SEL[2] shift_registerC_0/COL_SEL[30]
+ shift_registerC_0/COL_SEL[31] shift_registerC_0/COL_SEL[32] shift_registerC_0/COL_SEL[33]
+ shift_registerC_0/COL_SEL[34] shift_registerC_0/COL_SEL[35] shift_registerC_0/COL_SEL[36]
+ shift_registerC_0/COL_SEL[37] shift_registerC_0/COL_SEL[38] shift_registerC_0/COL_SEL[39]
+ shift_registerC_0/COL_SEL[3] shift_registerC_0/COL_SEL[40] shift_registerC_0/COL_SEL[41]
+ shift_registerC_0/COL_SEL[42] shift_registerC_0/COL_SEL[43] shift_registerC_0/COL_SEL[44]
+ shift_registerC_0/COL_SEL[45] shift_registerC_0/COL_SEL[46] shift_registerC_0/COL_SEL[47]
+ shift_registerC_0/COL_SEL[48] shift_registerC_0/COL_SEL[49] shift_registerC_0/COL_SEL[4]
+ shift_registerC_0/COL_SEL[50] shift_registerC_0/COL_SEL[51] shift_registerC_0/COL_SEL[52]
+ shift_registerC_0/COL_SEL[53] shift_registerC_0/COL_SEL[54] shift_registerC_0/COL_SEL[55]
+ shift_registerC_0/COL_SEL[56] shift_registerC_0/COL_SEL[57] shift_registerC_0/COL_SEL[58]
+ shift_registerC_0/COL_SEL[59] shift_registerC_0/COL_SEL[5] shift_registerC_0/COL_SEL[60]
+ shift_registerC_0/COL_SEL[61] shift_registerC_0/COL_SEL[62] shift_registerC_0/COL_SEL[63]
+ shift_registerC_0/COL_SEL[64] shift_registerC_0/COL_SEL[65] shift_registerC_0/COL_SEL[66]
+ shift_registerC_0/COL_SEL[67] shift_registerC_0/COL_SEL[68] shift_registerC_0/COL_SEL[69]
+ shift_registerC_0/COL_SEL[6] shift_registerC_0/COL_SEL[70] shift_registerC_0/COL_SEL[71]
+ shift_registerC_0/COL_SEL[72] shift_registerC_0/COL_SEL[73] shift_registerC_0/COL_SEL[74]
+ shift_registerC_0/COL_SEL[75] shift_registerC_0/COL_SEL[76] shift_registerC_0/COL_SEL[77]
+ shift_registerC_0/COL_SEL[78] shift_registerC_0/COL_SEL[79] shift_registerC_0/COL_SEL[7]
+ shift_registerC_0/COL_SEL[80] shift_registerC_0/COL_SEL[81] shift_registerC_0/COL_SEL[82]
+ shift_registerC_0/COL_SEL[83] shift_registerC_0/COL_SEL[84] shift_registerC_0/COL_SEL[85]
+ shift_registerC_0/COL_SEL[86] shift_registerC_0/COL_SEL[87] shift_registerC_0/COL_SEL[88]
+ shift_registerC_0/COL_SEL[89] shift_registerC_0/COL_SEL[8] shift_registerC_0/COL_SEL[90]
+ shift_registerC_0/COL_SEL[91] shift_registerC_0/COL_SEL[92] shift_registerC_0/COL_SEL[93]
+ shift_registerC_0/COL_SEL[94] shift_registerC_0/COL_SEL[95] shift_registerC_0/COL_SEL[96]
+ shift_registerC_0/COL_SEL[97] shift_registerC_0/COL_SEL[98] shift_registerC_0/COL_SEL[99]
+ shift_registerC_0/COL_SEL[9] COL_CLK COL_DIN COL_DOUT COL_ENA COL_RST VDD GND shift_registerC
Xshift_registerC_1 shift_registerC_1/COL_SEL[0] shift_registerC_1/COL_SEL[10] shift_registerC_1/COL_SEL[11]
+ shift_registerC_1/COL_SEL[12] shift_registerC_1/COL_SEL[13] shift_registerC_1/COL_SEL[14]
+ shift_registerC_1/COL_SEL[15] shift_registerC_1/COL_SEL[16] shift_registerC_1/COL_SEL[17]
+ shift_registerC_1/COL_SEL[18] shift_registerC_1/COL_SEL[19] shift_registerC_1/COL_SEL[1]
+ shift_registerC_1/COL_SEL[20] shift_registerC_1/COL_SEL[21] shift_registerC_1/COL_SEL[22]
+ shift_registerC_1/COL_SEL[23] shift_registerC_1/COL_SEL[24] shift_registerC_1/COL_SEL[25]
+ shift_registerC_1/COL_SEL[26] shift_registerC_1/COL_SEL[27] shift_registerC_1/COL_SEL[28]
+ shift_registerC_1/COL_SEL[29] shift_registerC_1/COL_SEL[2] shift_registerC_1/COL_SEL[30]
+ shift_registerC_1/COL_SEL[31] shift_registerC_1/COL_SEL[32] shift_registerC_1/COL_SEL[33]
+ shift_registerC_1/COL_SEL[34] shift_registerC_1/COL_SEL[35] shift_registerC_1/COL_SEL[36]
+ shift_registerC_1/COL_SEL[37] shift_registerC_1/COL_SEL[38] shift_registerC_1/COL_SEL[39]
+ shift_registerC_1/COL_SEL[3] shift_registerC_1/COL_SEL[40] shift_registerC_1/COL_SEL[41]
+ shift_registerC_1/COL_SEL[42] shift_registerC_1/COL_SEL[43] shift_registerC_1/COL_SEL[44]
+ shift_registerC_1/COL_SEL[45] shift_registerC_1/COL_SEL[46] shift_registerC_1/COL_SEL[47]
+ shift_registerC_1/COL_SEL[48] shift_registerC_1/COL_SEL[49] shift_registerC_1/COL_SEL[4]
+ shift_registerC_1/COL_SEL[50] shift_registerC_1/COL_SEL[51] shift_registerC_1/COL_SEL[52]
+ shift_registerC_1/COL_SEL[53] shift_registerC_1/COL_SEL[54] shift_registerC_1/COL_SEL[55]
+ shift_registerC_1/COL_SEL[56] shift_registerC_1/COL_SEL[57] shift_registerC_1/COL_SEL[58]
+ shift_registerC_1/COL_SEL[59] shift_registerC_1/COL_SEL[5] shift_registerC_1/COL_SEL[60]
+ shift_registerC_1/COL_SEL[61] shift_registerC_1/COL_SEL[62] shift_registerC_1/COL_SEL[63]
+ shift_registerC_1/COL_SEL[64] shift_registerC_1/COL_SEL[65] shift_registerC_1/COL_SEL[66]
+ shift_registerC_1/COL_SEL[67] shift_registerC_1/COL_SEL[68] shift_registerC_1/COL_SEL[69]
+ shift_registerC_1/COL_SEL[6] shift_registerC_1/COL_SEL[70] shift_registerC_1/COL_SEL[71]
+ shift_registerC_1/COL_SEL[72] shift_registerC_1/COL_SEL[73] shift_registerC_1/COL_SEL[74]
+ shift_registerC_1/COL_SEL[75] shift_registerC_1/COL_SEL[76] shift_registerC_1/COL_SEL[77]
+ shift_registerC_1/COL_SEL[78] shift_registerC_1/COL_SEL[79] shift_registerC_1/COL_SEL[7]
+ shift_registerC_1/COL_SEL[80] shift_registerC_1/COL_SEL[81] shift_registerC_1/COL_SEL[82]
+ shift_registerC_1/COL_SEL[83] shift_registerC_1/COL_SEL[84] shift_registerC_1/COL_SEL[85]
+ shift_registerC_1/COL_SEL[86] shift_registerC_1/COL_SEL[87] shift_registerC_1/COL_SEL[88]
+ shift_registerC_1/COL_SEL[89] shift_registerC_1/COL_SEL[8] shift_registerC_1/COL_SEL[90]
+ shift_registerC_1/COL_SEL[91] shift_registerC_1/COL_SEL[92] shift_registerC_1/COL_SEL[93]
+ shift_registerC_1/COL_SEL[94] shift_registerC_1/COL_SEL[95] shift_registerC_1/COL_SEL[96]
+ shift_registerC_1/COL_SEL[97] shift_registerC_1/COL_SEL[98] shift_registerC_1/COL_SEL[99]
+ shift_registerC_1/COL_SEL[9] ROW_CLK ROW_DIN shift_registerC_1/data_out ROW_ENA
+ ROW_RST VDD GND shift_registerC
.ends

.subckt sky130_fd_pr__pfet_01v8_YT7TV5 a_n505_21# a_n387_21# a_384_118# w_n1642_n937#
+ a_n623_21# a_620_118# a_n387_n815# a_n1150_118# a_n33_n815# a_n741_21# a_321_n815#
+ a_n560_n718# a_675_n815# a_1092_n718# a_n1331_n815# a_n1449_21# a_n914_n718# a_1446_n718#
+ a_1029_n815# a_n151_21# a_n560_118# a_1092_118# a_n269_n815# a_620_n718# a_1328_118#
+ a_30_118# a_203_n815# a_974_n718# a_n442_n718# a_557_n815# a_n796_n718# a_439_21#
+ a_n1213_n815# a_n1213_21# a_n1095_21# a_557_21# a_1328_n718# a_n1331_21# a_n206_118#
+ a_675_21# a_738_118# a_911_21# a_n1268_118# a_793_21# a_n1504_118# a_502_n718# a_n1095_n815#
+ a_856_n718# a_85_n815# a_n324_n718# a_439_n815# a_203_21# a_n678_n718# a_148_118#
+ a_n1449_n815# a_321_21# a_n678_118# a_n33_21# a_n914_118# a_1446_118# a_384_n718#
+ a_1029_21# a_n741_n815# a_30_n718# a_1147_21# a_738_n718# a_n206_n718# a_n324_118#
+ a_1265_21# a_n1150_n718# a_856_118# a_1383_n815# a_1383_21# a_n1386_118# a_n1504_n718#
+ a_266_n718# a_n88_118# a_266_118# a_n623_n815# a_n977_n815# a_502_118# a_n796_118#
+ a_n88_n718# a_n1032_118# a_911_n815# a_n1032_n718# a_1265_n815# a_n1386_n718# a_n151_n815#
+ a_n859_21# a_148_n718# a_n442_118# a_974_118# a_n505_n815# a_n977_21# a_1210_118#
+ a_793_n815# a_n859_n815# a_85_21# a_1210_n718# a_n269_21# a_1147_n815# a_n1268_n718#
X0 a_1446_118# a_1383_21# a_1328_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X1 a_n1032_n718# a_n1095_n815# a_n1150_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_n796_118# a_n859_21# a_n914_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_384_118# a_321_21# a_266_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_384_n718# a_321_n815# a_266_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_n88_n718# a_n151_n815# a_n206_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 a_1328_118# a_1265_21# a_1210_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X7 a_n1150_n718# a_n1213_n815# a_n1268_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_n678_118# a_n741_21# a_n796_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 a_1210_n718# a_1147_n815# a_1092_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_266_118# a_203_21# a_148_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_30_n718# a_n33_n815# a_n88_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_1210_118# a_1147_21# a_1092_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X13 a_n914_n718# a_n977_n815# a_n1032_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_n560_n718# a_n623_n815# a_n678_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 a_1446_n718# a_1383_n815# a_1328_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X16 a_n560_118# a_n623_21# a_n678_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 a_266_n718# a_203_n815# a_148_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X18 a_620_n718# a_557_n815# a_502_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 a_n1386_118# a_n1449_21# a_n1504_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X20 a_n324_118# a_n387_21# a_n442_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 a_856_118# a_793_21# a_738_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 a_1092_118# a_1029_21# a_974_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 a_n324_n718# a_n387_n815# a_n442_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 a_n442_118# a_n505_21# a_n560_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X25 a_148_118# a_85_21# a_30_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 a_n1386_n718# a_n1449_n815# a_n1504_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X27 a_856_n718# a_793_n815# a_738_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 a_974_118# a_911_21# a_856_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 a_1092_n718# a_1029_n815# a_974_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X30 a_n1268_118# a_n1331_21# a_n1386_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X31 a_n206_118# a_n269_21# a_n324_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X32 a_738_118# a_675_21# a_620_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X33 a_n796_n718# a_n859_n815# a_n914_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X34 a_n1032_118# a_n1095_21# a_n1150_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X35 a_148_n718# a_85_n815# a_30_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X36 a_1328_n718# a_1265_n815# a_1210_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X37 a_n88_118# a_n151_21# a_n206_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X38 a_30_118# a_n33_21# a_n88_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X39 a_620_118# a_557_21# a_502_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X40 a_502_n718# a_439_n815# a_384_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X41 a_n1150_118# a_n1213_21# a_n1268_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X42 a_n206_n718# a_n269_n815# a_n324_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X43 a_738_n718# a_675_n815# a_620_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X44 a_n1268_n718# a_n1331_n815# a_n1386_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X45 a_n914_118# a_n977_21# a_n1032_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X46 a_n442_n718# a_n505_n815# a_n560_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X47 a_502_118# a_439_21# a_384_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X48 a_974_n718# a_911_n815# a_856_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X49 a_n678_n718# a_n741_n815# a_n796_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_8HUREQ a_384_n709# a_557_n797# a_203_n797# a_n387_21#
+ a_n505_21# a_30_n709# a_n623_21# a_738_n709# a_n206_n709# a_n741_21# a_n324_109#
+ a_856_109# a_85_n797# a_n151_21# a_266_n709# a_439_n797# a_n88_109# a_266_109# a_n88_n709#
+ a_502_109# a_n796_109# a_439_21# a_n741_n797# a_557_21# a_148_n709# a_675_21# a_n442_109#
+ a_793_21# a_203_21# a_n623_n797# a_321_21# a_620_109# a_384_109# a_n33_21# a_n560_n709#
+ a_n151_n797# a_n914_n709# a_n1016_n883# a_793_n797# a_n505_n797# a_n859_n797# a_n560_109#
+ a_620_n709# a_n442_n709# a_30_109# a_n796_n709# a_n387_n797# a_321_n797# a_n33_n797#
+ a_n206_109# a_675_n797# a_738_109# a_502_n709# a_n859_21# a_856_n709# a_n324_n709#
+ a_n678_n709# a_148_109# a_85_21# a_n269_n797# a_n678_109# a_n914_109# a_n269_21#
X0 a_n678_109# a_n741_21# a_n796_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X1 a_266_109# a_203_21# a_148_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_30_n709# a_n33_n797# a_n88_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_n560_n709# a_n623_n797# a_n678_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_n560_109# a_n623_21# a_n678_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_n324_109# a_n387_21# a_n442_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 a_266_n709# a_203_n797# a_148_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X7 a_620_n709# a_557_n797# a_502_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_856_109# a_793_21# a_738_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X9 a_n324_n709# a_n387_n797# a_n442_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_n442_109# a_n505_21# a_n560_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_148_109# a_85_21# a_30_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_856_n709# a_793_n797# a_738_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X13 a_n206_109# a_n269_21# a_n324_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_738_109# a_675_21# a_620_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 a_n796_n709# a_n859_n797# a_n914_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X16 a_148_n709# a_85_n797# a_30_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 a_620_109# a_557_21# a_502_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X18 a_n88_109# a_n151_21# a_n206_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 a_30_109# a_n33_21# a_n88_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X20 a_502_n709# a_439_n797# a_384_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 a_n206_n709# a_n269_n797# a_n324_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 a_738_n709# a_675_n797# a_620_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 a_n442_n709# a_n505_n797# a_n560_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 a_502_109# a_439_21# a_384_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X25 a_n678_n709# a_n741_n797# a_n796_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 a_n796_109# a_n859_21# a_n914_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X27 a_384_109# a_321_21# a_266_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 a_384_n709# a_321_n797# a_266_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 a_n88_n709# a_n151_n797# a_n206_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_BLS9H9 m3_n1941_n1600# c1_n1841_n1500#
X0 c1_n1841_n1500# m3_n1941_n1600# sky130_fd_pr__cap_mim_m3_1 l=15 w=17.55
.ends

.subckt sky130_fd_pr__pfet_01v8_YC9MKB a_856_n300# a_n324_n300# a_n505_n397# a_n678_n300#
+ a_793_n397# a_n859_n397# a_384_n300# a_n387_n397# a_30_n300# a_321_n397# a_n33_n397#
+ a_738_n300# a_n206_n300# a_675_n397# a_266_n300# a_n269_n397# a_n88_n300# a_203_n397#
+ a_557_n397# a_148_n300# a_439_n397# a_85_n397# w_n1052_n519# a_n560_n300# a_n741_n397#
+ a_n914_n300# a_620_n300# a_n442_n300# a_n796_n300# a_n623_n397# a_n151_n397# a_502_n300#
X0 a_n560_n300# a_n623_n397# a_n678_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X1 a_30_n300# a_n33_n397# a_n88_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_266_n300# a_203_n397# a_148_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_620_n300# a_557_n397# a_502_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_n324_n300# a_n387_n397# a_n442_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_856_n300# a_793_n397# a_738_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X6 a_n796_n300# a_n859_n397# a_n914_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X7 a_148_n300# a_85_n397# a_30_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_502_n300# a_439_n397# a_384_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 a_n206_n300# a_n269_n397# a_n324_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_738_n300# a_675_n397# a_620_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_n442_n300# a_n505_n397# a_n560_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_n678_n300# a_n741_n397# a_n796_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X13 a_384_n300# a_321_n397# a_266_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_n88_n300# a_n151_n397# a_n206_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_GQFJAV a_15_n75# a_n69_97# a_n175_n249# a_n73_n75#
X0 a_15_n75# a_n69_97# a_n73_n75# a_n175_n249# sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_YCMRKB a_n1390_n815# a_89_n718# a_1678_21# a_915_118#
+ a_1151_n718# a_1914_21# a_n2216_21# a_734_n815# a_n2153_n718# a_380_21# a_n2098_21#
+ a_2032_n815# a_n973_n718# a_n1445_118# a_1796_21# a_1977_118# a_n92_21# a_2386_n815#
+ a_n1744_n815# a_1088_n815# a_n2334_21# w_n3117_n937# a_2803_n718# a_1206_21# a_1505_n718#
+ a_n2507_n718# a_n1209_n718# a_1088_21# a_1859_n718# a_2213_118# a_n2452_21# a_325_118#
+ a_1324_21# a_262_n815# a_n855_118# a_n2743_118# a_n2570_21# a_n328_n815# a_1387_118#
+ a_1442_21# a_1623_118# a_n2570_n815# a_n1272_n815# a_n501_n718# a_1033_n718# a_2331_n718#
+ a_1560_21# a_616_n815# a_n2035_n718# a_89_118# a_n855_n718# a_2685_n718# a_1387_n718#
+ a_2268_n815# a_n2389_n718# a_n2924_n815# a_n1626_n815# a_2685_118# a_n265_118# a_n2153_118#
+ a_797_118# a_n501_118# a_2921_118# a_1033_118# a_2858_21# a_561_n718# a_144_n815#
+ a_n1563_118# a_n383_n718# a_498_n815# a_n2452_n815# a_n1154_n815# a_915_n718# a_2095_118#
+ a_2213_n718# a_2268_21# a_n918_21# a_2331_118# a_n737_n718# a_2567_n718# a_1269_n718#
+ a_443_118# a_n2806_n815# a_2504_21# a_n1508_n815# a_n1681_n718# a_2386_21# a_26_21#
+ a_1560_n815# a_n973_118# a_n2861_118# a_2622_21# a_1741_118# a_1914_n815# a_443_n718#
+ a_n328_21# a_2740_21# a_797_n718# a_n1209_118# a_n800_n815# a_n265_n718# a_2095_n718#
+ a_n446_21# a_n2334_n815# a_n1036_n815# a_n383_118# a_n2271_118# a_n2688_n815# a_2032_21#
+ a_26_n815# a_1151_118# a_n564_21# a_n619_n718# a_2449_n718# a_2150_21# a_n800_21#
+ a_2740_n815# a_n2861_n718# a_n1563_n718# a_1442_n815# a_n619_118# a_n1681_118# a_n682_21#
+ a_n2507_118# a_1796_n815# a_n1508_21# a_n682_n815# a_n1917_n718# a_325_n718# a_n1626_21#
+ a_679_n718# a_n1917_118# a_n210_21# a_n147_n718# a_561_118# a_n2216_n815# a_970_n815#
+ a_n1744_21# a_n1091_n718# a_n1091_118# a_2449_118# a_n1980_n815# a_n1862_21# a_1741_n718#
+ a_n2979_118# a_n1036_21# a_2622_n815# a_n2743_n718# a_n1445_n718# a_1324_n815# a_1859_118#
+ a_n1327_118# a_n1980_21# a_1678_n815# a_n1799_n718# a_n1154_21# a_n210_n815# a_n564_n815#
+ a_207_n718# a_616_21# a_n2098_n815# a_n1272_21# a_n29_118# a_498_21# a_207_118#
+ a_n2389_118# a_734_21# a_852_n815# a_n2271_n718# a_n1390_21# a_n918_n815# a_2150_n815#
+ a_n737_118# a_n2625_118# a_n29_n718# a_1269_118# a_n1862_n815# a_1505_118# a_852_21#
+ a_2921_n718# a_1623_n718# a_n1799_118# a_2504_n815# a_n2625_n718# a_n1327_n718#
+ a_1206_n815# a_1977_n718# a_970_21# a_n2806_21# a_n2979_n718# a_n2688_21# a_2858_n815#
+ a_144_21# a_n92_n815# a_380_n815# a_n147_118# a_n2035_118# a_n2924_21# a_n446_n815#
+ a_2567_118# a_2803_118# a_679_118# a_262_21#
X0 a_561_n718# a_498_n815# a_443_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X1 a_n383_118# a_n446_21# a_n501_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_n265_n718# a_n328_n815# a_n383_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_n1445_118# a_n1508_21# a_n1563_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_915_118# a_852_21# a_797_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_n2625_n718# a_n2688_n815# a_n2743_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 a_1151_n718# a_1088_n815# a_1033_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X7 a_n2153_118# a_n2216_21# a_n2271_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_797_n718# a_734_n815# a_679_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 a_2803_118# a_2740_21# a_2685_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_2331_n718# a_2268_n815# a_2213_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_n29_118# a_n92_21# a_n147_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_n1681_n718# a_n1744_n815# a_n1799_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X13 a_n1209_118# a_n1272_21# a_n1327_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_1859_118# a_1796_21# a_1741_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 a_n2861_n718# a_n2924_n815# a_n2979_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X16 a_n265_118# a_n328_21# a_n383_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 a_n1917_n718# a_n1980_n815# a_n2035_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X18 a_n2035_n718# a_n2098_n815# a_n2153_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 a_797_118# a_734_21# a_679_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X20 a_1977_118# a_1914_21# a_1859_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 a_1269_n718# a_1206_n815# a_1151_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 a_1623_n718# a_1560_n815# a_1505_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 a_207_n718# a_144_n815# a_89_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 a_89_n718# a_26_n815# a_n29_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X25 a_n1091_118# a_n1154_21# a_n1209_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 a_2685_118# a_2622_21# a_2567_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X27 a_1741_118# a_1678_21# a_1623_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 a_2803_n718# a_2740_n815# a_2685_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 a_n1091_n718# a_n1154_n815# a_n1209_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X30 a_89_118# a_26_21# a_n29_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X31 a_n2271_n718# a_n2334_n815# a_n2389_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X32 a_1859_n718# a_1796_n815# a_1741_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X33 a_2449_118# a_2386_21# a_2331_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X34 a_n1327_n718# a_n1390_n815# a_n1445_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X35 a_n147_118# a_n210_21# a_n265_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X36 a_n147_n718# a_n210_n815# a_n265_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X37 a_n2861_118# a_n2924_21# a_n2979_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X38 a_n501_n718# a_n564_n815# a_n619_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X39 a_n2507_n718# a_n2570_n815# a_n2625_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X40 a_679_118# a_616_21# a_561_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X41 a_443_118# a_380_21# a_325_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X42 a_n973_118# a_n1036_21# a_n1091_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X43 a_n1917_118# a_n1980_21# a_n2035_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X44 a_679_n718# a_616_n815# a_561_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X45 a_1623_118# a_1560_21# a_1505_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X46 a_2213_n718# a_2150_n815# a_2095_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X47 a_2567_118# a_2504_21# a_2449_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X48 a_1033_n718# a_970_n815# a_915_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X49 a_n2625_118# a_n2688_21# a_n2743_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X50 a_n1563_n718# a_n1626_n815# a_n1681_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X51 a_n737_n718# a_n800_n815# a_n855_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X52 a_2331_118# a_2268_21# a_2213_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X53 a_n2743_n718# a_n2806_n815# a_n2861_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X54 a_2449_n718# a_2386_n815# a_2331_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X55 a_561_118# a_498_21# a_443_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X56 a_n1799_n718# a_n1862_n815# a_n1917_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X57 a_n2743_118# a_n2806_21# a_n2861_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X58 a_n737_118# a_n800_21# a_n855_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X59 a_1505_n718# a_1442_n815# a_1387_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X60 a_n1799_118# a_n1862_21# a_n1917_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X61 a_325_118# a_262_21# a_207_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X62 a_443_n718# a_380_n815# a_325_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X63 a_1505_118# a_1442_21# a_1387_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X64 a_2685_n718# a_2622_n815# a_2567_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X65 a_n973_n718# a_n1036_n815# a_n1091_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X66 a_n2507_118# a_n2570_21# a_n2625_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X67 a_n2153_n718# a_n2216_n815# a_n2271_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X68 a_2213_118# a_2150_21# a_2095_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X69 a_n855_118# a_n918_21# a_n973_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X70 a_n1209_n718# a_n1272_n815# a_n1327_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X71 a_n383_n718# a_n446_n815# a_n501_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X72 a_n2389_n718# a_n2452_n815# a_n2507_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X73 a_n1681_118# a_n1744_21# a_n1799_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X74 a_n619_118# a_n682_21# a_n737_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X75 a_1977_n718# a_1914_n815# a_1859_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X76 a_207_118# a_144_21# a_89_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X77 a_2095_n718# a_2032_n815# a_1977_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X78 a_1387_118# a_1324_21# a_1269_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X79 a_915_n718# a_852_n815# a_797_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X80 a_n29_n718# a_n92_n815# a_n147_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X81 a_n1445_n718# a_n1508_n815# a_n1563_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X82 a_n619_n718# a_n682_n815# a_n737_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X83 a_n2389_118# a_n2452_21# a_n2507_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X84 a_2095_118# a_2032_21# a_1977_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X85 a_1151_118# a_1088_21# a_1033_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X86 a_n501_118# a_n564_21# a_n619_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X87 a_1033_118# a_970_21# a_915_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X88 a_n1563_118# a_n1626_21# a_n1681_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X89 a_n855_n718# a_n918_n815# a_n973_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X90 a_1387_n718# a_1324_n815# a_1269_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X91 a_n2271_118# a_n2334_21# a_n2389_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X92 a_1741_n718# a_1678_n815# a_1623_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X93 a_325_n718# a_262_n815# a_207_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X94 a_2921_118# a_2858_21# a_2803_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X95 a_1269_118# a_1206_21# a_1151_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X96 a_2567_n718# a_2504_n815# a_2449_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X97 a_2921_n718# a_2858_n815# a_2803_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X98 a_n1327_118# a_n1390_21# a_n1445_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X99 a_n2035_118# a_n2098_21# a_n2153_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_8JUMX6 a_2117_109# a_n399_n1009# a_1879_n1097# a_5225_109#
+ a_3301_109# a_3803_21# a_547_21# a_785_n1009# a_1377_n1009# a_n193_21# a_n2027_109#
+ a_n3301_21# a_n3597_n1097# a_n3211_109# a_n5135_109# a_2767_n1097# a_4189_n1009#
+ a_3893_109# a_4395_21# a_n1673_n1097# a_2265_n1009# a_4691_n1097# a_n103_109# a_637_n1009#
+ a_n4485_n1097# a_4247_21# a_1229_n1009# a_3655_n1097# a_5077_n1009# a_n2561_n1097#
+ a_785_109# a_3655_21# a_399_21# a_n251_n1009# a_1731_n1097# a_n3449_n1097# a_1969_109#
+ a_2619_n1097# a_3153_n1009# a_n1525_n1097# a_n695_109# a_n3153_21# a_2117_n1009#
+ a_n5373_n1097# a_4543_n1097# a_3507_21# a_n2561_21# a_n4929_21# a_n1879_109# a_n4337_n1097#
+ a_5077_109# a_n4987_109# a_2915_21# a_n3005_21# a_3507_n1097# a_4041_n1009# a_3153_109#
+ a_n1583_n1009# a_n103_n1009# a_n2413_n1097# a_4099_21# a_n2413_21# a_3005_n1009#
+ a_n933_n1097# a_5431_n1097# a_n1821_21# a_n5225_n1097# a_n4395_n1009# a_n3063_109#
+ a_1969_n1009# a_399_n1097# a_n3301_n1097# a_n2471_n1009# a_1229_109# a_n3359_n1009#
+ a_n991_n1009# a_4337_109# a_2413_109# a_3359_21# a_3893_n1009# a_5521_109# a_n1435_n1009#
+ a_2767_21# a_n5283_n1009# a_2857_n1009# a_n1139_109# a_n2265_21# a_n4247_n1009#
+ a_n2323_109# a_n4247_109# a_n5431_109# a_2619_21# a_n1673_21# a_n2323_n1009# a_4781_n1009#
+ a_n843_n1009# a_n2117_21# a_3745_n1009# a_n45_n1097# a_n1525_21# a_n5135_n1009#
+ a_1821_n1009# a_251_n1097# a_45_109# a_2709_n1009# a_n193_n1097# a_1081_109# a_n3211_n1009#
+ a_n3507_109# a_n4929_n1097# a_4633_n1009# a_n991_109# a_n5521_21# a_103_n1097# a_4189_109#
+ a_1879_21# a_251_21# a_n4987_n1009# a_2265_109# a_5521_n1009# a_5373_109# a_n1377_21#
+ a_489_n1009# a_103_21# a_n4099_109# a_n2175_109# a_991_n1097# a_n5283_109# a_n45_21#
+ a_n1229_21# a_1583_n1097# a_341_109# a_n3951_n1009# a_n1377_n1097# a_3449_109# a_1525_109#
+ a_n4839_n1009# a_1081_n1009# a_4633_109# a_n933_21# a_n5373_21# a_n251_109# a_4395_n1097#
+ a_n2915_n1009# a_n4781_21# a_n4189_n1097# a_3359_n1097# a_2471_n1097# a_n1435_109#
+ a_n3359_109# a_n5225_21# a_843_n1097# a_n2265_n1097# a_n4543_109# a_1435_n1097#
+ a_n785_n1097# a_3211_21# a_n4633_21# a_5283_n1097# a_n3803_n1009# a_2709_109# a_341_n1009#
+ a_n1229_n1097# a_n5077_n1097# a_4247_n1097# a_n3153_n1097# a_n785_21# a_2323_n1097#
+ a_n2619_109# a_n2117_n1097# a_n1287_n1009# a_n637_n1097# a_n3803_109# a_4987_21#
+ a_n5077_21# a_5135_n1097# a_n637_21# a_n4041_n1097# a_193_109# a_3063_21# a_n4485_21#
+ a_3211_n1097# a_n4099_n1009# a_n3005_n1097# a_1377_109# a_2471_21# a_n3893_21# a_n2175_n1009#
+ a_4485_109# a_2561_109# a_4839_21# a_n695_n1009# a_n1139_n1009# a_45_n1009# a_3597_n1009#
+ a_n4337_21# a_n1969_n1097# a_2323_21# a_1673_n1009# a_n1287_109# a_n3745_21# a_4987_n1097#
+ a_n2471_109# a_n4395_109# a_1731_21# a_n5681_n1183# a_n3063_n1009# a_n3893_n1097#
+ a_n489_21# a_4485_n1009# a_n2027_n1009# a_3745_109# a_n547_n1009# a_2561_n1009#
+ a_n2857_n1097# a_1821_109# a_3449_n1009# a_933_n1009# a_1525_n1009# a_n4781_n1097#
+ a_3951_n1097# a_4839_n1097# a_5373_n1009# a_n3655_109# a_n5579_109# a_n4189_21#
+ a_n3745_n1097# a_637_109# a_n1731_109# a_2175_21# a_2915_n1097# a_n3597_21# a_4337_n1009#
+ a_n1821_n1097# a_4929_109# a_1583_21# a_n1879_n1009# a_n2709_n1097# a_n547_109#
+ a_2413_n1009# a_2027_21# a_n1081_21# a_n3449_21# a_n4633_n1097# a_3803_n1097# a_5225_n1009#
+ a_n4839_109# a_1435_21# a_n2857_21# a_3005_109# a_n2915_109# a_n2767_n1009# a_3301_n1009#
+ a_n4691_n1009# a_n5521_n1097# a_n2709_21# a_n5579_n1009# a_695_n1097# a_1287_n1097#
+ a_3597_109# a_1673_109# a_5431_21# a_n3655_n1009# a_193_n1009# a_4781_109# a_4099_n1097#
+ a_n2619_n1009# a_n1731_n1009# a_1287_21# a_991_21# a_2175_n1097# a_489_109# a_n1583_109#
+ a_n1081_n1097# a_n4691_109# a_n4543_n1009# a_547_n1097# a_1139_n1097# a_n489_n1097#
+ a_2857_109# a_n399_109# a_1139_21# a_843_21# a_n3507_n1009# a_3063_n1097# a_4929_n1009#
+ a_5283_21# a_n1969_21# a_n5431_n1009# a_n2767_109# a_4691_21# a_2027_n1097# a_n341_21#
+ a_4041_109# a_933_109# a_n3951_109# a_5135_21# a_n843_109# a_4543_21# a_695_21#
+ a_3951_21# a_n4041_21# a_n341_n1097#
X0 a_n4099_109# a_n4189_21# a_n4247_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X1 a_489_n1009# a_399_n1097# a_341_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X2 a_n843_n1009# a_n933_n1097# a_n991_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X3 a_n1731_n1009# a_n1821_n1097# a_n1879_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X4 a_3597_109# a_3507_21# a_3449_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X5 a_n1287_109# a_n1377_21# a_n1435_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X6 a_4633_109# a_4543_21# a_4485_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X7 a_4485_n1009# a_4395_n1097# a_4337_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X8 a_489_109# a_399_21# a_341_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X9 a_2709_109# a_2619_21# a_2561_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X10 a_1821_109# a_1731_21# a_1673_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X11 a_n2027_n1009# a_n2117_n1097# a_n2175_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X12 a_n547_n1009# a_n637_n1097# a_n695_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X13 a_n1435_n1009# a_n1525_n1097# a_n1583_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X14 a_3745_109# a_3655_21# a_3597_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X15 a_4781_109# a_4691_21# a_4633_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X16 a_4189_n1009# a_4099_n1097# a_4041_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X17 a_2857_109# a_2767_21# a_2709_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X18 a_n4839_109# a_n4929_21# a_n4987_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X19 a_5077_n1009# a_4987_n1097# a_4929_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X20 a_n1139_n1009# a_n1229_n1097# a_n1287_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X21 a_1969_109# a_1879_21# a_1821_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X22 a_n2619_n1009# a_n2709_n1097# a_n2767_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X23 a_193_n1009# a_103_n1097# a_45_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X24 a_n3951_n1009# a_n4041_n1097# a_n4099_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X25 a_n5431_n1009# a_n5521_n1097# a_n5579_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=0.45
X26 a_n547_109# a_n637_21# a_n695_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X27 a_45_109# a_n45_21# a_n103_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X28 a_2117_109# a_2027_21# a_1969_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X29 a_3153_109# a_3063_21# a_3005_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X30 a_n3211_109# a_n3301_21# a_n3359_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X31 a_45_n1009# a_n45_n1097# a_n103_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X32 a_n5135_n1009# a_n5225_n1097# a_n5283_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X33 a_n103_n1009# a_n193_n1097# a_n251_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X34 a_n991_n1009# a_n1081_n1097# a_n1139_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X35 a_n3063_n1009# a_n3153_n1097# a_n3211_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X36 a_n5135_109# a_n5225_21# a_n5283_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X37 a_1229_109# a_1139_21# a_1081_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X38 a_n2471_n1009# a_n2561_n1097# a_n2619_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X39 a_n4543_n1009# a_n4633_n1097# a_n4691_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X40 a_n695_109# a_n785_21# a_n843_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X41 a_3301_n1009# a_3211_n1097# a_3153_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X42 a_2265_109# a_2175_21# a_2117_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X43 a_n2323_109# a_n2413_21# a_n2471_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X44 a_4189_109# a_4099_21# a_4041_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X45 a_n4247_109# a_n4337_21# a_n4395_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X46 a_n5283_109# a_n5373_21# a_n5431_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X47 a_1377_109# a_1287_21# a_1229_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X48 a_n4247_n1009# a_n4337_n1097# a_n4395_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X49 a_n1435_109# a_n1525_21# a_n1583_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X50 a_n2175_n1009# a_n2265_n1097# a_n2323_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X51 a_n3359_109# a_n3449_21# a_n3507_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X52 a_n3655_n1009# a_n3745_n1097# a_n3803_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X53 a_n2471_109# a_n2561_21# a_n2619_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X54 a_n695_n1009# a_n785_n1097# a_n843_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X55 a_n1583_n1009# a_n1673_n1097# a_n1731_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X56 a_637_109# a_547_21# a_489_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X57 a_2413_n1009# a_2323_n1097# a_2265_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X58 a_n4395_109# a_n4485_21# a_n4543_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X59 a_3893_n1009# a_3803_n1097# a_3745_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X60 a_1821_n1009# a_1731_n1097# a_1673_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X61 a_3893_109# a_3803_21# a_3745_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X62 a_n1583_109# a_n1673_21# a_n1731_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X63 a_n3507_109# a_n3597_21# a_n3655_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X64 a_785_109# a_695_21# a_637_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X65 a_n3359_n1009# a_n3449_n1097# a_n3507_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X66 a_3005_109# a_2915_21# a_2857_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X67 a_n399_n1009# a_n489_n1097# a_n547_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X68 a_n1287_n1009# a_n1377_n1097# a_n1435_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X69 a_n4839_n1009# a_n4929_n1097# a_n4987_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X70 a_2117_n1009# a_2027_n1097# a_1969_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X71 a_341_n1009# a_251_n1097# a_193_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X72 a_n2767_n1009# a_n2857_n1097# a_n2915_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X73 a_4929_109# a_4839_21# a_4781_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X74 a_4041_109# a_3951_21# a_3893_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X75 a_n103_109# a_n193_21# a_n251_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X76 a_3597_n1009# a_3507_n1097# a_3449_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X77 a_1525_n1009# a_1435_n1097# a_1377_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X78 a_3005_n1009# a_2915_n1097# a_2857_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X79 a_5077_109# a_4987_21# a_4929_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X80 a_1229_n1009# a_1139_n1097# a_1081_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X81 a_n1879_n1009# a_n1969_n1097# a_n2027_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X82 a_2709_n1009# a_2619_n1097# a_2561_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X83 a_n5283_n1009# a_n5373_n1097# a_n5431_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X84 a_933_n1009# a_843_n1097# a_785_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X85 a_n4691_n1009# a_n4781_n1097# a_n4839_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X86 a_5521_n1009# a_5431_n1097# a_5373_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=0.45
X87 a_3301_109# a_3211_21# a_3153_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X88 a_5225_109# a_5135_21# a_5077_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X89 a_n991_109# a_n1081_21# a_n1139_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X90 a_n843_109# a_n933_21# a_n991_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X91 a_2413_109# a_2323_21# a_2265_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X92 a_n4987_n1009# a_n5077_n1097# a_n5135_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X93 a_637_n1009# a_547_n1097# a_489_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X94 a_4337_109# a_4247_21# a_4189_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X95 a_n4395_n1009# a_n4485_n1097# a_n4543_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X96 a_5225_n1009# a_5135_n1097# a_5077_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X97 a_3153_n1009# a_3063_n1097# a_3005_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X98 a_n3803_n1009# a_n3893_n1097# a_n3951_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X99 a_5373_109# a_5283_21# a_5225_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X100 a_n5431_109# a_n5521_21# a_n5579_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=0.45
X101 a_1525_109# a_1435_21# a_1377_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X102 a_4633_n1009# a_4543_n1097# a_4485_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X103 a_2561_n1009# a_2471_n1097# a_2413_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X104 a_4041_n1009# a_3951_n1097# a_3893_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X105 a_3449_109# a_3359_21# a_3301_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X106 a_2561_109# a_2471_21# a_2413_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X107 a_4485_109# a_4395_21# a_4337_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X108 a_n4543_109# a_n4633_21# a_n4691_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X109 a_n4099_n1009# a_n4189_n1097# a_n4247_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X110 a_1673_109# a_1583_21# a_1525_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X111 a_n3507_n1009# a_n3597_n1097# a_n3655_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X112 a_n2619_109# a_n2709_21# a_n2767_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X113 a_n1731_109# a_n1821_21# a_n1879_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X114 a_4337_n1009# a_4247_n1097# a_4189_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X115 a_2265_n1009# a_2175_n1097# a_2117_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X116 a_n3655_109# a_n3745_21# a_n3803_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X117 a_3745_n1009# a_3655_n1097# a_3597_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X118 a_933_109# a_843_21# a_785_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X119 a_1673_n1009# a_1583_n1097# a_1525_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X120 a_n4691_109# a_n4781_21# a_n4839_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X121 a_n251_109# a_n341_21# a_n399_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X122 a_n2767_109# a_n2857_21# a_n2915_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X123 a_n3803_109# a_n3893_21# a_n3951_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X124 a_1081_109# a_991_21# a_933_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X125 a_3449_n1009# a_3359_n1097# a_3301_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X126 a_4929_n1009# a_4839_n1097# a_4781_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X127 a_1377_n1009# a_1287_n1097# a_1229_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X128 a_n1879_109# a_n1969_21# a_n2027_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X129 a_2857_n1009# a_2767_n1097# a_2709_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X130 a_1081_n1009# a_991_n1097# a_933_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X131 a_n2915_109# a_n3005_21# a_n3063_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X132 a_193_109# a_103_21# a_45_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X133 a_n3951_109# a_n4041_21# a_n4099_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X134 a_n399_109# a_n489_21# a_n547_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X135 a_n3211_n1009# a_n3301_n1097# a_n3359_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X136 a_n251_n1009# a_n341_n1097# a_n399_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X137 a_n2027_109# a_n2117_21# a_n2175_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X138 a_785_n1009# a_695_n1097# a_637_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X139 a_1969_n1009# a_1879_n1097# a_1821_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X140 a_n3063_109# a_n3153_21# a_n3211_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X141 a_5373_n1009# a_5283_n1097# a_5225_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X142 a_341_109# a_251_21# a_193_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X143 a_n4987_109# a_n5077_21# a_n5135_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X144 a_4781_n1009# a_4691_n1097# a_4633_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X145 a_n1139_109# a_n1229_21# a_n1287_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X146 a_n2915_n1009# a_n3005_n1097# a_n3063_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X147 a_n2175_109# a_n2265_21# a_n2323_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X148 a_5521_109# a_5431_21# a_5373_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=0.45
X149 a_n2323_n1009# a_n2413_n1097# a_n2471_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
.ends

.subckt opamp_v1 iref vin_n vin_p vout vdd vss a_4019_n9933#
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[0] iref iref vdd vdd iref vdd iref vout iref iref
+ iref vdd iref vdd iref iref vout vout iref iref vdd vdd iref vdd vdd vout iref vout
+ vout iref vdd iref iref iref iref iref vdd iref vout iref vout iref vdd iref vdd
+ vout iref vdd iref vdd iref iref vout vdd iref iref vout iref vout vout vdd iref
+ iref vout iref vout vout vdd iref vout vdd iref iref vout vdd vout vdd vout iref
+ iref vout vdd vdd vdd iref vdd iref vout iref iref vdd vout vout iref iref vout
+ iref iref iref vout iref iref vdd sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[1] iref iref vdd vdd iref vdd iref vout iref iref
+ iref vdd iref vdd iref iref vout vout iref iref vdd vdd iref vdd vdd vout iref vout
+ vout iref vdd iref iref iref iref iref vdd iref vout iref vout iref vdd iref vdd
+ vout iref vdd iref vdd iref iref vout vdd iref iref vout iref vout vout vdd iref
+ iref vout iref vout vout vdd iref vout vdd iref iref vout vdd vout vdd vout iref
+ iref vout vdd vdd vdd iref vdd iref vout iref iref vdd vout vout iref iref vout
+ iref iref iref vout iref iref vdd sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[2] iref iref vdd vdd iref vdd iref vout iref iref
+ iref vdd iref vdd iref iref vout vout iref iref vdd vdd iref vdd vdd vout iref vout
+ vout iref vdd iref iref iref iref iref vdd iref vout iref vout iref vdd iref vdd
+ vout iref vdd iref vdd iref iref vout vdd iref iref vout iref vout vout vdd iref
+ iref vout iref vout vout vdd iref vout vdd iref iref vout vdd vout vdd vout iref
+ iref vout vdd vdd vdd iref vdd iref vout iref iref vdd vout vout iref iref vout
+ iref iref iref vout iref iref vdd sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__nfet_01v8_8HUREQ_0 vbn vbn vbn vbn vbn vss vbn vss vss vbn vbn vbn
+ vbn vbn vss vbn vbn vss vbn vss vbn vbn vbn vbn vbn vbn vss vbn vbn vbn vbn vbn
+ vbn vbn vbn vbn vss vss vbn vbn vbn vbn vbn vss vss vbn vbn vbn vbn vss vbn vss
+ vss vbn vbn vbn vss vbn vbn vbn vss vss vbn sky130_fd_pr__nfet_01v8_8HUREQ
Xsky130_fd_pr__nfet_01v8_8HUREQ_1 voe1 vbn vbn vbn vbn vss vbn vss vss vbn voe1 voe1
+ vbn vbn vss vbn voe1 vss voe1 vss voe1 vbn vbn vbn voe1 vbn vss vbn vbn vbn vbn
+ voe1 voe1 vbn voe1 vbn vss vss vbn vbn vbn voe1 voe1 vss vss voe1 vbn vbn vbn vss
+ vbn vss vss vbn voe1 voe1 vss voe1 vbn vbn vss vss vbn sky130_fd_pr__nfet_01v8_8HUREQ
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_0 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_1 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_2 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_YC9MKB_1 w_4660_n6791# w_4660_n6791# iref vdd iref iref w_4660_n6791#
+ iref vdd iref iref vdd vdd iref vdd iref w_4660_n6791# iref iref w_4660_n6791# iref
+ iref vdd w_4660_n6791# iref vdd w_4660_n6791# vdd w_4660_n6791# iref iref vdd sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__pfet_01v8_YC9MKB_0 iref iref iref vdd iref iref iref iref vdd iref
+ iref vdd vdd iref vdd iref iref iref iref iref iref iref vdd iref iref vdd iref
+ vdd iref iref iref vdd sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_3 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_YC9MKB_2 w_4660_n6791# w_4660_n6791# iref vdd iref iref w_4660_n6791#
+ iref vdd iref iref vdd vdd iref vdd iref w_4660_n6791# iref iref w_4660_n6791# iref
+ iref vdd w_4660_n6791# iref vdd w_4660_n6791# vdd w_4660_n6791# iref iref vdd sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_4 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_5 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__nfet_01v8_GQFJAV_0 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_1 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_2 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_3 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_4 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_5 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__pfet_01v8_YCMRKB_0 vin_p w_4660_n6791# vin_p voe1 voe1 vin_p vin_p
+ vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791# vin_p vin_p vin_p vin_p
+ vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 w_4660_n6791#
+ vin_p w_4660_n6791# vin_p vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p voe1 vin_p
+ voe1 vin_p vin_p voe1 w_4660_n6791# voe1 vin_p vin_p w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 vin_p vin_p w_4660_n6791# voe1 voe1
+ w_4660_n6791# voe1 w_4660_n6791# w_4660_n6791# vin_p w_4660_n6791# vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 voe1 w_4660_n6791# vin_p vin_p voe1 voe1 voe1
+ w_4660_n6791# voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791#
+ vin_p voe1 vin_p vin_p w_4660_n6791# voe1 vin_p voe1 voe1 vin_p vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p voe1 voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p
+ vin_p vin_p w_4660_n6791# w_4660_n6791# w_4660_n6791# vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p w_4660_n6791# voe1 vin_p voe1 w_4660_n6791# vin_p vin_p
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 vin_p voe1 voe1 vin_p
+ vin_p w_4660_n6791# vin_p vin_p vin_p voe1 voe1 voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p w_4660_n6791# voe1 w_4660_n6791# vin_p voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p vin_p w_4660_n6791# vin_p vin_p vin_p vin_p vin_p w_4660_n6791# w_4660_n6791#
+ vin_p vin_p voe1 voe1 voe1 vin_p sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__pfet_01v8_YCMRKB_1 vin_n w_4660_n6791# vin_n vbn vbn vin_n vin_n vin_n
+ vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vin_n vin_n vin_n vin_n
+ w_4660_n6791# vbn vin_n w_4660_n6791# w_4660_n6791# vbn vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vin_n
+ vbn vin_n vin_n vbn w_4660_n6791# vbn vin_n vin_n w_4660_n6791# w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# vbn vin_n vbn vin_n vin_n w_4660_n6791# vbn vbn w_4660_n6791# vbn
+ w_4660_n6791# w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vbn w_4660_n6791# vin_n vin_n vbn vbn vbn w_4660_n6791# vbn
+ vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vbn vin_n
+ vin_n w_4660_n6791# vbn vin_n vbn vbn vin_n vin_n vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vbn vin_n w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n vbn vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n
+ w_4660_n6791# vbn vin_n vbn w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vin_n vin_n vin_n vbn vin_n vbn vbn vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vbn vbn w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# vbn w_4660_n6791#
+ vin_n vbn w_4660_n6791# vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vbn vbn vin_n sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__pfet_01v8_YCMRKB_2 vin_n w_4660_n6791# vin_n vbn vbn vin_n vin_n vin_n
+ vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vin_n vin_n vin_n vin_n
+ w_4660_n6791# vbn vin_n w_4660_n6791# w_4660_n6791# vbn vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vin_n
+ vbn vin_n vin_n vbn w_4660_n6791# vbn vin_n vin_n w_4660_n6791# w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# vbn vin_n vbn vin_n vin_n w_4660_n6791# vbn vbn w_4660_n6791# vbn
+ w_4660_n6791# w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vbn w_4660_n6791# vin_n vin_n vbn vbn vbn w_4660_n6791# vbn
+ vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vbn vin_n
+ vin_n w_4660_n6791# vbn vin_n vbn vbn vin_n vin_n vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vbn vin_n w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n vbn vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n
+ w_4660_n6791# vbn vin_n vbn w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vin_n vin_n vin_n vbn vin_n vbn vbn vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vbn vbn w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# vbn w_4660_n6791#
+ vin_n vbn w_4660_n6791# vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vbn vbn vin_n sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__nfet_01v8_8JUMX6_0 vss vout voe1 vout vss voe1 voe1 vout vout voe1
+ vss voe1 voe1 vss vout voe1 vss vss voe1 voe1 vout voe1 vout vss voe1 voe1 vss voe1
+ vss voe1 vout voe1 voe1 vss voe1 voe1 vout voe1 vout voe1 vout voe1 vss voe1 voe1
+ voe1 voe1 voe1 vout voe1 vss vss voe1 voe1 voe1 vout vout vout vout voe1 voe1 voe1
+ vss voe1 voe1 voe1 voe1 vss vout vout voe1 voe1 vout vss vout vout vout vss voe1
+ vss vout vss voe1 vss vout vss voe1 vout vss vout vout voe1 voe1 vss vss vss voe1
+ vout voe1 voe1 vout vss voe1 vss vss voe1 vout vss vss voe1 vout vout voe1 voe1
+ vss voe1 voe1 vss vout vout vss voe1 vout voe1 vss vout voe1 vss voe1 voe1 voe1
+ vss vout voe1 vout vss vout vout vout voe1 voe1 vss voe1 vss voe1 voe1 voe1 voe1
+ vss vout voe1 voe1 voe1 vout voe1 voe1 voe1 voe1 voe1 vss vss vss voe1 voe1 voe1
+ voe1 voe1 voe1 vss voe1 vout voe1 vss voe1 voe1 voe1 voe1 voe1 vout voe1 voe1 voe1
+ vss voe1 vout voe1 voe1 vout vss vout voe1 vout vss vss vss voe1 voe1 voe1 vout
+ vout voe1 voe1 vout vss voe1 vss vout voe1 voe1 vss vss vout vss vout voe1 vss vout
+ vss vss voe1 voe1 voe1 vss vout vss voe1 voe1 vss vss voe1 voe1 voe1 vout voe1 vout
+ voe1 vout voe1 vss vss voe1 voe1 voe1 voe1 voe1 vout vout voe1 voe1 vss vss vout
+ vss vss voe1 voe1 vss voe1 voe1 vss vout voe1 vout vout vss voe1 vss vss voe1 voe1
+ voe1 vout vout voe1 vss vout voe1 voe1 voe1 vout vout voe1 voe1 vss voe1 vout voe1
+ voe1 vout vout voe1 voe1 voe1 vout vss vout voe1 vss voe1 voe1 voe1 voe1 voe1 sky130_fd_pr__nfet_01v8_8JUMX6
Xsky130_fd_pr__pfet_01v8_YCMRKB_3 vin_p w_4660_n6791# vin_p voe1 voe1 vin_p vin_p
+ vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791# vin_p vin_p vin_p vin_p
+ vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 w_4660_n6791#
+ vin_p w_4660_n6791# vin_p vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p voe1 vin_p
+ voe1 vin_p vin_p voe1 w_4660_n6791# voe1 vin_p vin_p w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 vin_p vin_p w_4660_n6791# voe1 voe1
+ w_4660_n6791# voe1 w_4660_n6791# w_4660_n6791# vin_p w_4660_n6791# vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 voe1 w_4660_n6791# vin_p vin_p voe1 voe1 voe1
+ w_4660_n6791# voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791#
+ vin_p voe1 vin_p vin_p w_4660_n6791# voe1 vin_p voe1 voe1 vin_p vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p voe1 voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p
+ vin_p vin_p w_4660_n6791# w_4660_n6791# w_4660_n6791# vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p w_4660_n6791# voe1 vin_p voe1 w_4660_n6791# vin_p vin_p
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 vin_p voe1 voe1 vin_p
+ vin_p w_4660_n6791# vin_p vin_p vin_p voe1 voe1 voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p w_4660_n6791# voe1 w_4660_n6791# vin_p voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p vin_p w_4660_n6791# vin_p vin_p vin_p vin_p vin_p w_4660_n6791# w_4660_n6791#
+ vin_p vin_p voe1 voe1 voe1 vin_p sky130_fd_pr__pfet_01v8_YCMRKB
.ends

.subckt opamp_wrapper AOUT OUT_IB AMP_IB ARRAY_OUT VSS VDD
Xopamp_v1_0 opamp_v1_0/iref AOUT ARRAY_OUT AOUT VDD VSS VSS opamp_v1
X0 ARRAY_OUT OUT_IB VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=31.9 pd=27 as=11.5 ps=22.3 w=10 l=0.15
X1 opamp_v1_0/iref AMP_IB VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=34.4 pd=27.7 as=11.5 ps=22.3 w=10 l=0.15
.ends

.subckt bias VDD NB1 NB2 OUT_IB AMP_IB GND SF_IB
X0 NB1 NB1 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.35 ps=2.7 w=1 l=1.2
X1 NB2 NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.35 ps=2.7 w=1 l=1.2
X2 AMP_IB AMP_IB GND GND sky130_fd_pr__nfet_01v8_lvt ad=5.6 pd=17.4 as=5.2 ps=17.3 w=8 l=2
X3 OUT_IB OUT_IB GND GND sky130_fd_pr__nfet_01v8_lvt ad=5.6 pd=17.4 as=5.2 ps=17.3 w=8 l=2
X4 SF_IB SF_IB VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.55 pd=3.1 as=0.45 ps=2.9 w=1 l=1
.ends

.subckt sky130_fd_pr__res_generic_m3_3NNQKJ m3_n50_n107# m3_n50_50#
R0 m3_n50_50# m3_n50_n107# sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xpixel_array_0 io_analog[7] io_analog[8] io_analog[4] io_analog[6] io_analog[9] io_analog[5]
+ io_in[20] io_in[21] io_in[22] pixel_array_0/PIX0_IN io_analog[10] pixel_array_0/PIX1_IN
+ pixel_array_0/PIX2_IN pixel_array_0/PIX3_IN pixel_array_0/PIX4_IN pixel_array_0/PIX5_IN
+ pixel_array_0/PIX6_IN pixel_array_0/PIX_OUT0 pixel_array_0/PIX7_IN pixel_array_0/PIX_OUT1
+ pixel_array_0/PIX8_IN pixel_array_0/PIX_OUT2 pixel_array_0/ARRAY_OUT io_in[23] io_in[24]
+ io_in[15] vccd1 vssd1 pixel_array
Xarray_SR_0 io_in[7] io_in[8] io_in[9] io_in[6] array_SR_0/COL_DOUT io_analog[9] array_SR_0/ARRAY_OUT
+ io_analog[5] io_analog[4] io_analog[7] io_analog[8] io_analog[6] io_in[19] io_in[16]
+ io_in[18] io_analog[10] io_in[17] vccd1 vssd1 array_SR
Xopamp_wrapper_0 io_analog[0] io_analog[3] io_analog[2] array_SR_0/ARRAY_OUT vssd1
+ vccd1 opamp_wrapper
Xopamp_wrapper_1 io_analog[1] io_analog[3] io_analog[2] pixel_array_0/ARRAY_OUT vssd1
+ vccd1 opamp_wrapper
Xbias_0 vccd1 io_analog[5] io_analog[4] io_analog[3] io_analog[2] vssd1 io_analog[6]
+ bias
Xsky130_fd_pr__res_generic_m3_3NNQKJ_0 vssd1 io_oeb[9] sky130_fd_pr__res_generic_m3_3NNQKJ
Xsky130_fd_pr__res_generic_m3_3NNQKJ_1 io_oeb[15] vssd1 sky130_fd_pr__res_generic_m3_3NNQKJ
R0 io_oeb[21] vssd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R1 vssd1 io_oeb[6] sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R2 vssd1 io_oeb[8] sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R3 io_oeb[19] vssd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R4 io_oeb[17] vssd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R5 io_oeb[24] vssd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R6 vssd1 io_oeb[7] sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R7 io_oeb[23] vssd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R8 io_oeb[16] vssd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R9 io_oeb[20] vssd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R10 io_oeb[22] vssd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R11 io_oeb[18] vssd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
.ends

