* NGSPICE file created from pixel_array100x100.ext - technology: sky130A

.subckt pixel gring VDD GND VREF ROW_SEL NB1 VBIAS NB2 AMP_IN SF_IB PIX_OUT CSA_VREF
X0 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5 pd=7.5 as=25.284374 ps=56.25 w=2 l=2
X1 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.2925 pd=2.2 as=1.57 ps=12.3 w=0.65 l=0.65
X2 a_4120_n520# VBIAS a_4120_n750# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.995 ps=8.8 w=1 l=0.8
X3 a_5720_n730# a_4600_n810# GND VDD sky130_fd_pr__pfet_01v8_lvt ad=0.25 pd=1.5 as=0.35 ps=2.7 w=1 l=1
X4 VDD SF_IB a_5720_n730# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.25 ps=1.5 w=1 l=1
X5 a_5460_10# a_4350_10# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X6 a_3860_n520# VBIAS a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.76 ps=8.8 w=1 l=0.8
X7 VDD a_4120_n520# a_4600_n810# GND sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=1
X8 a_4350_10# a_3860_n520# a_3860_n520# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X9 a_4120_n750# AMP_IN a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=1.995 pd=8.8 as=1.4 ps=7.4 w=7 l=0.15
X10 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.119375 pd=7.15 as=0 ps=0 w=2 l=3.35
X11 a_4120_n520# a_3860_n520# a_5460_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X12 GND NB1 a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0.42 pd=3.1 as=0.42 ps=3.1 w=1.2 l=1
X13 a_5750_n920# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=0.6 pd=2.95 as=5.4 ps=9.4 w=2 l=1
X14 a_4050_n2590# VREF a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=1.4 pd=7.4 as=1.76 ps=8.8 w=7 l=0.15
X15 a_4600_n810# NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1.15
X16 AMP_IN a_4600_n810# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VDD a_4350_10# a_4350_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X18 VDD a_5720_n730# a_5750_n920# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.6 ps=2.95 w=1 l=0.15
X19 AMP_IN CSA_VREF a_4600_n810# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.294 pd=2.24 as=0.273 ps=2.14 w=0.42 l=8
X20 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=10.715 pd=15.9 as=0 ps=0 w=2.6 l=0.35
.ends

.subckt pixel_array100x100 VBIAS VREF NB2 VDD NB1 ROW_SEL[0] GRING GND ROW_SEL[1]
+ ROW_SEL[2] ROW_SEL[3] ROW_SEL[4] ROW_SEL[5] ROW_SEL[6] ROW_SEL[7] ROW_SEL[8] ROW_SEL[9]
+ ROW_SEL[10] ROW_SEL[11] ROW_SEL[12] ROW_SEL[13] ROW_SEL[14] ROW_SEL[15] ROW_SEL[16]
+ ROW_SEL[17] ROW_SEL[18] ROW_SEL[19] ROW_SEL[20] ROW_SEL[21] ROW_SEL[22] ROW_SEL[23]
+ ROW_SEL[24] ROW_SEL[25] ROW_SEL[26] ROW_SEL[27] ROW_SEL[28] ROW_SEL[29] ROW_SEL[30]
+ ROW_SEL[31] ROW_SEL[32] ROW_SEL[33] ROW_SEL[34] ROW_SEL[35] ROW_SEL[36] ROW_SEL[37]
+ ROW_SEL[38] ROW_SEL[39] ROW_SEL[40] ROW_SEL[41] ROW_SEL[42] ROW_SEL[43] ROW_SEL[44]
+ ROW_SEL[45] ROW_SEL[46] ROW_SEL[47] ROW_SEL[48] ROW_SEL[49] ROW_SEL[50] ROW_SEL[51]
+ ROW_SEL[52] ROW_SEL[53] ROW_SEL[54] ROW_SEL[55] ROW_SEL[56] ROW_SEL[57] ROW_SEL[58]
+ ROW_SEL[59] ROW_SEL[60] ROW_SEL[61] ROW_SEL[62] ROW_SEL[63] ROW_SEL[64] ROW_SEL[65]
+ ROW_SEL[66] ROW_SEL[67] ROW_SEL[68] ROW_SEL[69] ROW_SEL[70] ROW_SEL[71] ROW_SEL[72]
+ ROW_SEL[73] ROW_SEL[74] ROW_SEL[75] ROW_SEL[76] ROW_SEL[77] ROW_SEL[78] ROW_SEL[79]
+ ROW_SEL[80] ROW_SEL[81] ROW_SEL[82] ROW_SEL[83] ROW_SEL[84] ROW_SEL[85] ROW_SEL[86]
+ ROW_SEL[87] ROW_SEL[88] ROW_SEL[89] ROW_SEL[90] ROW_SEL[91] ROW_SEL[92] ROW_SEL[93]
+ ROW_SEL[94] ROW_SEL[95] ROW_SEL[96] ROW_SEL[97] ROW_SEL[98] PIX_OUT0 COL_SEL[0]
+ CSA_VREF ROW_SEL[99] PIX_OUT1 COL_SEL[1] PIX_OUT2 COL_SEL[2] PIX_OUT3 COL_SEL[3]
+ PIX_OUT4 COL_SEL[4] PIX_OUT5 COL_SEL[5] PIX_OUT6 COL_SEL[6] PIX_OUT7 COL_SEL[7]
+ PIX_OUT8 COL_SEL[8] PIX_OUT9 COL_SEL[9] PIX_OUT10 COL_SEL[10] PIX_OUT11 COL_SEL[11]
+ PIX_OUT12 COL_SEL[12] PIX_OUT13 COL_SEL[13] PIX_OUT14 COL_SEL[14] PIX_OUT15 COL_SEL[15]
+ PIX_OUT16 COL_SEL[16] PIX_OUT17 COL_SEL[17] PIX_OUT18 COL_SEL[18] PIX_OUT19 COL_SEL[19]
+ PIX_OUT20 COL_SEL[20] PIX_OUT21 COL_SEL[21] PIX_OUT22 COL_SEL[22] PIX_OUT23 COL_SEL[23]
+ PIX_OUT24 COL_SEL[24] PIX_OUT25 COL_SEL[25] PIX_OUT26 COL_SEL[26] PIX_OUT27 COL_SEL[27]
+ PIX_OUT28 COL_SEL[28] PIX_OUT29 COL_SEL[29] PIX_OUT30 COL_SEL[30] PIX_OUT31 COL_SEL[31]
+ PIX_OUT32 COL_SEL[32] PIX_OUT33 COL_SEL[33] PIX_OUT34 COL_SEL[34] PIX_OUT35 COL_SEL[35]
+ PIX_OUT36 COL_SEL[36] PIX_OUT37 COL_SEL[37] PIX_OUT38 COL_SEL[38] PIX_OUT39 COL_SEL[39]
+ PIX_OUT40 COL_SEL[40] PIX_OUT41 COL_SEL[41] PIX_OUT42 COL_SEL[42] PIX_OUT43 COL_SEL[43]
+ PIX_OUT44 COL_SEL[44] PIX_OUT45 COL_SEL[45] PIX_OUT46 COL_SEL[46] PIX_OUT47 COL_SEL[47]
+ PIX_OUT48 COL_SEL[48] PIX_OUT49 COL_SEL[49] PIX_OUT50 COL_SEL[50] PIX_OUT51 COL_SEL[51]
+ PIX_OUT52 COL_SEL[52] PIX_OUT53 COL_SEL[53] PIX_OUT54 COL_SEL[54] PIX_OUT55 COL_SEL[55]
+ PIX_OUT56 COL_SEL[56] PIX_OUT57 COL_SEL[57] PIX_OUT58 COL_SEL[58] PIX_OUT59 COL_SEL[59]
+ PIX_OUT60 COL_SEL[60] PIX_OUT61 COL_SEL[61] PIX_OUT62 COL_SEL[62] PIX_OUT63 COL_SEL[63]
+ PIX_OUT64 COL_SEL[64] PIX_OUT65 COL_SEL[65] PIX_OUT66 COL_SEL[66] PIX_OUT67 COL_SEL[67]
+ PIX_OUT68 COL_SEL[68] PIX_OUT69 COL_SEL[69] PIX_OUT70 COL_SEL[70] PIX_OUT71 COL_SEL[71]
+ PIX_OUT72 COL_SEL[72] PIX_OUT73 COL_SEL[73] PIX_OUT74 COL_SEL[74] PIX_OUT75 COL_SEL[75]
+ PIX_OUT76 COL_SEL[76] PIX_OUT77 COL_SEL[77] PIX_OUT78 COL_SEL[78] PIX_OUT79 COL_SEL[79]
+ PIX_OUT80 COL_SEL[80] PIX_OUT81 COL_SEL[81] PIX_OUT82 COL_SEL[82] PIX_OUT83 COL_SEL[83]
+ PIX_OUT84 COL_SEL[84] PIX_OUT85 COL_SEL[85] PIX_OUT86 COL_SEL[86] PIX_OUT87 COL_SEL[87]
+ PIX_OUT88 COL_SEL[88] PIX_OUT89 COL_SEL[89] PIX_OUT90 COL_SEL[90] PIX_OUT91 COL_SEL[91]
+ PIX_OUT92 COL_SEL[92] PIX_OUT93 COL_SEL[93] PIX_OUT94 COL_SEL[94] PIX_OUT95 COL_SEL[95]
+ PIX_OUT96 COL_SEL[96] PIX_OUT97 COL_SEL[97] PIX_OUT98 COL_SEL[98] PIX_OUT99 ARRAY_OUT
+ COL_SEL[99] SF_IB
Xpixel_9273 pixel_9273/gring pixel_9273/VDD pixel_9273/GND pixel_9273/VREF pixel_9273/ROW_SEL
+ pixel_9273/NB1 pixel_9273/VBIAS pixel_9273/NB2 pixel_9273/AMP_IN pixel_9273/SF_IB
+ pixel_9273/PIX_OUT pixel_9273/CSA_VREF pixel
Xpixel_9262 pixel_9262/gring pixel_9262/VDD pixel_9262/GND pixel_9262/VREF pixel_9262/ROW_SEL
+ pixel_9262/NB1 pixel_9262/VBIAS pixel_9262/NB2 pixel_9262/AMP_IN pixel_9262/SF_IB
+ pixel_9262/PIX_OUT pixel_9262/CSA_VREF pixel
Xpixel_9251 pixel_9251/gring pixel_9251/VDD pixel_9251/GND pixel_9251/VREF pixel_9251/ROW_SEL
+ pixel_9251/NB1 pixel_9251/VBIAS pixel_9251/NB2 pixel_9251/AMP_IN pixel_9251/SF_IB
+ pixel_9251/PIX_OUT pixel_9251/CSA_VREF pixel
Xpixel_8572 pixel_8572/gring pixel_8572/VDD pixel_8572/GND pixel_8572/VREF pixel_8572/ROW_SEL
+ pixel_8572/NB1 pixel_8572/VBIAS pixel_8572/NB2 pixel_8572/AMP_IN pixel_8572/SF_IB
+ pixel_8572/PIX_OUT pixel_8572/CSA_VREF pixel
Xpixel_8561 pixel_8561/gring pixel_8561/VDD pixel_8561/GND pixel_8561/VREF pixel_8561/ROW_SEL
+ pixel_8561/NB1 pixel_8561/VBIAS pixel_8561/NB2 pixel_8561/AMP_IN pixel_8561/SF_IB
+ pixel_8561/PIX_OUT pixel_8561/CSA_VREF pixel
Xpixel_8550 pixel_8550/gring pixel_8550/VDD pixel_8550/GND pixel_8550/VREF pixel_8550/ROW_SEL
+ pixel_8550/NB1 pixel_8550/VBIAS pixel_8550/NB2 pixel_8550/AMP_IN pixel_8550/SF_IB
+ pixel_8550/PIX_OUT pixel_8550/CSA_VREF pixel
Xpixel_9295 pixel_9295/gring pixel_9295/VDD pixel_9295/GND pixel_9295/VREF pixel_9295/ROW_SEL
+ pixel_9295/NB1 pixel_9295/VBIAS pixel_9295/NB2 pixel_9295/AMP_IN pixel_9295/SF_IB
+ pixel_9295/PIX_OUT pixel_9295/CSA_VREF pixel
Xpixel_9284 pixel_9284/gring pixel_9284/VDD pixel_9284/GND pixel_9284/VREF pixel_9284/ROW_SEL
+ pixel_9284/NB1 pixel_9284/VBIAS pixel_9284/NB2 pixel_9284/AMP_IN pixel_9284/SF_IB
+ pixel_9284/PIX_OUT pixel_9284/CSA_VREF pixel
Xpixel_8594 pixel_8594/gring pixel_8594/VDD pixel_8594/GND pixel_8594/VREF pixel_8594/ROW_SEL
+ pixel_8594/NB1 pixel_8594/VBIAS pixel_8594/NB2 pixel_8594/AMP_IN pixel_8594/SF_IB
+ pixel_8594/PIX_OUT pixel_8594/CSA_VREF pixel
Xpixel_8583 pixel_8583/gring pixel_8583/VDD pixel_8583/GND pixel_8583/VREF pixel_8583/ROW_SEL
+ pixel_8583/NB1 pixel_8583/VBIAS pixel_8583/NB2 pixel_8583/AMP_IN pixel_8583/SF_IB
+ pixel_8583/PIX_OUT pixel_8583/CSA_VREF pixel
Xpixel_7860 pixel_7860/gring pixel_7860/VDD pixel_7860/GND pixel_7860/VREF pixel_7860/ROW_SEL
+ pixel_7860/NB1 pixel_7860/VBIAS pixel_7860/NB2 pixel_7860/AMP_IN pixel_7860/SF_IB
+ pixel_7860/PIX_OUT pixel_7860/CSA_VREF pixel
Xpixel_7871 pixel_7871/gring pixel_7871/VDD pixel_7871/GND pixel_7871/VREF pixel_7871/ROW_SEL
+ pixel_7871/NB1 pixel_7871/VBIAS pixel_7871/NB2 pixel_7871/AMP_IN pixel_7871/SF_IB
+ pixel_7871/PIX_OUT pixel_7871/CSA_VREF pixel
Xpixel_7882 pixel_7882/gring pixel_7882/VDD pixel_7882/GND pixel_7882/VREF pixel_7882/ROW_SEL
+ pixel_7882/NB1 pixel_7882/VBIAS pixel_7882/NB2 pixel_7882/AMP_IN pixel_7882/SF_IB
+ pixel_7882/PIX_OUT pixel_7882/CSA_VREF pixel
Xpixel_7893 pixel_7893/gring pixel_7893/VDD pixel_7893/GND pixel_7893/VREF pixel_7893/ROW_SEL
+ pixel_7893/NB1 pixel_7893/VBIAS pixel_7893/NB2 pixel_7893/AMP_IN pixel_7893/SF_IB
+ pixel_7893/PIX_OUT pixel_7893/CSA_VREF pixel
Xpixel_5209 pixel_5209/gring pixel_5209/VDD pixel_5209/GND pixel_5209/VREF pixel_5209/ROW_SEL
+ pixel_5209/NB1 pixel_5209/VBIAS pixel_5209/NB2 pixel_5209/AMP_IN pixel_5209/SF_IB
+ pixel_5209/PIX_OUT pixel_5209/CSA_VREF pixel
Xpixel_514 pixel_514/gring pixel_514/VDD pixel_514/GND pixel_514/VREF pixel_514/ROW_SEL
+ pixel_514/NB1 pixel_514/VBIAS pixel_514/NB2 pixel_514/AMP_IN pixel_514/SF_IB pixel_514/PIX_OUT
+ pixel_514/CSA_VREF pixel
Xpixel_503 pixel_503/gring pixel_503/VDD pixel_503/GND pixel_503/VREF pixel_503/ROW_SEL
+ pixel_503/NB1 pixel_503/VBIAS pixel_503/NB2 pixel_503/AMP_IN pixel_503/SF_IB pixel_503/PIX_OUT
+ pixel_503/CSA_VREF pixel
Xpixel_4508 pixel_4508/gring pixel_4508/VDD pixel_4508/GND pixel_4508/VREF pixel_4508/ROW_SEL
+ pixel_4508/NB1 pixel_4508/VBIAS pixel_4508/NB2 pixel_4508/AMP_IN pixel_4508/SF_IB
+ pixel_4508/PIX_OUT pixel_4508/CSA_VREF pixel
Xpixel_4519 pixel_4519/gring pixel_4519/VDD pixel_4519/GND pixel_4519/VREF pixel_4519/ROW_SEL
+ pixel_4519/NB1 pixel_4519/VBIAS pixel_4519/NB2 pixel_4519/AMP_IN pixel_4519/SF_IB
+ pixel_4519/PIX_OUT pixel_4519/CSA_VREF pixel
Xpixel_547 pixel_547/gring pixel_547/VDD pixel_547/GND pixel_547/VREF pixel_547/ROW_SEL
+ pixel_547/NB1 pixel_547/VBIAS pixel_547/NB2 pixel_547/AMP_IN pixel_547/SF_IB pixel_547/PIX_OUT
+ pixel_547/CSA_VREF pixel
Xpixel_536 pixel_536/gring pixel_536/VDD pixel_536/GND pixel_536/VREF pixel_536/ROW_SEL
+ pixel_536/NB1 pixel_536/VBIAS pixel_536/NB2 pixel_536/AMP_IN pixel_536/SF_IB pixel_536/PIX_OUT
+ pixel_536/CSA_VREF pixel
Xpixel_525 pixel_525/gring pixel_525/VDD pixel_525/GND pixel_525/VREF pixel_525/ROW_SEL
+ pixel_525/NB1 pixel_525/VBIAS pixel_525/NB2 pixel_525/AMP_IN pixel_525/SF_IB pixel_525/PIX_OUT
+ pixel_525/CSA_VREF pixel
Xpixel_3807 pixel_3807/gring pixel_3807/VDD pixel_3807/GND pixel_3807/VREF pixel_3807/ROW_SEL
+ pixel_3807/NB1 pixel_3807/VBIAS pixel_3807/NB2 pixel_3807/AMP_IN pixel_3807/SF_IB
+ pixel_3807/PIX_OUT pixel_3807/CSA_VREF pixel
Xpixel_569 pixel_569/gring pixel_569/VDD pixel_569/GND pixel_569/VREF pixel_569/ROW_SEL
+ pixel_569/NB1 pixel_569/VBIAS pixel_569/NB2 pixel_569/AMP_IN pixel_569/SF_IB pixel_569/PIX_OUT
+ pixel_569/CSA_VREF pixel
Xpixel_558 pixel_558/gring pixel_558/VDD pixel_558/GND pixel_558/VREF pixel_558/ROW_SEL
+ pixel_558/NB1 pixel_558/VBIAS pixel_558/NB2 pixel_558/AMP_IN pixel_558/SF_IB pixel_558/PIX_OUT
+ pixel_558/CSA_VREF pixel
Xpixel_3818 pixel_3818/gring pixel_3818/VDD pixel_3818/GND pixel_3818/VREF pixel_3818/ROW_SEL
+ pixel_3818/NB1 pixel_3818/VBIAS pixel_3818/NB2 pixel_3818/AMP_IN pixel_3818/SF_IB
+ pixel_3818/PIX_OUT pixel_3818/CSA_VREF pixel
Xpixel_3829 pixel_3829/gring pixel_3829/VDD pixel_3829/GND pixel_3829/VREF pixel_3829/ROW_SEL
+ pixel_3829/NB1 pixel_3829/VBIAS pixel_3829/NB2 pixel_3829/AMP_IN pixel_3829/SF_IB
+ pixel_3829/PIX_OUT pixel_3829/CSA_VREF pixel
Xpixel_7101 pixel_7101/gring pixel_7101/VDD pixel_7101/GND pixel_7101/VREF pixel_7101/ROW_SEL
+ pixel_7101/NB1 pixel_7101/VBIAS pixel_7101/NB2 pixel_7101/AMP_IN pixel_7101/SF_IB
+ pixel_7101/PIX_OUT pixel_7101/CSA_VREF pixel
Xpixel_7112 pixel_7112/gring pixel_7112/VDD pixel_7112/GND pixel_7112/VREF pixel_7112/ROW_SEL
+ pixel_7112/NB1 pixel_7112/VBIAS pixel_7112/NB2 pixel_7112/AMP_IN pixel_7112/SF_IB
+ pixel_7112/PIX_OUT pixel_7112/CSA_VREF pixel
Xpixel_7123 pixel_7123/gring pixel_7123/VDD pixel_7123/GND pixel_7123/VREF pixel_7123/ROW_SEL
+ pixel_7123/NB1 pixel_7123/VBIAS pixel_7123/NB2 pixel_7123/AMP_IN pixel_7123/SF_IB
+ pixel_7123/PIX_OUT pixel_7123/CSA_VREF pixel
Xpixel_7134 pixel_7134/gring pixel_7134/VDD pixel_7134/GND pixel_7134/VREF pixel_7134/ROW_SEL
+ pixel_7134/NB1 pixel_7134/VBIAS pixel_7134/NB2 pixel_7134/AMP_IN pixel_7134/SF_IB
+ pixel_7134/PIX_OUT pixel_7134/CSA_VREF pixel
Xpixel_7145 pixel_7145/gring pixel_7145/VDD pixel_7145/GND pixel_7145/VREF pixel_7145/ROW_SEL
+ pixel_7145/NB1 pixel_7145/VBIAS pixel_7145/NB2 pixel_7145/AMP_IN pixel_7145/SF_IB
+ pixel_7145/PIX_OUT pixel_7145/CSA_VREF pixel
Xpixel_7156 pixel_7156/gring pixel_7156/VDD pixel_7156/GND pixel_7156/VREF pixel_7156/ROW_SEL
+ pixel_7156/NB1 pixel_7156/VBIAS pixel_7156/NB2 pixel_7156/AMP_IN pixel_7156/SF_IB
+ pixel_7156/PIX_OUT pixel_7156/CSA_VREF pixel
Xpixel_6400 pixel_6400/gring pixel_6400/VDD pixel_6400/GND pixel_6400/VREF pixel_6400/ROW_SEL
+ pixel_6400/NB1 pixel_6400/VBIAS pixel_6400/NB2 pixel_6400/AMP_IN pixel_6400/SF_IB
+ pixel_6400/PIX_OUT pixel_6400/CSA_VREF pixel
Xpixel_6411 pixel_6411/gring pixel_6411/VDD pixel_6411/GND pixel_6411/VREF pixel_6411/ROW_SEL
+ pixel_6411/NB1 pixel_6411/VBIAS pixel_6411/NB2 pixel_6411/AMP_IN pixel_6411/SF_IB
+ pixel_6411/PIX_OUT pixel_6411/CSA_VREF pixel
Xpixel_7167 pixel_7167/gring pixel_7167/VDD pixel_7167/GND pixel_7167/VREF pixel_7167/ROW_SEL
+ pixel_7167/NB1 pixel_7167/VBIAS pixel_7167/NB2 pixel_7167/AMP_IN pixel_7167/SF_IB
+ pixel_7167/PIX_OUT pixel_7167/CSA_VREF pixel
Xpixel_7178 pixel_7178/gring pixel_7178/VDD pixel_7178/GND pixel_7178/VREF pixel_7178/ROW_SEL
+ pixel_7178/NB1 pixel_7178/VBIAS pixel_7178/NB2 pixel_7178/AMP_IN pixel_7178/SF_IB
+ pixel_7178/PIX_OUT pixel_7178/CSA_VREF pixel
Xpixel_7189 pixel_7189/gring pixel_7189/VDD pixel_7189/GND pixel_7189/VREF pixel_7189/ROW_SEL
+ pixel_7189/NB1 pixel_7189/VBIAS pixel_7189/NB2 pixel_7189/AMP_IN pixel_7189/SF_IB
+ pixel_7189/PIX_OUT pixel_7189/CSA_VREF pixel
Xpixel_6422 pixel_6422/gring pixel_6422/VDD pixel_6422/GND pixel_6422/VREF pixel_6422/ROW_SEL
+ pixel_6422/NB1 pixel_6422/VBIAS pixel_6422/NB2 pixel_6422/AMP_IN pixel_6422/SF_IB
+ pixel_6422/PIX_OUT pixel_6422/CSA_VREF pixel
Xpixel_6433 pixel_6433/gring pixel_6433/VDD pixel_6433/GND pixel_6433/VREF pixel_6433/ROW_SEL
+ pixel_6433/NB1 pixel_6433/VBIAS pixel_6433/NB2 pixel_6433/AMP_IN pixel_6433/SF_IB
+ pixel_6433/PIX_OUT pixel_6433/CSA_VREF pixel
Xpixel_6444 pixel_6444/gring pixel_6444/VDD pixel_6444/GND pixel_6444/VREF pixel_6444/ROW_SEL
+ pixel_6444/NB1 pixel_6444/VBIAS pixel_6444/NB2 pixel_6444/AMP_IN pixel_6444/SF_IB
+ pixel_6444/PIX_OUT pixel_6444/CSA_VREF pixel
Xpixel_6455 pixel_6455/gring pixel_6455/VDD pixel_6455/GND pixel_6455/VREF pixel_6455/ROW_SEL
+ pixel_6455/NB1 pixel_6455/VBIAS pixel_6455/NB2 pixel_6455/AMP_IN pixel_6455/SF_IB
+ pixel_6455/PIX_OUT pixel_6455/CSA_VREF pixel
Xpixel_6466 pixel_6466/gring pixel_6466/VDD pixel_6466/GND pixel_6466/VREF pixel_6466/ROW_SEL
+ pixel_6466/NB1 pixel_6466/VBIAS pixel_6466/NB2 pixel_6466/AMP_IN pixel_6466/SF_IB
+ pixel_6466/PIX_OUT pixel_6466/CSA_VREF pixel
Xpixel_6477 pixel_6477/gring pixel_6477/VDD pixel_6477/GND pixel_6477/VREF pixel_6477/ROW_SEL
+ pixel_6477/NB1 pixel_6477/VBIAS pixel_6477/NB2 pixel_6477/AMP_IN pixel_6477/SF_IB
+ pixel_6477/PIX_OUT pixel_6477/CSA_VREF pixel
Xpixel_5710 pixel_5710/gring pixel_5710/VDD pixel_5710/GND pixel_5710/VREF pixel_5710/ROW_SEL
+ pixel_5710/NB1 pixel_5710/VBIAS pixel_5710/NB2 pixel_5710/AMP_IN pixel_5710/SF_IB
+ pixel_5710/PIX_OUT pixel_5710/CSA_VREF pixel
Xpixel_5721 pixel_5721/gring pixel_5721/VDD pixel_5721/GND pixel_5721/VREF pixel_5721/ROW_SEL
+ pixel_5721/NB1 pixel_5721/VBIAS pixel_5721/NB2 pixel_5721/AMP_IN pixel_5721/SF_IB
+ pixel_5721/PIX_OUT pixel_5721/CSA_VREF pixel
Xpixel_5732 pixel_5732/gring pixel_5732/VDD pixel_5732/GND pixel_5732/VREF pixel_5732/ROW_SEL
+ pixel_5732/NB1 pixel_5732/VBIAS pixel_5732/NB2 pixel_5732/AMP_IN pixel_5732/SF_IB
+ pixel_5732/PIX_OUT pixel_5732/CSA_VREF pixel
Xpixel_5743 pixel_5743/gring pixel_5743/VDD pixel_5743/GND pixel_5743/VREF pixel_5743/ROW_SEL
+ pixel_5743/NB1 pixel_5743/VBIAS pixel_5743/NB2 pixel_5743/AMP_IN pixel_5743/SF_IB
+ pixel_5743/PIX_OUT pixel_5743/CSA_VREF pixel
Xpixel_6488 pixel_6488/gring pixel_6488/VDD pixel_6488/GND pixel_6488/VREF pixel_6488/ROW_SEL
+ pixel_6488/NB1 pixel_6488/VBIAS pixel_6488/NB2 pixel_6488/AMP_IN pixel_6488/SF_IB
+ pixel_6488/PIX_OUT pixel_6488/CSA_VREF pixel
Xpixel_6499 pixel_6499/gring pixel_6499/VDD pixel_6499/GND pixel_6499/VREF pixel_6499/ROW_SEL
+ pixel_6499/NB1 pixel_6499/VBIAS pixel_6499/NB2 pixel_6499/AMP_IN pixel_6499/SF_IB
+ pixel_6499/PIX_OUT pixel_6499/CSA_VREF pixel
Xpixel_5754 pixel_5754/gring pixel_5754/VDD pixel_5754/GND pixel_5754/VREF pixel_5754/ROW_SEL
+ pixel_5754/NB1 pixel_5754/VBIAS pixel_5754/NB2 pixel_5754/AMP_IN pixel_5754/SF_IB
+ pixel_5754/PIX_OUT pixel_5754/CSA_VREF pixel
Xpixel_5765 pixel_5765/gring pixel_5765/VDD pixel_5765/GND pixel_5765/VREF pixel_5765/ROW_SEL
+ pixel_5765/NB1 pixel_5765/VBIAS pixel_5765/NB2 pixel_5765/AMP_IN pixel_5765/SF_IB
+ pixel_5765/PIX_OUT pixel_5765/CSA_VREF pixel
Xpixel_5776 pixel_5776/gring pixel_5776/VDD pixel_5776/GND pixel_5776/VREF pixel_5776/ROW_SEL
+ pixel_5776/NB1 pixel_5776/VBIAS pixel_5776/NB2 pixel_5776/AMP_IN pixel_5776/SF_IB
+ pixel_5776/PIX_OUT pixel_5776/CSA_VREF pixel
Xpixel_5787 pixel_5787/gring pixel_5787/VDD pixel_5787/GND pixel_5787/VREF pixel_5787/ROW_SEL
+ pixel_5787/NB1 pixel_5787/VBIAS pixel_5787/NB2 pixel_5787/AMP_IN pixel_5787/SF_IB
+ pixel_5787/PIX_OUT pixel_5787/CSA_VREF pixel
Xpixel_5798 pixel_5798/gring pixel_5798/VDD pixel_5798/GND pixel_5798/VREF pixel_5798/ROW_SEL
+ pixel_5798/NB1 pixel_5798/VBIAS pixel_5798/NB2 pixel_5798/AMP_IN pixel_5798/SF_IB
+ pixel_5798/PIX_OUT pixel_5798/CSA_VREF pixel
Xpixel_9081 pixel_9081/gring pixel_9081/VDD pixel_9081/GND pixel_9081/VREF pixel_9081/ROW_SEL
+ pixel_9081/NB1 pixel_9081/VBIAS pixel_9081/NB2 pixel_9081/AMP_IN pixel_9081/SF_IB
+ pixel_9081/PIX_OUT pixel_9081/CSA_VREF pixel
Xpixel_9070 pixel_9070/gring pixel_9070/VDD pixel_9070/GND pixel_9070/VREF pixel_9070/ROW_SEL
+ pixel_9070/NB1 pixel_9070/VBIAS pixel_9070/NB2 pixel_9070/AMP_IN pixel_9070/SF_IB
+ pixel_9070/PIX_OUT pixel_9070/CSA_VREF pixel
Xpixel_9092 pixel_9092/gring pixel_9092/VDD pixel_9092/GND pixel_9092/VREF pixel_9092/ROW_SEL
+ pixel_9092/NB1 pixel_9092/VBIAS pixel_9092/NB2 pixel_9092/AMP_IN pixel_9092/SF_IB
+ pixel_9092/PIX_OUT pixel_9092/CSA_VREF pixel
Xpixel_8380 pixel_8380/gring pixel_8380/VDD pixel_8380/GND pixel_8380/VREF pixel_8380/ROW_SEL
+ pixel_8380/NB1 pixel_8380/VBIAS pixel_8380/NB2 pixel_8380/AMP_IN pixel_8380/SF_IB
+ pixel_8380/PIX_OUT pixel_8380/CSA_VREF pixel
Xpixel_8391 pixel_8391/gring pixel_8391/VDD pixel_8391/GND pixel_8391/VREF pixel_8391/ROW_SEL
+ pixel_8391/NB1 pixel_8391/VBIAS pixel_8391/NB2 pixel_8391/AMP_IN pixel_8391/SF_IB
+ pixel_8391/PIX_OUT pixel_8391/CSA_VREF pixel
Xpixel_7690 pixel_7690/gring pixel_7690/VDD pixel_7690/GND pixel_7690/VREF pixel_7690/ROW_SEL
+ pixel_7690/NB1 pixel_7690/VBIAS pixel_7690/NB2 pixel_7690/AMP_IN pixel_7690/SF_IB
+ pixel_7690/PIX_OUT pixel_7690/CSA_VREF pixel
Xpixel_81 pixel_81/gring pixel_81/VDD pixel_81/GND pixel_81/VREF pixel_81/ROW_SEL
+ pixel_81/NB1 pixel_81/VBIAS pixel_81/NB2 pixel_81/AMP_IN pixel_81/SF_IB pixel_81/PIX_OUT
+ pixel_81/CSA_VREF pixel
Xpixel_70 pixel_70/gring pixel_70/VDD pixel_70/GND pixel_70/VREF pixel_70/ROW_SEL
+ pixel_70/NB1 pixel_70/VBIAS pixel_70/NB2 pixel_70/AMP_IN pixel_70/SF_IB pixel_70/PIX_OUT
+ pixel_70/CSA_VREF pixel
Xpixel_92 pixel_92/gring pixel_92/VDD pixel_92/GND pixel_92/VREF pixel_92/ROW_SEL
+ pixel_92/NB1 pixel_92/VBIAS pixel_92/NB2 pixel_92/AMP_IN pixel_92/SF_IB pixel_92/PIX_OUT
+ pixel_92/CSA_VREF pixel
Xpixel_5006 pixel_5006/gring pixel_5006/VDD pixel_5006/GND pixel_5006/VREF pixel_5006/ROW_SEL
+ pixel_5006/NB1 pixel_5006/VBIAS pixel_5006/NB2 pixel_5006/AMP_IN pixel_5006/SF_IB
+ pixel_5006/PIX_OUT pixel_5006/CSA_VREF pixel
Xpixel_5017 pixel_5017/gring pixel_5017/VDD pixel_5017/GND pixel_5017/VREF pixel_5017/ROW_SEL
+ pixel_5017/NB1 pixel_5017/VBIAS pixel_5017/NB2 pixel_5017/AMP_IN pixel_5017/SF_IB
+ pixel_5017/PIX_OUT pixel_5017/CSA_VREF pixel
Xpixel_5028 pixel_5028/gring pixel_5028/VDD pixel_5028/GND pixel_5028/VREF pixel_5028/ROW_SEL
+ pixel_5028/NB1 pixel_5028/VBIAS pixel_5028/NB2 pixel_5028/AMP_IN pixel_5028/SF_IB
+ pixel_5028/PIX_OUT pixel_5028/CSA_VREF pixel
Xpixel_322 pixel_322/gring pixel_322/VDD pixel_322/GND pixel_322/VREF pixel_322/ROW_SEL
+ pixel_322/NB1 pixel_322/VBIAS pixel_322/NB2 pixel_322/AMP_IN pixel_322/SF_IB pixel_322/PIX_OUT
+ pixel_322/CSA_VREF pixel
Xpixel_311 pixel_311/gring pixel_311/VDD pixel_311/GND pixel_311/VREF pixel_311/ROW_SEL
+ pixel_311/NB1 pixel_311/VBIAS pixel_311/NB2 pixel_311/AMP_IN pixel_311/SF_IB pixel_311/PIX_OUT
+ pixel_311/CSA_VREF pixel
Xpixel_300 pixel_300/gring pixel_300/VDD pixel_300/GND pixel_300/VREF pixel_300/ROW_SEL
+ pixel_300/NB1 pixel_300/VBIAS pixel_300/NB2 pixel_300/AMP_IN pixel_300/SF_IB pixel_300/PIX_OUT
+ pixel_300/CSA_VREF pixel
Xpixel_5039 pixel_5039/gring pixel_5039/VDD pixel_5039/GND pixel_5039/VREF pixel_5039/ROW_SEL
+ pixel_5039/NB1 pixel_5039/VBIAS pixel_5039/NB2 pixel_5039/AMP_IN pixel_5039/SF_IB
+ pixel_5039/PIX_OUT pixel_5039/CSA_VREF pixel
Xpixel_4305 pixel_4305/gring pixel_4305/VDD pixel_4305/GND pixel_4305/VREF pixel_4305/ROW_SEL
+ pixel_4305/NB1 pixel_4305/VBIAS pixel_4305/NB2 pixel_4305/AMP_IN pixel_4305/SF_IB
+ pixel_4305/PIX_OUT pixel_4305/CSA_VREF pixel
Xpixel_4316 pixel_4316/gring pixel_4316/VDD pixel_4316/GND pixel_4316/VREF pixel_4316/ROW_SEL
+ pixel_4316/NB1 pixel_4316/VBIAS pixel_4316/NB2 pixel_4316/AMP_IN pixel_4316/SF_IB
+ pixel_4316/PIX_OUT pixel_4316/CSA_VREF pixel
Xpixel_4327 pixel_4327/gring pixel_4327/VDD pixel_4327/GND pixel_4327/VREF pixel_4327/ROW_SEL
+ pixel_4327/NB1 pixel_4327/VBIAS pixel_4327/NB2 pixel_4327/AMP_IN pixel_4327/SF_IB
+ pixel_4327/PIX_OUT pixel_4327/CSA_VREF pixel
Xpixel_355 pixel_355/gring pixel_355/VDD pixel_355/GND pixel_355/VREF pixel_355/ROW_SEL
+ pixel_355/NB1 pixel_355/VBIAS pixel_355/NB2 pixel_355/AMP_IN pixel_355/SF_IB pixel_355/PIX_OUT
+ pixel_355/CSA_VREF pixel
Xpixel_344 pixel_344/gring pixel_344/VDD pixel_344/GND pixel_344/VREF pixel_344/ROW_SEL
+ pixel_344/NB1 pixel_344/VBIAS pixel_344/NB2 pixel_344/AMP_IN pixel_344/SF_IB pixel_344/PIX_OUT
+ pixel_344/CSA_VREF pixel
Xpixel_333 pixel_333/gring pixel_333/VDD pixel_333/GND pixel_333/VREF pixel_333/ROW_SEL
+ pixel_333/NB1 pixel_333/VBIAS pixel_333/NB2 pixel_333/AMP_IN pixel_333/SF_IB pixel_333/PIX_OUT
+ pixel_333/CSA_VREF pixel
Xpixel_3615 pixel_3615/gring pixel_3615/VDD pixel_3615/GND pixel_3615/VREF pixel_3615/ROW_SEL
+ pixel_3615/NB1 pixel_3615/VBIAS pixel_3615/NB2 pixel_3615/AMP_IN pixel_3615/SF_IB
+ pixel_3615/PIX_OUT pixel_3615/CSA_VREF pixel
Xpixel_3604 pixel_3604/gring pixel_3604/VDD pixel_3604/GND pixel_3604/VREF pixel_3604/ROW_SEL
+ pixel_3604/NB1 pixel_3604/VBIAS pixel_3604/NB2 pixel_3604/AMP_IN pixel_3604/SF_IB
+ pixel_3604/PIX_OUT pixel_3604/CSA_VREF pixel
Xpixel_4338 pixel_4338/gring pixel_4338/VDD pixel_4338/GND pixel_4338/VREF pixel_4338/ROW_SEL
+ pixel_4338/NB1 pixel_4338/VBIAS pixel_4338/NB2 pixel_4338/AMP_IN pixel_4338/SF_IB
+ pixel_4338/PIX_OUT pixel_4338/CSA_VREF pixel
Xpixel_4349 pixel_4349/gring pixel_4349/VDD pixel_4349/GND pixel_4349/VREF pixel_4349/ROW_SEL
+ pixel_4349/NB1 pixel_4349/VBIAS pixel_4349/NB2 pixel_4349/AMP_IN pixel_4349/SF_IB
+ pixel_4349/PIX_OUT pixel_4349/CSA_VREF pixel
Xpixel_399 pixel_399/gring pixel_399/VDD pixel_399/GND pixel_399/VREF pixel_399/ROW_SEL
+ pixel_399/NB1 pixel_399/VBIAS pixel_399/NB2 pixel_399/AMP_IN pixel_399/SF_IB pixel_399/PIX_OUT
+ pixel_399/CSA_VREF pixel
Xpixel_388 pixel_388/gring pixel_388/VDD pixel_388/GND pixel_388/VREF pixel_388/ROW_SEL
+ pixel_388/NB1 pixel_388/VBIAS pixel_388/NB2 pixel_388/AMP_IN pixel_388/SF_IB pixel_388/PIX_OUT
+ pixel_388/CSA_VREF pixel
Xpixel_377 pixel_377/gring pixel_377/VDD pixel_377/GND pixel_377/VREF pixel_377/ROW_SEL
+ pixel_377/NB1 pixel_377/VBIAS pixel_377/NB2 pixel_377/AMP_IN pixel_377/SF_IB pixel_377/PIX_OUT
+ pixel_377/CSA_VREF pixel
Xpixel_366 pixel_366/gring pixel_366/VDD pixel_366/GND pixel_366/VREF pixel_366/ROW_SEL
+ pixel_366/NB1 pixel_366/VBIAS pixel_366/NB2 pixel_366/AMP_IN pixel_366/SF_IB pixel_366/PIX_OUT
+ pixel_366/CSA_VREF pixel
Xpixel_2914 pixel_2914/gring pixel_2914/VDD pixel_2914/GND pixel_2914/VREF pixel_2914/ROW_SEL
+ pixel_2914/NB1 pixel_2914/VBIAS pixel_2914/NB2 pixel_2914/AMP_IN pixel_2914/SF_IB
+ pixel_2914/PIX_OUT pixel_2914/CSA_VREF pixel
Xpixel_2903 pixel_2903/gring pixel_2903/VDD pixel_2903/GND pixel_2903/VREF pixel_2903/ROW_SEL
+ pixel_2903/NB1 pixel_2903/VBIAS pixel_2903/NB2 pixel_2903/AMP_IN pixel_2903/SF_IB
+ pixel_2903/PIX_OUT pixel_2903/CSA_VREF pixel
Xpixel_3648 pixel_3648/gring pixel_3648/VDD pixel_3648/GND pixel_3648/VREF pixel_3648/ROW_SEL
+ pixel_3648/NB1 pixel_3648/VBIAS pixel_3648/NB2 pixel_3648/AMP_IN pixel_3648/SF_IB
+ pixel_3648/PIX_OUT pixel_3648/CSA_VREF pixel
Xpixel_3637 pixel_3637/gring pixel_3637/VDD pixel_3637/GND pixel_3637/VREF pixel_3637/ROW_SEL
+ pixel_3637/NB1 pixel_3637/VBIAS pixel_3637/NB2 pixel_3637/AMP_IN pixel_3637/SF_IB
+ pixel_3637/PIX_OUT pixel_3637/CSA_VREF pixel
Xpixel_3626 pixel_3626/gring pixel_3626/VDD pixel_3626/GND pixel_3626/VREF pixel_3626/ROW_SEL
+ pixel_3626/NB1 pixel_3626/VBIAS pixel_3626/NB2 pixel_3626/AMP_IN pixel_3626/SF_IB
+ pixel_3626/PIX_OUT pixel_3626/CSA_VREF pixel
Xpixel_2947 pixel_2947/gring pixel_2947/VDD pixel_2947/GND pixel_2947/VREF pixel_2947/ROW_SEL
+ pixel_2947/NB1 pixel_2947/VBIAS pixel_2947/NB2 pixel_2947/AMP_IN pixel_2947/SF_IB
+ pixel_2947/PIX_OUT pixel_2947/CSA_VREF pixel
Xpixel_2936 pixel_2936/gring pixel_2936/VDD pixel_2936/GND pixel_2936/VREF pixel_2936/ROW_SEL
+ pixel_2936/NB1 pixel_2936/VBIAS pixel_2936/NB2 pixel_2936/AMP_IN pixel_2936/SF_IB
+ pixel_2936/PIX_OUT pixel_2936/CSA_VREF pixel
Xpixel_2925 pixel_2925/gring pixel_2925/VDD pixel_2925/GND pixel_2925/VREF pixel_2925/ROW_SEL
+ pixel_2925/NB1 pixel_2925/VBIAS pixel_2925/NB2 pixel_2925/AMP_IN pixel_2925/SF_IB
+ pixel_2925/PIX_OUT pixel_2925/CSA_VREF pixel
Xpixel_3659 pixel_3659/gring pixel_3659/VDD pixel_3659/GND pixel_3659/VREF pixel_3659/ROW_SEL
+ pixel_3659/NB1 pixel_3659/VBIAS pixel_3659/NB2 pixel_3659/AMP_IN pixel_3659/SF_IB
+ pixel_3659/PIX_OUT pixel_3659/CSA_VREF pixel
Xpixel_2969 pixel_2969/gring pixel_2969/VDD pixel_2969/GND pixel_2969/VREF pixel_2969/ROW_SEL
+ pixel_2969/NB1 pixel_2969/VBIAS pixel_2969/NB2 pixel_2969/AMP_IN pixel_2969/SF_IB
+ pixel_2969/PIX_OUT pixel_2969/CSA_VREF pixel
Xpixel_2958 pixel_2958/gring pixel_2958/VDD pixel_2958/GND pixel_2958/VREF pixel_2958/ROW_SEL
+ pixel_2958/NB1 pixel_2958/VBIAS pixel_2958/NB2 pixel_2958/AMP_IN pixel_2958/SF_IB
+ pixel_2958/PIX_OUT pixel_2958/CSA_VREF pixel
Xpixel_6230 pixel_6230/gring pixel_6230/VDD pixel_6230/GND pixel_6230/VREF pixel_6230/ROW_SEL
+ pixel_6230/NB1 pixel_6230/VBIAS pixel_6230/NB2 pixel_6230/AMP_IN pixel_6230/SF_IB
+ pixel_6230/PIX_OUT pixel_6230/CSA_VREF pixel
Xpixel_6241 pixel_6241/gring pixel_6241/VDD pixel_6241/GND pixel_6241/VREF pixel_6241/ROW_SEL
+ pixel_6241/NB1 pixel_6241/VBIAS pixel_6241/NB2 pixel_6241/AMP_IN pixel_6241/SF_IB
+ pixel_6241/PIX_OUT pixel_6241/CSA_VREF pixel
Xpixel_6252 pixel_6252/gring pixel_6252/VDD pixel_6252/GND pixel_6252/VREF pixel_6252/ROW_SEL
+ pixel_6252/NB1 pixel_6252/VBIAS pixel_6252/NB2 pixel_6252/AMP_IN pixel_6252/SF_IB
+ pixel_6252/PIX_OUT pixel_6252/CSA_VREF pixel
Xpixel_6263 pixel_6263/gring pixel_6263/VDD pixel_6263/GND pixel_6263/VREF pixel_6263/ROW_SEL
+ pixel_6263/NB1 pixel_6263/VBIAS pixel_6263/NB2 pixel_6263/AMP_IN pixel_6263/SF_IB
+ pixel_6263/PIX_OUT pixel_6263/CSA_VREF pixel
Xpixel_6274 pixel_6274/gring pixel_6274/VDD pixel_6274/GND pixel_6274/VREF pixel_6274/ROW_SEL
+ pixel_6274/NB1 pixel_6274/VBIAS pixel_6274/NB2 pixel_6274/AMP_IN pixel_6274/SF_IB
+ pixel_6274/PIX_OUT pixel_6274/CSA_VREF pixel
Xpixel_6285 pixel_6285/gring pixel_6285/VDD pixel_6285/GND pixel_6285/VREF pixel_6285/ROW_SEL
+ pixel_6285/NB1 pixel_6285/VBIAS pixel_6285/NB2 pixel_6285/AMP_IN pixel_6285/SF_IB
+ pixel_6285/PIX_OUT pixel_6285/CSA_VREF pixel
Xpixel_6296 pixel_6296/gring pixel_6296/VDD pixel_6296/GND pixel_6296/VREF pixel_6296/ROW_SEL
+ pixel_6296/NB1 pixel_6296/VBIAS pixel_6296/NB2 pixel_6296/AMP_IN pixel_6296/SF_IB
+ pixel_6296/PIX_OUT pixel_6296/CSA_VREF pixel
Xpixel_5540 pixel_5540/gring pixel_5540/VDD pixel_5540/GND pixel_5540/VREF pixel_5540/ROW_SEL
+ pixel_5540/NB1 pixel_5540/VBIAS pixel_5540/NB2 pixel_5540/AMP_IN pixel_5540/SF_IB
+ pixel_5540/PIX_OUT pixel_5540/CSA_VREF pixel
Xpixel_5551 pixel_5551/gring pixel_5551/VDD pixel_5551/GND pixel_5551/VREF pixel_5551/ROW_SEL
+ pixel_5551/NB1 pixel_5551/VBIAS pixel_5551/NB2 pixel_5551/AMP_IN pixel_5551/SF_IB
+ pixel_5551/PIX_OUT pixel_5551/CSA_VREF pixel
Xpixel_5562 pixel_5562/gring pixel_5562/VDD pixel_5562/GND pixel_5562/VREF pixel_5562/ROW_SEL
+ pixel_5562/NB1 pixel_5562/VBIAS pixel_5562/NB2 pixel_5562/AMP_IN pixel_5562/SF_IB
+ pixel_5562/PIX_OUT pixel_5562/CSA_VREF pixel
Xpixel_5573 pixel_5573/gring pixel_5573/VDD pixel_5573/GND pixel_5573/VREF pixel_5573/ROW_SEL
+ pixel_5573/NB1 pixel_5573/VBIAS pixel_5573/NB2 pixel_5573/AMP_IN pixel_5573/SF_IB
+ pixel_5573/PIX_OUT pixel_5573/CSA_VREF pixel
Xpixel_5584 pixel_5584/gring pixel_5584/VDD pixel_5584/GND pixel_5584/VREF pixel_5584/ROW_SEL
+ pixel_5584/NB1 pixel_5584/VBIAS pixel_5584/NB2 pixel_5584/AMP_IN pixel_5584/SF_IB
+ pixel_5584/PIX_OUT pixel_5584/CSA_VREF pixel
Xpixel_5595 pixel_5595/gring pixel_5595/VDD pixel_5595/GND pixel_5595/VREF pixel_5595/ROW_SEL
+ pixel_5595/NB1 pixel_5595/VBIAS pixel_5595/NB2 pixel_5595/AMP_IN pixel_5595/SF_IB
+ pixel_5595/PIX_OUT pixel_5595/CSA_VREF pixel
Xpixel_4850 pixel_4850/gring pixel_4850/VDD pixel_4850/GND pixel_4850/VREF pixel_4850/ROW_SEL
+ pixel_4850/NB1 pixel_4850/VBIAS pixel_4850/NB2 pixel_4850/AMP_IN pixel_4850/SF_IB
+ pixel_4850/PIX_OUT pixel_4850/CSA_VREF pixel
Xpixel_4861 pixel_4861/gring pixel_4861/VDD pixel_4861/GND pixel_4861/VREF pixel_4861/ROW_SEL
+ pixel_4861/NB1 pixel_4861/VBIAS pixel_4861/NB2 pixel_4861/AMP_IN pixel_4861/SF_IB
+ pixel_4861/PIX_OUT pixel_4861/CSA_VREF pixel
Xpixel_4872 pixel_4872/gring pixel_4872/VDD pixel_4872/GND pixel_4872/VREF pixel_4872/ROW_SEL
+ pixel_4872/NB1 pixel_4872/VBIAS pixel_4872/NB2 pixel_4872/AMP_IN pixel_4872/SF_IB
+ pixel_4872/PIX_OUT pixel_4872/CSA_VREF pixel
Xpixel_4883 pixel_4883/gring pixel_4883/VDD pixel_4883/GND pixel_4883/VREF pixel_4883/ROW_SEL
+ pixel_4883/NB1 pixel_4883/VBIAS pixel_4883/NB2 pixel_4883/AMP_IN pixel_4883/SF_IB
+ pixel_4883/PIX_OUT pixel_4883/CSA_VREF pixel
Xpixel_4894 pixel_4894/gring pixel_4894/VDD pixel_4894/GND pixel_4894/VREF pixel_4894/ROW_SEL
+ pixel_4894/NB1 pixel_4894/VBIAS pixel_4894/NB2 pixel_4894/AMP_IN pixel_4894/SF_IB
+ pixel_4894/PIX_OUT pixel_4894/CSA_VREF pixel
Xpixel_1509 pixel_1509/gring pixel_1509/VDD pixel_1509/GND pixel_1509/VREF pixel_1509/ROW_SEL
+ pixel_1509/NB1 pixel_1509/VBIAS pixel_1509/NB2 pixel_1509/AMP_IN pixel_1509/SF_IB
+ pixel_1509/PIX_OUT pixel_1509/CSA_VREF pixel
Xpixel_9806 pixel_9806/gring pixel_9806/VDD pixel_9806/GND pixel_9806/VREF pixel_9806/ROW_SEL
+ pixel_9806/NB1 pixel_9806/VBIAS pixel_9806/NB2 pixel_9806/AMP_IN pixel_9806/SF_IB
+ pixel_9806/PIX_OUT pixel_9806/CSA_VREF pixel
Xpixel_9839 pixel_9839/gring pixel_9839/VDD pixel_9839/GND pixel_9839/VREF pixel_9839/ROW_SEL
+ pixel_9839/NB1 pixel_9839/VBIAS pixel_9839/NB2 pixel_9839/AMP_IN pixel_9839/SF_IB
+ pixel_9839/PIX_OUT pixel_9839/CSA_VREF pixel
Xpixel_9828 pixel_9828/gring pixel_9828/VDD pixel_9828/GND pixel_9828/VREF pixel_9828/ROW_SEL
+ pixel_9828/NB1 pixel_9828/VBIAS pixel_9828/NB2 pixel_9828/AMP_IN pixel_9828/SF_IB
+ pixel_9828/PIX_OUT pixel_9828/CSA_VREF pixel
Xpixel_9817 pixel_9817/gring pixel_9817/VDD pixel_9817/GND pixel_9817/VREF pixel_9817/ROW_SEL
+ pixel_9817/NB1 pixel_9817/VBIAS pixel_9817/NB2 pixel_9817/AMP_IN pixel_9817/SF_IB
+ pixel_9817/PIX_OUT pixel_9817/CSA_VREF pixel
Xpixel_4102 pixel_4102/gring pixel_4102/VDD pixel_4102/GND pixel_4102/VREF pixel_4102/ROW_SEL
+ pixel_4102/NB1 pixel_4102/VBIAS pixel_4102/NB2 pixel_4102/AMP_IN pixel_4102/SF_IB
+ pixel_4102/PIX_OUT pixel_4102/CSA_VREF pixel
Xpixel_130 pixel_130/gring pixel_130/VDD pixel_130/GND pixel_130/VREF pixel_130/ROW_SEL
+ pixel_130/NB1 pixel_130/VBIAS pixel_130/NB2 pixel_130/AMP_IN pixel_130/SF_IB pixel_130/PIX_OUT
+ pixel_130/CSA_VREF pixel
Xpixel_4113 pixel_4113/gring pixel_4113/VDD pixel_4113/GND pixel_4113/VREF pixel_4113/ROW_SEL
+ pixel_4113/NB1 pixel_4113/VBIAS pixel_4113/NB2 pixel_4113/AMP_IN pixel_4113/SF_IB
+ pixel_4113/PIX_OUT pixel_4113/CSA_VREF pixel
Xpixel_4124 pixel_4124/gring pixel_4124/VDD pixel_4124/GND pixel_4124/VREF pixel_4124/ROW_SEL
+ pixel_4124/NB1 pixel_4124/VBIAS pixel_4124/NB2 pixel_4124/AMP_IN pixel_4124/SF_IB
+ pixel_4124/PIX_OUT pixel_4124/CSA_VREF pixel
Xpixel_4135 pixel_4135/gring pixel_4135/VDD pixel_4135/GND pixel_4135/VREF pixel_4135/ROW_SEL
+ pixel_4135/NB1 pixel_4135/VBIAS pixel_4135/NB2 pixel_4135/AMP_IN pixel_4135/SF_IB
+ pixel_4135/PIX_OUT pixel_4135/CSA_VREF pixel
Xpixel_163 pixel_163/gring pixel_163/VDD pixel_163/GND pixel_163/VREF pixel_163/ROW_SEL
+ pixel_163/NB1 pixel_163/VBIAS pixel_163/NB2 pixel_163/AMP_IN pixel_163/SF_IB pixel_163/PIX_OUT
+ pixel_163/CSA_VREF pixel
Xpixel_152 pixel_152/gring pixel_152/VDD pixel_152/GND pixel_152/VREF pixel_152/ROW_SEL
+ pixel_152/NB1 pixel_152/VBIAS pixel_152/NB2 pixel_152/AMP_IN pixel_152/SF_IB pixel_152/PIX_OUT
+ pixel_152/CSA_VREF pixel
Xpixel_141 pixel_141/gring pixel_141/VDD pixel_141/GND pixel_141/VREF pixel_141/ROW_SEL
+ pixel_141/NB1 pixel_141/VBIAS pixel_141/NB2 pixel_141/AMP_IN pixel_141/SF_IB pixel_141/PIX_OUT
+ pixel_141/CSA_VREF pixel
Xpixel_3423 pixel_3423/gring pixel_3423/VDD pixel_3423/GND pixel_3423/VREF pixel_3423/ROW_SEL
+ pixel_3423/NB1 pixel_3423/VBIAS pixel_3423/NB2 pixel_3423/AMP_IN pixel_3423/SF_IB
+ pixel_3423/PIX_OUT pixel_3423/CSA_VREF pixel
Xpixel_3412 pixel_3412/gring pixel_3412/VDD pixel_3412/GND pixel_3412/VREF pixel_3412/ROW_SEL
+ pixel_3412/NB1 pixel_3412/VBIAS pixel_3412/NB2 pixel_3412/AMP_IN pixel_3412/SF_IB
+ pixel_3412/PIX_OUT pixel_3412/CSA_VREF pixel
Xpixel_3401 pixel_3401/gring pixel_3401/VDD pixel_3401/GND pixel_3401/VREF pixel_3401/ROW_SEL
+ pixel_3401/NB1 pixel_3401/VBIAS pixel_3401/NB2 pixel_3401/AMP_IN pixel_3401/SF_IB
+ pixel_3401/PIX_OUT pixel_3401/CSA_VREF pixel
Xpixel_4146 pixel_4146/gring pixel_4146/VDD pixel_4146/GND pixel_4146/VREF pixel_4146/ROW_SEL
+ pixel_4146/NB1 pixel_4146/VBIAS pixel_4146/NB2 pixel_4146/AMP_IN pixel_4146/SF_IB
+ pixel_4146/PIX_OUT pixel_4146/CSA_VREF pixel
Xpixel_4157 pixel_4157/gring pixel_4157/VDD pixel_4157/GND pixel_4157/VREF pixel_4157/ROW_SEL
+ pixel_4157/NB1 pixel_4157/VBIAS pixel_4157/NB2 pixel_4157/AMP_IN pixel_4157/SF_IB
+ pixel_4157/PIX_OUT pixel_4157/CSA_VREF pixel
Xpixel_4168 pixel_4168/gring pixel_4168/VDD pixel_4168/GND pixel_4168/VREF pixel_4168/ROW_SEL
+ pixel_4168/NB1 pixel_4168/VBIAS pixel_4168/NB2 pixel_4168/AMP_IN pixel_4168/SF_IB
+ pixel_4168/PIX_OUT pixel_4168/CSA_VREF pixel
Xpixel_196 pixel_196/gring pixel_196/VDD pixel_196/GND pixel_196/VREF pixel_196/ROW_SEL
+ pixel_196/NB1 pixel_196/VBIAS pixel_196/NB2 pixel_196/AMP_IN pixel_196/SF_IB pixel_196/PIX_OUT
+ pixel_196/CSA_VREF pixel
Xpixel_185 pixel_185/gring pixel_185/VDD pixel_185/GND pixel_185/VREF pixel_185/ROW_SEL
+ pixel_185/NB1 pixel_185/VBIAS pixel_185/NB2 pixel_185/AMP_IN pixel_185/SF_IB pixel_185/PIX_OUT
+ pixel_185/CSA_VREF pixel
Xpixel_174 pixel_174/gring pixel_174/VDD pixel_174/GND pixel_174/VREF pixel_174/ROW_SEL
+ pixel_174/NB1 pixel_174/VBIAS pixel_174/NB2 pixel_174/AMP_IN pixel_174/SF_IB pixel_174/PIX_OUT
+ pixel_174/CSA_VREF pixel
Xpixel_2722 pixel_2722/gring pixel_2722/VDD pixel_2722/GND pixel_2722/VREF pixel_2722/ROW_SEL
+ pixel_2722/NB1 pixel_2722/VBIAS pixel_2722/NB2 pixel_2722/AMP_IN pixel_2722/SF_IB
+ pixel_2722/PIX_OUT pixel_2722/CSA_VREF pixel
Xpixel_2711 pixel_2711/gring pixel_2711/VDD pixel_2711/GND pixel_2711/VREF pixel_2711/ROW_SEL
+ pixel_2711/NB1 pixel_2711/VBIAS pixel_2711/NB2 pixel_2711/AMP_IN pixel_2711/SF_IB
+ pixel_2711/PIX_OUT pixel_2711/CSA_VREF pixel
Xpixel_2700 pixel_2700/gring pixel_2700/VDD pixel_2700/GND pixel_2700/VREF pixel_2700/ROW_SEL
+ pixel_2700/NB1 pixel_2700/VBIAS pixel_2700/NB2 pixel_2700/AMP_IN pixel_2700/SF_IB
+ pixel_2700/PIX_OUT pixel_2700/CSA_VREF pixel
Xpixel_3467 pixel_3467/gring pixel_3467/VDD pixel_3467/GND pixel_3467/VREF pixel_3467/ROW_SEL
+ pixel_3467/NB1 pixel_3467/VBIAS pixel_3467/NB2 pixel_3467/AMP_IN pixel_3467/SF_IB
+ pixel_3467/PIX_OUT pixel_3467/CSA_VREF pixel
Xpixel_3456 pixel_3456/gring pixel_3456/VDD pixel_3456/GND pixel_3456/VREF pixel_3456/ROW_SEL
+ pixel_3456/NB1 pixel_3456/VBIAS pixel_3456/NB2 pixel_3456/AMP_IN pixel_3456/SF_IB
+ pixel_3456/PIX_OUT pixel_3456/CSA_VREF pixel
Xpixel_3445 pixel_3445/gring pixel_3445/VDD pixel_3445/GND pixel_3445/VREF pixel_3445/ROW_SEL
+ pixel_3445/NB1 pixel_3445/VBIAS pixel_3445/NB2 pixel_3445/AMP_IN pixel_3445/SF_IB
+ pixel_3445/PIX_OUT pixel_3445/CSA_VREF pixel
Xpixel_3434 pixel_3434/gring pixel_3434/VDD pixel_3434/GND pixel_3434/VREF pixel_3434/ROW_SEL
+ pixel_3434/NB1 pixel_3434/VBIAS pixel_3434/NB2 pixel_3434/AMP_IN pixel_3434/SF_IB
+ pixel_3434/PIX_OUT pixel_3434/CSA_VREF pixel
Xpixel_4179 pixel_4179/gring pixel_4179/VDD pixel_4179/GND pixel_4179/VREF pixel_4179/ROW_SEL
+ pixel_4179/NB1 pixel_4179/VBIAS pixel_4179/NB2 pixel_4179/AMP_IN pixel_4179/SF_IB
+ pixel_4179/PIX_OUT pixel_4179/CSA_VREF pixel
Xpixel_2755 pixel_2755/gring pixel_2755/VDD pixel_2755/GND pixel_2755/VREF pixel_2755/ROW_SEL
+ pixel_2755/NB1 pixel_2755/VBIAS pixel_2755/NB2 pixel_2755/AMP_IN pixel_2755/SF_IB
+ pixel_2755/PIX_OUT pixel_2755/CSA_VREF pixel
Xpixel_2744 pixel_2744/gring pixel_2744/VDD pixel_2744/GND pixel_2744/VREF pixel_2744/ROW_SEL
+ pixel_2744/NB1 pixel_2744/VBIAS pixel_2744/NB2 pixel_2744/AMP_IN pixel_2744/SF_IB
+ pixel_2744/PIX_OUT pixel_2744/CSA_VREF pixel
Xpixel_2733 pixel_2733/gring pixel_2733/VDD pixel_2733/GND pixel_2733/VREF pixel_2733/ROW_SEL
+ pixel_2733/NB1 pixel_2733/VBIAS pixel_2733/NB2 pixel_2733/AMP_IN pixel_2733/SF_IB
+ pixel_2733/PIX_OUT pixel_2733/CSA_VREF pixel
Xpixel_3489 pixel_3489/gring pixel_3489/VDD pixel_3489/GND pixel_3489/VREF pixel_3489/ROW_SEL
+ pixel_3489/NB1 pixel_3489/VBIAS pixel_3489/NB2 pixel_3489/AMP_IN pixel_3489/SF_IB
+ pixel_3489/PIX_OUT pixel_3489/CSA_VREF pixel
Xpixel_3478 pixel_3478/gring pixel_3478/VDD pixel_3478/GND pixel_3478/VREF pixel_3478/ROW_SEL
+ pixel_3478/NB1 pixel_3478/VBIAS pixel_3478/NB2 pixel_3478/AMP_IN pixel_3478/SF_IB
+ pixel_3478/PIX_OUT pixel_3478/CSA_VREF pixel
Xpixel_2788 pixel_2788/gring pixel_2788/VDD pixel_2788/GND pixel_2788/VREF pixel_2788/ROW_SEL
+ pixel_2788/NB1 pixel_2788/VBIAS pixel_2788/NB2 pixel_2788/AMP_IN pixel_2788/SF_IB
+ pixel_2788/PIX_OUT pixel_2788/CSA_VREF pixel
Xpixel_2777 pixel_2777/gring pixel_2777/VDD pixel_2777/GND pixel_2777/VREF pixel_2777/ROW_SEL
+ pixel_2777/NB1 pixel_2777/VBIAS pixel_2777/NB2 pixel_2777/AMP_IN pixel_2777/SF_IB
+ pixel_2777/PIX_OUT pixel_2777/CSA_VREF pixel
Xpixel_2766 pixel_2766/gring pixel_2766/VDD pixel_2766/GND pixel_2766/VREF pixel_2766/ROW_SEL
+ pixel_2766/NB1 pixel_2766/VBIAS pixel_2766/NB2 pixel_2766/AMP_IN pixel_2766/SF_IB
+ pixel_2766/PIX_OUT pixel_2766/CSA_VREF pixel
Xpixel_2799 pixel_2799/gring pixel_2799/VDD pixel_2799/GND pixel_2799/VREF pixel_2799/ROW_SEL
+ pixel_2799/NB1 pixel_2799/VBIAS pixel_2799/NB2 pixel_2799/AMP_IN pixel_2799/SF_IB
+ pixel_2799/PIX_OUT pixel_2799/CSA_VREF pixel
Xpixel_6060 pixel_6060/gring pixel_6060/VDD pixel_6060/GND pixel_6060/VREF pixel_6060/ROW_SEL
+ pixel_6060/NB1 pixel_6060/VBIAS pixel_6060/NB2 pixel_6060/AMP_IN pixel_6060/SF_IB
+ pixel_6060/PIX_OUT pixel_6060/CSA_VREF pixel
Xpixel_6071 pixel_6071/gring pixel_6071/VDD pixel_6071/GND pixel_6071/VREF pixel_6071/ROW_SEL
+ pixel_6071/NB1 pixel_6071/VBIAS pixel_6071/NB2 pixel_6071/AMP_IN pixel_6071/SF_IB
+ pixel_6071/PIX_OUT pixel_6071/CSA_VREF pixel
Xpixel_6082 pixel_6082/gring pixel_6082/VDD pixel_6082/GND pixel_6082/VREF pixel_6082/ROW_SEL
+ pixel_6082/NB1 pixel_6082/VBIAS pixel_6082/NB2 pixel_6082/AMP_IN pixel_6082/SF_IB
+ pixel_6082/PIX_OUT pixel_6082/CSA_VREF pixel
Xpixel_6093 pixel_6093/gring pixel_6093/VDD pixel_6093/GND pixel_6093/VREF pixel_6093/ROW_SEL
+ pixel_6093/NB1 pixel_6093/VBIAS pixel_6093/NB2 pixel_6093/AMP_IN pixel_6093/SF_IB
+ pixel_6093/PIX_OUT pixel_6093/CSA_VREF pixel
Xpixel_5370 pixel_5370/gring pixel_5370/VDD pixel_5370/GND pixel_5370/VREF pixel_5370/ROW_SEL
+ pixel_5370/NB1 pixel_5370/VBIAS pixel_5370/NB2 pixel_5370/AMP_IN pixel_5370/SF_IB
+ pixel_5370/PIX_OUT pixel_5370/CSA_VREF pixel
Xpixel_5381 pixel_5381/gring pixel_5381/VDD pixel_5381/GND pixel_5381/VREF pixel_5381/ROW_SEL
+ pixel_5381/NB1 pixel_5381/VBIAS pixel_5381/NB2 pixel_5381/AMP_IN pixel_5381/SF_IB
+ pixel_5381/PIX_OUT pixel_5381/CSA_VREF pixel
Xpixel_5392 pixel_5392/gring pixel_5392/VDD pixel_5392/GND pixel_5392/VREF pixel_5392/ROW_SEL
+ pixel_5392/NB1 pixel_5392/VBIAS pixel_5392/NB2 pixel_5392/AMP_IN pixel_5392/SF_IB
+ pixel_5392/PIX_OUT pixel_5392/CSA_VREF pixel
Xpixel_4680 pixel_4680/gring pixel_4680/VDD pixel_4680/GND pixel_4680/VREF pixel_4680/ROW_SEL
+ pixel_4680/NB1 pixel_4680/VBIAS pixel_4680/NB2 pixel_4680/AMP_IN pixel_4680/SF_IB
+ pixel_4680/PIX_OUT pixel_4680/CSA_VREF pixel
Xpixel_4691 pixel_4691/gring pixel_4691/VDD pixel_4691/GND pixel_4691/VREF pixel_4691/ROW_SEL
+ pixel_4691/NB1 pixel_4691/VBIAS pixel_4691/NB2 pixel_4691/AMP_IN pixel_4691/SF_IB
+ pixel_4691/PIX_OUT pixel_4691/CSA_VREF pixel
Xpixel_3990 pixel_3990/gring pixel_3990/VDD pixel_3990/GND pixel_3990/VREF pixel_3990/ROW_SEL
+ pixel_3990/NB1 pixel_3990/VBIAS pixel_3990/NB2 pixel_3990/AMP_IN pixel_3990/SF_IB
+ pixel_3990/PIX_OUT pixel_3990/CSA_VREF pixel
Xpixel_0 pixel_0/gring pixel_0/VDD pixel_0/GND pixel_0/VREF pixel_0/ROW_SEL pixel_0/NB1
+ pixel_0/VBIAS pixel_0/NB2 pixel_0/AMP_IN pixel_0/SF_IB pixel_0/PIX_OUT pixel_0/CSA_VREF
+ pixel
Xpixel_2018 pixel_2018/gring pixel_2018/VDD pixel_2018/GND pixel_2018/VREF pixel_2018/ROW_SEL
+ pixel_2018/NB1 pixel_2018/VBIAS pixel_2018/NB2 pixel_2018/AMP_IN pixel_2018/SF_IB
+ pixel_2018/PIX_OUT pixel_2018/CSA_VREF pixel
Xpixel_2007 pixel_2007/gring pixel_2007/VDD pixel_2007/GND pixel_2007/VREF pixel_2007/ROW_SEL
+ pixel_2007/NB1 pixel_2007/VBIAS pixel_2007/NB2 pixel_2007/AMP_IN pixel_2007/SF_IB
+ pixel_2007/PIX_OUT pixel_2007/CSA_VREF pixel
Xpixel_1306 pixel_1306/gring pixel_1306/VDD pixel_1306/GND pixel_1306/VREF pixel_1306/ROW_SEL
+ pixel_1306/NB1 pixel_1306/VBIAS pixel_1306/NB2 pixel_1306/AMP_IN pixel_1306/SF_IB
+ pixel_1306/PIX_OUT pixel_1306/CSA_VREF pixel
Xpixel_2029 pixel_2029/gring pixel_2029/VDD pixel_2029/GND pixel_2029/VREF pixel_2029/ROW_SEL
+ pixel_2029/NB1 pixel_2029/VBIAS pixel_2029/NB2 pixel_2029/AMP_IN pixel_2029/SF_IB
+ pixel_2029/PIX_OUT pixel_2029/CSA_VREF pixel
Xpixel_1339 pixel_1339/gring pixel_1339/VDD pixel_1339/GND pixel_1339/VREF pixel_1339/ROW_SEL
+ pixel_1339/NB1 pixel_1339/VBIAS pixel_1339/NB2 pixel_1339/AMP_IN pixel_1339/SF_IB
+ pixel_1339/PIX_OUT pixel_1339/CSA_VREF pixel
Xpixel_1328 pixel_1328/gring pixel_1328/VDD pixel_1328/GND pixel_1328/VREF pixel_1328/ROW_SEL
+ pixel_1328/NB1 pixel_1328/VBIAS pixel_1328/NB2 pixel_1328/AMP_IN pixel_1328/SF_IB
+ pixel_1328/PIX_OUT pixel_1328/CSA_VREF pixel
Xpixel_1317 pixel_1317/gring pixel_1317/VDD pixel_1317/GND pixel_1317/VREF pixel_1317/ROW_SEL
+ pixel_1317/NB1 pixel_1317/VBIAS pixel_1317/NB2 pixel_1317/AMP_IN pixel_1317/SF_IB
+ pixel_1317/PIX_OUT pixel_1317/CSA_VREF pixel
Xpixel_9603 pixel_9603/gring pixel_9603/VDD pixel_9603/GND pixel_9603/VREF pixel_9603/ROW_SEL
+ pixel_9603/NB1 pixel_9603/VBIAS pixel_9603/NB2 pixel_9603/AMP_IN pixel_9603/SF_IB
+ pixel_9603/PIX_OUT pixel_9603/CSA_VREF pixel
Xpixel_9614 pixel_9614/gring pixel_9614/VDD pixel_9614/GND pixel_9614/VREF pixel_9614/ROW_SEL
+ pixel_9614/NB1 pixel_9614/VBIAS pixel_9614/NB2 pixel_9614/AMP_IN pixel_9614/SF_IB
+ pixel_9614/PIX_OUT pixel_9614/CSA_VREF pixel
Xpixel_8902 pixel_8902/gring pixel_8902/VDD pixel_8902/GND pixel_8902/VREF pixel_8902/ROW_SEL
+ pixel_8902/NB1 pixel_8902/VBIAS pixel_8902/NB2 pixel_8902/AMP_IN pixel_8902/SF_IB
+ pixel_8902/PIX_OUT pixel_8902/CSA_VREF pixel
Xpixel_9625 pixel_9625/gring pixel_9625/VDD pixel_9625/GND pixel_9625/VREF pixel_9625/ROW_SEL
+ pixel_9625/NB1 pixel_9625/VBIAS pixel_9625/NB2 pixel_9625/AMP_IN pixel_9625/SF_IB
+ pixel_9625/PIX_OUT pixel_9625/CSA_VREF pixel
Xpixel_9636 pixel_9636/gring pixel_9636/VDD pixel_9636/GND pixel_9636/VREF pixel_9636/ROW_SEL
+ pixel_9636/NB1 pixel_9636/VBIAS pixel_9636/NB2 pixel_9636/AMP_IN pixel_9636/SF_IB
+ pixel_9636/PIX_OUT pixel_9636/CSA_VREF pixel
Xpixel_9647 pixel_9647/gring pixel_9647/VDD pixel_9647/GND pixel_9647/VREF pixel_9647/ROW_SEL
+ pixel_9647/NB1 pixel_9647/VBIAS pixel_9647/NB2 pixel_9647/AMP_IN pixel_9647/SF_IB
+ pixel_9647/PIX_OUT pixel_9647/CSA_VREF pixel
Xpixel_8946 pixel_8946/gring pixel_8946/VDD pixel_8946/GND pixel_8946/VREF pixel_8946/ROW_SEL
+ pixel_8946/NB1 pixel_8946/VBIAS pixel_8946/NB2 pixel_8946/AMP_IN pixel_8946/SF_IB
+ pixel_8946/PIX_OUT pixel_8946/CSA_VREF pixel
Xpixel_8935 pixel_8935/gring pixel_8935/VDD pixel_8935/GND pixel_8935/VREF pixel_8935/ROW_SEL
+ pixel_8935/NB1 pixel_8935/VBIAS pixel_8935/NB2 pixel_8935/AMP_IN pixel_8935/SF_IB
+ pixel_8935/PIX_OUT pixel_8935/CSA_VREF pixel
Xpixel_8924 pixel_8924/gring pixel_8924/VDD pixel_8924/GND pixel_8924/VREF pixel_8924/ROW_SEL
+ pixel_8924/NB1 pixel_8924/VBIAS pixel_8924/NB2 pixel_8924/AMP_IN pixel_8924/SF_IB
+ pixel_8924/PIX_OUT pixel_8924/CSA_VREF pixel
Xpixel_8913 pixel_8913/gring pixel_8913/VDD pixel_8913/GND pixel_8913/VREF pixel_8913/ROW_SEL
+ pixel_8913/NB1 pixel_8913/VBIAS pixel_8913/NB2 pixel_8913/AMP_IN pixel_8913/SF_IB
+ pixel_8913/PIX_OUT pixel_8913/CSA_VREF pixel
Xpixel_9658 pixel_9658/gring pixel_9658/VDD pixel_9658/GND pixel_9658/VREF pixel_9658/ROW_SEL
+ pixel_9658/NB1 pixel_9658/VBIAS pixel_9658/NB2 pixel_9658/AMP_IN pixel_9658/SF_IB
+ pixel_9658/PIX_OUT pixel_9658/CSA_VREF pixel
Xpixel_9669 pixel_9669/gring pixel_9669/VDD pixel_9669/GND pixel_9669/VREF pixel_9669/ROW_SEL
+ pixel_9669/NB1 pixel_9669/VBIAS pixel_9669/NB2 pixel_9669/AMP_IN pixel_9669/SF_IB
+ pixel_9669/PIX_OUT pixel_9669/CSA_VREF pixel
Xpixel_8979 pixel_8979/gring pixel_8979/VDD pixel_8979/GND pixel_8979/VREF pixel_8979/ROW_SEL
+ pixel_8979/NB1 pixel_8979/VBIAS pixel_8979/NB2 pixel_8979/AMP_IN pixel_8979/SF_IB
+ pixel_8979/PIX_OUT pixel_8979/CSA_VREF pixel
Xpixel_8968 pixel_8968/gring pixel_8968/VDD pixel_8968/GND pixel_8968/VREF pixel_8968/ROW_SEL
+ pixel_8968/NB1 pixel_8968/VBIAS pixel_8968/NB2 pixel_8968/AMP_IN pixel_8968/SF_IB
+ pixel_8968/PIX_OUT pixel_8968/CSA_VREF pixel
Xpixel_8957 pixel_8957/gring pixel_8957/VDD pixel_8957/GND pixel_8957/VREF pixel_8957/ROW_SEL
+ pixel_8957/NB1 pixel_8957/VBIAS pixel_8957/NB2 pixel_8957/AMP_IN pixel_8957/SF_IB
+ pixel_8957/PIX_OUT pixel_8957/CSA_VREF pixel
Xpixel_3242 pixel_3242/gring pixel_3242/VDD pixel_3242/GND pixel_3242/VREF pixel_3242/ROW_SEL
+ pixel_3242/NB1 pixel_3242/VBIAS pixel_3242/NB2 pixel_3242/AMP_IN pixel_3242/SF_IB
+ pixel_3242/PIX_OUT pixel_3242/CSA_VREF pixel
Xpixel_3231 pixel_3231/gring pixel_3231/VDD pixel_3231/GND pixel_3231/VREF pixel_3231/ROW_SEL
+ pixel_3231/NB1 pixel_3231/VBIAS pixel_3231/NB2 pixel_3231/AMP_IN pixel_3231/SF_IB
+ pixel_3231/PIX_OUT pixel_3231/CSA_VREF pixel
Xpixel_3220 pixel_3220/gring pixel_3220/VDD pixel_3220/GND pixel_3220/VREF pixel_3220/ROW_SEL
+ pixel_3220/NB1 pixel_3220/VBIAS pixel_3220/NB2 pixel_3220/AMP_IN pixel_3220/SF_IB
+ pixel_3220/PIX_OUT pixel_3220/CSA_VREF pixel
Xpixel_2530 pixel_2530/gring pixel_2530/VDD pixel_2530/GND pixel_2530/VREF pixel_2530/ROW_SEL
+ pixel_2530/NB1 pixel_2530/VBIAS pixel_2530/NB2 pixel_2530/AMP_IN pixel_2530/SF_IB
+ pixel_2530/PIX_OUT pixel_2530/CSA_VREF pixel
Xpixel_3275 pixel_3275/gring pixel_3275/VDD pixel_3275/GND pixel_3275/VREF pixel_3275/ROW_SEL
+ pixel_3275/NB1 pixel_3275/VBIAS pixel_3275/NB2 pixel_3275/AMP_IN pixel_3275/SF_IB
+ pixel_3275/PIX_OUT pixel_3275/CSA_VREF pixel
Xpixel_3264 pixel_3264/gring pixel_3264/VDD pixel_3264/GND pixel_3264/VREF pixel_3264/ROW_SEL
+ pixel_3264/NB1 pixel_3264/VBIAS pixel_3264/NB2 pixel_3264/AMP_IN pixel_3264/SF_IB
+ pixel_3264/PIX_OUT pixel_3264/CSA_VREF pixel
Xpixel_3253 pixel_3253/gring pixel_3253/VDD pixel_3253/GND pixel_3253/VREF pixel_3253/ROW_SEL
+ pixel_3253/NB1 pixel_3253/VBIAS pixel_3253/NB2 pixel_3253/AMP_IN pixel_3253/SF_IB
+ pixel_3253/PIX_OUT pixel_3253/CSA_VREF pixel
Xpixel_2563 pixel_2563/gring pixel_2563/VDD pixel_2563/GND pixel_2563/VREF pixel_2563/ROW_SEL
+ pixel_2563/NB1 pixel_2563/VBIAS pixel_2563/NB2 pixel_2563/AMP_IN pixel_2563/SF_IB
+ pixel_2563/PIX_OUT pixel_2563/CSA_VREF pixel
Xpixel_2552 pixel_2552/gring pixel_2552/VDD pixel_2552/GND pixel_2552/VREF pixel_2552/ROW_SEL
+ pixel_2552/NB1 pixel_2552/VBIAS pixel_2552/NB2 pixel_2552/AMP_IN pixel_2552/SF_IB
+ pixel_2552/PIX_OUT pixel_2552/CSA_VREF pixel
Xpixel_2541 pixel_2541/gring pixel_2541/VDD pixel_2541/GND pixel_2541/VREF pixel_2541/ROW_SEL
+ pixel_2541/NB1 pixel_2541/VBIAS pixel_2541/NB2 pixel_2541/AMP_IN pixel_2541/SF_IB
+ pixel_2541/PIX_OUT pixel_2541/CSA_VREF pixel
Xpixel_3297 pixel_3297/gring pixel_3297/VDD pixel_3297/GND pixel_3297/VREF pixel_3297/ROW_SEL
+ pixel_3297/NB1 pixel_3297/VBIAS pixel_3297/NB2 pixel_3297/AMP_IN pixel_3297/SF_IB
+ pixel_3297/PIX_OUT pixel_3297/CSA_VREF pixel
Xpixel_3286 pixel_3286/gring pixel_3286/VDD pixel_3286/GND pixel_3286/VREF pixel_3286/ROW_SEL
+ pixel_3286/NB1 pixel_3286/VBIAS pixel_3286/NB2 pixel_3286/AMP_IN pixel_3286/SF_IB
+ pixel_3286/PIX_OUT pixel_3286/CSA_VREF pixel
Xpixel_1862 pixel_1862/gring pixel_1862/VDD pixel_1862/GND pixel_1862/VREF pixel_1862/ROW_SEL
+ pixel_1862/NB1 pixel_1862/VBIAS pixel_1862/NB2 pixel_1862/AMP_IN pixel_1862/SF_IB
+ pixel_1862/PIX_OUT pixel_1862/CSA_VREF pixel
Xpixel_1851 pixel_1851/gring pixel_1851/VDD pixel_1851/GND pixel_1851/VREF pixel_1851/ROW_SEL
+ pixel_1851/NB1 pixel_1851/VBIAS pixel_1851/NB2 pixel_1851/AMP_IN pixel_1851/SF_IB
+ pixel_1851/PIX_OUT pixel_1851/CSA_VREF pixel
Xpixel_1840 pixel_1840/gring pixel_1840/VDD pixel_1840/GND pixel_1840/VREF pixel_1840/ROW_SEL
+ pixel_1840/NB1 pixel_1840/VBIAS pixel_1840/NB2 pixel_1840/AMP_IN pixel_1840/SF_IB
+ pixel_1840/PIX_OUT pixel_1840/CSA_VREF pixel
Xpixel_2596 pixel_2596/gring pixel_2596/VDD pixel_2596/GND pixel_2596/VREF pixel_2596/ROW_SEL
+ pixel_2596/NB1 pixel_2596/VBIAS pixel_2596/NB2 pixel_2596/AMP_IN pixel_2596/SF_IB
+ pixel_2596/PIX_OUT pixel_2596/CSA_VREF pixel
Xpixel_2585 pixel_2585/gring pixel_2585/VDD pixel_2585/GND pixel_2585/VREF pixel_2585/ROW_SEL
+ pixel_2585/NB1 pixel_2585/VBIAS pixel_2585/NB2 pixel_2585/AMP_IN pixel_2585/SF_IB
+ pixel_2585/PIX_OUT pixel_2585/CSA_VREF pixel
Xpixel_2574 pixel_2574/gring pixel_2574/VDD pixel_2574/GND pixel_2574/VREF pixel_2574/ROW_SEL
+ pixel_2574/NB1 pixel_2574/VBIAS pixel_2574/NB2 pixel_2574/AMP_IN pixel_2574/SF_IB
+ pixel_2574/PIX_OUT pixel_2574/CSA_VREF pixel
Xpixel_1895 pixel_1895/gring pixel_1895/VDD pixel_1895/GND pixel_1895/VREF pixel_1895/ROW_SEL
+ pixel_1895/NB1 pixel_1895/VBIAS pixel_1895/NB2 pixel_1895/AMP_IN pixel_1895/SF_IB
+ pixel_1895/PIX_OUT pixel_1895/CSA_VREF pixel
Xpixel_1884 pixel_1884/gring pixel_1884/VDD pixel_1884/GND pixel_1884/VREF pixel_1884/ROW_SEL
+ pixel_1884/NB1 pixel_1884/VBIAS pixel_1884/NB2 pixel_1884/AMP_IN pixel_1884/SF_IB
+ pixel_1884/PIX_OUT pixel_1884/CSA_VREF pixel
Xpixel_1873 pixel_1873/gring pixel_1873/VDD pixel_1873/GND pixel_1873/VREF pixel_1873/ROW_SEL
+ pixel_1873/NB1 pixel_1873/VBIAS pixel_1873/NB2 pixel_1873/AMP_IN pixel_1873/SF_IB
+ pixel_1873/PIX_OUT pixel_1873/CSA_VREF pixel
Xpixel_8209 pixel_8209/gring pixel_8209/VDD pixel_8209/GND pixel_8209/VREF pixel_8209/ROW_SEL
+ pixel_8209/NB1 pixel_8209/VBIAS pixel_8209/NB2 pixel_8209/AMP_IN pixel_8209/SF_IB
+ pixel_8209/PIX_OUT pixel_8209/CSA_VREF pixel
Xpixel_7508 pixel_7508/gring pixel_7508/VDD pixel_7508/GND pixel_7508/VREF pixel_7508/ROW_SEL
+ pixel_7508/NB1 pixel_7508/VBIAS pixel_7508/NB2 pixel_7508/AMP_IN pixel_7508/SF_IB
+ pixel_7508/PIX_OUT pixel_7508/CSA_VREF pixel
Xpixel_7519 pixel_7519/gring pixel_7519/VDD pixel_7519/GND pixel_7519/VREF pixel_7519/ROW_SEL
+ pixel_7519/NB1 pixel_7519/VBIAS pixel_7519/NB2 pixel_7519/AMP_IN pixel_7519/SF_IB
+ pixel_7519/PIX_OUT pixel_7519/CSA_VREF pixel
Xpixel_6807 pixel_6807/gring pixel_6807/VDD pixel_6807/GND pixel_6807/VREF pixel_6807/ROW_SEL
+ pixel_6807/NB1 pixel_6807/VBIAS pixel_6807/NB2 pixel_6807/AMP_IN pixel_6807/SF_IB
+ pixel_6807/PIX_OUT pixel_6807/CSA_VREF pixel
Xpixel_6818 pixel_6818/gring pixel_6818/VDD pixel_6818/GND pixel_6818/VREF pixel_6818/ROW_SEL
+ pixel_6818/NB1 pixel_6818/VBIAS pixel_6818/NB2 pixel_6818/AMP_IN pixel_6818/SF_IB
+ pixel_6818/PIX_OUT pixel_6818/CSA_VREF pixel
Xpixel_6829 pixel_6829/gring pixel_6829/VDD pixel_6829/GND pixel_6829/VREF pixel_6829/ROW_SEL
+ pixel_6829/NB1 pixel_6829/VBIAS pixel_6829/NB2 pixel_6829/AMP_IN pixel_6829/SF_IB
+ pixel_6829/PIX_OUT pixel_6829/CSA_VREF pixel
Xpixel_1114 pixel_1114/gring pixel_1114/VDD pixel_1114/GND pixel_1114/VREF pixel_1114/ROW_SEL
+ pixel_1114/NB1 pixel_1114/VBIAS pixel_1114/NB2 pixel_1114/AMP_IN pixel_1114/SF_IB
+ pixel_1114/PIX_OUT pixel_1114/CSA_VREF pixel
Xpixel_1103 pixel_1103/gring pixel_1103/VDD pixel_1103/GND pixel_1103/VREF pixel_1103/ROW_SEL
+ pixel_1103/NB1 pixel_1103/VBIAS pixel_1103/NB2 pixel_1103/AMP_IN pixel_1103/SF_IB
+ pixel_1103/PIX_OUT pixel_1103/CSA_VREF pixel
Xpixel_1147 pixel_1147/gring pixel_1147/VDD pixel_1147/GND pixel_1147/VREF pixel_1147/ROW_SEL
+ pixel_1147/NB1 pixel_1147/VBIAS pixel_1147/NB2 pixel_1147/AMP_IN pixel_1147/SF_IB
+ pixel_1147/PIX_OUT pixel_1147/CSA_VREF pixel
Xpixel_1136 pixel_1136/gring pixel_1136/VDD pixel_1136/GND pixel_1136/VREF pixel_1136/ROW_SEL
+ pixel_1136/NB1 pixel_1136/VBIAS pixel_1136/NB2 pixel_1136/AMP_IN pixel_1136/SF_IB
+ pixel_1136/PIX_OUT pixel_1136/CSA_VREF pixel
Xpixel_1125 pixel_1125/gring pixel_1125/VDD pixel_1125/GND pixel_1125/VREF pixel_1125/ROW_SEL
+ pixel_1125/NB1 pixel_1125/VBIAS pixel_1125/NB2 pixel_1125/AMP_IN pixel_1125/SF_IB
+ pixel_1125/PIX_OUT pixel_1125/CSA_VREF pixel
Xpixel_1169 pixel_1169/gring pixel_1169/VDD pixel_1169/GND pixel_1169/VREF pixel_1169/ROW_SEL
+ pixel_1169/NB1 pixel_1169/VBIAS pixel_1169/NB2 pixel_1169/AMP_IN pixel_1169/SF_IB
+ pixel_1169/PIX_OUT pixel_1169/CSA_VREF pixel
Xpixel_1158 pixel_1158/gring pixel_1158/VDD pixel_1158/GND pixel_1158/VREF pixel_1158/ROW_SEL
+ pixel_1158/NB1 pixel_1158/VBIAS pixel_1158/NB2 pixel_1158/AMP_IN pixel_1158/SF_IB
+ pixel_1158/PIX_OUT pixel_1158/CSA_VREF pixel
Xpixel_9422 pixel_9422/gring pixel_9422/VDD pixel_9422/GND pixel_9422/VREF pixel_9422/ROW_SEL
+ pixel_9422/NB1 pixel_9422/VBIAS pixel_9422/NB2 pixel_9422/AMP_IN pixel_9422/SF_IB
+ pixel_9422/PIX_OUT pixel_9422/CSA_VREF pixel
Xpixel_9411 pixel_9411/gring pixel_9411/VDD pixel_9411/GND pixel_9411/VREF pixel_9411/ROW_SEL
+ pixel_9411/NB1 pixel_9411/VBIAS pixel_9411/NB2 pixel_9411/AMP_IN pixel_9411/SF_IB
+ pixel_9411/PIX_OUT pixel_9411/CSA_VREF pixel
Xpixel_9400 pixel_9400/gring pixel_9400/VDD pixel_9400/GND pixel_9400/VREF pixel_9400/ROW_SEL
+ pixel_9400/NB1 pixel_9400/VBIAS pixel_9400/NB2 pixel_9400/AMP_IN pixel_9400/SF_IB
+ pixel_9400/PIX_OUT pixel_9400/CSA_VREF pixel
Xpixel_8721 pixel_8721/gring pixel_8721/VDD pixel_8721/GND pixel_8721/VREF pixel_8721/ROW_SEL
+ pixel_8721/NB1 pixel_8721/VBIAS pixel_8721/NB2 pixel_8721/AMP_IN pixel_8721/SF_IB
+ pixel_8721/PIX_OUT pixel_8721/CSA_VREF pixel
Xpixel_8710 pixel_8710/gring pixel_8710/VDD pixel_8710/GND pixel_8710/VREF pixel_8710/ROW_SEL
+ pixel_8710/NB1 pixel_8710/VBIAS pixel_8710/NB2 pixel_8710/AMP_IN pixel_8710/SF_IB
+ pixel_8710/PIX_OUT pixel_8710/CSA_VREF pixel
Xpixel_9455 pixel_9455/gring pixel_9455/VDD pixel_9455/GND pixel_9455/VREF pixel_9455/ROW_SEL
+ pixel_9455/NB1 pixel_9455/VBIAS pixel_9455/NB2 pixel_9455/AMP_IN pixel_9455/SF_IB
+ pixel_9455/PIX_OUT pixel_9455/CSA_VREF pixel
Xpixel_9444 pixel_9444/gring pixel_9444/VDD pixel_9444/GND pixel_9444/VREF pixel_9444/ROW_SEL
+ pixel_9444/NB1 pixel_9444/VBIAS pixel_9444/NB2 pixel_9444/AMP_IN pixel_9444/SF_IB
+ pixel_9444/PIX_OUT pixel_9444/CSA_VREF pixel
Xpixel_9433 pixel_9433/gring pixel_9433/VDD pixel_9433/GND pixel_9433/VREF pixel_9433/ROW_SEL
+ pixel_9433/NB1 pixel_9433/VBIAS pixel_9433/NB2 pixel_9433/AMP_IN pixel_9433/SF_IB
+ pixel_9433/PIX_OUT pixel_9433/CSA_VREF pixel
Xpixel_8754 pixel_8754/gring pixel_8754/VDD pixel_8754/GND pixel_8754/VREF pixel_8754/ROW_SEL
+ pixel_8754/NB1 pixel_8754/VBIAS pixel_8754/NB2 pixel_8754/AMP_IN pixel_8754/SF_IB
+ pixel_8754/PIX_OUT pixel_8754/CSA_VREF pixel
Xpixel_8743 pixel_8743/gring pixel_8743/VDD pixel_8743/GND pixel_8743/VREF pixel_8743/ROW_SEL
+ pixel_8743/NB1 pixel_8743/VBIAS pixel_8743/NB2 pixel_8743/AMP_IN pixel_8743/SF_IB
+ pixel_8743/PIX_OUT pixel_8743/CSA_VREF pixel
Xpixel_8732 pixel_8732/gring pixel_8732/VDD pixel_8732/GND pixel_8732/VREF pixel_8732/ROW_SEL
+ pixel_8732/NB1 pixel_8732/VBIAS pixel_8732/NB2 pixel_8732/AMP_IN pixel_8732/SF_IB
+ pixel_8732/PIX_OUT pixel_8732/CSA_VREF pixel
Xpixel_9499 pixel_9499/gring pixel_9499/VDD pixel_9499/GND pixel_9499/VREF pixel_9499/ROW_SEL
+ pixel_9499/NB1 pixel_9499/VBIAS pixel_9499/NB2 pixel_9499/AMP_IN pixel_9499/SF_IB
+ pixel_9499/PIX_OUT pixel_9499/CSA_VREF pixel
Xpixel_9488 pixel_9488/gring pixel_9488/VDD pixel_9488/GND pixel_9488/VREF pixel_9488/ROW_SEL
+ pixel_9488/NB1 pixel_9488/VBIAS pixel_9488/NB2 pixel_9488/AMP_IN pixel_9488/SF_IB
+ pixel_9488/PIX_OUT pixel_9488/CSA_VREF pixel
Xpixel_9477 pixel_9477/gring pixel_9477/VDD pixel_9477/GND pixel_9477/VREF pixel_9477/ROW_SEL
+ pixel_9477/NB1 pixel_9477/VBIAS pixel_9477/NB2 pixel_9477/AMP_IN pixel_9477/SF_IB
+ pixel_9477/PIX_OUT pixel_9477/CSA_VREF pixel
Xpixel_9466 pixel_9466/gring pixel_9466/VDD pixel_9466/GND pixel_9466/VREF pixel_9466/ROW_SEL
+ pixel_9466/NB1 pixel_9466/VBIAS pixel_9466/NB2 pixel_9466/AMP_IN pixel_9466/SF_IB
+ pixel_9466/PIX_OUT pixel_9466/CSA_VREF pixel
Xpixel_8787 pixel_8787/gring pixel_8787/VDD pixel_8787/GND pixel_8787/VREF pixel_8787/ROW_SEL
+ pixel_8787/NB1 pixel_8787/VBIAS pixel_8787/NB2 pixel_8787/AMP_IN pixel_8787/SF_IB
+ pixel_8787/PIX_OUT pixel_8787/CSA_VREF pixel
Xpixel_8776 pixel_8776/gring pixel_8776/VDD pixel_8776/GND pixel_8776/VREF pixel_8776/ROW_SEL
+ pixel_8776/NB1 pixel_8776/VBIAS pixel_8776/NB2 pixel_8776/AMP_IN pixel_8776/SF_IB
+ pixel_8776/PIX_OUT pixel_8776/CSA_VREF pixel
Xpixel_8765 pixel_8765/gring pixel_8765/VDD pixel_8765/GND pixel_8765/VREF pixel_8765/ROW_SEL
+ pixel_8765/NB1 pixel_8765/VBIAS pixel_8765/NB2 pixel_8765/AMP_IN pixel_8765/SF_IB
+ pixel_8765/PIX_OUT pixel_8765/CSA_VREF pixel
Xpixel_8798 pixel_8798/gring pixel_8798/VDD pixel_8798/GND pixel_8798/VREF pixel_8798/ROW_SEL
+ pixel_8798/NB1 pixel_8798/VBIAS pixel_8798/NB2 pixel_8798/AMP_IN pixel_8798/SF_IB
+ pixel_8798/PIX_OUT pixel_8798/CSA_VREF pixel
Xpixel_3050 pixel_3050/gring pixel_3050/VDD pixel_3050/GND pixel_3050/VREF pixel_3050/ROW_SEL
+ pixel_3050/NB1 pixel_3050/VBIAS pixel_3050/NB2 pixel_3050/AMP_IN pixel_3050/SF_IB
+ pixel_3050/PIX_OUT pixel_3050/CSA_VREF pixel
Xpixel_3083 pixel_3083/gring pixel_3083/VDD pixel_3083/GND pixel_3083/VREF pixel_3083/ROW_SEL
+ pixel_3083/NB1 pixel_3083/VBIAS pixel_3083/NB2 pixel_3083/AMP_IN pixel_3083/SF_IB
+ pixel_3083/PIX_OUT pixel_3083/CSA_VREF pixel
Xpixel_3072 pixel_3072/gring pixel_3072/VDD pixel_3072/GND pixel_3072/VREF pixel_3072/ROW_SEL
+ pixel_3072/NB1 pixel_3072/VBIAS pixel_3072/NB2 pixel_3072/AMP_IN pixel_3072/SF_IB
+ pixel_3072/PIX_OUT pixel_3072/CSA_VREF pixel
Xpixel_3061 pixel_3061/gring pixel_3061/VDD pixel_3061/GND pixel_3061/VREF pixel_3061/ROW_SEL
+ pixel_3061/NB1 pixel_3061/VBIAS pixel_3061/NB2 pixel_3061/AMP_IN pixel_3061/SF_IB
+ pixel_3061/PIX_OUT pixel_3061/CSA_VREF pixel
Xpixel_2382 pixel_2382/gring pixel_2382/VDD pixel_2382/GND pixel_2382/VREF pixel_2382/ROW_SEL
+ pixel_2382/NB1 pixel_2382/VBIAS pixel_2382/NB2 pixel_2382/AMP_IN pixel_2382/SF_IB
+ pixel_2382/PIX_OUT pixel_2382/CSA_VREF pixel
Xpixel_2371 pixel_2371/gring pixel_2371/VDD pixel_2371/GND pixel_2371/VREF pixel_2371/ROW_SEL
+ pixel_2371/NB1 pixel_2371/VBIAS pixel_2371/NB2 pixel_2371/AMP_IN pixel_2371/SF_IB
+ pixel_2371/PIX_OUT pixel_2371/CSA_VREF pixel
Xpixel_2360 pixel_2360/gring pixel_2360/VDD pixel_2360/GND pixel_2360/VREF pixel_2360/ROW_SEL
+ pixel_2360/NB1 pixel_2360/VBIAS pixel_2360/NB2 pixel_2360/AMP_IN pixel_2360/SF_IB
+ pixel_2360/PIX_OUT pixel_2360/CSA_VREF pixel
Xpixel_3094 pixel_3094/gring pixel_3094/VDD pixel_3094/GND pixel_3094/VREF pixel_3094/ROW_SEL
+ pixel_3094/NB1 pixel_3094/VBIAS pixel_3094/NB2 pixel_3094/AMP_IN pixel_3094/SF_IB
+ pixel_3094/PIX_OUT pixel_3094/CSA_VREF pixel
Xpixel_1670 pixel_1670/gring pixel_1670/VDD pixel_1670/GND pixel_1670/VREF pixel_1670/ROW_SEL
+ pixel_1670/NB1 pixel_1670/VBIAS pixel_1670/NB2 pixel_1670/AMP_IN pixel_1670/SF_IB
+ pixel_1670/PIX_OUT pixel_1670/CSA_VREF pixel
Xpixel_2393 pixel_2393/gring pixel_2393/VDD pixel_2393/GND pixel_2393/VREF pixel_2393/ROW_SEL
+ pixel_2393/NB1 pixel_2393/VBIAS pixel_2393/NB2 pixel_2393/AMP_IN pixel_2393/SF_IB
+ pixel_2393/PIX_OUT pixel_2393/CSA_VREF pixel
Xpixel_1692 pixel_1692/gring pixel_1692/VDD pixel_1692/GND pixel_1692/VREF pixel_1692/ROW_SEL
+ pixel_1692/NB1 pixel_1692/VBIAS pixel_1692/NB2 pixel_1692/AMP_IN pixel_1692/SF_IB
+ pixel_1692/PIX_OUT pixel_1692/CSA_VREF pixel
Xpixel_1681 pixel_1681/gring pixel_1681/VDD pixel_1681/GND pixel_1681/VREF pixel_1681/ROW_SEL
+ pixel_1681/NB1 pixel_1681/VBIAS pixel_1681/NB2 pixel_1681/AMP_IN pixel_1681/SF_IB
+ pixel_1681/PIX_OUT pixel_1681/CSA_VREF pixel
Xpixel_729 pixel_729/gring pixel_729/VDD pixel_729/GND pixel_729/VREF pixel_729/ROW_SEL
+ pixel_729/NB1 pixel_729/VBIAS pixel_729/NB2 pixel_729/AMP_IN pixel_729/SF_IB pixel_729/PIX_OUT
+ pixel_729/CSA_VREF pixel
Xpixel_718 pixel_718/gring pixel_718/VDD pixel_718/GND pixel_718/VREF pixel_718/ROW_SEL
+ pixel_718/NB1 pixel_718/VBIAS pixel_718/NB2 pixel_718/AMP_IN pixel_718/SF_IB pixel_718/PIX_OUT
+ pixel_718/CSA_VREF pixel
Xpixel_707 pixel_707/gring pixel_707/VDD pixel_707/GND pixel_707/VREF pixel_707/ROW_SEL
+ pixel_707/NB1 pixel_707/VBIAS pixel_707/NB2 pixel_707/AMP_IN pixel_707/SF_IB pixel_707/PIX_OUT
+ pixel_707/CSA_VREF pixel
Xpixel_8006 pixel_8006/gring pixel_8006/VDD pixel_8006/GND pixel_8006/VREF pixel_8006/ROW_SEL
+ pixel_8006/NB1 pixel_8006/VBIAS pixel_8006/NB2 pixel_8006/AMP_IN pixel_8006/SF_IB
+ pixel_8006/PIX_OUT pixel_8006/CSA_VREF pixel
Xpixel_8017 pixel_8017/gring pixel_8017/VDD pixel_8017/GND pixel_8017/VREF pixel_8017/ROW_SEL
+ pixel_8017/NB1 pixel_8017/VBIAS pixel_8017/NB2 pixel_8017/AMP_IN pixel_8017/SF_IB
+ pixel_8017/PIX_OUT pixel_8017/CSA_VREF pixel
Xpixel_8028 pixel_8028/gring pixel_8028/VDD pixel_8028/GND pixel_8028/VREF pixel_8028/ROW_SEL
+ pixel_8028/NB1 pixel_8028/VBIAS pixel_8028/NB2 pixel_8028/AMP_IN pixel_8028/SF_IB
+ pixel_8028/PIX_OUT pixel_8028/CSA_VREF pixel
Xpixel_8039 pixel_8039/gring pixel_8039/VDD pixel_8039/GND pixel_8039/VREF pixel_8039/ROW_SEL
+ pixel_8039/NB1 pixel_8039/VBIAS pixel_8039/NB2 pixel_8039/AMP_IN pixel_8039/SF_IB
+ pixel_8039/PIX_OUT pixel_8039/CSA_VREF pixel
Xpixel_7305 pixel_7305/gring pixel_7305/VDD pixel_7305/GND pixel_7305/VREF pixel_7305/ROW_SEL
+ pixel_7305/NB1 pixel_7305/VBIAS pixel_7305/NB2 pixel_7305/AMP_IN pixel_7305/SF_IB
+ pixel_7305/PIX_OUT pixel_7305/CSA_VREF pixel
Xpixel_7316 pixel_7316/gring pixel_7316/VDD pixel_7316/GND pixel_7316/VREF pixel_7316/ROW_SEL
+ pixel_7316/NB1 pixel_7316/VBIAS pixel_7316/NB2 pixel_7316/AMP_IN pixel_7316/SF_IB
+ pixel_7316/PIX_OUT pixel_7316/CSA_VREF pixel
Xpixel_7327 pixel_7327/gring pixel_7327/VDD pixel_7327/GND pixel_7327/VREF pixel_7327/ROW_SEL
+ pixel_7327/NB1 pixel_7327/VBIAS pixel_7327/NB2 pixel_7327/AMP_IN pixel_7327/SF_IB
+ pixel_7327/PIX_OUT pixel_7327/CSA_VREF pixel
Xpixel_7338 pixel_7338/gring pixel_7338/VDD pixel_7338/GND pixel_7338/VREF pixel_7338/ROW_SEL
+ pixel_7338/NB1 pixel_7338/VBIAS pixel_7338/NB2 pixel_7338/AMP_IN pixel_7338/SF_IB
+ pixel_7338/PIX_OUT pixel_7338/CSA_VREF pixel
Xpixel_7349 pixel_7349/gring pixel_7349/VDD pixel_7349/GND pixel_7349/VREF pixel_7349/ROW_SEL
+ pixel_7349/NB1 pixel_7349/VBIAS pixel_7349/NB2 pixel_7349/AMP_IN pixel_7349/SF_IB
+ pixel_7349/PIX_OUT pixel_7349/CSA_VREF pixel
Xpixel_6604 pixel_6604/gring pixel_6604/VDD pixel_6604/GND pixel_6604/VREF pixel_6604/ROW_SEL
+ pixel_6604/NB1 pixel_6604/VBIAS pixel_6604/NB2 pixel_6604/AMP_IN pixel_6604/SF_IB
+ pixel_6604/PIX_OUT pixel_6604/CSA_VREF pixel
Xpixel_6615 pixel_6615/gring pixel_6615/VDD pixel_6615/GND pixel_6615/VREF pixel_6615/ROW_SEL
+ pixel_6615/NB1 pixel_6615/VBIAS pixel_6615/NB2 pixel_6615/AMP_IN pixel_6615/SF_IB
+ pixel_6615/PIX_OUT pixel_6615/CSA_VREF pixel
Xpixel_6626 pixel_6626/gring pixel_6626/VDD pixel_6626/GND pixel_6626/VREF pixel_6626/ROW_SEL
+ pixel_6626/NB1 pixel_6626/VBIAS pixel_6626/NB2 pixel_6626/AMP_IN pixel_6626/SF_IB
+ pixel_6626/PIX_OUT pixel_6626/CSA_VREF pixel
Xpixel_6637 pixel_6637/gring pixel_6637/VDD pixel_6637/GND pixel_6637/VREF pixel_6637/ROW_SEL
+ pixel_6637/NB1 pixel_6637/VBIAS pixel_6637/NB2 pixel_6637/AMP_IN pixel_6637/SF_IB
+ pixel_6637/PIX_OUT pixel_6637/CSA_VREF pixel
Xpixel_6648 pixel_6648/gring pixel_6648/VDD pixel_6648/GND pixel_6648/VREF pixel_6648/ROW_SEL
+ pixel_6648/NB1 pixel_6648/VBIAS pixel_6648/NB2 pixel_6648/AMP_IN pixel_6648/SF_IB
+ pixel_6648/PIX_OUT pixel_6648/CSA_VREF pixel
Xpixel_6659 pixel_6659/gring pixel_6659/VDD pixel_6659/GND pixel_6659/VREF pixel_6659/ROW_SEL
+ pixel_6659/NB1 pixel_6659/VBIAS pixel_6659/NB2 pixel_6659/AMP_IN pixel_6659/SF_IB
+ pixel_6659/PIX_OUT pixel_6659/CSA_VREF pixel
Xpixel_5903 pixel_5903/gring pixel_5903/VDD pixel_5903/GND pixel_5903/VREF pixel_5903/ROW_SEL
+ pixel_5903/NB1 pixel_5903/VBIAS pixel_5903/NB2 pixel_5903/AMP_IN pixel_5903/SF_IB
+ pixel_5903/PIX_OUT pixel_5903/CSA_VREF pixel
Xpixel_5914 pixel_5914/gring pixel_5914/VDD pixel_5914/GND pixel_5914/VREF pixel_5914/ROW_SEL
+ pixel_5914/NB1 pixel_5914/VBIAS pixel_5914/NB2 pixel_5914/AMP_IN pixel_5914/SF_IB
+ pixel_5914/PIX_OUT pixel_5914/CSA_VREF pixel
Xpixel_5925 pixel_5925/gring pixel_5925/VDD pixel_5925/GND pixel_5925/VREF pixel_5925/ROW_SEL
+ pixel_5925/NB1 pixel_5925/VBIAS pixel_5925/NB2 pixel_5925/AMP_IN pixel_5925/SF_IB
+ pixel_5925/PIX_OUT pixel_5925/CSA_VREF pixel
Xpixel_5936 pixel_5936/gring pixel_5936/VDD pixel_5936/GND pixel_5936/VREF pixel_5936/ROW_SEL
+ pixel_5936/NB1 pixel_5936/VBIAS pixel_5936/NB2 pixel_5936/AMP_IN pixel_5936/SF_IB
+ pixel_5936/PIX_OUT pixel_5936/CSA_VREF pixel
Xpixel_5947 pixel_5947/gring pixel_5947/VDD pixel_5947/GND pixel_5947/VREF pixel_5947/ROW_SEL
+ pixel_5947/NB1 pixel_5947/VBIAS pixel_5947/NB2 pixel_5947/AMP_IN pixel_5947/SF_IB
+ pixel_5947/PIX_OUT pixel_5947/CSA_VREF pixel
Xpixel_5958 pixel_5958/gring pixel_5958/VDD pixel_5958/GND pixel_5958/VREF pixel_5958/ROW_SEL
+ pixel_5958/NB1 pixel_5958/VBIAS pixel_5958/NB2 pixel_5958/AMP_IN pixel_5958/SF_IB
+ pixel_5958/PIX_OUT pixel_5958/CSA_VREF pixel
Xpixel_5969 pixel_5969/gring pixel_5969/VDD pixel_5969/GND pixel_5969/VREF pixel_5969/ROW_SEL
+ pixel_5969/NB1 pixel_5969/VBIAS pixel_5969/NB2 pixel_5969/AMP_IN pixel_5969/SF_IB
+ pixel_5969/PIX_OUT pixel_5969/CSA_VREF pixel
Xpixel_9230 pixel_9230/gring pixel_9230/VDD pixel_9230/GND pixel_9230/VREF pixel_9230/ROW_SEL
+ pixel_9230/NB1 pixel_9230/VBIAS pixel_9230/NB2 pixel_9230/AMP_IN pixel_9230/SF_IB
+ pixel_9230/PIX_OUT pixel_9230/CSA_VREF pixel
Xpixel_9274 pixel_9274/gring pixel_9274/VDD pixel_9274/GND pixel_9274/VREF pixel_9274/ROW_SEL
+ pixel_9274/NB1 pixel_9274/VBIAS pixel_9274/NB2 pixel_9274/AMP_IN pixel_9274/SF_IB
+ pixel_9274/PIX_OUT pixel_9274/CSA_VREF pixel
Xpixel_9263 pixel_9263/gring pixel_9263/VDD pixel_9263/GND pixel_9263/VREF pixel_9263/ROW_SEL
+ pixel_9263/NB1 pixel_9263/VBIAS pixel_9263/NB2 pixel_9263/AMP_IN pixel_9263/SF_IB
+ pixel_9263/PIX_OUT pixel_9263/CSA_VREF pixel
Xpixel_9252 pixel_9252/gring pixel_9252/VDD pixel_9252/GND pixel_9252/VREF pixel_9252/ROW_SEL
+ pixel_9252/NB1 pixel_9252/VBIAS pixel_9252/NB2 pixel_9252/AMP_IN pixel_9252/SF_IB
+ pixel_9252/PIX_OUT pixel_9252/CSA_VREF pixel
Xpixel_9241 pixel_9241/gring pixel_9241/VDD pixel_9241/GND pixel_9241/VREF pixel_9241/ROW_SEL
+ pixel_9241/NB1 pixel_9241/VBIAS pixel_9241/NB2 pixel_9241/AMP_IN pixel_9241/SF_IB
+ pixel_9241/PIX_OUT pixel_9241/CSA_VREF pixel
Xpixel_8562 pixel_8562/gring pixel_8562/VDD pixel_8562/GND pixel_8562/VREF pixel_8562/ROW_SEL
+ pixel_8562/NB1 pixel_8562/VBIAS pixel_8562/NB2 pixel_8562/AMP_IN pixel_8562/SF_IB
+ pixel_8562/PIX_OUT pixel_8562/CSA_VREF pixel
Xpixel_8551 pixel_8551/gring pixel_8551/VDD pixel_8551/GND pixel_8551/VREF pixel_8551/ROW_SEL
+ pixel_8551/NB1 pixel_8551/VBIAS pixel_8551/NB2 pixel_8551/AMP_IN pixel_8551/SF_IB
+ pixel_8551/PIX_OUT pixel_8551/CSA_VREF pixel
Xpixel_8540 pixel_8540/gring pixel_8540/VDD pixel_8540/GND pixel_8540/VREF pixel_8540/ROW_SEL
+ pixel_8540/NB1 pixel_8540/VBIAS pixel_8540/NB2 pixel_8540/AMP_IN pixel_8540/SF_IB
+ pixel_8540/PIX_OUT pixel_8540/CSA_VREF pixel
Xpixel_9296 pixel_9296/gring pixel_9296/VDD pixel_9296/GND pixel_9296/VREF pixel_9296/ROW_SEL
+ pixel_9296/NB1 pixel_9296/VBIAS pixel_9296/NB2 pixel_9296/AMP_IN pixel_9296/SF_IB
+ pixel_9296/PIX_OUT pixel_9296/CSA_VREF pixel
Xpixel_9285 pixel_9285/gring pixel_9285/VDD pixel_9285/GND pixel_9285/VREF pixel_9285/ROW_SEL
+ pixel_9285/NB1 pixel_9285/VBIAS pixel_9285/NB2 pixel_9285/AMP_IN pixel_9285/SF_IB
+ pixel_9285/PIX_OUT pixel_9285/CSA_VREF pixel
Xpixel_8595 pixel_8595/gring pixel_8595/VDD pixel_8595/GND pixel_8595/VREF pixel_8595/ROW_SEL
+ pixel_8595/NB1 pixel_8595/VBIAS pixel_8595/NB2 pixel_8595/AMP_IN pixel_8595/SF_IB
+ pixel_8595/PIX_OUT pixel_8595/CSA_VREF pixel
Xpixel_8584 pixel_8584/gring pixel_8584/VDD pixel_8584/GND pixel_8584/VREF pixel_8584/ROW_SEL
+ pixel_8584/NB1 pixel_8584/VBIAS pixel_8584/NB2 pixel_8584/AMP_IN pixel_8584/SF_IB
+ pixel_8584/PIX_OUT pixel_8584/CSA_VREF pixel
Xpixel_8573 pixel_8573/gring pixel_8573/VDD pixel_8573/GND pixel_8573/VREF pixel_8573/ROW_SEL
+ pixel_8573/NB1 pixel_8573/VBIAS pixel_8573/NB2 pixel_8573/AMP_IN pixel_8573/SF_IB
+ pixel_8573/PIX_OUT pixel_8573/CSA_VREF pixel
Xpixel_7850 pixel_7850/gring pixel_7850/VDD pixel_7850/GND pixel_7850/VREF pixel_7850/ROW_SEL
+ pixel_7850/NB1 pixel_7850/VBIAS pixel_7850/NB2 pixel_7850/AMP_IN pixel_7850/SF_IB
+ pixel_7850/PIX_OUT pixel_7850/CSA_VREF pixel
Xpixel_7861 pixel_7861/gring pixel_7861/VDD pixel_7861/GND pixel_7861/VREF pixel_7861/ROW_SEL
+ pixel_7861/NB1 pixel_7861/VBIAS pixel_7861/NB2 pixel_7861/AMP_IN pixel_7861/SF_IB
+ pixel_7861/PIX_OUT pixel_7861/CSA_VREF pixel
Xpixel_7872 pixel_7872/gring pixel_7872/VDD pixel_7872/GND pixel_7872/VREF pixel_7872/ROW_SEL
+ pixel_7872/NB1 pixel_7872/VBIAS pixel_7872/NB2 pixel_7872/AMP_IN pixel_7872/SF_IB
+ pixel_7872/PIX_OUT pixel_7872/CSA_VREF pixel
Xpixel_7883 pixel_7883/gring pixel_7883/VDD pixel_7883/GND pixel_7883/VREF pixel_7883/ROW_SEL
+ pixel_7883/NB1 pixel_7883/VBIAS pixel_7883/NB2 pixel_7883/AMP_IN pixel_7883/SF_IB
+ pixel_7883/PIX_OUT pixel_7883/CSA_VREF pixel
Xpixel_7894 pixel_7894/gring pixel_7894/VDD pixel_7894/GND pixel_7894/VREF pixel_7894/ROW_SEL
+ pixel_7894/NB1 pixel_7894/VBIAS pixel_7894/NB2 pixel_7894/AMP_IN pixel_7894/SF_IB
+ pixel_7894/PIX_OUT pixel_7894/CSA_VREF pixel
Xpixel_2190 pixel_2190/gring pixel_2190/VDD pixel_2190/GND pixel_2190/VREF pixel_2190/ROW_SEL
+ pixel_2190/NB1 pixel_2190/VBIAS pixel_2190/NB2 pixel_2190/AMP_IN pixel_2190/SF_IB
+ pixel_2190/PIX_OUT pixel_2190/CSA_VREF pixel
Xpixel_504 pixel_504/gring pixel_504/VDD pixel_504/GND pixel_504/VREF pixel_504/ROW_SEL
+ pixel_504/NB1 pixel_504/VBIAS pixel_504/NB2 pixel_504/AMP_IN pixel_504/SF_IB pixel_504/PIX_OUT
+ pixel_504/CSA_VREF pixel
Xpixel_4509 pixel_4509/gring pixel_4509/VDD pixel_4509/GND pixel_4509/VREF pixel_4509/ROW_SEL
+ pixel_4509/NB1 pixel_4509/VBIAS pixel_4509/NB2 pixel_4509/AMP_IN pixel_4509/SF_IB
+ pixel_4509/PIX_OUT pixel_4509/CSA_VREF pixel
Xpixel_548 pixel_548/gring pixel_548/VDD pixel_548/GND pixel_548/VREF pixel_548/ROW_SEL
+ pixel_548/NB1 pixel_548/VBIAS pixel_548/NB2 pixel_548/AMP_IN pixel_548/SF_IB pixel_548/PIX_OUT
+ pixel_548/CSA_VREF pixel
Xpixel_537 pixel_537/gring pixel_537/VDD pixel_537/GND pixel_537/VREF pixel_537/ROW_SEL
+ pixel_537/NB1 pixel_537/VBIAS pixel_537/NB2 pixel_537/AMP_IN pixel_537/SF_IB pixel_537/PIX_OUT
+ pixel_537/CSA_VREF pixel
Xpixel_526 pixel_526/gring pixel_526/VDD pixel_526/GND pixel_526/VREF pixel_526/ROW_SEL
+ pixel_526/NB1 pixel_526/VBIAS pixel_526/NB2 pixel_526/AMP_IN pixel_526/SF_IB pixel_526/PIX_OUT
+ pixel_526/CSA_VREF pixel
Xpixel_515 pixel_515/gring pixel_515/VDD pixel_515/GND pixel_515/VREF pixel_515/ROW_SEL
+ pixel_515/NB1 pixel_515/VBIAS pixel_515/NB2 pixel_515/AMP_IN pixel_515/SF_IB pixel_515/PIX_OUT
+ pixel_515/CSA_VREF pixel
Xpixel_559 pixel_559/gring pixel_559/VDD pixel_559/GND pixel_559/VREF pixel_559/ROW_SEL
+ pixel_559/NB1 pixel_559/VBIAS pixel_559/NB2 pixel_559/AMP_IN pixel_559/SF_IB pixel_559/PIX_OUT
+ pixel_559/CSA_VREF pixel
Xpixel_3808 pixel_3808/gring pixel_3808/VDD pixel_3808/GND pixel_3808/VREF pixel_3808/ROW_SEL
+ pixel_3808/NB1 pixel_3808/VBIAS pixel_3808/NB2 pixel_3808/AMP_IN pixel_3808/SF_IB
+ pixel_3808/PIX_OUT pixel_3808/CSA_VREF pixel
Xpixel_3819 pixel_3819/gring pixel_3819/VDD pixel_3819/GND pixel_3819/VREF pixel_3819/ROW_SEL
+ pixel_3819/NB1 pixel_3819/VBIAS pixel_3819/NB2 pixel_3819/AMP_IN pixel_3819/SF_IB
+ pixel_3819/PIX_OUT pixel_3819/CSA_VREF pixel
Xpixel_7102 pixel_7102/gring pixel_7102/VDD pixel_7102/GND pixel_7102/VREF pixel_7102/ROW_SEL
+ pixel_7102/NB1 pixel_7102/VBIAS pixel_7102/NB2 pixel_7102/AMP_IN pixel_7102/SF_IB
+ pixel_7102/PIX_OUT pixel_7102/CSA_VREF pixel
Xpixel_7113 pixel_7113/gring pixel_7113/VDD pixel_7113/GND pixel_7113/VREF pixel_7113/ROW_SEL
+ pixel_7113/NB1 pixel_7113/VBIAS pixel_7113/NB2 pixel_7113/AMP_IN pixel_7113/SF_IB
+ pixel_7113/PIX_OUT pixel_7113/CSA_VREF pixel
Xpixel_7124 pixel_7124/gring pixel_7124/VDD pixel_7124/GND pixel_7124/VREF pixel_7124/ROW_SEL
+ pixel_7124/NB1 pixel_7124/VBIAS pixel_7124/NB2 pixel_7124/AMP_IN pixel_7124/SF_IB
+ pixel_7124/PIX_OUT pixel_7124/CSA_VREF pixel
Xpixel_7135 pixel_7135/gring pixel_7135/VDD pixel_7135/GND pixel_7135/VREF pixel_7135/ROW_SEL
+ pixel_7135/NB1 pixel_7135/VBIAS pixel_7135/NB2 pixel_7135/AMP_IN pixel_7135/SF_IB
+ pixel_7135/PIX_OUT pixel_7135/CSA_VREF pixel
Xpixel_7146 pixel_7146/gring pixel_7146/VDD pixel_7146/GND pixel_7146/VREF pixel_7146/ROW_SEL
+ pixel_7146/NB1 pixel_7146/VBIAS pixel_7146/NB2 pixel_7146/AMP_IN pixel_7146/SF_IB
+ pixel_7146/PIX_OUT pixel_7146/CSA_VREF pixel
Xpixel_6401 pixel_6401/gring pixel_6401/VDD pixel_6401/GND pixel_6401/VREF pixel_6401/ROW_SEL
+ pixel_6401/NB1 pixel_6401/VBIAS pixel_6401/NB2 pixel_6401/AMP_IN pixel_6401/SF_IB
+ pixel_6401/PIX_OUT pixel_6401/CSA_VREF pixel
Xpixel_7157 pixel_7157/gring pixel_7157/VDD pixel_7157/GND pixel_7157/VREF pixel_7157/ROW_SEL
+ pixel_7157/NB1 pixel_7157/VBIAS pixel_7157/NB2 pixel_7157/AMP_IN pixel_7157/SF_IB
+ pixel_7157/PIX_OUT pixel_7157/CSA_VREF pixel
Xpixel_7168 pixel_7168/gring pixel_7168/VDD pixel_7168/GND pixel_7168/VREF pixel_7168/ROW_SEL
+ pixel_7168/NB1 pixel_7168/VBIAS pixel_7168/NB2 pixel_7168/AMP_IN pixel_7168/SF_IB
+ pixel_7168/PIX_OUT pixel_7168/CSA_VREF pixel
Xpixel_7179 pixel_7179/gring pixel_7179/VDD pixel_7179/GND pixel_7179/VREF pixel_7179/ROW_SEL
+ pixel_7179/NB1 pixel_7179/VBIAS pixel_7179/NB2 pixel_7179/AMP_IN pixel_7179/SF_IB
+ pixel_7179/PIX_OUT pixel_7179/CSA_VREF pixel
Xpixel_6412 pixel_6412/gring pixel_6412/VDD pixel_6412/GND pixel_6412/VREF pixel_6412/ROW_SEL
+ pixel_6412/NB1 pixel_6412/VBIAS pixel_6412/NB2 pixel_6412/AMP_IN pixel_6412/SF_IB
+ pixel_6412/PIX_OUT pixel_6412/CSA_VREF pixel
Xpixel_6423 pixel_6423/gring pixel_6423/VDD pixel_6423/GND pixel_6423/VREF pixel_6423/ROW_SEL
+ pixel_6423/NB1 pixel_6423/VBIAS pixel_6423/NB2 pixel_6423/AMP_IN pixel_6423/SF_IB
+ pixel_6423/PIX_OUT pixel_6423/CSA_VREF pixel
Xpixel_6434 pixel_6434/gring pixel_6434/VDD pixel_6434/GND pixel_6434/VREF pixel_6434/ROW_SEL
+ pixel_6434/NB1 pixel_6434/VBIAS pixel_6434/NB2 pixel_6434/AMP_IN pixel_6434/SF_IB
+ pixel_6434/PIX_OUT pixel_6434/CSA_VREF pixel
Xpixel_6445 pixel_6445/gring pixel_6445/VDD pixel_6445/GND pixel_6445/VREF pixel_6445/ROW_SEL
+ pixel_6445/NB1 pixel_6445/VBIAS pixel_6445/NB2 pixel_6445/AMP_IN pixel_6445/SF_IB
+ pixel_6445/PIX_OUT pixel_6445/CSA_VREF pixel
Xpixel_5700 pixel_5700/gring pixel_5700/VDD pixel_5700/GND pixel_5700/VREF pixel_5700/ROW_SEL
+ pixel_5700/NB1 pixel_5700/VBIAS pixel_5700/NB2 pixel_5700/AMP_IN pixel_5700/SF_IB
+ pixel_5700/PIX_OUT pixel_5700/CSA_VREF pixel
Xpixel_6456 pixel_6456/gring pixel_6456/VDD pixel_6456/GND pixel_6456/VREF pixel_6456/ROW_SEL
+ pixel_6456/NB1 pixel_6456/VBIAS pixel_6456/NB2 pixel_6456/AMP_IN pixel_6456/SF_IB
+ pixel_6456/PIX_OUT pixel_6456/CSA_VREF pixel
Xpixel_6467 pixel_6467/gring pixel_6467/VDD pixel_6467/GND pixel_6467/VREF pixel_6467/ROW_SEL
+ pixel_6467/NB1 pixel_6467/VBIAS pixel_6467/NB2 pixel_6467/AMP_IN pixel_6467/SF_IB
+ pixel_6467/PIX_OUT pixel_6467/CSA_VREF pixel
Xpixel_6478 pixel_6478/gring pixel_6478/VDD pixel_6478/GND pixel_6478/VREF pixel_6478/ROW_SEL
+ pixel_6478/NB1 pixel_6478/VBIAS pixel_6478/NB2 pixel_6478/AMP_IN pixel_6478/SF_IB
+ pixel_6478/PIX_OUT pixel_6478/CSA_VREF pixel
Xpixel_5711 pixel_5711/gring pixel_5711/VDD pixel_5711/GND pixel_5711/VREF pixel_5711/ROW_SEL
+ pixel_5711/NB1 pixel_5711/VBIAS pixel_5711/NB2 pixel_5711/AMP_IN pixel_5711/SF_IB
+ pixel_5711/PIX_OUT pixel_5711/CSA_VREF pixel
Xpixel_5722 pixel_5722/gring pixel_5722/VDD pixel_5722/GND pixel_5722/VREF pixel_5722/ROW_SEL
+ pixel_5722/NB1 pixel_5722/VBIAS pixel_5722/NB2 pixel_5722/AMP_IN pixel_5722/SF_IB
+ pixel_5722/PIX_OUT pixel_5722/CSA_VREF pixel
Xpixel_5733 pixel_5733/gring pixel_5733/VDD pixel_5733/GND pixel_5733/VREF pixel_5733/ROW_SEL
+ pixel_5733/NB1 pixel_5733/VBIAS pixel_5733/NB2 pixel_5733/AMP_IN pixel_5733/SF_IB
+ pixel_5733/PIX_OUT pixel_5733/CSA_VREF pixel
Xpixel_6489 pixel_6489/gring pixel_6489/VDD pixel_6489/GND pixel_6489/VREF pixel_6489/ROW_SEL
+ pixel_6489/NB1 pixel_6489/VBIAS pixel_6489/NB2 pixel_6489/AMP_IN pixel_6489/SF_IB
+ pixel_6489/PIX_OUT pixel_6489/CSA_VREF pixel
Xpixel_5744 pixel_5744/gring pixel_5744/VDD pixel_5744/GND pixel_5744/VREF pixel_5744/ROW_SEL
+ pixel_5744/NB1 pixel_5744/VBIAS pixel_5744/NB2 pixel_5744/AMP_IN pixel_5744/SF_IB
+ pixel_5744/PIX_OUT pixel_5744/CSA_VREF pixel
Xpixel_5755 pixel_5755/gring pixel_5755/VDD pixel_5755/GND pixel_5755/VREF pixel_5755/ROW_SEL
+ pixel_5755/NB1 pixel_5755/VBIAS pixel_5755/NB2 pixel_5755/AMP_IN pixel_5755/SF_IB
+ pixel_5755/PIX_OUT pixel_5755/CSA_VREF pixel
Xpixel_5766 pixel_5766/gring pixel_5766/VDD pixel_5766/GND pixel_5766/VREF pixel_5766/ROW_SEL
+ pixel_5766/NB1 pixel_5766/VBIAS pixel_5766/NB2 pixel_5766/AMP_IN pixel_5766/SF_IB
+ pixel_5766/PIX_OUT pixel_5766/CSA_VREF pixel
Xpixel_5777 pixel_5777/gring pixel_5777/VDD pixel_5777/GND pixel_5777/VREF pixel_5777/ROW_SEL
+ pixel_5777/NB1 pixel_5777/VBIAS pixel_5777/NB2 pixel_5777/AMP_IN pixel_5777/SF_IB
+ pixel_5777/PIX_OUT pixel_5777/CSA_VREF pixel
Xpixel_5788 pixel_5788/gring pixel_5788/VDD pixel_5788/GND pixel_5788/VREF pixel_5788/ROW_SEL
+ pixel_5788/NB1 pixel_5788/VBIAS pixel_5788/NB2 pixel_5788/AMP_IN pixel_5788/SF_IB
+ pixel_5788/PIX_OUT pixel_5788/CSA_VREF pixel
Xpixel_5799 pixel_5799/gring pixel_5799/VDD pixel_5799/GND pixel_5799/VREF pixel_5799/ROW_SEL
+ pixel_5799/NB1 pixel_5799/VBIAS pixel_5799/NB2 pixel_5799/AMP_IN pixel_5799/SF_IB
+ pixel_5799/PIX_OUT pixel_5799/CSA_VREF pixel
Xpixel_9082 pixel_9082/gring pixel_9082/VDD pixel_9082/GND pixel_9082/VREF pixel_9082/ROW_SEL
+ pixel_9082/NB1 pixel_9082/VBIAS pixel_9082/NB2 pixel_9082/AMP_IN pixel_9082/SF_IB
+ pixel_9082/PIX_OUT pixel_9082/CSA_VREF pixel
Xpixel_9071 pixel_9071/gring pixel_9071/VDD pixel_9071/GND pixel_9071/VREF pixel_9071/ROW_SEL
+ pixel_9071/NB1 pixel_9071/VBIAS pixel_9071/NB2 pixel_9071/AMP_IN pixel_9071/SF_IB
+ pixel_9071/PIX_OUT pixel_9071/CSA_VREF pixel
Xpixel_9060 pixel_9060/gring pixel_9060/VDD pixel_9060/GND pixel_9060/VREF pixel_9060/ROW_SEL
+ pixel_9060/NB1 pixel_9060/VBIAS pixel_9060/NB2 pixel_9060/AMP_IN pixel_9060/SF_IB
+ pixel_9060/PIX_OUT pixel_9060/CSA_VREF pixel
Xpixel_9093 pixel_9093/gring pixel_9093/VDD pixel_9093/GND pixel_9093/VREF pixel_9093/ROW_SEL
+ pixel_9093/NB1 pixel_9093/VBIAS pixel_9093/NB2 pixel_9093/AMP_IN pixel_9093/SF_IB
+ pixel_9093/PIX_OUT pixel_9093/CSA_VREF pixel
Xpixel_8370 pixel_8370/gring pixel_8370/VDD pixel_8370/GND pixel_8370/VREF pixel_8370/ROW_SEL
+ pixel_8370/NB1 pixel_8370/VBIAS pixel_8370/NB2 pixel_8370/AMP_IN pixel_8370/SF_IB
+ pixel_8370/PIX_OUT pixel_8370/CSA_VREF pixel
Xpixel_8381 pixel_8381/gring pixel_8381/VDD pixel_8381/GND pixel_8381/VREF pixel_8381/ROW_SEL
+ pixel_8381/NB1 pixel_8381/VBIAS pixel_8381/NB2 pixel_8381/AMP_IN pixel_8381/SF_IB
+ pixel_8381/PIX_OUT pixel_8381/CSA_VREF pixel
Xpixel_8392 pixel_8392/gring pixel_8392/VDD pixel_8392/GND pixel_8392/VREF pixel_8392/ROW_SEL
+ pixel_8392/NB1 pixel_8392/VBIAS pixel_8392/NB2 pixel_8392/AMP_IN pixel_8392/SF_IB
+ pixel_8392/PIX_OUT pixel_8392/CSA_VREF pixel
Xpixel_7680 pixel_7680/gring pixel_7680/VDD pixel_7680/GND pixel_7680/VREF pixel_7680/ROW_SEL
+ pixel_7680/NB1 pixel_7680/VBIAS pixel_7680/NB2 pixel_7680/AMP_IN pixel_7680/SF_IB
+ pixel_7680/PIX_OUT pixel_7680/CSA_VREF pixel
Xpixel_7691 pixel_7691/gring pixel_7691/VDD pixel_7691/GND pixel_7691/VREF pixel_7691/ROW_SEL
+ pixel_7691/NB1 pixel_7691/VBIAS pixel_7691/NB2 pixel_7691/AMP_IN pixel_7691/SF_IB
+ pixel_7691/PIX_OUT pixel_7691/CSA_VREF pixel
Xpixel_6990 pixel_6990/gring pixel_6990/VDD pixel_6990/GND pixel_6990/VREF pixel_6990/ROW_SEL
+ pixel_6990/NB1 pixel_6990/VBIAS pixel_6990/NB2 pixel_6990/AMP_IN pixel_6990/SF_IB
+ pixel_6990/PIX_OUT pixel_6990/CSA_VREF pixel
Xpixel_82 pixel_82/gring pixel_82/VDD pixel_82/GND pixel_82/VREF pixel_82/ROW_SEL
+ pixel_82/NB1 pixel_82/VBIAS pixel_82/NB2 pixel_82/AMP_IN pixel_82/SF_IB pixel_82/PIX_OUT
+ pixel_82/CSA_VREF pixel
Xpixel_71 pixel_71/gring pixel_71/VDD pixel_71/GND pixel_71/VREF pixel_71/ROW_SEL
+ pixel_71/NB1 pixel_71/VBIAS pixel_71/NB2 pixel_71/AMP_IN pixel_71/SF_IB pixel_71/PIX_OUT
+ pixel_71/CSA_VREF pixel
Xpixel_60 pixel_60/gring pixel_60/VDD pixel_60/GND pixel_60/VREF pixel_60/ROW_SEL
+ pixel_60/NB1 pixel_60/VBIAS pixel_60/NB2 pixel_60/AMP_IN pixel_60/SF_IB pixel_60/PIX_OUT
+ pixel_60/CSA_VREF pixel
Xpixel_93 pixel_93/gring pixel_93/VDD pixel_93/GND pixel_93/VREF pixel_93/ROW_SEL
+ pixel_93/NB1 pixel_93/VBIAS pixel_93/NB2 pixel_93/AMP_IN pixel_93/SF_IB pixel_93/PIX_OUT
+ pixel_93/CSA_VREF pixel
Xpixel_5007 pixel_5007/gring pixel_5007/VDD pixel_5007/GND pixel_5007/VREF pixel_5007/ROW_SEL
+ pixel_5007/NB1 pixel_5007/VBIAS pixel_5007/NB2 pixel_5007/AMP_IN pixel_5007/SF_IB
+ pixel_5007/PIX_OUT pixel_5007/CSA_VREF pixel
Xpixel_5018 pixel_5018/gring pixel_5018/VDD pixel_5018/GND pixel_5018/VREF pixel_5018/ROW_SEL
+ pixel_5018/NB1 pixel_5018/VBIAS pixel_5018/NB2 pixel_5018/AMP_IN pixel_5018/SF_IB
+ pixel_5018/PIX_OUT pixel_5018/CSA_VREF pixel
Xpixel_5029 pixel_5029/gring pixel_5029/VDD pixel_5029/GND pixel_5029/VREF pixel_5029/ROW_SEL
+ pixel_5029/NB1 pixel_5029/VBIAS pixel_5029/NB2 pixel_5029/AMP_IN pixel_5029/SF_IB
+ pixel_5029/PIX_OUT pixel_5029/CSA_VREF pixel
Xpixel_312 pixel_312/gring pixel_312/VDD pixel_312/GND pixel_312/VREF pixel_312/ROW_SEL
+ pixel_312/NB1 pixel_312/VBIAS pixel_312/NB2 pixel_312/AMP_IN pixel_312/SF_IB pixel_312/PIX_OUT
+ pixel_312/CSA_VREF pixel
Xpixel_301 pixel_301/gring pixel_301/VDD pixel_301/GND pixel_301/VREF pixel_301/ROW_SEL
+ pixel_301/NB1 pixel_301/VBIAS pixel_301/NB2 pixel_301/AMP_IN pixel_301/SF_IB pixel_301/PIX_OUT
+ pixel_301/CSA_VREF pixel
Xpixel_4306 pixel_4306/gring pixel_4306/VDD pixel_4306/GND pixel_4306/VREF pixel_4306/ROW_SEL
+ pixel_4306/NB1 pixel_4306/VBIAS pixel_4306/NB2 pixel_4306/AMP_IN pixel_4306/SF_IB
+ pixel_4306/PIX_OUT pixel_4306/CSA_VREF pixel
Xpixel_4317 pixel_4317/gring pixel_4317/VDD pixel_4317/GND pixel_4317/VREF pixel_4317/ROW_SEL
+ pixel_4317/NB1 pixel_4317/VBIAS pixel_4317/NB2 pixel_4317/AMP_IN pixel_4317/SF_IB
+ pixel_4317/PIX_OUT pixel_4317/CSA_VREF pixel
Xpixel_356 pixel_356/gring pixel_356/VDD pixel_356/GND pixel_356/VREF pixel_356/ROW_SEL
+ pixel_356/NB1 pixel_356/VBIAS pixel_356/NB2 pixel_356/AMP_IN pixel_356/SF_IB pixel_356/PIX_OUT
+ pixel_356/CSA_VREF pixel
Xpixel_345 pixel_345/gring pixel_345/VDD pixel_345/GND pixel_345/VREF pixel_345/ROW_SEL
+ pixel_345/NB1 pixel_345/VBIAS pixel_345/NB2 pixel_345/AMP_IN pixel_345/SF_IB pixel_345/PIX_OUT
+ pixel_345/CSA_VREF pixel
Xpixel_334 pixel_334/gring pixel_334/VDD pixel_334/GND pixel_334/VREF pixel_334/ROW_SEL
+ pixel_334/NB1 pixel_334/VBIAS pixel_334/NB2 pixel_334/AMP_IN pixel_334/SF_IB pixel_334/PIX_OUT
+ pixel_334/CSA_VREF pixel
Xpixel_323 pixel_323/gring pixel_323/VDD pixel_323/GND pixel_323/VREF pixel_323/ROW_SEL
+ pixel_323/NB1 pixel_323/VBIAS pixel_323/NB2 pixel_323/AMP_IN pixel_323/SF_IB pixel_323/PIX_OUT
+ pixel_323/CSA_VREF pixel
Xpixel_3616 pixel_3616/gring pixel_3616/VDD pixel_3616/GND pixel_3616/VREF pixel_3616/ROW_SEL
+ pixel_3616/NB1 pixel_3616/VBIAS pixel_3616/NB2 pixel_3616/AMP_IN pixel_3616/SF_IB
+ pixel_3616/PIX_OUT pixel_3616/CSA_VREF pixel
Xpixel_3605 pixel_3605/gring pixel_3605/VDD pixel_3605/GND pixel_3605/VREF pixel_3605/ROW_SEL
+ pixel_3605/NB1 pixel_3605/VBIAS pixel_3605/NB2 pixel_3605/AMP_IN pixel_3605/SF_IB
+ pixel_3605/PIX_OUT pixel_3605/CSA_VREF pixel
Xpixel_4328 pixel_4328/gring pixel_4328/VDD pixel_4328/GND pixel_4328/VREF pixel_4328/ROW_SEL
+ pixel_4328/NB1 pixel_4328/VBIAS pixel_4328/NB2 pixel_4328/AMP_IN pixel_4328/SF_IB
+ pixel_4328/PIX_OUT pixel_4328/CSA_VREF pixel
Xpixel_4339 pixel_4339/gring pixel_4339/VDD pixel_4339/GND pixel_4339/VREF pixel_4339/ROW_SEL
+ pixel_4339/NB1 pixel_4339/VBIAS pixel_4339/NB2 pixel_4339/AMP_IN pixel_4339/SF_IB
+ pixel_4339/PIX_OUT pixel_4339/CSA_VREF pixel
Xpixel_389 pixel_389/gring pixel_389/VDD pixel_389/GND pixel_389/VREF pixel_389/ROW_SEL
+ pixel_389/NB1 pixel_389/VBIAS pixel_389/NB2 pixel_389/AMP_IN pixel_389/SF_IB pixel_389/PIX_OUT
+ pixel_389/CSA_VREF pixel
Xpixel_378 pixel_378/gring pixel_378/VDD pixel_378/GND pixel_378/VREF pixel_378/ROW_SEL
+ pixel_378/NB1 pixel_378/VBIAS pixel_378/NB2 pixel_378/AMP_IN pixel_378/SF_IB pixel_378/PIX_OUT
+ pixel_378/CSA_VREF pixel
Xpixel_367 pixel_367/gring pixel_367/VDD pixel_367/GND pixel_367/VREF pixel_367/ROW_SEL
+ pixel_367/NB1 pixel_367/VBIAS pixel_367/NB2 pixel_367/AMP_IN pixel_367/SF_IB pixel_367/PIX_OUT
+ pixel_367/CSA_VREF pixel
Xpixel_2904 pixel_2904/gring pixel_2904/VDD pixel_2904/GND pixel_2904/VREF pixel_2904/ROW_SEL
+ pixel_2904/NB1 pixel_2904/VBIAS pixel_2904/NB2 pixel_2904/AMP_IN pixel_2904/SF_IB
+ pixel_2904/PIX_OUT pixel_2904/CSA_VREF pixel
Xpixel_3649 pixel_3649/gring pixel_3649/VDD pixel_3649/GND pixel_3649/VREF pixel_3649/ROW_SEL
+ pixel_3649/NB1 pixel_3649/VBIAS pixel_3649/NB2 pixel_3649/AMP_IN pixel_3649/SF_IB
+ pixel_3649/PIX_OUT pixel_3649/CSA_VREF pixel
Xpixel_3638 pixel_3638/gring pixel_3638/VDD pixel_3638/GND pixel_3638/VREF pixel_3638/ROW_SEL
+ pixel_3638/NB1 pixel_3638/VBIAS pixel_3638/NB2 pixel_3638/AMP_IN pixel_3638/SF_IB
+ pixel_3638/PIX_OUT pixel_3638/CSA_VREF pixel
Xpixel_3627 pixel_3627/gring pixel_3627/VDD pixel_3627/GND pixel_3627/VREF pixel_3627/ROW_SEL
+ pixel_3627/NB1 pixel_3627/VBIAS pixel_3627/NB2 pixel_3627/AMP_IN pixel_3627/SF_IB
+ pixel_3627/PIX_OUT pixel_3627/CSA_VREF pixel
Xpixel_2937 pixel_2937/gring pixel_2937/VDD pixel_2937/GND pixel_2937/VREF pixel_2937/ROW_SEL
+ pixel_2937/NB1 pixel_2937/VBIAS pixel_2937/NB2 pixel_2937/AMP_IN pixel_2937/SF_IB
+ pixel_2937/PIX_OUT pixel_2937/CSA_VREF pixel
Xpixel_2926 pixel_2926/gring pixel_2926/VDD pixel_2926/GND pixel_2926/VREF pixel_2926/ROW_SEL
+ pixel_2926/NB1 pixel_2926/VBIAS pixel_2926/NB2 pixel_2926/AMP_IN pixel_2926/SF_IB
+ pixel_2926/PIX_OUT pixel_2926/CSA_VREF pixel
Xpixel_2915 pixel_2915/gring pixel_2915/VDD pixel_2915/GND pixel_2915/VREF pixel_2915/ROW_SEL
+ pixel_2915/NB1 pixel_2915/VBIAS pixel_2915/NB2 pixel_2915/AMP_IN pixel_2915/SF_IB
+ pixel_2915/PIX_OUT pixel_2915/CSA_VREF pixel
Xpixel_2959 pixel_2959/gring pixel_2959/VDD pixel_2959/GND pixel_2959/VREF pixel_2959/ROW_SEL
+ pixel_2959/NB1 pixel_2959/VBIAS pixel_2959/NB2 pixel_2959/AMP_IN pixel_2959/SF_IB
+ pixel_2959/PIX_OUT pixel_2959/CSA_VREF pixel
Xpixel_2948 pixel_2948/gring pixel_2948/VDD pixel_2948/GND pixel_2948/VREF pixel_2948/ROW_SEL
+ pixel_2948/NB1 pixel_2948/VBIAS pixel_2948/NB2 pixel_2948/AMP_IN pixel_2948/SF_IB
+ pixel_2948/PIX_OUT pixel_2948/CSA_VREF pixel
Xpixel_6220 pixel_6220/gring pixel_6220/VDD pixel_6220/GND pixel_6220/VREF pixel_6220/ROW_SEL
+ pixel_6220/NB1 pixel_6220/VBIAS pixel_6220/NB2 pixel_6220/AMP_IN pixel_6220/SF_IB
+ pixel_6220/PIX_OUT pixel_6220/CSA_VREF pixel
Xpixel_6231 pixel_6231/gring pixel_6231/VDD pixel_6231/GND pixel_6231/VREF pixel_6231/ROW_SEL
+ pixel_6231/NB1 pixel_6231/VBIAS pixel_6231/NB2 pixel_6231/AMP_IN pixel_6231/SF_IB
+ pixel_6231/PIX_OUT pixel_6231/CSA_VREF pixel
Xpixel_6242 pixel_6242/gring pixel_6242/VDD pixel_6242/GND pixel_6242/VREF pixel_6242/ROW_SEL
+ pixel_6242/NB1 pixel_6242/VBIAS pixel_6242/NB2 pixel_6242/AMP_IN pixel_6242/SF_IB
+ pixel_6242/PIX_OUT pixel_6242/CSA_VREF pixel
Xpixel_6253 pixel_6253/gring pixel_6253/VDD pixel_6253/GND pixel_6253/VREF pixel_6253/ROW_SEL
+ pixel_6253/NB1 pixel_6253/VBIAS pixel_6253/NB2 pixel_6253/AMP_IN pixel_6253/SF_IB
+ pixel_6253/PIX_OUT pixel_6253/CSA_VREF pixel
Xpixel_6264 pixel_6264/gring pixel_6264/VDD pixel_6264/GND pixel_6264/VREF pixel_6264/ROW_SEL
+ pixel_6264/NB1 pixel_6264/VBIAS pixel_6264/NB2 pixel_6264/AMP_IN pixel_6264/SF_IB
+ pixel_6264/PIX_OUT pixel_6264/CSA_VREF pixel
Xpixel_6275 pixel_6275/gring pixel_6275/VDD pixel_6275/GND pixel_6275/VREF pixel_6275/ROW_SEL
+ pixel_6275/NB1 pixel_6275/VBIAS pixel_6275/NB2 pixel_6275/AMP_IN pixel_6275/SF_IB
+ pixel_6275/PIX_OUT pixel_6275/CSA_VREF pixel
Xpixel_6286 pixel_6286/gring pixel_6286/VDD pixel_6286/GND pixel_6286/VREF pixel_6286/ROW_SEL
+ pixel_6286/NB1 pixel_6286/VBIAS pixel_6286/NB2 pixel_6286/AMP_IN pixel_6286/SF_IB
+ pixel_6286/PIX_OUT pixel_6286/CSA_VREF pixel
Xpixel_5530 pixel_5530/gring pixel_5530/VDD pixel_5530/GND pixel_5530/VREF pixel_5530/ROW_SEL
+ pixel_5530/NB1 pixel_5530/VBIAS pixel_5530/NB2 pixel_5530/AMP_IN pixel_5530/SF_IB
+ pixel_5530/PIX_OUT pixel_5530/CSA_VREF pixel
Xpixel_5541 pixel_5541/gring pixel_5541/VDD pixel_5541/GND pixel_5541/VREF pixel_5541/ROW_SEL
+ pixel_5541/NB1 pixel_5541/VBIAS pixel_5541/NB2 pixel_5541/AMP_IN pixel_5541/SF_IB
+ pixel_5541/PIX_OUT pixel_5541/CSA_VREF pixel
Xpixel_6297 pixel_6297/gring pixel_6297/VDD pixel_6297/GND pixel_6297/VREF pixel_6297/ROW_SEL
+ pixel_6297/NB1 pixel_6297/VBIAS pixel_6297/NB2 pixel_6297/AMP_IN pixel_6297/SF_IB
+ pixel_6297/PIX_OUT pixel_6297/CSA_VREF pixel
Xpixel_5552 pixel_5552/gring pixel_5552/VDD pixel_5552/GND pixel_5552/VREF pixel_5552/ROW_SEL
+ pixel_5552/NB1 pixel_5552/VBIAS pixel_5552/NB2 pixel_5552/AMP_IN pixel_5552/SF_IB
+ pixel_5552/PIX_OUT pixel_5552/CSA_VREF pixel
Xpixel_5563 pixel_5563/gring pixel_5563/VDD pixel_5563/GND pixel_5563/VREF pixel_5563/ROW_SEL
+ pixel_5563/NB1 pixel_5563/VBIAS pixel_5563/NB2 pixel_5563/AMP_IN pixel_5563/SF_IB
+ pixel_5563/PIX_OUT pixel_5563/CSA_VREF pixel
Xpixel_5574 pixel_5574/gring pixel_5574/VDD pixel_5574/GND pixel_5574/VREF pixel_5574/ROW_SEL
+ pixel_5574/NB1 pixel_5574/VBIAS pixel_5574/NB2 pixel_5574/AMP_IN pixel_5574/SF_IB
+ pixel_5574/PIX_OUT pixel_5574/CSA_VREF pixel
Xpixel_5585 pixel_5585/gring pixel_5585/VDD pixel_5585/GND pixel_5585/VREF pixel_5585/ROW_SEL
+ pixel_5585/NB1 pixel_5585/VBIAS pixel_5585/NB2 pixel_5585/AMP_IN pixel_5585/SF_IB
+ pixel_5585/PIX_OUT pixel_5585/CSA_VREF pixel
Xpixel_4840 pixel_4840/gring pixel_4840/VDD pixel_4840/GND pixel_4840/VREF pixel_4840/ROW_SEL
+ pixel_4840/NB1 pixel_4840/VBIAS pixel_4840/NB2 pixel_4840/AMP_IN pixel_4840/SF_IB
+ pixel_4840/PIX_OUT pixel_4840/CSA_VREF pixel
Xpixel_5596 pixel_5596/gring pixel_5596/VDD pixel_5596/GND pixel_5596/VREF pixel_5596/ROW_SEL
+ pixel_5596/NB1 pixel_5596/VBIAS pixel_5596/NB2 pixel_5596/AMP_IN pixel_5596/SF_IB
+ pixel_5596/PIX_OUT pixel_5596/CSA_VREF pixel
Xpixel_4851 pixel_4851/gring pixel_4851/VDD pixel_4851/GND pixel_4851/VREF pixel_4851/ROW_SEL
+ pixel_4851/NB1 pixel_4851/VBIAS pixel_4851/NB2 pixel_4851/AMP_IN pixel_4851/SF_IB
+ pixel_4851/PIX_OUT pixel_4851/CSA_VREF pixel
Xpixel_4862 pixel_4862/gring pixel_4862/VDD pixel_4862/GND pixel_4862/VREF pixel_4862/ROW_SEL
+ pixel_4862/NB1 pixel_4862/VBIAS pixel_4862/NB2 pixel_4862/AMP_IN pixel_4862/SF_IB
+ pixel_4862/PIX_OUT pixel_4862/CSA_VREF pixel
Xpixel_4873 pixel_4873/gring pixel_4873/VDD pixel_4873/GND pixel_4873/VREF pixel_4873/ROW_SEL
+ pixel_4873/NB1 pixel_4873/VBIAS pixel_4873/NB2 pixel_4873/AMP_IN pixel_4873/SF_IB
+ pixel_4873/PIX_OUT pixel_4873/CSA_VREF pixel
Xpixel_890 pixel_890/gring pixel_890/VDD pixel_890/GND pixel_890/VREF pixel_890/ROW_SEL
+ pixel_890/NB1 pixel_890/VBIAS pixel_890/NB2 pixel_890/AMP_IN pixel_890/SF_IB pixel_890/PIX_OUT
+ pixel_890/CSA_VREF pixel
Xpixel_4884 pixel_4884/gring pixel_4884/VDD pixel_4884/GND pixel_4884/VREF pixel_4884/ROW_SEL
+ pixel_4884/NB1 pixel_4884/VBIAS pixel_4884/NB2 pixel_4884/AMP_IN pixel_4884/SF_IB
+ pixel_4884/PIX_OUT pixel_4884/CSA_VREF pixel
Xpixel_4895 pixel_4895/gring pixel_4895/VDD pixel_4895/GND pixel_4895/VREF pixel_4895/ROW_SEL
+ pixel_4895/NB1 pixel_4895/VBIAS pixel_4895/NB2 pixel_4895/AMP_IN pixel_4895/SF_IB
+ pixel_4895/PIX_OUT pixel_4895/CSA_VREF pixel
Xpixel_9829 pixel_9829/gring pixel_9829/VDD pixel_9829/GND pixel_9829/VREF pixel_9829/ROW_SEL
+ pixel_9829/NB1 pixel_9829/VBIAS pixel_9829/NB2 pixel_9829/AMP_IN pixel_9829/SF_IB
+ pixel_9829/PIX_OUT pixel_9829/CSA_VREF pixel
Xpixel_9818 pixel_9818/gring pixel_9818/VDD pixel_9818/GND pixel_9818/VREF pixel_9818/ROW_SEL
+ pixel_9818/NB1 pixel_9818/VBIAS pixel_9818/NB2 pixel_9818/AMP_IN pixel_9818/SF_IB
+ pixel_9818/PIX_OUT pixel_9818/CSA_VREF pixel
Xpixel_9807 pixel_9807/gring pixel_9807/VDD pixel_9807/GND pixel_9807/VREF pixel_9807/ROW_SEL
+ pixel_9807/NB1 pixel_9807/VBIAS pixel_9807/NB2 pixel_9807/AMP_IN pixel_9807/SF_IB
+ pixel_9807/PIX_OUT pixel_9807/CSA_VREF pixel
Xpixel_131 pixel_131/gring pixel_131/VDD pixel_131/GND pixel_131/VREF pixel_131/ROW_SEL
+ pixel_131/NB1 pixel_131/VBIAS pixel_131/NB2 pixel_131/AMP_IN pixel_131/SF_IB pixel_131/PIX_OUT
+ pixel_131/CSA_VREF pixel
Xpixel_120 pixel_120/gring pixel_120/VDD pixel_120/GND pixel_120/VREF pixel_120/ROW_SEL
+ pixel_120/NB1 pixel_120/VBIAS pixel_120/NB2 pixel_120/AMP_IN pixel_120/SF_IB pixel_120/PIX_OUT
+ pixel_120/CSA_VREF pixel
Xpixel_4103 pixel_4103/gring pixel_4103/VDD pixel_4103/GND pixel_4103/VREF pixel_4103/ROW_SEL
+ pixel_4103/NB1 pixel_4103/VBIAS pixel_4103/NB2 pixel_4103/AMP_IN pixel_4103/SF_IB
+ pixel_4103/PIX_OUT pixel_4103/CSA_VREF pixel
Xpixel_4114 pixel_4114/gring pixel_4114/VDD pixel_4114/GND pixel_4114/VREF pixel_4114/ROW_SEL
+ pixel_4114/NB1 pixel_4114/VBIAS pixel_4114/NB2 pixel_4114/AMP_IN pixel_4114/SF_IB
+ pixel_4114/PIX_OUT pixel_4114/CSA_VREF pixel
Xpixel_4125 pixel_4125/gring pixel_4125/VDD pixel_4125/GND pixel_4125/VREF pixel_4125/ROW_SEL
+ pixel_4125/NB1 pixel_4125/VBIAS pixel_4125/NB2 pixel_4125/AMP_IN pixel_4125/SF_IB
+ pixel_4125/PIX_OUT pixel_4125/CSA_VREF pixel
Xpixel_164 pixel_164/gring pixel_164/VDD pixel_164/GND pixel_164/VREF pixel_164/ROW_SEL
+ pixel_164/NB1 pixel_164/VBIAS pixel_164/NB2 pixel_164/AMP_IN pixel_164/SF_IB pixel_164/PIX_OUT
+ pixel_164/CSA_VREF pixel
Xpixel_153 pixel_153/gring pixel_153/VDD pixel_153/GND pixel_153/VREF pixel_153/ROW_SEL
+ pixel_153/NB1 pixel_153/VBIAS pixel_153/NB2 pixel_153/AMP_IN pixel_153/SF_IB pixel_153/PIX_OUT
+ pixel_153/CSA_VREF pixel
Xpixel_142 pixel_142/gring pixel_142/VDD pixel_142/GND pixel_142/VREF pixel_142/ROW_SEL
+ pixel_142/NB1 pixel_142/VBIAS pixel_142/NB2 pixel_142/AMP_IN pixel_142/SF_IB pixel_142/PIX_OUT
+ pixel_142/CSA_VREF pixel
Xpixel_3424 pixel_3424/gring pixel_3424/VDD pixel_3424/GND pixel_3424/VREF pixel_3424/ROW_SEL
+ pixel_3424/NB1 pixel_3424/VBIAS pixel_3424/NB2 pixel_3424/AMP_IN pixel_3424/SF_IB
+ pixel_3424/PIX_OUT pixel_3424/CSA_VREF pixel
Xpixel_3413 pixel_3413/gring pixel_3413/VDD pixel_3413/GND pixel_3413/VREF pixel_3413/ROW_SEL
+ pixel_3413/NB1 pixel_3413/VBIAS pixel_3413/NB2 pixel_3413/AMP_IN pixel_3413/SF_IB
+ pixel_3413/PIX_OUT pixel_3413/CSA_VREF pixel
Xpixel_3402 pixel_3402/gring pixel_3402/VDD pixel_3402/GND pixel_3402/VREF pixel_3402/ROW_SEL
+ pixel_3402/NB1 pixel_3402/VBIAS pixel_3402/NB2 pixel_3402/AMP_IN pixel_3402/SF_IB
+ pixel_3402/PIX_OUT pixel_3402/CSA_VREF pixel
Xpixel_4136 pixel_4136/gring pixel_4136/VDD pixel_4136/GND pixel_4136/VREF pixel_4136/ROW_SEL
+ pixel_4136/NB1 pixel_4136/VBIAS pixel_4136/NB2 pixel_4136/AMP_IN pixel_4136/SF_IB
+ pixel_4136/PIX_OUT pixel_4136/CSA_VREF pixel
Xpixel_4147 pixel_4147/gring pixel_4147/VDD pixel_4147/GND pixel_4147/VREF pixel_4147/ROW_SEL
+ pixel_4147/NB1 pixel_4147/VBIAS pixel_4147/NB2 pixel_4147/AMP_IN pixel_4147/SF_IB
+ pixel_4147/PIX_OUT pixel_4147/CSA_VREF pixel
Xpixel_4158 pixel_4158/gring pixel_4158/VDD pixel_4158/GND pixel_4158/VREF pixel_4158/ROW_SEL
+ pixel_4158/NB1 pixel_4158/VBIAS pixel_4158/NB2 pixel_4158/AMP_IN pixel_4158/SF_IB
+ pixel_4158/PIX_OUT pixel_4158/CSA_VREF pixel
Xpixel_4169 pixel_4169/gring pixel_4169/VDD pixel_4169/GND pixel_4169/VREF pixel_4169/ROW_SEL
+ pixel_4169/NB1 pixel_4169/VBIAS pixel_4169/NB2 pixel_4169/AMP_IN pixel_4169/SF_IB
+ pixel_4169/PIX_OUT pixel_4169/CSA_VREF pixel
Xpixel_197 pixel_197/gring pixel_197/VDD pixel_197/GND pixel_197/VREF pixel_197/ROW_SEL
+ pixel_197/NB1 pixel_197/VBIAS pixel_197/NB2 pixel_197/AMP_IN pixel_197/SF_IB pixel_197/PIX_OUT
+ pixel_197/CSA_VREF pixel
Xpixel_186 pixel_186/gring pixel_186/VDD pixel_186/GND pixel_186/VREF pixel_186/ROW_SEL
+ pixel_186/NB1 pixel_186/VBIAS pixel_186/NB2 pixel_186/AMP_IN pixel_186/SF_IB pixel_186/PIX_OUT
+ pixel_186/CSA_VREF pixel
Xpixel_175 pixel_175/gring pixel_175/VDD pixel_175/GND pixel_175/VREF pixel_175/ROW_SEL
+ pixel_175/NB1 pixel_175/VBIAS pixel_175/NB2 pixel_175/AMP_IN pixel_175/SF_IB pixel_175/PIX_OUT
+ pixel_175/CSA_VREF pixel
Xpixel_2712 pixel_2712/gring pixel_2712/VDD pixel_2712/GND pixel_2712/VREF pixel_2712/ROW_SEL
+ pixel_2712/NB1 pixel_2712/VBIAS pixel_2712/NB2 pixel_2712/AMP_IN pixel_2712/SF_IB
+ pixel_2712/PIX_OUT pixel_2712/CSA_VREF pixel
Xpixel_2701 pixel_2701/gring pixel_2701/VDD pixel_2701/GND pixel_2701/VREF pixel_2701/ROW_SEL
+ pixel_2701/NB1 pixel_2701/VBIAS pixel_2701/NB2 pixel_2701/AMP_IN pixel_2701/SF_IB
+ pixel_2701/PIX_OUT pixel_2701/CSA_VREF pixel
Xpixel_3457 pixel_3457/gring pixel_3457/VDD pixel_3457/GND pixel_3457/VREF pixel_3457/ROW_SEL
+ pixel_3457/NB1 pixel_3457/VBIAS pixel_3457/NB2 pixel_3457/AMP_IN pixel_3457/SF_IB
+ pixel_3457/PIX_OUT pixel_3457/CSA_VREF pixel
Xpixel_3446 pixel_3446/gring pixel_3446/VDD pixel_3446/GND pixel_3446/VREF pixel_3446/ROW_SEL
+ pixel_3446/NB1 pixel_3446/VBIAS pixel_3446/NB2 pixel_3446/AMP_IN pixel_3446/SF_IB
+ pixel_3446/PIX_OUT pixel_3446/CSA_VREF pixel
Xpixel_3435 pixel_3435/gring pixel_3435/VDD pixel_3435/GND pixel_3435/VREF pixel_3435/ROW_SEL
+ pixel_3435/NB1 pixel_3435/VBIAS pixel_3435/NB2 pixel_3435/AMP_IN pixel_3435/SF_IB
+ pixel_3435/PIX_OUT pixel_3435/CSA_VREF pixel
Xpixel_2756 pixel_2756/gring pixel_2756/VDD pixel_2756/GND pixel_2756/VREF pixel_2756/ROW_SEL
+ pixel_2756/NB1 pixel_2756/VBIAS pixel_2756/NB2 pixel_2756/AMP_IN pixel_2756/SF_IB
+ pixel_2756/PIX_OUT pixel_2756/CSA_VREF pixel
Xpixel_2745 pixel_2745/gring pixel_2745/VDD pixel_2745/GND pixel_2745/VREF pixel_2745/ROW_SEL
+ pixel_2745/NB1 pixel_2745/VBIAS pixel_2745/NB2 pixel_2745/AMP_IN pixel_2745/SF_IB
+ pixel_2745/PIX_OUT pixel_2745/CSA_VREF pixel
Xpixel_2734 pixel_2734/gring pixel_2734/VDD pixel_2734/GND pixel_2734/VREF pixel_2734/ROW_SEL
+ pixel_2734/NB1 pixel_2734/VBIAS pixel_2734/NB2 pixel_2734/AMP_IN pixel_2734/SF_IB
+ pixel_2734/PIX_OUT pixel_2734/CSA_VREF pixel
Xpixel_2723 pixel_2723/gring pixel_2723/VDD pixel_2723/GND pixel_2723/VREF pixel_2723/ROW_SEL
+ pixel_2723/NB1 pixel_2723/VBIAS pixel_2723/NB2 pixel_2723/AMP_IN pixel_2723/SF_IB
+ pixel_2723/PIX_OUT pixel_2723/CSA_VREF pixel
Xpixel_3479 pixel_3479/gring pixel_3479/VDD pixel_3479/GND pixel_3479/VREF pixel_3479/ROW_SEL
+ pixel_3479/NB1 pixel_3479/VBIAS pixel_3479/NB2 pixel_3479/AMP_IN pixel_3479/SF_IB
+ pixel_3479/PIX_OUT pixel_3479/CSA_VREF pixel
Xpixel_3468 pixel_3468/gring pixel_3468/VDD pixel_3468/GND pixel_3468/VREF pixel_3468/ROW_SEL
+ pixel_3468/NB1 pixel_3468/VBIAS pixel_3468/NB2 pixel_3468/AMP_IN pixel_3468/SF_IB
+ pixel_3468/PIX_OUT pixel_3468/CSA_VREF pixel
Xpixel_2789 pixel_2789/gring pixel_2789/VDD pixel_2789/GND pixel_2789/VREF pixel_2789/ROW_SEL
+ pixel_2789/NB1 pixel_2789/VBIAS pixel_2789/NB2 pixel_2789/AMP_IN pixel_2789/SF_IB
+ pixel_2789/PIX_OUT pixel_2789/CSA_VREF pixel
Xpixel_2778 pixel_2778/gring pixel_2778/VDD pixel_2778/GND pixel_2778/VREF pixel_2778/ROW_SEL
+ pixel_2778/NB1 pixel_2778/VBIAS pixel_2778/NB2 pixel_2778/AMP_IN pixel_2778/SF_IB
+ pixel_2778/PIX_OUT pixel_2778/CSA_VREF pixel
Xpixel_2767 pixel_2767/gring pixel_2767/VDD pixel_2767/GND pixel_2767/VREF pixel_2767/ROW_SEL
+ pixel_2767/NB1 pixel_2767/VBIAS pixel_2767/NB2 pixel_2767/AMP_IN pixel_2767/SF_IB
+ pixel_2767/PIX_OUT pixel_2767/CSA_VREF pixel
Xpixel_6050 pixel_6050/gring pixel_6050/VDD pixel_6050/GND pixel_6050/VREF pixel_6050/ROW_SEL
+ pixel_6050/NB1 pixel_6050/VBIAS pixel_6050/NB2 pixel_6050/AMP_IN pixel_6050/SF_IB
+ pixel_6050/PIX_OUT pixel_6050/CSA_VREF pixel
Xpixel_6061 pixel_6061/gring pixel_6061/VDD pixel_6061/GND pixel_6061/VREF pixel_6061/ROW_SEL
+ pixel_6061/NB1 pixel_6061/VBIAS pixel_6061/NB2 pixel_6061/AMP_IN pixel_6061/SF_IB
+ pixel_6061/PIX_OUT pixel_6061/CSA_VREF pixel
Xpixel_6072 pixel_6072/gring pixel_6072/VDD pixel_6072/GND pixel_6072/VREF pixel_6072/ROW_SEL
+ pixel_6072/NB1 pixel_6072/VBIAS pixel_6072/NB2 pixel_6072/AMP_IN pixel_6072/SF_IB
+ pixel_6072/PIX_OUT pixel_6072/CSA_VREF pixel
Xpixel_6083 pixel_6083/gring pixel_6083/VDD pixel_6083/GND pixel_6083/VREF pixel_6083/ROW_SEL
+ pixel_6083/NB1 pixel_6083/VBIAS pixel_6083/NB2 pixel_6083/AMP_IN pixel_6083/SF_IB
+ pixel_6083/PIX_OUT pixel_6083/CSA_VREF pixel
Xpixel_6094 pixel_6094/gring pixel_6094/VDD pixel_6094/GND pixel_6094/VREF pixel_6094/ROW_SEL
+ pixel_6094/NB1 pixel_6094/VBIAS pixel_6094/NB2 pixel_6094/AMP_IN pixel_6094/SF_IB
+ pixel_6094/PIX_OUT pixel_6094/CSA_VREF pixel
Xpixel_5360 pixel_5360/gring pixel_5360/VDD pixel_5360/GND pixel_5360/VREF pixel_5360/ROW_SEL
+ pixel_5360/NB1 pixel_5360/VBIAS pixel_5360/NB2 pixel_5360/AMP_IN pixel_5360/SF_IB
+ pixel_5360/PIX_OUT pixel_5360/CSA_VREF pixel
Xpixel_5371 pixel_5371/gring pixel_5371/VDD pixel_5371/GND pixel_5371/VREF pixel_5371/ROW_SEL
+ pixel_5371/NB1 pixel_5371/VBIAS pixel_5371/NB2 pixel_5371/AMP_IN pixel_5371/SF_IB
+ pixel_5371/PIX_OUT pixel_5371/CSA_VREF pixel
Xpixel_5382 pixel_5382/gring pixel_5382/VDD pixel_5382/GND pixel_5382/VREF pixel_5382/ROW_SEL
+ pixel_5382/NB1 pixel_5382/VBIAS pixel_5382/NB2 pixel_5382/AMP_IN pixel_5382/SF_IB
+ pixel_5382/PIX_OUT pixel_5382/CSA_VREF pixel
Xpixel_5393 pixel_5393/gring pixel_5393/VDD pixel_5393/GND pixel_5393/VREF pixel_5393/ROW_SEL
+ pixel_5393/NB1 pixel_5393/VBIAS pixel_5393/NB2 pixel_5393/AMP_IN pixel_5393/SF_IB
+ pixel_5393/PIX_OUT pixel_5393/CSA_VREF pixel
Xpixel_4670 pixel_4670/gring pixel_4670/VDD pixel_4670/GND pixel_4670/VREF pixel_4670/ROW_SEL
+ pixel_4670/NB1 pixel_4670/VBIAS pixel_4670/NB2 pixel_4670/AMP_IN pixel_4670/SF_IB
+ pixel_4670/PIX_OUT pixel_4670/CSA_VREF pixel
Xpixel_4681 pixel_4681/gring pixel_4681/VDD pixel_4681/GND pixel_4681/VREF pixel_4681/ROW_SEL
+ pixel_4681/NB1 pixel_4681/VBIAS pixel_4681/NB2 pixel_4681/AMP_IN pixel_4681/SF_IB
+ pixel_4681/PIX_OUT pixel_4681/CSA_VREF pixel
Xpixel_4692 pixel_4692/gring pixel_4692/VDD pixel_4692/GND pixel_4692/VREF pixel_4692/ROW_SEL
+ pixel_4692/NB1 pixel_4692/VBIAS pixel_4692/NB2 pixel_4692/AMP_IN pixel_4692/SF_IB
+ pixel_4692/PIX_OUT pixel_4692/CSA_VREF pixel
Xpixel_3980 pixel_3980/gring pixel_3980/VDD pixel_3980/GND pixel_3980/VREF pixel_3980/ROW_SEL
+ pixel_3980/NB1 pixel_3980/VBIAS pixel_3980/NB2 pixel_3980/AMP_IN pixel_3980/SF_IB
+ pixel_3980/PIX_OUT pixel_3980/CSA_VREF pixel
Xpixel_3991 pixel_3991/gring pixel_3991/VDD pixel_3991/GND pixel_3991/VREF pixel_3991/ROW_SEL
+ pixel_3991/NB1 pixel_3991/VBIAS pixel_3991/NB2 pixel_3991/AMP_IN pixel_3991/SF_IB
+ pixel_3991/PIX_OUT pixel_3991/CSA_VREF pixel
Xpixel_1 pixel_1/gring pixel_1/VDD pixel_1/GND pixel_1/VREF pixel_1/ROW_SEL pixel_1/NB1
+ pixel_1/VBIAS pixel_1/NB2 pixel_1/AMP_IN pixel_1/SF_IB pixel_1/PIX_OUT pixel_1/CSA_VREF
+ pixel
Xpixel_2008 pixel_2008/gring pixel_2008/VDD pixel_2008/GND pixel_2008/VREF pixel_2008/ROW_SEL
+ pixel_2008/NB1 pixel_2008/VBIAS pixel_2008/NB2 pixel_2008/AMP_IN pixel_2008/SF_IB
+ pixel_2008/PIX_OUT pixel_2008/CSA_VREF pixel
Xpixel_2019 pixel_2019/gring pixel_2019/VDD pixel_2019/GND pixel_2019/VREF pixel_2019/ROW_SEL
+ pixel_2019/NB1 pixel_2019/VBIAS pixel_2019/NB2 pixel_2019/AMP_IN pixel_2019/SF_IB
+ pixel_2019/PIX_OUT pixel_2019/CSA_VREF pixel
Xpixel_1329 pixel_1329/gring pixel_1329/VDD pixel_1329/GND pixel_1329/VREF pixel_1329/ROW_SEL
+ pixel_1329/NB1 pixel_1329/VBIAS pixel_1329/NB2 pixel_1329/AMP_IN pixel_1329/SF_IB
+ pixel_1329/PIX_OUT pixel_1329/CSA_VREF pixel
Xpixel_1318 pixel_1318/gring pixel_1318/VDD pixel_1318/GND pixel_1318/VREF pixel_1318/ROW_SEL
+ pixel_1318/NB1 pixel_1318/VBIAS pixel_1318/NB2 pixel_1318/AMP_IN pixel_1318/SF_IB
+ pixel_1318/PIX_OUT pixel_1318/CSA_VREF pixel
Xpixel_1307 pixel_1307/gring pixel_1307/VDD pixel_1307/GND pixel_1307/VREF pixel_1307/ROW_SEL
+ pixel_1307/NB1 pixel_1307/VBIAS pixel_1307/NB2 pixel_1307/AMP_IN pixel_1307/SF_IB
+ pixel_1307/PIX_OUT pixel_1307/CSA_VREF pixel
Xpixel_9604 pixel_9604/gring pixel_9604/VDD pixel_9604/GND pixel_9604/VREF pixel_9604/ROW_SEL
+ pixel_9604/NB1 pixel_9604/VBIAS pixel_9604/NB2 pixel_9604/AMP_IN pixel_9604/SF_IB
+ pixel_9604/PIX_OUT pixel_9604/CSA_VREF pixel
Xpixel_8903 pixel_8903/gring pixel_8903/VDD pixel_8903/GND pixel_8903/VREF pixel_8903/ROW_SEL
+ pixel_8903/NB1 pixel_8903/VBIAS pixel_8903/NB2 pixel_8903/AMP_IN pixel_8903/SF_IB
+ pixel_8903/PIX_OUT pixel_8903/CSA_VREF pixel
Xpixel_9615 pixel_9615/gring pixel_9615/VDD pixel_9615/GND pixel_9615/VREF pixel_9615/ROW_SEL
+ pixel_9615/NB1 pixel_9615/VBIAS pixel_9615/NB2 pixel_9615/AMP_IN pixel_9615/SF_IB
+ pixel_9615/PIX_OUT pixel_9615/CSA_VREF pixel
Xpixel_9626 pixel_9626/gring pixel_9626/VDD pixel_9626/GND pixel_9626/VREF pixel_9626/ROW_SEL
+ pixel_9626/NB1 pixel_9626/VBIAS pixel_9626/NB2 pixel_9626/AMP_IN pixel_9626/SF_IB
+ pixel_9626/PIX_OUT pixel_9626/CSA_VREF pixel
Xpixel_9637 pixel_9637/gring pixel_9637/VDD pixel_9637/GND pixel_9637/VREF pixel_9637/ROW_SEL
+ pixel_9637/NB1 pixel_9637/VBIAS pixel_9637/NB2 pixel_9637/AMP_IN pixel_9637/SF_IB
+ pixel_9637/PIX_OUT pixel_9637/CSA_VREF pixel
Xpixel_9648 pixel_9648/gring pixel_9648/VDD pixel_9648/GND pixel_9648/VREF pixel_9648/ROW_SEL
+ pixel_9648/NB1 pixel_9648/VBIAS pixel_9648/NB2 pixel_9648/AMP_IN pixel_9648/SF_IB
+ pixel_9648/PIX_OUT pixel_9648/CSA_VREF pixel
Xpixel_8936 pixel_8936/gring pixel_8936/VDD pixel_8936/GND pixel_8936/VREF pixel_8936/ROW_SEL
+ pixel_8936/NB1 pixel_8936/VBIAS pixel_8936/NB2 pixel_8936/AMP_IN pixel_8936/SF_IB
+ pixel_8936/PIX_OUT pixel_8936/CSA_VREF pixel
Xpixel_8925 pixel_8925/gring pixel_8925/VDD pixel_8925/GND pixel_8925/VREF pixel_8925/ROW_SEL
+ pixel_8925/NB1 pixel_8925/VBIAS pixel_8925/NB2 pixel_8925/AMP_IN pixel_8925/SF_IB
+ pixel_8925/PIX_OUT pixel_8925/CSA_VREF pixel
Xpixel_8914 pixel_8914/gring pixel_8914/VDD pixel_8914/GND pixel_8914/VREF pixel_8914/ROW_SEL
+ pixel_8914/NB1 pixel_8914/VBIAS pixel_8914/NB2 pixel_8914/AMP_IN pixel_8914/SF_IB
+ pixel_8914/PIX_OUT pixel_8914/CSA_VREF pixel
Xpixel_9659 pixel_9659/gring pixel_9659/VDD pixel_9659/GND pixel_9659/VREF pixel_9659/ROW_SEL
+ pixel_9659/NB1 pixel_9659/VBIAS pixel_9659/NB2 pixel_9659/AMP_IN pixel_9659/SF_IB
+ pixel_9659/PIX_OUT pixel_9659/CSA_VREF pixel
Xpixel_8969 pixel_8969/gring pixel_8969/VDD pixel_8969/GND pixel_8969/VREF pixel_8969/ROW_SEL
+ pixel_8969/NB1 pixel_8969/VBIAS pixel_8969/NB2 pixel_8969/AMP_IN pixel_8969/SF_IB
+ pixel_8969/PIX_OUT pixel_8969/CSA_VREF pixel
Xpixel_8958 pixel_8958/gring pixel_8958/VDD pixel_8958/GND pixel_8958/VREF pixel_8958/ROW_SEL
+ pixel_8958/NB1 pixel_8958/VBIAS pixel_8958/NB2 pixel_8958/AMP_IN pixel_8958/SF_IB
+ pixel_8958/PIX_OUT pixel_8958/CSA_VREF pixel
Xpixel_8947 pixel_8947/gring pixel_8947/VDD pixel_8947/GND pixel_8947/VREF pixel_8947/ROW_SEL
+ pixel_8947/NB1 pixel_8947/VBIAS pixel_8947/NB2 pixel_8947/AMP_IN pixel_8947/SF_IB
+ pixel_8947/PIX_OUT pixel_8947/CSA_VREF pixel
Xpixel_3232 pixel_3232/gring pixel_3232/VDD pixel_3232/GND pixel_3232/VREF pixel_3232/ROW_SEL
+ pixel_3232/NB1 pixel_3232/VBIAS pixel_3232/NB2 pixel_3232/AMP_IN pixel_3232/SF_IB
+ pixel_3232/PIX_OUT pixel_3232/CSA_VREF pixel
Xpixel_3221 pixel_3221/gring pixel_3221/VDD pixel_3221/GND pixel_3221/VREF pixel_3221/ROW_SEL
+ pixel_3221/NB1 pixel_3221/VBIAS pixel_3221/NB2 pixel_3221/AMP_IN pixel_3221/SF_IB
+ pixel_3221/PIX_OUT pixel_3221/CSA_VREF pixel
Xpixel_3210 pixel_3210/gring pixel_3210/VDD pixel_3210/GND pixel_3210/VREF pixel_3210/ROW_SEL
+ pixel_3210/NB1 pixel_3210/VBIAS pixel_3210/NB2 pixel_3210/AMP_IN pixel_3210/SF_IB
+ pixel_3210/PIX_OUT pixel_3210/CSA_VREF pixel
Xpixel_2531 pixel_2531/gring pixel_2531/VDD pixel_2531/GND pixel_2531/VREF pixel_2531/ROW_SEL
+ pixel_2531/NB1 pixel_2531/VBIAS pixel_2531/NB2 pixel_2531/AMP_IN pixel_2531/SF_IB
+ pixel_2531/PIX_OUT pixel_2531/CSA_VREF pixel
Xpixel_2520 pixel_2520/gring pixel_2520/VDD pixel_2520/GND pixel_2520/VREF pixel_2520/ROW_SEL
+ pixel_2520/NB1 pixel_2520/VBIAS pixel_2520/NB2 pixel_2520/AMP_IN pixel_2520/SF_IB
+ pixel_2520/PIX_OUT pixel_2520/CSA_VREF pixel
Xpixel_3265 pixel_3265/gring pixel_3265/VDD pixel_3265/GND pixel_3265/VREF pixel_3265/ROW_SEL
+ pixel_3265/NB1 pixel_3265/VBIAS pixel_3265/NB2 pixel_3265/AMP_IN pixel_3265/SF_IB
+ pixel_3265/PIX_OUT pixel_3265/CSA_VREF pixel
Xpixel_3254 pixel_3254/gring pixel_3254/VDD pixel_3254/GND pixel_3254/VREF pixel_3254/ROW_SEL
+ pixel_3254/NB1 pixel_3254/VBIAS pixel_3254/NB2 pixel_3254/AMP_IN pixel_3254/SF_IB
+ pixel_3254/PIX_OUT pixel_3254/CSA_VREF pixel
Xpixel_3243 pixel_3243/gring pixel_3243/VDD pixel_3243/GND pixel_3243/VREF pixel_3243/ROW_SEL
+ pixel_3243/NB1 pixel_3243/VBIAS pixel_3243/NB2 pixel_3243/AMP_IN pixel_3243/SF_IB
+ pixel_3243/PIX_OUT pixel_3243/CSA_VREF pixel
Xpixel_2564 pixel_2564/gring pixel_2564/VDD pixel_2564/GND pixel_2564/VREF pixel_2564/ROW_SEL
+ pixel_2564/NB1 pixel_2564/VBIAS pixel_2564/NB2 pixel_2564/AMP_IN pixel_2564/SF_IB
+ pixel_2564/PIX_OUT pixel_2564/CSA_VREF pixel
Xpixel_2553 pixel_2553/gring pixel_2553/VDD pixel_2553/GND pixel_2553/VREF pixel_2553/ROW_SEL
+ pixel_2553/NB1 pixel_2553/VBIAS pixel_2553/NB2 pixel_2553/AMP_IN pixel_2553/SF_IB
+ pixel_2553/PIX_OUT pixel_2553/CSA_VREF pixel
Xpixel_2542 pixel_2542/gring pixel_2542/VDD pixel_2542/GND pixel_2542/VREF pixel_2542/ROW_SEL
+ pixel_2542/NB1 pixel_2542/VBIAS pixel_2542/NB2 pixel_2542/AMP_IN pixel_2542/SF_IB
+ pixel_2542/PIX_OUT pixel_2542/CSA_VREF pixel
Xpixel_3298 pixel_3298/gring pixel_3298/VDD pixel_3298/GND pixel_3298/VREF pixel_3298/ROW_SEL
+ pixel_3298/NB1 pixel_3298/VBIAS pixel_3298/NB2 pixel_3298/AMP_IN pixel_3298/SF_IB
+ pixel_3298/PIX_OUT pixel_3298/CSA_VREF pixel
Xpixel_3287 pixel_3287/gring pixel_3287/VDD pixel_3287/GND pixel_3287/VREF pixel_3287/ROW_SEL
+ pixel_3287/NB1 pixel_3287/VBIAS pixel_3287/NB2 pixel_3287/AMP_IN pixel_3287/SF_IB
+ pixel_3287/PIX_OUT pixel_3287/CSA_VREF pixel
Xpixel_3276 pixel_3276/gring pixel_3276/VDD pixel_3276/GND pixel_3276/VREF pixel_3276/ROW_SEL
+ pixel_3276/NB1 pixel_3276/VBIAS pixel_3276/NB2 pixel_3276/AMP_IN pixel_3276/SF_IB
+ pixel_3276/PIX_OUT pixel_3276/CSA_VREF pixel
Xpixel_1852 pixel_1852/gring pixel_1852/VDD pixel_1852/GND pixel_1852/VREF pixel_1852/ROW_SEL
+ pixel_1852/NB1 pixel_1852/VBIAS pixel_1852/NB2 pixel_1852/AMP_IN pixel_1852/SF_IB
+ pixel_1852/PIX_OUT pixel_1852/CSA_VREF pixel
Xpixel_1841 pixel_1841/gring pixel_1841/VDD pixel_1841/GND pixel_1841/VREF pixel_1841/ROW_SEL
+ pixel_1841/NB1 pixel_1841/VBIAS pixel_1841/NB2 pixel_1841/AMP_IN pixel_1841/SF_IB
+ pixel_1841/PIX_OUT pixel_1841/CSA_VREF pixel
Xpixel_1830 pixel_1830/gring pixel_1830/VDD pixel_1830/GND pixel_1830/VREF pixel_1830/ROW_SEL
+ pixel_1830/NB1 pixel_1830/VBIAS pixel_1830/NB2 pixel_1830/AMP_IN pixel_1830/SF_IB
+ pixel_1830/PIX_OUT pixel_1830/CSA_VREF pixel
Xpixel_2597 pixel_2597/gring pixel_2597/VDD pixel_2597/GND pixel_2597/VREF pixel_2597/ROW_SEL
+ pixel_2597/NB1 pixel_2597/VBIAS pixel_2597/NB2 pixel_2597/AMP_IN pixel_2597/SF_IB
+ pixel_2597/PIX_OUT pixel_2597/CSA_VREF pixel
Xpixel_2586 pixel_2586/gring pixel_2586/VDD pixel_2586/GND pixel_2586/VREF pixel_2586/ROW_SEL
+ pixel_2586/NB1 pixel_2586/VBIAS pixel_2586/NB2 pixel_2586/AMP_IN pixel_2586/SF_IB
+ pixel_2586/PIX_OUT pixel_2586/CSA_VREF pixel
Xpixel_2575 pixel_2575/gring pixel_2575/VDD pixel_2575/GND pixel_2575/VREF pixel_2575/ROW_SEL
+ pixel_2575/NB1 pixel_2575/VBIAS pixel_2575/NB2 pixel_2575/AMP_IN pixel_2575/SF_IB
+ pixel_2575/PIX_OUT pixel_2575/CSA_VREF pixel
Xpixel_1896 pixel_1896/gring pixel_1896/VDD pixel_1896/GND pixel_1896/VREF pixel_1896/ROW_SEL
+ pixel_1896/NB1 pixel_1896/VBIAS pixel_1896/NB2 pixel_1896/AMP_IN pixel_1896/SF_IB
+ pixel_1896/PIX_OUT pixel_1896/CSA_VREF pixel
Xpixel_1885 pixel_1885/gring pixel_1885/VDD pixel_1885/GND pixel_1885/VREF pixel_1885/ROW_SEL
+ pixel_1885/NB1 pixel_1885/VBIAS pixel_1885/NB2 pixel_1885/AMP_IN pixel_1885/SF_IB
+ pixel_1885/PIX_OUT pixel_1885/CSA_VREF pixel
Xpixel_1874 pixel_1874/gring pixel_1874/VDD pixel_1874/GND pixel_1874/VREF pixel_1874/ROW_SEL
+ pixel_1874/NB1 pixel_1874/VBIAS pixel_1874/NB2 pixel_1874/AMP_IN pixel_1874/SF_IB
+ pixel_1874/PIX_OUT pixel_1874/CSA_VREF pixel
Xpixel_1863 pixel_1863/gring pixel_1863/VDD pixel_1863/GND pixel_1863/VREF pixel_1863/ROW_SEL
+ pixel_1863/NB1 pixel_1863/VBIAS pixel_1863/NB2 pixel_1863/AMP_IN pixel_1863/SF_IB
+ pixel_1863/PIX_OUT pixel_1863/CSA_VREF pixel
Xpixel_5190 pixel_5190/gring pixel_5190/VDD pixel_5190/GND pixel_5190/VREF pixel_5190/ROW_SEL
+ pixel_5190/NB1 pixel_5190/VBIAS pixel_5190/NB2 pixel_5190/AMP_IN pixel_5190/SF_IB
+ pixel_5190/PIX_OUT pixel_5190/CSA_VREF pixel
Xpixel_7509 pixel_7509/gring pixel_7509/VDD pixel_7509/GND pixel_7509/VREF pixel_7509/ROW_SEL
+ pixel_7509/NB1 pixel_7509/VBIAS pixel_7509/NB2 pixel_7509/AMP_IN pixel_7509/SF_IB
+ pixel_7509/PIX_OUT pixel_7509/CSA_VREF pixel
Xpixel_6808 pixel_6808/gring pixel_6808/VDD pixel_6808/GND pixel_6808/VREF pixel_6808/ROW_SEL
+ pixel_6808/NB1 pixel_6808/VBIAS pixel_6808/NB2 pixel_6808/AMP_IN pixel_6808/SF_IB
+ pixel_6808/PIX_OUT pixel_6808/CSA_VREF pixel
Xpixel_6819 pixel_6819/gring pixel_6819/VDD pixel_6819/GND pixel_6819/VREF pixel_6819/ROW_SEL
+ pixel_6819/NB1 pixel_6819/VBIAS pixel_6819/NB2 pixel_6819/AMP_IN pixel_6819/SF_IB
+ pixel_6819/PIX_OUT pixel_6819/CSA_VREF pixel
Xpixel_1115 pixel_1115/gring pixel_1115/VDD pixel_1115/GND pixel_1115/VREF pixel_1115/ROW_SEL
+ pixel_1115/NB1 pixel_1115/VBIAS pixel_1115/NB2 pixel_1115/AMP_IN pixel_1115/SF_IB
+ pixel_1115/PIX_OUT pixel_1115/CSA_VREF pixel
Xpixel_1104 pixel_1104/gring pixel_1104/VDD pixel_1104/GND pixel_1104/VREF pixel_1104/ROW_SEL
+ pixel_1104/NB1 pixel_1104/VBIAS pixel_1104/NB2 pixel_1104/AMP_IN pixel_1104/SF_IB
+ pixel_1104/PIX_OUT pixel_1104/CSA_VREF pixel
Xpixel_1148 pixel_1148/gring pixel_1148/VDD pixel_1148/GND pixel_1148/VREF pixel_1148/ROW_SEL
+ pixel_1148/NB1 pixel_1148/VBIAS pixel_1148/NB2 pixel_1148/AMP_IN pixel_1148/SF_IB
+ pixel_1148/PIX_OUT pixel_1148/CSA_VREF pixel
Xpixel_1137 pixel_1137/gring pixel_1137/VDD pixel_1137/GND pixel_1137/VREF pixel_1137/ROW_SEL
+ pixel_1137/NB1 pixel_1137/VBIAS pixel_1137/NB2 pixel_1137/AMP_IN pixel_1137/SF_IB
+ pixel_1137/PIX_OUT pixel_1137/CSA_VREF pixel
Xpixel_1126 pixel_1126/gring pixel_1126/VDD pixel_1126/GND pixel_1126/VREF pixel_1126/ROW_SEL
+ pixel_1126/NB1 pixel_1126/VBIAS pixel_1126/NB2 pixel_1126/AMP_IN pixel_1126/SF_IB
+ pixel_1126/PIX_OUT pixel_1126/CSA_VREF pixel
Xpixel_1159 pixel_1159/gring pixel_1159/VDD pixel_1159/GND pixel_1159/VREF pixel_1159/ROW_SEL
+ pixel_1159/NB1 pixel_1159/VBIAS pixel_1159/NB2 pixel_1159/AMP_IN pixel_1159/SF_IB
+ pixel_1159/PIX_OUT pixel_1159/CSA_VREF pixel
Xpixel_9423 pixel_9423/gring pixel_9423/VDD pixel_9423/GND pixel_9423/VREF pixel_9423/ROW_SEL
+ pixel_9423/NB1 pixel_9423/VBIAS pixel_9423/NB2 pixel_9423/AMP_IN pixel_9423/SF_IB
+ pixel_9423/PIX_OUT pixel_9423/CSA_VREF pixel
Xpixel_9412 pixel_9412/gring pixel_9412/VDD pixel_9412/GND pixel_9412/VREF pixel_9412/ROW_SEL
+ pixel_9412/NB1 pixel_9412/VBIAS pixel_9412/NB2 pixel_9412/AMP_IN pixel_9412/SF_IB
+ pixel_9412/PIX_OUT pixel_9412/CSA_VREF pixel
Xpixel_9401 pixel_9401/gring pixel_9401/VDD pixel_9401/GND pixel_9401/VREF pixel_9401/ROW_SEL
+ pixel_9401/NB1 pixel_9401/VBIAS pixel_9401/NB2 pixel_9401/AMP_IN pixel_9401/SF_IB
+ pixel_9401/PIX_OUT pixel_9401/CSA_VREF pixel
Xpixel_8711 pixel_8711/gring pixel_8711/VDD pixel_8711/GND pixel_8711/VREF pixel_8711/ROW_SEL
+ pixel_8711/NB1 pixel_8711/VBIAS pixel_8711/NB2 pixel_8711/AMP_IN pixel_8711/SF_IB
+ pixel_8711/PIX_OUT pixel_8711/CSA_VREF pixel
Xpixel_8700 pixel_8700/gring pixel_8700/VDD pixel_8700/GND pixel_8700/VREF pixel_8700/ROW_SEL
+ pixel_8700/NB1 pixel_8700/VBIAS pixel_8700/NB2 pixel_8700/AMP_IN pixel_8700/SF_IB
+ pixel_8700/PIX_OUT pixel_8700/CSA_VREF pixel
Xpixel_9456 pixel_9456/gring pixel_9456/VDD pixel_9456/GND pixel_9456/VREF pixel_9456/ROW_SEL
+ pixel_9456/NB1 pixel_9456/VBIAS pixel_9456/NB2 pixel_9456/AMP_IN pixel_9456/SF_IB
+ pixel_9456/PIX_OUT pixel_9456/CSA_VREF pixel
Xpixel_9445 pixel_9445/gring pixel_9445/VDD pixel_9445/GND pixel_9445/VREF pixel_9445/ROW_SEL
+ pixel_9445/NB1 pixel_9445/VBIAS pixel_9445/NB2 pixel_9445/AMP_IN pixel_9445/SF_IB
+ pixel_9445/PIX_OUT pixel_9445/CSA_VREF pixel
Xpixel_9434 pixel_9434/gring pixel_9434/VDD pixel_9434/GND pixel_9434/VREF pixel_9434/ROW_SEL
+ pixel_9434/NB1 pixel_9434/VBIAS pixel_9434/NB2 pixel_9434/AMP_IN pixel_9434/SF_IB
+ pixel_9434/PIX_OUT pixel_9434/CSA_VREF pixel
Xpixel_8744 pixel_8744/gring pixel_8744/VDD pixel_8744/GND pixel_8744/VREF pixel_8744/ROW_SEL
+ pixel_8744/NB1 pixel_8744/VBIAS pixel_8744/NB2 pixel_8744/AMP_IN pixel_8744/SF_IB
+ pixel_8744/PIX_OUT pixel_8744/CSA_VREF pixel
Xpixel_8733 pixel_8733/gring pixel_8733/VDD pixel_8733/GND pixel_8733/VREF pixel_8733/ROW_SEL
+ pixel_8733/NB1 pixel_8733/VBIAS pixel_8733/NB2 pixel_8733/AMP_IN pixel_8733/SF_IB
+ pixel_8733/PIX_OUT pixel_8733/CSA_VREF pixel
Xpixel_8722 pixel_8722/gring pixel_8722/VDD pixel_8722/GND pixel_8722/VREF pixel_8722/ROW_SEL
+ pixel_8722/NB1 pixel_8722/VBIAS pixel_8722/NB2 pixel_8722/AMP_IN pixel_8722/SF_IB
+ pixel_8722/PIX_OUT pixel_8722/CSA_VREF pixel
Xpixel_9489 pixel_9489/gring pixel_9489/VDD pixel_9489/GND pixel_9489/VREF pixel_9489/ROW_SEL
+ pixel_9489/NB1 pixel_9489/VBIAS pixel_9489/NB2 pixel_9489/AMP_IN pixel_9489/SF_IB
+ pixel_9489/PIX_OUT pixel_9489/CSA_VREF pixel
Xpixel_9478 pixel_9478/gring pixel_9478/VDD pixel_9478/GND pixel_9478/VREF pixel_9478/ROW_SEL
+ pixel_9478/NB1 pixel_9478/VBIAS pixel_9478/NB2 pixel_9478/AMP_IN pixel_9478/SF_IB
+ pixel_9478/PIX_OUT pixel_9478/CSA_VREF pixel
Xpixel_9467 pixel_9467/gring pixel_9467/VDD pixel_9467/GND pixel_9467/VREF pixel_9467/ROW_SEL
+ pixel_9467/NB1 pixel_9467/VBIAS pixel_9467/NB2 pixel_9467/AMP_IN pixel_9467/SF_IB
+ pixel_9467/PIX_OUT pixel_9467/CSA_VREF pixel
Xpixel_8788 pixel_8788/gring pixel_8788/VDD pixel_8788/GND pixel_8788/VREF pixel_8788/ROW_SEL
+ pixel_8788/NB1 pixel_8788/VBIAS pixel_8788/NB2 pixel_8788/AMP_IN pixel_8788/SF_IB
+ pixel_8788/PIX_OUT pixel_8788/CSA_VREF pixel
Xpixel_8777 pixel_8777/gring pixel_8777/VDD pixel_8777/GND pixel_8777/VREF pixel_8777/ROW_SEL
+ pixel_8777/NB1 pixel_8777/VBIAS pixel_8777/NB2 pixel_8777/AMP_IN pixel_8777/SF_IB
+ pixel_8777/PIX_OUT pixel_8777/CSA_VREF pixel
Xpixel_8766 pixel_8766/gring pixel_8766/VDD pixel_8766/GND pixel_8766/VREF pixel_8766/ROW_SEL
+ pixel_8766/NB1 pixel_8766/VBIAS pixel_8766/NB2 pixel_8766/AMP_IN pixel_8766/SF_IB
+ pixel_8766/PIX_OUT pixel_8766/CSA_VREF pixel
Xpixel_8755 pixel_8755/gring pixel_8755/VDD pixel_8755/GND pixel_8755/VREF pixel_8755/ROW_SEL
+ pixel_8755/NB1 pixel_8755/VBIAS pixel_8755/NB2 pixel_8755/AMP_IN pixel_8755/SF_IB
+ pixel_8755/PIX_OUT pixel_8755/CSA_VREF pixel
Xpixel_8799 pixel_8799/gring pixel_8799/VDD pixel_8799/GND pixel_8799/VREF pixel_8799/ROW_SEL
+ pixel_8799/NB1 pixel_8799/VBIAS pixel_8799/NB2 pixel_8799/AMP_IN pixel_8799/SF_IB
+ pixel_8799/PIX_OUT pixel_8799/CSA_VREF pixel
Xpixel_3040 pixel_3040/gring pixel_3040/VDD pixel_3040/GND pixel_3040/VREF pixel_3040/ROW_SEL
+ pixel_3040/NB1 pixel_3040/VBIAS pixel_3040/NB2 pixel_3040/AMP_IN pixel_3040/SF_IB
+ pixel_3040/PIX_OUT pixel_3040/CSA_VREF pixel
Xpixel_3084 pixel_3084/gring pixel_3084/VDD pixel_3084/GND pixel_3084/VREF pixel_3084/ROW_SEL
+ pixel_3084/NB1 pixel_3084/VBIAS pixel_3084/NB2 pixel_3084/AMP_IN pixel_3084/SF_IB
+ pixel_3084/PIX_OUT pixel_3084/CSA_VREF pixel
Xpixel_3073 pixel_3073/gring pixel_3073/VDD pixel_3073/GND pixel_3073/VREF pixel_3073/ROW_SEL
+ pixel_3073/NB1 pixel_3073/VBIAS pixel_3073/NB2 pixel_3073/AMP_IN pixel_3073/SF_IB
+ pixel_3073/PIX_OUT pixel_3073/CSA_VREF pixel
Xpixel_3062 pixel_3062/gring pixel_3062/VDD pixel_3062/GND pixel_3062/VREF pixel_3062/ROW_SEL
+ pixel_3062/NB1 pixel_3062/VBIAS pixel_3062/NB2 pixel_3062/AMP_IN pixel_3062/SF_IB
+ pixel_3062/PIX_OUT pixel_3062/CSA_VREF pixel
Xpixel_3051 pixel_3051/gring pixel_3051/VDD pixel_3051/GND pixel_3051/VREF pixel_3051/ROW_SEL
+ pixel_3051/NB1 pixel_3051/VBIAS pixel_3051/NB2 pixel_3051/AMP_IN pixel_3051/SF_IB
+ pixel_3051/PIX_OUT pixel_3051/CSA_VREF pixel
Xpixel_2372 pixel_2372/gring pixel_2372/VDD pixel_2372/GND pixel_2372/VREF pixel_2372/ROW_SEL
+ pixel_2372/NB1 pixel_2372/VBIAS pixel_2372/NB2 pixel_2372/AMP_IN pixel_2372/SF_IB
+ pixel_2372/PIX_OUT pixel_2372/CSA_VREF pixel
Xpixel_2361 pixel_2361/gring pixel_2361/VDD pixel_2361/GND pixel_2361/VREF pixel_2361/ROW_SEL
+ pixel_2361/NB1 pixel_2361/VBIAS pixel_2361/NB2 pixel_2361/AMP_IN pixel_2361/SF_IB
+ pixel_2361/PIX_OUT pixel_2361/CSA_VREF pixel
Xpixel_2350 pixel_2350/gring pixel_2350/VDD pixel_2350/GND pixel_2350/VREF pixel_2350/ROW_SEL
+ pixel_2350/NB1 pixel_2350/VBIAS pixel_2350/NB2 pixel_2350/AMP_IN pixel_2350/SF_IB
+ pixel_2350/PIX_OUT pixel_2350/CSA_VREF pixel
Xpixel_3095 pixel_3095/gring pixel_3095/VDD pixel_3095/GND pixel_3095/VREF pixel_3095/ROW_SEL
+ pixel_3095/NB1 pixel_3095/VBIAS pixel_3095/NB2 pixel_3095/AMP_IN pixel_3095/SF_IB
+ pixel_3095/PIX_OUT pixel_3095/CSA_VREF pixel
Xpixel_1660 pixel_1660/gring pixel_1660/VDD pixel_1660/GND pixel_1660/VREF pixel_1660/ROW_SEL
+ pixel_1660/NB1 pixel_1660/VBIAS pixel_1660/NB2 pixel_1660/AMP_IN pixel_1660/SF_IB
+ pixel_1660/PIX_OUT pixel_1660/CSA_VREF pixel
Xpixel_2394 pixel_2394/gring pixel_2394/VDD pixel_2394/GND pixel_2394/VREF pixel_2394/ROW_SEL
+ pixel_2394/NB1 pixel_2394/VBIAS pixel_2394/NB2 pixel_2394/AMP_IN pixel_2394/SF_IB
+ pixel_2394/PIX_OUT pixel_2394/CSA_VREF pixel
Xpixel_2383 pixel_2383/gring pixel_2383/VDD pixel_2383/GND pixel_2383/VREF pixel_2383/ROW_SEL
+ pixel_2383/NB1 pixel_2383/VBIAS pixel_2383/NB2 pixel_2383/AMP_IN pixel_2383/SF_IB
+ pixel_2383/PIX_OUT pixel_2383/CSA_VREF pixel
Xpixel_1693 pixel_1693/gring pixel_1693/VDD pixel_1693/GND pixel_1693/VREF pixel_1693/ROW_SEL
+ pixel_1693/NB1 pixel_1693/VBIAS pixel_1693/NB2 pixel_1693/AMP_IN pixel_1693/SF_IB
+ pixel_1693/PIX_OUT pixel_1693/CSA_VREF pixel
Xpixel_1682 pixel_1682/gring pixel_1682/VDD pixel_1682/GND pixel_1682/VREF pixel_1682/ROW_SEL
+ pixel_1682/NB1 pixel_1682/VBIAS pixel_1682/NB2 pixel_1682/AMP_IN pixel_1682/SF_IB
+ pixel_1682/PIX_OUT pixel_1682/CSA_VREF pixel
Xpixel_1671 pixel_1671/gring pixel_1671/VDD pixel_1671/GND pixel_1671/VREF pixel_1671/ROW_SEL
+ pixel_1671/NB1 pixel_1671/VBIAS pixel_1671/NB2 pixel_1671/AMP_IN pixel_1671/SF_IB
+ pixel_1671/PIX_OUT pixel_1671/CSA_VREF pixel
Xpixel_9990 pixel_9990/gring pixel_9990/VDD pixel_9990/GND pixel_9990/VREF pixel_9990/ROW_SEL
+ pixel_9990/NB1 pixel_9990/VBIAS pixel_9990/NB2 pixel_9990/AMP_IN pixel_9990/SF_IB
+ pixel_9990/PIX_OUT pixel_9990/CSA_VREF pixel
Xpixel_719 pixel_719/gring pixel_719/VDD pixel_719/GND pixel_719/VREF pixel_719/ROW_SEL
+ pixel_719/NB1 pixel_719/VBIAS pixel_719/NB2 pixel_719/AMP_IN pixel_719/SF_IB pixel_719/PIX_OUT
+ pixel_719/CSA_VREF pixel
Xpixel_708 pixel_708/gring pixel_708/VDD pixel_708/GND pixel_708/VREF pixel_708/ROW_SEL
+ pixel_708/NB1 pixel_708/VBIAS pixel_708/NB2 pixel_708/AMP_IN pixel_708/SF_IB pixel_708/PIX_OUT
+ pixel_708/CSA_VREF pixel
Xpixel_8007 pixel_8007/gring pixel_8007/VDD pixel_8007/GND pixel_8007/VREF pixel_8007/ROW_SEL
+ pixel_8007/NB1 pixel_8007/VBIAS pixel_8007/NB2 pixel_8007/AMP_IN pixel_8007/SF_IB
+ pixel_8007/PIX_OUT pixel_8007/CSA_VREF pixel
Xpixel_8018 pixel_8018/gring pixel_8018/VDD pixel_8018/GND pixel_8018/VREF pixel_8018/ROW_SEL
+ pixel_8018/NB1 pixel_8018/VBIAS pixel_8018/NB2 pixel_8018/AMP_IN pixel_8018/SF_IB
+ pixel_8018/PIX_OUT pixel_8018/CSA_VREF pixel
Xpixel_8029 pixel_8029/gring pixel_8029/VDD pixel_8029/GND pixel_8029/VREF pixel_8029/ROW_SEL
+ pixel_8029/NB1 pixel_8029/VBIAS pixel_8029/NB2 pixel_8029/AMP_IN pixel_8029/SF_IB
+ pixel_8029/PIX_OUT pixel_8029/CSA_VREF pixel
Xpixel_7306 pixel_7306/gring pixel_7306/VDD pixel_7306/GND pixel_7306/VREF pixel_7306/ROW_SEL
+ pixel_7306/NB1 pixel_7306/VBIAS pixel_7306/NB2 pixel_7306/AMP_IN pixel_7306/SF_IB
+ pixel_7306/PIX_OUT pixel_7306/CSA_VREF pixel
Xpixel_7317 pixel_7317/gring pixel_7317/VDD pixel_7317/GND pixel_7317/VREF pixel_7317/ROW_SEL
+ pixel_7317/NB1 pixel_7317/VBIAS pixel_7317/NB2 pixel_7317/AMP_IN pixel_7317/SF_IB
+ pixel_7317/PIX_OUT pixel_7317/CSA_VREF pixel
Xpixel_7328 pixel_7328/gring pixel_7328/VDD pixel_7328/GND pixel_7328/VREF pixel_7328/ROW_SEL
+ pixel_7328/NB1 pixel_7328/VBIAS pixel_7328/NB2 pixel_7328/AMP_IN pixel_7328/SF_IB
+ pixel_7328/PIX_OUT pixel_7328/CSA_VREF pixel
Xpixel_7339 pixel_7339/gring pixel_7339/VDD pixel_7339/GND pixel_7339/VREF pixel_7339/ROW_SEL
+ pixel_7339/NB1 pixel_7339/VBIAS pixel_7339/NB2 pixel_7339/AMP_IN pixel_7339/SF_IB
+ pixel_7339/PIX_OUT pixel_7339/CSA_VREF pixel
Xpixel_6605 pixel_6605/gring pixel_6605/VDD pixel_6605/GND pixel_6605/VREF pixel_6605/ROW_SEL
+ pixel_6605/NB1 pixel_6605/VBIAS pixel_6605/NB2 pixel_6605/AMP_IN pixel_6605/SF_IB
+ pixel_6605/PIX_OUT pixel_6605/CSA_VREF pixel
Xpixel_6616 pixel_6616/gring pixel_6616/VDD pixel_6616/GND pixel_6616/VREF pixel_6616/ROW_SEL
+ pixel_6616/NB1 pixel_6616/VBIAS pixel_6616/NB2 pixel_6616/AMP_IN pixel_6616/SF_IB
+ pixel_6616/PIX_OUT pixel_6616/CSA_VREF pixel
Xpixel_6627 pixel_6627/gring pixel_6627/VDD pixel_6627/GND pixel_6627/VREF pixel_6627/ROW_SEL
+ pixel_6627/NB1 pixel_6627/VBIAS pixel_6627/NB2 pixel_6627/AMP_IN pixel_6627/SF_IB
+ pixel_6627/PIX_OUT pixel_6627/CSA_VREF pixel
Xpixel_6638 pixel_6638/gring pixel_6638/VDD pixel_6638/GND pixel_6638/VREF pixel_6638/ROW_SEL
+ pixel_6638/NB1 pixel_6638/VBIAS pixel_6638/NB2 pixel_6638/AMP_IN pixel_6638/SF_IB
+ pixel_6638/PIX_OUT pixel_6638/CSA_VREF pixel
Xpixel_6649 pixel_6649/gring pixel_6649/VDD pixel_6649/GND pixel_6649/VREF pixel_6649/ROW_SEL
+ pixel_6649/NB1 pixel_6649/VBIAS pixel_6649/NB2 pixel_6649/AMP_IN pixel_6649/SF_IB
+ pixel_6649/PIX_OUT pixel_6649/CSA_VREF pixel
Xpixel_5904 pixel_5904/gring pixel_5904/VDD pixel_5904/GND pixel_5904/VREF pixel_5904/ROW_SEL
+ pixel_5904/NB1 pixel_5904/VBIAS pixel_5904/NB2 pixel_5904/AMP_IN pixel_5904/SF_IB
+ pixel_5904/PIX_OUT pixel_5904/CSA_VREF pixel
Xpixel_5915 pixel_5915/gring pixel_5915/VDD pixel_5915/GND pixel_5915/VREF pixel_5915/ROW_SEL
+ pixel_5915/NB1 pixel_5915/VBIAS pixel_5915/NB2 pixel_5915/AMP_IN pixel_5915/SF_IB
+ pixel_5915/PIX_OUT pixel_5915/CSA_VREF pixel
Xpixel_5926 pixel_5926/gring pixel_5926/VDD pixel_5926/GND pixel_5926/VREF pixel_5926/ROW_SEL
+ pixel_5926/NB1 pixel_5926/VBIAS pixel_5926/NB2 pixel_5926/AMP_IN pixel_5926/SF_IB
+ pixel_5926/PIX_OUT pixel_5926/CSA_VREF pixel
Xpixel_5937 pixel_5937/gring pixel_5937/VDD pixel_5937/GND pixel_5937/VREF pixel_5937/ROW_SEL
+ pixel_5937/NB1 pixel_5937/VBIAS pixel_5937/NB2 pixel_5937/AMP_IN pixel_5937/SF_IB
+ pixel_5937/PIX_OUT pixel_5937/CSA_VREF pixel
Xpixel_5948 pixel_5948/gring pixel_5948/VDD pixel_5948/GND pixel_5948/VREF pixel_5948/ROW_SEL
+ pixel_5948/NB1 pixel_5948/VBIAS pixel_5948/NB2 pixel_5948/AMP_IN pixel_5948/SF_IB
+ pixel_5948/PIX_OUT pixel_5948/CSA_VREF pixel
Xpixel_5959 pixel_5959/gring pixel_5959/VDD pixel_5959/GND pixel_5959/VREF pixel_5959/ROW_SEL
+ pixel_5959/NB1 pixel_5959/VBIAS pixel_5959/NB2 pixel_5959/AMP_IN pixel_5959/SF_IB
+ pixel_5959/PIX_OUT pixel_5959/CSA_VREF pixel
Xpixel_9231 pixel_9231/gring pixel_9231/VDD pixel_9231/GND pixel_9231/VREF pixel_9231/ROW_SEL
+ pixel_9231/NB1 pixel_9231/VBIAS pixel_9231/NB2 pixel_9231/AMP_IN pixel_9231/SF_IB
+ pixel_9231/PIX_OUT pixel_9231/CSA_VREF pixel
Xpixel_9220 pixel_9220/gring pixel_9220/VDD pixel_9220/GND pixel_9220/VREF pixel_9220/ROW_SEL
+ pixel_9220/NB1 pixel_9220/VBIAS pixel_9220/NB2 pixel_9220/AMP_IN pixel_9220/SF_IB
+ pixel_9220/PIX_OUT pixel_9220/CSA_VREF pixel
Xpixel_9264 pixel_9264/gring pixel_9264/VDD pixel_9264/GND pixel_9264/VREF pixel_9264/ROW_SEL
+ pixel_9264/NB1 pixel_9264/VBIAS pixel_9264/NB2 pixel_9264/AMP_IN pixel_9264/SF_IB
+ pixel_9264/PIX_OUT pixel_9264/CSA_VREF pixel
Xpixel_9253 pixel_9253/gring pixel_9253/VDD pixel_9253/GND pixel_9253/VREF pixel_9253/ROW_SEL
+ pixel_9253/NB1 pixel_9253/VBIAS pixel_9253/NB2 pixel_9253/AMP_IN pixel_9253/SF_IB
+ pixel_9253/PIX_OUT pixel_9253/CSA_VREF pixel
Xpixel_9242 pixel_9242/gring pixel_9242/VDD pixel_9242/GND pixel_9242/VREF pixel_9242/ROW_SEL
+ pixel_9242/NB1 pixel_9242/VBIAS pixel_9242/NB2 pixel_9242/AMP_IN pixel_9242/SF_IB
+ pixel_9242/PIX_OUT pixel_9242/CSA_VREF pixel
Xpixel_8563 pixel_8563/gring pixel_8563/VDD pixel_8563/GND pixel_8563/VREF pixel_8563/ROW_SEL
+ pixel_8563/NB1 pixel_8563/VBIAS pixel_8563/NB2 pixel_8563/AMP_IN pixel_8563/SF_IB
+ pixel_8563/PIX_OUT pixel_8563/CSA_VREF pixel
Xpixel_8552 pixel_8552/gring pixel_8552/VDD pixel_8552/GND pixel_8552/VREF pixel_8552/ROW_SEL
+ pixel_8552/NB1 pixel_8552/VBIAS pixel_8552/NB2 pixel_8552/AMP_IN pixel_8552/SF_IB
+ pixel_8552/PIX_OUT pixel_8552/CSA_VREF pixel
Xpixel_8541 pixel_8541/gring pixel_8541/VDD pixel_8541/GND pixel_8541/VREF pixel_8541/ROW_SEL
+ pixel_8541/NB1 pixel_8541/VBIAS pixel_8541/NB2 pixel_8541/AMP_IN pixel_8541/SF_IB
+ pixel_8541/PIX_OUT pixel_8541/CSA_VREF pixel
Xpixel_8530 pixel_8530/gring pixel_8530/VDD pixel_8530/GND pixel_8530/VREF pixel_8530/ROW_SEL
+ pixel_8530/NB1 pixel_8530/VBIAS pixel_8530/NB2 pixel_8530/AMP_IN pixel_8530/SF_IB
+ pixel_8530/PIX_OUT pixel_8530/CSA_VREF pixel
Xpixel_9297 pixel_9297/gring pixel_9297/VDD pixel_9297/GND pixel_9297/VREF pixel_9297/ROW_SEL
+ pixel_9297/NB1 pixel_9297/VBIAS pixel_9297/NB2 pixel_9297/AMP_IN pixel_9297/SF_IB
+ pixel_9297/PIX_OUT pixel_9297/CSA_VREF pixel
Xpixel_9286 pixel_9286/gring pixel_9286/VDD pixel_9286/GND pixel_9286/VREF pixel_9286/ROW_SEL
+ pixel_9286/NB1 pixel_9286/VBIAS pixel_9286/NB2 pixel_9286/AMP_IN pixel_9286/SF_IB
+ pixel_9286/PIX_OUT pixel_9286/CSA_VREF pixel
Xpixel_9275 pixel_9275/gring pixel_9275/VDD pixel_9275/GND pixel_9275/VREF pixel_9275/ROW_SEL
+ pixel_9275/NB1 pixel_9275/VBIAS pixel_9275/NB2 pixel_9275/AMP_IN pixel_9275/SF_IB
+ pixel_9275/PIX_OUT pixel_9275/CSA_VREF pixel
Xpixel_8596 pixel_8596/gring pixel_8596/VDD pixel_8596/GND pixel_8596/VREF pixel_8596/ROW_SEL
+ pixel_8596/NB1 pixel_8596/VBIAS pixel_8596/NB2 pixel_8596/AMP_IN pixel_8596/SF_IB
+ pixel_8596/PIX_OUT pixel_8596/CSA_VREF pixel
Xpixel_8585 pixel_8585/gring pixel_8585/VDD pixel_8585/GND pixel_8585/VREF pixel_8585/ROW_SEL
+ pixel_8585/NB1 pixel_8585/VBIAS pixel_8585/NB2 pixel_8585/AMP_IN pixel_8585/SF_IB
+ pixel_8585/PIX_OUT pixel_8585/CSA_VREF pixel
Xpixel_8574 pixel_8574/gring pixel_8574/VDD pixel_8574/GND pixel_8574/VREF pixel_8574/ROW_SEL
+ pixel_8574/NB1 pixel_8574/VBIAS pixel_8574/NB2 pixel_8574/AMP_IN pixel_8574/SF_IB
+ pixel_8574/PIX_OUT pixel_8574/CSA_VREF pixel
Xpixel_7840 pixel_7840/gring pixel_7840/VDD pixel_7840/GND pixel_7840/VREF pixel_7840/ROW_SEL
+ pixel_7840/NB1 pixel_7840/VBIAS pixel_7840/NB2 pixel_7840/AMP_IN pixel_7840/SF_IB
+ pixel_7840/PIX_OUT pixel_7840/CSA_VREF pixel
Xpixel_7851 pixel_7851/gring pixel_7851/VDD pixel_7851/GND pixel_7851/VREF pixel_7851/ROW_SEL
+ pixel_7851/NB1 pixel_7851/VBIAS pixel_7851/NB2 pixel_7851/AMP_IN pixel_7851/SF_IB
+ pixel_7851/PIX_OUT pixel_7851/CSA_VREF pixel
Xpixel_7862 pixel_7862/gring pixel_7862/VDD pixel_7862/GND pixel_7862/VREF pixel_7862/ROW_SEL
+ pixel_7862/NB1 pixel_7862/VBIAS pixel_7862/NB2 pixel_7862/AMP_IN pixel_7862/SF_IB
+ pixel_7862/PIX_OUT pixel_7862/CSA_VREF pixel
Xpixel_7873 pixel_7873/gring pixel_7873/VDD pixel_7873/GND pixel_7873/VREF pixel_7873/ROW_SEL
+ pixel_7873/NB1 pixel_7873/VBIAS pixel_7873/NB2 pixel_7873/AMP_IN pixel_7873/SF_IB
+ pixel_7873/PIX_OUT pixel_7873/CSA_VREF pixel
Xpixel_7884 pixel_7884/gring pixel_7884/VDD pixel_7884/GND pixel_7884/VREF pixel_7884/ROW_SEL
+ pixel_7884/NB1 pixel_7884/VBIAS pixel_7884/NB2 pixel_7884/AMP_IN pixel_7884/SF_IB
+ pixel_7884/PIX_OUT pixel_7884/CSA_VREF pixel
Xpixel_7895 pixel_7895/gring pixel_7895/VDD pixel_7895/GND pixel_7895/VREF pixel_7895/ROW_SEL
+ pixel_7895/NB1 pixel_7895/VBIAS pixel_7895/NB2 pixel_7895/AMP_IN pixel_7895/SF_IB
+ pixel_7895/PIX_OUT pixel_7895/CSA_VREF pixel
Xpixel_2180 pixel_2180/gring pixel_2180/VDD pixel_2180/GND pixel_2180/VREF pixel_2180/ROW_SEL
+ pixel_2180/NB1 pixel_2180/VBIAS pixel_2180/NB2 pixel_2180/AMP_IN pixel_2180/SF_IB
+ pixel_2180/PIX_OUT pixel_2180/CSA_VREF pixel
Xpixel_2191 pixel_2191/gring pixel_2191/VDD pixel_2191/GND pixel_2191/VREF pixel_2191/ROW_SEL
+ pixel_2191/NB1 pixel_2191/VBIAS pixel_2191/NB2 pixel_2191/AMP_IN pixel_2191/SF_IB
+ pixel_2191/PIX_OUT pixel_2191/CSA_VREF pixel
Xpixel_1490 pixel_1490/gring pixel_1490/VDD pixel_1490/GND pixel_1490/VREF pixel_1490/ROW_SEL
+ pixel_1490/NB1 pixel_1490/VBIAS pixel_1490/NB2 pixel_1490/AMP_IN pixel_1490/SF_IB
+ pixel_1490/PIX_OUT pixel_1490/CSA_VREF pixel
Xpixel_505 pixel_505/gring pixel_505/VDD pixel_505/GND pixel_505/VREF pixel_505/ROW_SEL
+ pixel_505/NB1 pixel_505/VBIAS pixel_505/NB2 pixel_505/AMP_IN pixel_505/SF_IB pixel_505/PIX_OUT
+ pixel_505/CSA_VREF pixel
Xpixel_538 pixel_538/gring pixel_538/VDD pixel_538/GND pixel_538/VREF pixel_538/ROW_SEL
+ pixel_538/NB1 pixel_538/VBIAS pixel_538/NB2 pixel_538/AMP_IN pixel_538/SF_IB pixel_538/PIX_OUT
+ pixel_538/CSA_VREF pixel
Xpixel_527 pixel_527/gring pixel_527/VDD pixel_527/GND pixel_527/VREF pixel_527/ROW_SEL
+ pixel_527/NB1 pixel_527/VBIAS pixel_527/NB2 pixel_527/AMP_IN pixel_527/SF_IB pixel_527/PIX_OUT
+ pixel_527/CSA_VREF pixel
Xpixel_516 pixel_516/gring pixel_516/VDD pixel_516/GND pixel_516/VREF pixel_516/ROW_SEL
+ pixel_516/NB1 pixel_516/VBIAS pixel_516/NB2 pixel_516/AMP_IN pixel_516/SF_IB pixel_516/PIX_OUT
+ pixel_516/CSA_VREF pixel
Xpixel_549 pixel_549/gring pixel_549/VDD pixel_549/GND pixel_549/VREF pixel_549/ROW_SEL
+ pixel_549/NB1 pixel_549/VBIAS pixel_549/NB2 pixel_549/AMP_IN pixel_549/SF_IB pixel_549/PIX_OUT
+ pixel_549/CSA_VREF pixel
Xpixel_3809 pixel_3809/gring pixel_3809/VDD pixel_3809/GND pixel_3809/VREF pixel_3809/ROW_SEL
+ pixel_3809/NB1 pixel_3809/VBIAS pixel_3809/NB2 pixel_3809/AMP_IN pixel_3809/SF_IB
+ pixel_3809/PIX_OUT pixel_3809/CSA_VREF pixel
Xpixel_7103 pixel_7103/gring pixel_7103/VDD pixel_7103/GND pixel_7103/VREF pixel_7103/ROW_SEL
+ pixel_7103/NB1 pixel_7103/VBIAS pixel_7103/NB2 pixel_7103/AMP_IN pixel_7103/SF_IB
+ pixel_7103/PIX_OUT pixel_7103/CSA_VREF pixel
Xpixel_7114 pixel_7114/gring pixel_7114/VDD pixel_7114/GND pixel_7114/VREF pixel_7114/ROW_SEL
+ pixel_7114/NB1 pixel_7114/VBIAS pixel_7114/NB2 pixel_7114/AMP_IN pixel_7114/SF_IB
+ pixel_7114/PIX_OUT pixel_7114/CSA_VREF pixel
Xpixel_7125 pixel_7125/gring pixel_7125/VDD pixel_7125/GND pixel_7125/VREF pixel_7125/ROW_SEL
+ pixel_7125/NB1 pixel_7125/VBIAS pixel_7125/NB2 pixel_7125/AMP_IN pixel_7125/SF_IB
+ pixel_7125/PIX_OUT pixel_7125/CSA_VREF pixel
Xpixel_7136 pixel_7136/gring pixel_7136/VDD pixel_7136/GND pixel_7136/VREF pixel_7136/ROW_SEL
+ pixel_7136/NB1 pixel_7136/VBIAS pixel_7136/NB2 pixel_7136/AMP_IN pixel_7136/SF_IB
+ pixel_7136/PIX_OUT pixel_7136/CSA_VREF pixel
Xpixel_7147 pixel_7147/gring pixel_7147/VDD pixel_7147/GND pixel_7147/VREF pixel_7147/ROW_SEL
+ pixel_7147/NB1 pixel_7147/VBIAS pixel_7147/NB2 pixel_7147/AMP_IN pixel_7147/SF_IB
+ pixel_7147/PIX_OUT pixel_7147/CSA_VREF pixel
Xpixel_6402 pixel_6402/gring pixel_6402/VDD pixel_6402/GND pixel_6402/VREF pixel_6402/ROW_SEL
+ pixel_6402/NB1 pixel_6402/VBIAS pixel_6402/NB2 pixel_6402/AMP_IN pixel_6402/SF_IB
+ pixel_6402/PIX_OUT pixel_6402/CSA_VREF pixel
Xpixel_7158 pixel_7158/gring pixel_7158/VDD pixel_7158/GND pixel_7158/VREF pixel_7158/ROW_SEL
+ pixel_7158/NB1 pixel_7158/VBIAS pixel_7158/NB2 pixel_7158/AMP_IN pixel_7158/SF_IB
+ pixel_7158/PIX_OUT pixel_7158/CSA_VREF pixel
Xpixel_7169 pixel_7169/gring pixel_7169/VDD pixel_7169/GND pixel_7169/VREF pixel_7169/ROW_SEL
+ pixel_7169/NB1 pixel_7169/VBIAS pixel_7169/NB2 pixel_7169/AMP_IN pixel_7169/SF_IB
+ pixel_7169/PIX_OUT pixel_7169/CSA_VREF pixel
Xpixel_6413 pixel_6413/gring pixel_6413/VDD pixel_6413/GND pixel_6413/VREF pixel_6413/ROW_SEL
+ pixel_6413/NB1 pixel_6413/VBIAS pixel_6413/NB2 pixel_6413/AMP_IN pixel_6413/SF_IB
+ pixel_6413/PIX_OUT pixel_6413/CSA_VREF pixel
Xpixel_6424 pixel_6424/gring pixel_6424/VDD pixel_6424/GND pixel_6424/VREF pixel_6424/ROW_SEL
+ pixel_6424/NB1 pixel_6424/VBIAS pixel_6424/NB2 pixel_6424/AMP_IN pixel_6424/SF_IB
+ pixel_6424/PIX_OUT pixel_6424/CSA_VREF pixel
Xpixel_6435 pixel_6435/gring pixel_6435/VDD pixel_6435/GND pixel_6435/VREF pixel_6435/ROW_SEL
+ pixel_6435/NB1 pixel_6435/VBIAS pixel_6435/NB2 pixel_6435/AMP_IN pixel_6435/SF_IB
+ pixel_6435/PIX_OUT pixel_6435/CSA_VREF pixel
Xpixel_6446 pixel_6446/gring pixel_6446/VDD pixel_6446/GND pixel_6446/VREF pixel_6446/ROW_SEL
+ pixel_6446/NB1 pixel_6446/VBIAS pixel_6446/NB2 pixel_6446/AMP_IN pixel_6446/SF_IB
+ pixel_6446/PIX_OUT pixel_6446/CSA_VREF pixel
Xpixel_6457 pixel_6457/gring pixel_6457/VDD pixel_6457/GND pixel_6457/VREF pixel_6457/ROW_SEL
+ pixel_6457/NB1 pixel_6457/VBIAS pixel_6457/NB2 pixel_6457/AMP_IN pixel_6457/SF_IB
+ pixel_6457/PIX_OUT pixel_6457/CSA_VREF pixel
Xpixel_6468 pixel_6468/gring pixel_6468/VDD pixel_6468/GND pixel_6468/VREF pixel_6468/ROW_SEL
+ pixel_6468/NB1 pixel_6468/VBIAS pixel_6468/NB2 pixel_6468/AMP_IN pixel_6468/SF_IB
+ pixel_6468/PIX_OUT pixel_6468/CSA_VREF pixel
Xpixel_5701 pixel_5701/gring pixel_5701/VDD pixel_5701/GND pixel_5701/VREF pixel_5701/ROW_SEL
+ pixel_5701/NB1 pixel_5701/VBIAS pixel_5701/NB2 pixel_5701/AMP_IN pixel_5701/SF_IB
+ pixel_5701/PIX_OUT pixel_5701/CSA_VREF pixel
Xpixel_5712 pixel_5712/gring pixel_5712/VDD pixel_5712/GND pixel_5712/VREF pixel_5712/ROW_SEL
+ pixel_5712/NB1 pixel_5712/VBIAS pixel_5712/NB2 pixel_5712/AMP_IN pixel_5712/SF_IB
+ pixel_5712/PIX_OUT pixel_5712/CSA_VREF pixel
Xpixel_5723 pixel_5723/gring pixel_5723/VDD pixel_5723/GND pixel_5723/VREF pixel_5723/ROW_SEL
+ pixel_5723/NB1 pixel_5723/VBIAS pixel_5723/NB2 pixel_5723/AMP_IN pixel_5723/SF_IB
+ pixel_5723/PIX_OUT pixel_5723/CSA_VREF pixel
Xpixel_5734 pixel_5734/gring pixel_5734/VDD pixel_5734/GND pixel_5734/VREF pixel_5734/ROW_SEL
+ pixel_5734/NB1 pixel_5734/VBIAS pixel_5734/NB2 pixel_5734/AMP_IN pixel_5734/SF_IB
+ pixel_5734/PIX_OUT pixel_5734/CSA_VREF pixel
Xpixel_6479 pixel_6479/gring pixel_6479/VDD pixel_6479/GND pixel_6479/VREF pixel_6479/ROW_SEL
+ pixel_6479/NB1 pixel_6479/VBIAS pixel_6479/NB2 pixel_6479/AMP_IN pixel_6479/SF_IB
+ pixel_6479/PIX_OUT pixel_6479/CSA_VREF pixel
Xpixel_5745 pixel_5745/gring pixel_5745/VDD pixel_5745/GND pixel_5745/VREF pixel_5745/ROW_SEL
+ pixel_5745/NB1 pixel_5745/VBIAS pixel_5745/NB2 pixel_5745/AMP_IN pixel_5745/SF_IB
+ pixel_5745/PIX_OUT pixel_5745/CSA_VREF pixel
Xpixel_5756 pixel_5756/gring pixel_5756/VDD pixel_5756/GND pixel_5756/VREF pixel_5756/ROW_SEL
+ pixel_5756/NB1 pixel_5756/VBIAS pixel_5756/NB2 pixel_5756/AMP_IN pixel_5756/SF_IB
+ pixel_5756/PIX_OUT pixel_5756/CSA_VREF pixel
Xpixel_5767 pixel_5767/gring pixel_5767/VDD pixel_5767/GND pixel_5767/VREF pixel_5767/ROW_SEL
+ pixel_5767/NB1 pixel_5767/VBIAS pixel_5767/NB2 pixel_5767/AMP_IN pixel_5767/SF_IB
+ pixel_5767/PIX_OUT pixel_5767/CSA_VREF pixel
Xpixel_5778 pixel_5778/gring pixel_5778/VDD pixel_5778/GND pixel_5778/VREF pixel_5778/ROW_SEL
+ pixel_5778/NB1 pixel_5778/VBIAS pixel_5778/NB2 pixel_5778/AMP_IN pixel_5778/SF_IB
+ pixel_5778/PIX_OUT pixel_5778/CSA_VREF pixel
Xpixel_5789 pixel_5789/gring pixel_5789/VDD pixel_5789/GND pixel_5789/VREF pixel_5789/ROW_SEL
+ pixel_5789/NB1 pixel_5789/VBIAS pixel_5789/NB2 pixel_5789/AMP_IN pixel_5789/SF_IB
+ pixel_5789/PIX_OUT pixel_5789/CSA_VREF pixel
Xpixel_9072 pixel_9072/gring pixel_9072/VDD pixel_9072/GND pixel_9072/VREF pixel_9072/ROW_SEL
+ pixel_9072/NB1 pixel_9072/VBIAS pixel_9072/NB2 pixel_9072/AMP_IN pixel_9072/SF_IB
+ pixel_9072/PIX_OUT pixel_9072/CSA_VREF pixel
Xpixel_9061 pixel_9061/gring pixel_9061/VDD pixel_9061/GND pixel_9061/VREF pixel_9061/ROW_SEL
+ pixel_9061/NB1 pixel_9061/VBIAS pixel_9061/NB2 pixel_9061/AMP_IN pixel_9061/SF_IB
+ pixel_9061/PIX_OUT pixel_9061/CSA_VREF pixel
Xpixel_9050 pixel_9050/gring pixel_9050/VDD pixel_9050/GND pixel_9050/VREF pixel_9050/ROW_SEL
+ pixel_9050/NB1 pixel_9050/VBIAS pixel_9050/NB2 pixel_9050/AMP_IN pixel_9050/SF_IB
+ pixel_9050/PIX_OUT pixel_9050/CSA_VREF pixel
Xpixel_9094 pixel_9094/gring pixel_9094/VDD pixel_9094/GND pixel_9094/VREF pixel_9094/ROW_SEL
+ pixel_9094/NB1 pixel_9094/VBIAS pixel_9094/NB2 pixel_9094/AMP_IN pixel_9094/SF_IB
+ pixel_9094/PIX_OUT pixel_9094/CSA_VREF pixel
Xpixel_9083 pixel_9083/gring pixel_9083/VDD pixel_9083/GND pixel_9083/VREF pixel_9083/ROW_SEL
+ pixel_9083/NB1 pixel_9083/VBIAS pixel_9083/NB2 pixel_9083/AMP_IN pixel_9083/SF_IB
+ pixel_9083/PIX_OUT pixel_9083/CSA_VREF pixel
Xpixel_8360 pixel_8360/gring pixel_8360/VDD pixel_8360/GND pixel_8360/VREF pixel_8360/ROW_SEL
+ pixel_8360/NB1 pixel_8360/VBIAS pixel_8360/NB2 pixel_8360/AMP_IN pixel_8360/SF_IB
+ pixel_8360/PIX_OUT pixel_8360/CSA_VREF pixel
Xpixel_8371 pixel_8371/gring pixel_8371/VDD pixel_8371/GND pixel_8371/VREF pixel_8371/ROW_SEL
+ pixel_8371/NB1 pixel_8371/VBIAS pixel_8371/NB2 pixel_8371/AMP_IN pixel_8371/SF_IB
+ pixel_8371/PIX_OUT pixel_8371/CSA_VREF pixel
Xpixel_8382 pixel_8382/gring pixel_8382/VDD pixel_8382/GND pixel_8382/VREF pixel_8382/ROW_SEL
+ pixel_8382/NB1 pixel_8382/VBIAS pixel_8382/NB2 pixel_8382/AMP_IN pixel_8382/SF_IB
+ pixel_8382/PIX_OUT pixel_8382/CSA_VREF pixel
Xpixel_8393 pixel_8393/gring pixel_8393/VDD pixel_8393/GND pixel_8393/VREF pixel_8393/ROW_SEL
+ pixel_8393/NB1 pixel_8393/VBIAS pixel_8393/NB2 pixel_8393/AMP_IN pixel_8393/SF_IB
+ pixel_8393/PIX_OUT pixel_8393/CSA_VREF pixel
Xpixel_7670 pixel_7670/gring pixel_7670/VDD pixel_7670/GND pixel_7670/VREF pixel_7670/ROW_SEL
+ pixel_7670/NB1 pixel_7670/VBIAS pixel_7670/NB2 pixel_7670/AMP_IN pixel_7670/SF_IB
+ pixel_7670/PIX_OUT pixel_7670/CSA_VREF pixel
Xpixel_7681 pixel_7681/gring pixel_7681/VDD pixel_7681/GND pixel_7681/VREF pixel_7681/ROW_SEL
+ pixel_7681/NB1 pixel_7681/VBIAS pixel_7681/NB2 pixel_7681/AMP_IN pixel_7681/SF_IB
+ pixel_7681/PIX_OUT pixel_7681/CSA_VREF pixel
Xpixel_7692 pixel_7692/gring pixel_7692/VDD pixel_7692/GND pixel_7692/VREF pixel_7692/ROW_SEL
+ pixel_7692/NB1 pixel_7692/VBIAS pixel_7692/NB2 pixel_7692/AMP_IN pixel_7692/SF_IB
+ pixel_7692/PIX_OUT pixel_7692/CSA_VREF pixel
Xpixel_6980 pixel_6980/gring pixel_6980/VDD pixel_6980/GND pixel_6980/VREF pixel_6980/ROW_SEL
+ pixel_6980/NB1 pixel_6980/VBIAS pixel_6980/NB2 pixel_6980/AMP_IN pixel_6980/SF_IB
+ pixel_6980/PIX_OUT pixel_6980/CSA_VREF pixel
Xpixel_6991 pixel_6991/gring pixel_6991/VDD pixel_6991/GND pixel_6991/VREF pixel_6991/ROW_SEL
+ pixel_6991/NB1 pixel_6991/VBIAS pixel_6991/NB2 pixel_6991/AMP_IN pixel_6991/SF_IB
+ pixel_6991/PIX_OUT pixel_6991/CSA_VREF pixel
Xpixel_72 pixel_72/gring pixel_72/VDD pixel_72/GND pixel_72/VREF pixel_72/ROW_SEL
+ pixel_72/NB1 pixel_72/VBIAS pixel_72/NB2 pixel_72/AMP_IN pixel_72/SF_IB pixel_72/PIX_OUT
+ pixel_72/CSA_VREF pixel
Xpixel_61 pixel_61/gring pixel_61/VDD pixel_61/GND pixel_61/VREF pixel_61/ROW_SEL
+ pixel_61/NB1 pixel_61/VBIAS pixel_61/NB2 pixel_61/AMP_IN pixel_61/SF_IB pixel_61/PIX_OUT
+ pixel_61/CSA_VREF pixel
Xpixel_50 pixel_50/gring pixel_50/VDD pixel_50/GND pixel_50/VREF pixel_50/ROW_SEL
+ pixel_50/NB1 pixel_50/VBIAS pixel_50/NB2 pixel_50/AMP_IN pixel_50/SF_IB pixel_50/PIX_OUT
+ pixel_50/CSA_VREF pixel
Xpixel_94 pixel_94/gring pixel_94/VDD pixel_94/GND pixel_94/VREF pixel_94/ROW_SEL
+ pixel_94/NB1 pixel_94/VBIAS pixel_94/NB2 pixel_94/AMP_IN pixel_94/SF_IB pixel_94/PIX_OUT
+ pixel_94/CSA_VREF pixel
Xpixel_83 pixel_83/gring pixel_83/VDD pixel_83/GND pixel_83/VREF pixel_83/ROW_SEL
+ pixel_83/NB1 pixel_83/VBIAS pixel_83/NB2 pixel_83/AMP_IN pixel_83/SF_IB pixel_83/PIX_OUT
+ pixel_83/CSA_VREF pixel
Xpixel_5008 pixel_5008/gring pixel_5008/VDD pixel_5008/GND pixel_5008/VREF pixel_5008/ROW_SEL
+ pixel_5008/NB1 pixel_5008/VBIAS pixel_5008/NB2 pixel_5008/AMP_IN pixel_5008/SF_IB
+ pixel_5008/PIX_OUT pixel_5008/CSA_VREF pixel
Xpixel_5019 pixel_5019/gring pixel_5019/VDD pixel_5019/GND pixel_5019/VREF pixel_5019/ROW_SEL
+ pixel_5019/NB1 pixel_5019/VBIAS pixel_5019/NB2 pixel_5019/AMP_IN pixel_5019/SF_IB
+ pixel_5019/PIX_OUT pixel_5019/CSA_VREF pixel
Xpixel_313 pixel_313/gring pixel_313/VDD pixel_313/GND pixel_313/VREF pixel_313/ROW_SEL
+ pixel_313/NB1 pixel_313/VBIAS pixel_313/NB2 pixel_313/AMP_IN pixel_313/SF_IB pixel_313/PIX_OUT
+ pixel_313/CSA_VREF pixel
Xpixel_302 pixel_302/gring pixel_302/VDD pixel_302/GND pixel_302/VREF pixel_302/ROW_SEL
+ pixel_302/NB1 pixel_302/VBIAS pixel_302/NB2 pixel_302/AMP_IN pixel_302/SF_IB pixel_302/PIX_OUT
+ pixel_302/CSA_VREF pixel
Xpixel_4307 pixel_4307/gring pixel_4307/VDD pixel_4307/GND pixel_4307/VREF pixel_4307/ROW_SEL
+ pixel_4307/NB1 pixel_4307/VBIAS pixel_4307/NB2 pixel_4307/AMP_IN pixel_4307/SF_IB
+ pixel_4307/PIX_OUT pixel_4307/CSA_VREF pixel
Xpixel_4318 pixel_4318/gring pixel_4318/VDD pixel_4318/GND pixel_4318/VREF pixel_4318/ROW_SEL
+ pixel_4318/NB1 pixel_4318/VBIAS pixel_4318/NB2 pixel_4318/AMP_IN pixel_4318/SF_IB
+ pixel_4318/PIX_OUT pixel_4318/CSA_VREF pixel
Xpixel_346 pixel_346/gring pixel_346/VDD pixel_346/GND pixel_346/VREF pixel_346/ROW_SEL
+ pixel_346/NB1 pixel_346/VBIAS pixel_346/NB2 pixel_346/AMP_IN pixel_346/SF_IB pixel_346/PIX_OUT
+ pixel_346/CSA_VREF pixel
Xpixel_335 pixel_335/gring pixel_335/VDD pixel_335/GND pixel_335/VREF pixel_335/ROW_SEL
+ pixel_335/NB1 pixel_335/VBIAS pixel_335/NB2 pixel_335/AMP_IN pixel_335/SF_IB pixel_335/PIX_OUT
+ pixel_335/CSA_VREF pixel
Xpixel_324 pixel_324/gring pixel_324/VDD pixel_324/GND pixel_324/VREF pixel_324/ROW_SEL
+ pixel_324/NB1 pixel_324/VBIAS pixel_324/NB2 pixel_324/AMP_IN pixel_324/SF_IB pixel_324/PIX_OUT
+ pixel_324/CSA_VREF pixel
Xpixel_3606 pixel_3606/gring pixel_3606/VDD pixel_3606/GND pixel_3606/VREF pixel_3606/ROW_SEL
+ pixel_3606/NB1 pixel_3606/VBIAS pixel_3606/NB2 pixel_3606/AMP_IN pixel_3606/SF_IB
+ pixel_3606/PIX_OUT pixel_3606/CSA_VREF pixel
Xpixel_4329 pixel_4329/gring pixel_4329/VDD pixel_4329/GND pixel_4329/VREF pixel_4329/ROW_SEL
+ pixel_4329/NB1 pixel_4329/VBIAS pixel_4329/NB2 pixel_4329/AMP_IN pixel_4329/SF_IB
+ pixel_4329/PIX_OUT pixel_4329/CSA_VREF pixel
Xpixel_379 pixel_379/gring pixel_379/VDD pixel_379/GND pixel_379/VREF pixel_379/ROW_SEL
+ pixel_379/NB1 pixel_379/VBIAS pixel_379/NB2 pixel_379/AMP_IN pixel_379/SF_IB pixel_379/PIX_OUT
+ pixel_379/CSA_VREF pixel
Xpixel_368 pixel_368/gring pixel_368/VDD pixel_368/GND pixel_368/VREF pixel_368/ROW_SEL
+ pixel_368/NB1 pixel_368/VBIAS pixel_368/NB2 pixel_368/AMP_IN pixel_368/SF_IB pixel_368/PIX_OUT
+ pixel_368/CSA_VREF pixel
Xpixel_357 pixel_357/gring pixel_357/VDD pixel_357/GND pixel_357/VREF pixel_357/ROW_SEL
+ pixel_357/NB1 pixel_357/VBIAS pixel_357/NB2 pixel_357/AMP_IN pixel_357/SF_IB pixel_357/PIX_OUT
+ pixel_357/CSA_VREF pixel
Xpixel_2905 pixel_2905/gring pixel_2905/VDD pixel_2905/GND pixel_2905/VREF pixel_2905/ROW_SEL
+ pixel_2905/NB1 pixel_2905/VBIAS pixel_2905/NB2 pixel_2905/AMP_IN pixel_2905/SF_IB
+ pixel_2905/PIX_OUT pixel_2905/CSA_VREF pixel
Xpixel_3639 pixel_3639/gring pixel_3639/VDD pixel_3639/GND pixel_3639/VREF pixel_3639/ROW_SEL
+ pixel_3639/NB1 pixel_3639/VBIAS pixel_3639/NB2 pixel_3639/AMP_IN pixel_3639/SF_IB
+ pixel_3639/PIX_OUT pixel_3639/CSA_VREF pixel
Xpixel_3628 pixel_3628/gring pixel_3628/VDD pixel_3628/GND pixel_3628/VREF pixel_3628/ROW_SEL
+ pixel_3628/NB1 pixel_3628/VBIAS pixel_3628/NB2 pixel_3628/AMP_IN pixel_3628/SF_IB
+ pixel_3628/PIX_OUT pixel_3628/CSA_VREF pixel
Xpixel_3617 pixel_3617/gring pixel_3617/VDD pixel_3617/GND pixel_3617/VREF pixel_3617/ROW_SEL
+ pixel_3617/NB1 pixel_3617/VBIAS pixel_3617/NB2 pixel_3617/AMP_IN pixel_3617/SF_IB
+ pixel_3617/PIX_OUT pixel_3617/CSA_VREF pixel
Xpixel_2938 pixel_2938/gring pixel_2938/VDD pixel_2938/GND pixel_2938/VREF pixel_2938/ROW_SEL
+ pixel_2938/NB1 pixel_2938/VBIAS pixel_2938/NB2 pixel_2938/AMP_IN pixel_2938/SF_IB
+ pixel_2938/PIX_OUT pixel_2938/CSA_VREF pixel
Xpixel_2927 pixel_2927/gring pixel_2927/VDD pixel_2927/GND pixel_2927/VREF pixel_2927/ROW_SEL
+ pixel_2927/NB1 pixel_2927/VBIAS pixel_2927/NB2 pixel_2927/AMP_IN pixel_2927/SF_IB
+ pixel_2927/PIX_OUT pixel_2927/CSA_VREF pixel
Xpixel_2916 pixel_2916/gring pixel_2916/VDD pixel_2916/GND pixel_2916/VREF pixel_2916/ROW_SEL
+ pixel_2916/NB1 pixel_2916/VBIAS pixel_2916/NB2 pixel_2916/AMP_IN pixel_2916/SF_IB
+ pixel_2916/PIX_OUT pixel_2916/CSA_VREF pixel
Xpixel_2949 pixel_2949/gring pixel_2949/VDD pixel_2949/GND pixel_2949/VREF pixel_2949/ROW_SEL
+ pixel_2949/NB1 pixel_2949/VBIAS pixel_2949/NB2 pixel_2949/AMP_IN pixel_2949/SF_IB
+ pixel_2949/PIX_OUT pixel_2949/CSA_VREF pixel
Xpixel_6210 pixel_6210/gring pixel_6210/VDD pixel_6210/GND pixel_6210/VREF pixel_6210/ROW_SEL
+ pixel_6210/NB1 pixel_6210/VBIAS pixel_6210/NB2 pixel_6210/AMP_IN pixel_6210/SF_IB
+ pixel_6210/PIX_OUT pixel_6210/CSA_VREF pixel
Xpixel_6221 pixel_6221/gring pixel_6221/VDD pixel_6221/GND pixel_6221/VREF pixel_6221/ROW_SEL
+ pixel_6221/NB1 pixel_6221/VBIAS pixel_6221/NB2 pixel_6221/AMP_IN pixel_6221/SF_IB
+ pixel_6221/PIX_OUT pixel_6221/CSA_VREF pixel
Xpixel_6232 pixel_6232/gring pixel_6232/VDD pixel_6232/GND pixel_6232/VREF pixel_6232/ROW_SEL
+ pixel_6232/NB1 pixel_6232/VBIAS pixel_6232/NB2 pixel_6232/AMP_IN pixel_6232/SF_IB
+ pixel_6232/PIX_OUT pixel_6232/CSA_VREF pixel
Xpixel_6243 pixel_6243/gring pixel_6243/VDD pixel_6243/GND pixel_6243/VREF pixel_6243/ROW_SEL
+ pixel_6243/NB1 pixel_6243/VBIAS pixel_6243/NB2 pixel_6243/AMP_IN pixel_6243/SF_IB
+ pixel_6243/PIX_OUT pixel_6243/CSA_VREF pixel
Xpixel_6254 pixel_6254/gring pixel_6254/VDD pixel_6254/GND pixel_6254/VREF pixel_6254/ROW_SEL
+ pixel_6254/NB1 pixel_6254/VBIAS pixel_6254/NB2 pixel_6254/AMP_IN pixel_6254/SF_IB
+ pixel_6254/PIX_OUT pixel_6254/CSA_VREF pixel
Xpixel_6265 pixel_6265/gring pixel_6265/VDD pixel_6265/GND pixel_6265/VREF pixel_6265/ROW_SEL
+ pixel_6265/NB1 pixel_6265/VBIAS pixel_6265/NB2 pixel_6265/AMP_IN pixel_6265/SF_IB
+ pixel_6265/PIX_OUT pixel_6265/CSA_VREF pixel
Xpixel_6276 pixel_6276/gring pixel_6276/VDD pixel_6276/GND pixel_6276/VREF pixel_6276/ROW_SEL
+ pixel_6276/NB1 pixel_6276/VBIAS pixel_6276/NB2 pixel_6276/AMP_IN pixel_6276/SF_IB
+ pixel_6276/PIX_OUT pixel_6276/CSA_VREF pixel
Xpixel_6287 pixel_6287/gring pixel_6287/VDD pixel_6287/GND pixel_6287/VREF pixel_6287/ROW_SEL
+ pixel_6287/NB1 pixel_6287/VBIAS pixel_6287/NB2 pixel_6287/AMP_IN pixel_6287/SF_IB
+ pixel_6287/PIX_OUT pixel_6287/CSA_VREF pixel
Xpixel_5520 pixel_5520/gring pixel_5520/VDD pixel_5520/GND pixel_5520/VREF pixel_5520/ROW_SEL
+ pixel_5520/NB1 pixel_5520/VBIAS pixel_5520/NB2 pixel_5520/AMP_IN pixel_5520/SF_IB
+ pixel_5520/PIX_OUT pixel_5520/CSA_VREF pixel
Xpixel_5531 pixel_5531/gring pixel_5531/VDD pixel_5531/GND pixel_5531/VREF pixel_5531/ROW_SEL
+ pixel_5531/NB1 pixel_5531/VBIAS pixel_5531/NB2 pixel_5531/AMP_IN pixel_5531/SF_IB
+ pixel_5531/PIX_OUT pixel_5531/CSA_VREF pixel
Xpixel_5542 pixel_5542/gring pixel_5542/VDD pixel_5542/GND pixel_5542/VREF pixel_5542/ROW_SEL
+ pixel_5542/NB1 pixel_5542/VBIAS pixel_5542/NB2 pixel_5542/AMP_IN pixel_5542/SF_IB
+ pixel_5542/PIX_OUT pixel_5542/CSA_VREF pixel
Xpixel_6298 pixel_6298/gring pixel_6298/VDD pixel_6298/GND pixel_6298/VREF pixel_6298/ROW_SEL
+ pixel_6298/NB1 pixel_6298/VBIAS pixel_6298/NB2 pixel_6298/AMP_IN pixel_6298/SF_IB
+ pixel_6298/PIX_OUT pixel_6298/CSA_VREF pixel
Xpixel_5553 pixel_5553/gring pixel_5553/VDD pixel_5553/GND pixel_5553/VREF pixel_5553/ROW_SEL
+ pixel_5553/NB1 pixel_5553/VBIAS pixel_5553/NB2 pixel_5553/AMP_IN pixel_5553/SF_IB
+ pixel_5553/PIX_OUT pixel_5553/CSA_VREF pixel
Xpixel_5564 pixel_5564/gring pixel_5564/VDD pixel_5564/GND pixel_5564/VREF pixel_5564/ROW_SEL
+ pixel_5564/NB1 pixel_5564/VBIAS pixel_5564/NB2 pixel_5564/AMP_IN pixel_5564/SF_IB
+ pixel_5564/PIX_OUT pixel_5564/CSA_VREF pixel
Xpixel_5575 pixel_5575/gring pixel_5575/VDD pixel_5575/GND pixel_5575/VREF pixel_5575/ROW_SEL
+ pixel_5575/NB1 pixel_5575/VBIAS pixel_5575/NB2 pixel_5575/AMP_IN pixel_5575/SF_IB
+ pixel_5575/PIX_OUT pixel_5575/CSA_VREF pixel
Xpixel_4830 pixel_4830/gring pixel_4830/VDD pixel_4830/GND pixel_4830/VREF pixel_4830/ROW_SEL
+ pixel_4830/NB1 pixel_4830/VBIAS pixel_4830/NB2 pixel_4830/AMP_IN pixel_4830/SF_IB
+ pixel_4830/PIX_OUT pixel_4830/CSA_VREF pixel
Xpixel_5586 pixel_5586/gring pixel_5586/VDD pixel_5586/GND pixel_5586/VREF pixel_5586/ROW_SEL
+ pixel_5586/NB1 pixel_5586/VBIAS pixel_5586/NB2 pixel_5586/AMP_IN pixel_5586/SF_IB
+ pixel_5586/PIX_OUT pixel_5586/CSA_VREF pixel
Xpixel_5597 pixel_5597/gring pixel_5597/VDD pixel_5597/GND pixel_5597/VREF pixel_5597/ROW_SEL
+ pixel_5597/NB1 pixel_5597/VBIAS pixel_5597/NB2 pixel_5597/AMP_IN pixel_5597/SF_IB
+ pixel_5597/PIX_OUT pixel_5597/CSA_VREF pixel
Xpixel_4841 pixel_4841/gring pixel_4841/VDD pixel_4841/GND pixel_4841/VREF pixel_4841/ROW_SEL
+ pixel_4841/NB1 pixel_4841/VBIAS pixel_4841/NB2 pixel_4841/AMP_IN pixel_4841/SF_IB
+ pixel_4841/PIX_OUT pixel_4841/CSA_VREF pixel
Xpixel_4852 pixel_4852/gring pixel_4852/VDD pixel_4852/GND pixel_4852/VREF pixel_4852/ROW_SEL
+ pixel_4852/NB1 pixel_4852/VBIAS pixel_4852/NB2 pixel_4852/AMP_IN pixel_4852/SF_IB
+ pixel_4852/PIX_OUT pixel_4852/CSA_VREF pixel
Xpixel_4863 pixel_4863/gring pixel_4863/VDD pixel_4863/GND pixel_4863/VREF pixel_4863/ROW_SEL
+ pixel_4863/NB1 pixel_4863/VBIAS pixel_4863/NB2 pixel_4863/AMP_IN pixel_4863/SF_IB
+ pixel_4863/PIX_OUT pixel_4863/CSA_VREF pixel
Xpixel_4874 pixel_4874/gring pixel_4874/VDD pixel_4874/GND pixel_4874/VREF pixel_4874/ROW_SEL
+ pixel_4874/NB1 pixel_4874/VBIAS pixel_4874/NB2 pixel_4874/AMP_IN pixel_4874/SF_IB
+ pixel_4874/PIX_OUT pixel_4874/CSA_VREF pixel
Xpixel_891 pixel_891/gring pixel_891/VDD pixel_891/GND pixel_891/VREF pixel_891/ROW_SEL
+ pixel_891/NB1 pixel_891/VBIAS pixel_891/NB2 pixel_891/AMP_IN pixel_891/SF_IB pixel_891/PIX_OUT
+ pixel_891/CSA_VREF pixel
Xpixel_880 pixel_880/gring pixel_880/VDD pixel_880/GND pixel_880/VREF pixel_880/ROW_SEL
+ pixel_880/NB1 pixel_880/VBIAS pixel_880/NB2 pixel_880/AMP_IN pixel_880/SF_IB pixel_880/PIX_OUT
+ pixel_880/CSA_VREF pixel
Xpixel_4885 pixel_4885/gring pixel_4885/VDD pixel_4885/GND pixel_4885/VREF pixel_4885/ROW_SEL
+ pixel_4885/NB1 pixel_4885/VBIAS pixel_4885/NB2 pixel_4885/AMP_IN pixel_4885/SF_IB
+ pixel_4885/PIX_OUT pixel_4885/CSA_VREF pixel
Xpixel_4896 pixel_4896/gring pixel_4896/VDD pixel_4896/GND pixel_4896/VREF pixel_4896/ROW_SEL
+ pixel_4896/NB1 pixel_4896/VBIAS pixel_4896/NB2 pixel_4896/AMP_IN pixel_4896/SF_IB
+ pixel_4896/PIX_OUT pixel_4896/CSA_VREF pixel
Xpixel_8190 pixel_8190/gring pixel_8190/VDD pixel_8190/GND pixel_8190/VREF pixel_8190/ROW_SEL
+ pixel_8190/NB1 pixel_8190/VBIAS pixel_8190/NB2 pixel_8190/AMP_IN pixel_8190/SF_IB
+ pixel_8190/PIX_OUT pixel_8190/CSA_VREF pixel
Xpixel_9819 pixel_9819/gring pixel_9819/VDD pixel_9819/GND pixel_9819/VREF pixel_9819/ROW_SEL
+ pixel_9819/NB1 pixel_9819/VBIAS pixel_9819/NB2 pixel_9819/AMP_IN pixel_9819/SF_IB
+ pixel_9819/PIX_OUT pixel_9819/CSA_VREF pixel
Xpixel_9808 pixel_9808/gring pixel_9808/VDD pixel_9808/GND pixel_9808/VREF pixel_9808/ROW_SEL
+ pixel_9808/NB1 pixel_9808/VBIAS pixel_9808/NB2 pixel_9808/AMP_IN pixel_9808/SF_IB
+ pixel_9808/PIX_OUT pixel_9808/CSA_VREF pixel
Xpixel_121 pixel_121/gring pixel_121/VDD pixel_121/GND pixel_121/VREF pixel_121/ROW_SEL
+ pixel_121/NB1 pixel_121/VBIAS pixel_121/NB2 pixel_121/AMP_IN pixel_121/SF_IB pixel_121/PIX_OUT
+ pixel_121/CSA_VREF pixel
Xpixel_110 pixel_110/gring pixel_110/VDD pixel_110/GND pixel_110/VREF pixel_110/ROW_SEL
+ pixel_110/NB1 pixel_110/VBIAS pixel_110/NB2 pixel_110/AMP_IN pixel_110/SF_IB pixel_110/PIX_OUT
+ pixel_110/CSA_VREF pixel
Xpixel_4104 pixel_4104/gring pixel_4104/VDD pixel_4104/GND pixel_4104/VREF pixel_4104/ROW_SEL
+ pixel_4104/NB1 pixel_4104/VBIAS pixel_4104/NB2 pixel_4104/AMP_IN pixel_4104/SF_IB
+ pixel_4104/PIX_OUT pixel_4104/CSA_VREF pixel
Xpixel_4115 pixel_4115/gring pixel_4115/VDD pixel_4115/GND pixel_4115/VREF pixel_4115/ROW_SEL
+ pixel_4115/NB1 pixel_4115/VBIAS pixel_4115/NB2 pixel_4115/AMP_IN pixel_4115/SF_IB
+ pixel_4115/PIX_OUT pixel_4115/CSA_VREF pixel
Xpixel_4126 pixel_4126/gring pixel_4126/VDD pixel_4126/GND pixel_4126/VREF pixel_4126/ROW_SEL
+ pixel_4126/NB1 pixel_4126/VBIAS pixel_4126/NB2 pixel_4126/AMP_IN pixel_4126/SF_IB
+ pixel_4126/PIX_OUT pixel_4126/CSA_VREF pixel
Xpixel_154 pixel_154/gring pixel_154/VDD pixel_154/GND pixel_154/VREF pixel_154/ROW_SEL
+ pixel_154/NB1 pixel_154/VBIAS pixel_154/NB2 pixel_154/AMP_IN pixel_154/SF_IB pixel_154/PIX_OUT
+ pixel_154/CSA_VREF pixel
Xpixel_143 pixel_143/gring pixel_143/VDD pixel_143/GND pixel_143/VREF pixel_143/ROW_SEL
+ pixel_143/NB1 pixel_143/VBIAS pixel_143/NB2 pixel_143/AMP_IN pixel_143/SF_IB pixel_143/PIX_OUT
+ pixel_143/CSA_VREF pixel
Xpixel_132 pixel_132/gring pixel_132/VDD pixel_132/GND pixel_132/VREF pixel_132/ROW_SEL
+ pixel_132/NB1 pixel_132/VBIAS pixel_132/NB2 pixel_132/AMP_IN pixel_132/SF_IB pixel_132/PIX_OUT
+ pixel_132/CSA_VREF pixel
Xpixel_3414 pixel_3414/gring pixel_3414/VDD pixel_3414/GND pixel_3414/VREF pixel_3414/ROW_SEL
+ pixel_3414/NB1 pixel_3414/VBIAS pixel_3414/NB2 pixel_3414/AMP_IN pixel_3414/SF_IB
+ pixel_3414/PIX_OUT pixel_3414/CSA_VREF pixel
Xpixel_3403 pixel_3403/gring pixel_3403/VDD pixel_3403/GND pixel_3403/VREF pixel_3403/ROW_SEL
+ pixel_3403/NB1 pixel_3403/VBIAS pixel_3403/NB2 pixel_3403/AMP_IN pixel_3403/SF_IB
+ pixel_3403/PIX_OUT pixel_3403/CSA_VREF pixel
Xpixel_4137 pixel_4137/gring pixel_4137/VDD pixel_4137/GND pixel_4137/VREF pixel_4137/ROW_SEL
+ pixel_4137/NB1 pixel_4137/VBIAS pixel_4137/NB2 pixel_4137/AMP_IN pixel_4137/SF_IB
+ pixel_4137/PIX_OUT pixel_4137/CSA_VREF pixel
Xpixel_4148 pixel_4148/gring pixel_4148/VDD pixel_4148/GND pixel_4148/VREF pixel_4148/ROW_SEL
+ pixel_4148/NB1 pixel_4148/VBIAS pixel_4148/NB2 pixel_4148/AMP_IN pixel_4148/SF_IB
+ pixel_4148/PIX_OUT pixel_4148/CSA_VREF pixel
Xpixel_4159 pixel_4159/gring pixel_4159/VDD pixel_4159/GND pixel_4159/VREF pixel_4159/ROW_SEL
+ pixel_4159/NB1 pixel_4159/VBIAS pixel_4159/NB2 pixel_4159/AMP_IN pixel_4159/SF_IB
+ pixel_4159/PIX_OUT pixel_4159/CSA_VREF pixel
Xpixel_198 pixel_198/gring pixel_198/VDD pixel_198/GND pixel_198/VREF pixel_198/ROW_SEL
+ pixel_198/NB1 pixel_198/VBIAS pixel_198/NB2 pixel_198/AMP_IN pixel_198/SF_IB pixel_198/PIX_OUT
+ pixel_198/CSA_VREF pixel
Xpixel_187 pixel_187/gring pixel_187/VDD pixel_187/GND pixel_187/VREF pixel_187/ROW_SEL
+ pixel_187/NB1 pixel_187/VBIAS pixel_187/NB2 pixel_187/AMP_IN pixel_187/SF_IB pixel_187/PIX_OUT
+ pixel_187/CSA_VREF pixel
Xpixel_176 pixel_176/gring pixel_176/VDD pixel_176/GND pixel_176/VREF pixel_176/ROW_SEL
+ pixel_176/NB1 pixel_176/VBIAS pixel_176/NB2 pixel_176/AMP_IN pixel_176/SF_IB pixel_176/PIX_OUT
+ pixel_176/CSA_VREF pixel
Xpixel_165 pixel_165/gring pixel_165/VDD pixel_165/GND pixel_165/VREF pixel_165/ROW_SEL
+ pixel_165/NB1 pixel_165/VBIAS pixel_165/NB2 pixel_165/AMP_IN pixel_165/SF_IB pixel_165/PIX_OUT
+ pixel_165/CSA_VREF pixel
Xpixel_2713 pixel_2713/gring pixel_2713/VDD pixel_2713/GND pixel_2713/VREF pixel_2713/ROW_SEL
+ pixel_2713/NB1 pixel_2713/VBIAS pixel_2713/NB2 pixel_2713/AMP_IN pixel_2713/SF_IB
+ pixel_2713/PIX_OUT pixel_2713/CSA_VREF pixel
Xpixel_2702 pixel_2702/gring pixel_2702/VDD pixel_2702/GND pixel_2702/VREF pixel_2702/ROW_SEL
+ pixel_2702/NB1 pixel_2702/VBIAS pixel_2702/NB2 pixel_2702/AMP_IN pixel_2702/SF_IB
+ pixel_2702/PIX_OUT pixel_2702/CSA_VREF pixel
Xpixel_3458 pixel_3458/gring pixel_3458/VDD pixel_3458/GND pixel_3458/VREF pixel_3458/ROW_SEL
+ pixel_3458/NB1 pixel_3458/VBIAS pixel_3458/NB2 pixel_3458/AMP_IN pixel_3458/SF_IB
+ pixel_3458/PIX_OUT pixel_3458/CSA_VREF pixel
Xpixel_3447 pixel_3447/gring pixel_3447/VDD pixel_3447/GND pixel_3447/VREF pixel_3447/ROW_SEL
+ pixel_3447/NB1 pixel_3447/VBIAS pixel_3447/NB2 pixel_3447/AMP_IN pixel_3447/SF_IB
+ pixel_3447/PIX_OUT pixel_3447/CSA_VREF pixel
Xpixel_3436 pixel_3436/gring pixel_3436/VDD pixel_3436/GND pixel_3436/VREF pixel_3436/ROW_SEL
+ pixel_3436/NB1 pixel_3436/VBIAS pixel_3436/NB2 pixel_3436/AMP_IN pixel_3436/SF_IB
+ pixel_3436/PIX_OUT pixel_3436/CSA_VREF pixel
Xpixel_3425 pixel_3425/gring pixel_3425/VDD pixel_3425/GND pixel_3425/VREF pixel_3425/ROW_SEL
+ pixel_3425/NB1 pixel_3425/VBIAS pixel_3425/NB2 pixel_3425/AMP_IN pixel_3425/SF_IB
+ pixel_3425/PIX_OUT pixel_3425/CSA_VREF pixel
Xpixel_2746 pixel_2746/gring pixel_2746/VDD pixel_2746/GND pixel_2746/VREF pixel_2746/ROW_SEL
+ pixel_2746/NB1 pixel_2746/VBIAS pixel_2746/NB2 pixel_2746/AMP_IN pixel_2746/SF_IB
+ pixel_2746/PIX_OUT pixel_2746/CSA_VREF pixel
Xpixel_2735 pixel_2735/gring pixel_2735/VDD pixel_2735/GND pixel_2735/VREF pixel_2735/ROW_SEL
+ pixel_2735/NB1 pixel_2735/VBIAS pixel_2735/NB2 pixel_2735/AMP_IN pixel_2735/SF_IB
+ pixel_2735/PIX_OUT pixel_2735/CSA_VREF pixel
Xpixel_2724 pixel_2724/gring pixel_2724/VDD pixel_2724/GND pixel_2724/VREF pixel_2724/ROW_SEL
+ pixel_2724/NB1 pixel_2724/VBIAS pixel_2724/NB2 pixel_2724/AMP_IN pixel_2724/SF_IB
+ pixel_2724/PIX_OUT pixel_2724/CSA_VREF pixel
Xpixel_3469 pixel_3469/gring pixel_3469/VDD pixel_3469/GND pixel_3469/VREF pixel_3469/ROW_SEL
+ pixel_3469/NB1 pixel_3469/VBIAS pixel_3469/NB2 pixel_3469/AMP_IN pixel_3469/SF_IB
+ pixel_3469/PIX_OUT pixel_3469/CSA_VREF pixel
Xpixel_2779 pixel_2779/gring pixel_2779/VDD pixel_2779/GND pixel_2779/VREF pixel_2779/ROW_SEL
+ pixel_2779/NB1 pixel_2779/VBIAS pixel_2779/NB2 pixel_2779/AMP_IN pixel_2779/SF_IB
+ pixel_2779/PIX_OUT pixel_2779/CSA_VREF pixel
Xpixel_2768 pixel_2768/gring pixel_2768/VDD pixel_2768/GND pixel_2768/VREF pixel_2768/ROW_SEL
+ pixel_2768/NB1 pixel_2768/VBIAS pixel_2768/NB2 pixel_2768/AMP_IN pixel_2768/SF_IB
+ pixel_2768/PIX_OUT pixel_2768/CSA_VREF pixel
Xpixel_2757 pixel_2757/gring pixel_2757/VDD pixel_2757/GND pixel_2757/VREF pixel_2757/ROW_SEL
+ pixel_2757/NB1 pixel_2757/VBIAS pixel_2757/NB2 pixel_2757/AMP_IN pixel_2757/SF_IB
+ pixel_2757/PIX_OUT pixel_2757/CSA_VREF pixel
Xpixel_6040 pixel_6040/gring pixel_6040/VDD pixel_6040/GND pixel_6040/VREF pixel_6040/ROW_SEL
+ pixel_6040/NB1 pixel_6040/VBIAS pixel_6040/NB2 pixel_6040/AMP_IN pixel_6040/SF_IB
+ pixel_6040/PIX_OUT pixel_6040/CSA_VREF pixel
Xpixel_6051 pixel_6051/gring pixel_6051/VDD pixel_6051/GND pixel_6051/VREF pixel_6051/ROW_SEL
+ pixel_6051/NB1 pixel_6051/VBIAS pixel_6051/NB2 pixel_6051/AMP_IN pixel_6051/SF_IB
+ pixel_6051/PIX_OUT pixel_6051/CSA_VREF pixel
Xpixel_6062 pixel_6062/gring pixel_6062/VDD pixel_6062/GND pixel_6062/VREF pixel_6062/ROW_SEL
+ pixel_6062/NB1 pixel_6062/VBIAS pixel_6062/NB2 pixel_6062/AMP_IN pixel_6062/SF_IB
+ pixel_6062/PIX_OUT pixel_6062/CSA_VREF pixel
Xpixel_6073 pixel_6073/gring pixel_6073/VDD pixel_6073/GND pixel_6073/VREF pixel_6073/ROW_SEL
+ pixel_6073/NB1 pixel_6073/VBIAS pixel_6073/NB2 pixel_6073/AMP_IN pixel_6073/SF_IB
+ pixel_6073/PIX_OUT pixel_6073/CSA_VREF pixel
Xpixel_6084 pixel_6084/gring pixel_6084/VDD pixel_6084/GND pixel_6084/VREF pixel_6084/ROW_SEL
+ pixel_6084/NB1 pixel_6084/VBIAS pixel_6084/NB2 pixel_6084/AMP_IN pixel_6084/SF_IB
+ pixel_6084/PIX_OUT pixel_6084/CSA_VREF pixel
Xpixel_6095 pixel_6095/gring pixel_6095/VDD pixel_6095/GND pixel_6095/VREF pixel_6095/ROW_SEL
+ pixel_6095/NB1 pixel_6095/VBIAS pixel_6095/NB2 pixel_6095/AMP_IN pixel_6095/SF_IB
+ pixel_6095/PIX_OUT pixel_6095/CSA_VREF pixel
Xpixel_5350 pixel_5350/gring pixel_5350/VDD pixel_5350/GND pixel_5350/VREF pixel_5350/ROW_SEL
+ pixel_5350/NB1 pixel_5350/VBIAS pixel_5350/NB2 pixel_5350/AMP_IN pixel_5350/SF_IB
+ pixel_5350/PIX_OUT pixel_5350/CSA_VREF pixel
Xpixel_5361 pixel_5361/gring pixel_5361/VDD pixel_5361/GND pixel_5361/VREF pixel_5361/ROW_SEL
+ pixel_5361/NB1 pixel_5361/VBIAS pixel_5361/NB2 pixel_5361/AMP_IN pixel_5361/SF_IB
+ pixel_5361/PIX_OUT pixel_5361/CSA_VREF pixel
Xpixel_5372 pixel_5372/gring pixel_5372/VDD pixel_5372/GND pixel_5372/VREF pixel_5372/ROW_SEL
+ pixel_5372/NB1 pixel_5372/VBIAS pixel_5372/NB2 pixel_5372/AMP_IN pixel_5372/SF_IB
+ pixel_5372/PIX_OUT pixel_5372/CSA_VREF pixel
Xpixel_5383 pixel_5383/gring pixel_5383/VDD pixel_5383/GND pixel_5383/VREF pixel_5383/ROW_SEL
+ pixel_5383/NB1 pixel_5383/VBIAS pixel_5383/NB2 pixel_5383/AMP_IN pixel_5383/SF_IB
+ pixel_5383/PIX_OUT pixel_5383/CSA_VREF pixel
Xpixel_5394 pixel_5394/gring pixel_5394/VDD pixel_5394/GND pixel_5394/VREF pixel_5394/ROW_SEL
+ pixel_5394/NB1 pixel_5394/VBIAS pixel_5394/NB2 pixel_5394/AMP_IN pixel_5394/SF_IB
+ pixel_5394/PIX_OUT pixel_5394/CSA_VREF pixel
Xpixel_4660 pixel_4660/gring pixel_4660/VDD pixel_4660/GND pixel_4660/VREF pixel_4660/ROW_SEL
+ pixel_4660/NB1 pixel_4660/VBIAS pixel_4660/NB2 pixel_4660/AMP_IN pixel_4660/SF_IB
+ pixel_4660/PIX_OUT pixel_4660/CSA_VREF pixel
Xpixel_4671 pixel_4671/gring pixel_4671/VDD pixel_4671/GND pixel_4671/VREF pixel_4671/ROW_SEL
+ pixel_4671/NB1 pixel_4671/VBIAS pixel_4671/NB2 pixel_4671/AMP_IN pixel_4671/SF_IB
+ pixel_4671/PIX_OUT pixel_4671/CSA_VREF pixel
Xpixel_4682 pixel_4682/gring pixel_4682/VDD pixel_4682/GND pixel_4682/VREF pixel_4682/ROW_SEL
+ pixel_4682/NB1 pixel_4682/VBIAS pixel_4682/NB2 pixel_4682/AMP_IN pixel_4682/SF_IB
+ pixel_4682/PIX_OUT pixel_4682/CSA_VREF pixel
Xpixel_4693 pixel_4693/gring pixel_4693/VDD pixel_4693/GND pixel_4693/VREF pixel_4693/ROW_SEL
+ pixel_4693/NB1 pixel_4693/VBIAS pixel_4693/NB2 pixel_4693/AMP_IN pixel_4693/SF_IB
+ pixel_4693/PIX_OUT pixel_4693/CSA_VREF pixel
Xpixel_3970 pixel_3970/gring pixel_3970/VDD pixel_3970/GND pixel_3970/VREF pixel_3970/ROW_SEL
+ pixel_3970/NB1 pixel_3970/VBIAS pixel_3970/NB2 pixel_3970/AMP_IN pixel_3970/SF_IB
+ pixel_3970/PIX_OUT pixel_3970/CSA_VREF pixel
Xpixel_3981 pixel_3981/gring pixel_3981/VDD pixel_3981/GND pixel_3981/VREF pixel_3981/ROW_SEL
+ pixel_3981/NB1 pixel_3981/VBIAS pixel_3981/NB2 pixel_3981/AMP_IN pixel_3981/SF_IB
+ pixel_3981/PIX_OUT pixel_3981/CSA_VREF pixel
Xpixel_3992 pixel_3992/gring pixel_3992/VDD pixel_3992/GND pixel_3992/VREF pixel_3992/ROW_SEL
+ pixel_3992/NB1 pixel_3992/VBIAS pixel_3992/NB2 pixel_3992/AMP_IN pixel_3992/SF_IB
+ pixel_3992/PIX_OUT pixel_3992/CSA_VREF pixel
Xpixel_2 pixel_2/gring pixel_2/VDD pixel_2/GND pixel_2/VREF pixel_2/ROW_SEL pixel_2/NB1
+ pixel_2/VBIAS pixel_2/NB2 pixel_2/AMP_IN pixel_2/SF_IB pixel_2/PIX_OUT pixel_2/CSA_VREF
+ pixel
Xpixel_2009 pixel_2009/gring pixel_2009/VDD pixel_2009/GND pixel_2009/VREF pixel_2009/ROW_SEL
+ pixel_2009/NB1 pixel_2009/VBIAS pixel_2009/NB2 pixel_2009/AMP_IN pixel_2009/SF_IB
+ pixel_2009/PIX_OUT pixel_2009/CSA_VREF pixel
Xpixel_1319 pixel_1319/gring pixel_1319/VDD pixel_1319/GND pixel_1319/VREF pixel_1319/ROW_SEL
+ pixel_1319/NB1 pixel_1319/VBIAS pixel_1319/NB2 pixel_1319/AMP_IN pixel_1319/SF_IB
+ pixel_1319/PIX_OUT pixel_1319/CSA_VREF pixel
Xpixel_1308 pixel_1308/gring pixel_1308/VDD pixel_1308/GND pixel_1308/VREF pixel_1308/ROW_SEL
+ pixel_1308/NB1 pixel_1308/VBIAS pixel_1308/NB2 pixel_1308/AMP_IN pixel_1308/SF_IB
+ pixel_1308/PIX_OUT pixel_1308/CSA_VREF pixel
Xpixel_9605 pixel_9605/gring pixel_9605/VDD pixel_9605/GND pixel_9605/VREF pixel_9605/ROW_SEL
+ pixel_9605/NB1 pixel_9605/VBIAS pixel_9605/NB2 pixel_9605/AMP_IN pixel_9605/SF_IB
+ pixel_9605/PIX_OUT pixel_9605/CSA_VREF pixel
Xpixel_9616 pixel_9616/gring pixel_9616/VDD pixel_9616/GND pixel_9616/VREF pixel_9616/ROW_SEL
+ pixel_9616/NB1 pixel_9616/VBIAS pixel_9616/NB2 pixel_9616/AMP_IN pixel_9616/SF_IB
+ pixel_9616/PIX_OUT pixel_9616/CSA_VREF pixel
Xpixel_9627 pixel_9627/gring pixel_9627/VDD pixel_9627/GND pixel_9627/VREF pixel_9627/ROW_SEL
+ pixel_9627/NB1 pixel_9627/VBIAS pixel_9627/NB2 pixel_9627/AMP_IN pixel_9627/SF_IB
+ pixel_9627/PIX_OUT pixel_9627/CSA_VREF pixel
Xpixel_9638 pixel_9638/gring pixel_9638/VDD pixel_9638/GND pixel_9638/VREF pixel_9638/ROW_SEL
+ pixel_9638/NB1 pixel_9638/VBIAS pixel_9638/NB2 pixel_9638/AMP_IN pixel_9638/SF_IB
+ pixel_9638/PIX_OUT pixel_9638/CSA_VREF pixel
Xpixel_8937 pixel_8937/gring pixel_8937/VDD pixel_8937/GND pixel_8937/VREF pixel_8937/ROW_SEL
+ pixel_8937/NB1 pixel_8937/VBIAS pixel_8937/NB2 pixel_8937/AMP_IN pixel_8937/SF_IB
+ pixel_8937/PIX_OUT pixel_8937/CSA_VREF pixel
Xpixel_8926 pixel_8926/gring pixel_8926/VDD pixel_8926/GND pixel_8926/VREF pixel_8926/ROW_SEL
+ pixel_8926/NB1 pixel_8926/VBIAS pixel_8926/NB2 pixel_8926/AMP_IN pixel_8926/SF_IB
+ pixel_8926/PIX_OUT pixel_8926/CSA_VREF pixel
Xpixel_8915 pixel_8915/gring pixel_8915/VDD pixel_8915/GND pixel_8915/VREF pixel_8915/ROW_SEL
+ pixel_8915/NB1 pixel_8915/VBIAS pixel_8915/NB2 pixel_8915/AMP_IN pixel_8915/SF_IB
+ pixel_8915/PIX_OUT pixel_8915/CSA_VREF pixel
Xpixel_8904 pixel_8904/gring pixel_8904/VDD pixel_8904/GND pixel_8904/VREF pixel_8904/ROW_SEL
+ pixel_8904/NB1 pixel_8904/VBIAS pixel_8904/NB2 pixel_8904/AMP_IN pixel_8904/SF_IB
+ pixel_8904/PIX_OUT pixel_8904/CSA_VREF pixel
Xpixel_9649 pixel_9649/gring pixel_9649/VDD pixel_9649/GND pixel_9649/VREF pixel_9649/ROW_SEL
+ pixel_9649/NB1 pixel_9649/VBIAS pixel_9649/NB2 pixel_9649/AMP_IN pixel_9649/SF_IB
+ pixel_9649/PIX_OUT pixel_9649/CSA_VREF pixel
Xpixel_8959 pixel_8959/gring pixel_8959/VDD pixel_8959/GND pixel_8959/VREF pixel_8959/ROW_SEL
+ pixel_8959/NB1 pixel_8959/VBIAS pixel_8959/NB2 pixel_8959/AMP_IN pixel_8959/SF_IB
+ pixel_8959/PIX_OUT pixel_8959/CSA_VREF pixel
Xpixel_8948 pixel_8948/gring pixel_8948/VDD pixel_8948/GND pixel_8948/VREF pixel_8948/ROW_SEL
+ pixel_8948/NB1 pixel_8948/VBIAS pixel_8948/NB2 pixel_8948/AMP_IN pixel_8948/SF_IB
+ pixel_8948/PIX_OUT pixel_8948/CSA_VREF pixel
Xpixel_3233 pixel_3233/gring pixel_3233/VDD pixel_3233/GND pixel_3233/VREF pixel_3233/ROW_SEL
+ pixel_3233/NB1 pixel_3233/VBIAS pixel_3233/NB2 pixel_3233/AMP_IN pixel_3233/SF_IB
+ pixel_3233/PIX_OUT pixel_3233/CSA_VREF pixel
Xpixel_3222 pixel_3222/gring pixel_3222/VDD pixel_3222/GND pixel_3222/VREF pixel_3222/ROW_SEL
+ pixel_3222/NB1 pixel_3222/VBIAS pixel_3222/NB2 pixel_3222/AMP_IN pixel_3222/SF_IB
+ pixel_3222/PIX_OUT pixel_3222/CSA_VREF pixel
Xpixel_3211 pixel_3211/gring pixel_3211/VDD pixel_3211/GND pixel_3211/VREF pixel_3211/ROW_SEL
+ pixel_3211/NB1 pixel_3211/VBIAS pixel_3211/NB2 pixel_3211/AMP_IN pixel_3211/SF_IB
+ pixel_3211/PIX_OUT pixel_3211/CSA_VREF pixel
Xpixel_3200 pixel_3200/gring pixel_3200/VDD pixel_3200/GND pixel_3200/VREF pixel_3200/ROW_SEL
+ pixel_3200/NB1 pixel_3200/VBIAS pixel_3200/NB2 pixel_3200/AMP_IN pixel_3200/SF_IB
+ pixel_3200/PIX_OUT pixel_3200/CSA_VREF pixel
Xpixel_2521 pixel_2521/gring pixel_2521/VDD pixel_2521/GND pixel_2521/VREF pixel_2521/ROW_SEL
+ pixel_2521/NB1 pixel_2521/VBIAS pixel_2521/NB2 pixel_2521/AMP_IN pixel_2521/SF_IB
+ pixel_2521/PIX_OUT pixel_2521/CSA_VREF pixel
Xpixel_2510 pixel_2510/gring pixel_2510/VDD pixel_2510/GND pixel_2510/VREF pixel_2510/ROW_SEL
+ pixel_2510/NB1 pixel_2510/VBIAS pixel_2510/NB2 pixel_2510/AMP_IN pixel_2510/SF_IB
+ pixel_2510/PIX_OUT pixel_2510/CSA_VREF pixel
Xpixel_3266 pixel_3266/gring pixel_3266/VDD pixel_3266/GND pixel_3266/VREF pixel_3266/ROW_SEL
+ pixel_3266/NB1 pixel_3266/VBIAS pixel_3266/NB2 pixel_3266/AMP_IN pixel_3266/SF_IB
+ pixel_3266/PIX_OUT pixel_3266/CSA_VREF pixel
Xpixel_3255 pixel_3255/gring pixel_3255/VDD pixel_3255/GND pixel_3255/VREF pixel_3255/ROW_SEL
+ pixel_3255/NB1 pixel_3255/VBIAS pixel_3255/NB2 pixel_3255/AMP_IN pixel_3255/SF_IB
+ pixel_3255/PIX_OUT pixel_3255/CSA_VREF pixel
Xpixel_3244 pixel_3244/gring pixel_3244/VDD pixel_3244/GND pixel_3244/VREF pixel_3244/ROW_SEL
+ pixel_3244/NB1 pixel_3244/VBIAS pixel_3244/NB2 pixel_3244/AMP_IN pixel_3244/SF_IB
+ pixel_3244/PIX_OUT pixel_3244/CSA_VREF pixel
Xpixel_2554 pixel_2554/gring pixel_2554/VDD pixel_2554/GND pixel_2554/VREF pixel_2554/ROW_SEL
+ pixel_2554/NB1 pixel_2554/VBIAS pixel_2554/NB2 pixel_2554/AMP_IN pixel_2554/SF_IB
+ pixel_2554/PIX_OUT pixel_2554/CSA_VREF pixel
Xpixel_2543 pixel_2543/gring pixel_2543/VDD pixel_2543/GND pixel_2543/VREF pixel_2543/ROW_SEL
+ pixel_2543/NB1 pixel_2543/VBIAS pixel_2543/NB2 pixel_2543/AMP_IN pixel_2543/SF_IB
+ pixel_2543/PIX_OUT pixel_2543/CSA_VREF pixel
Xpixel_2532 pixel_2532/gring pixel_2532/VDD pixel_2532/GND pixel_2532/VREF pixel_2532/ROW_SEL
+ pixel_2532/NB1 pixel_2532/VBIAS pixel_2532/NB2 pixel_2532/AMP_IN pixel_2532/SF_IB
+ pixel_2532/PIX_OUT pixel_2532/CSA_VREF pixel
Xpixel_3299 pixel_3299/gring pixel_3299/VDD pixel_3299/GND pixel_3299/VREF pixel_3299/ROW_SEL
+ pixel_3299/NB1 pixel_3299/VBIAS pixel_3299/NB2 pixel_3299/AMP_IN pixel_3299/SF_IB
+ pixel_3299/PIX_OUT pixel_3299/CSA_VREF pixel
Xpixel_3288 pixel_3288/gring pixel_3288/VDD pixel_3288/GND pixel_3288/VREF pixel_3288/ROW_SEL
+ pixel_3288/NB1 pixel_3288/VBIAS pixel_3288/NB2 pixel_3288/AMP_IN pixel_3288/SF_IB
+ pixel_3288/PIX_OUT pixel_3288/CSA_VREF pixel
Xpixel_3277 pixel_3277/gring pixel_3277/VDD pixel_3277/GND pixel_3277/VREF pixel_3277/ROW_SEL
+ pixel_3277/NB1 pixel_3277/VBIAS pixel_3277/NB2 pixel_3277/AMP_IN pixel_3277/SF_IB
+ pixel_3277/PIX_OUT pixel_3277/CSA_VREF pixel
Xpixel_1853 pixel_1853/gring pixel_1853/VDD pixel_1853/GND pixel_1853/VREF pixel_1853/ROW_SEL
+ pixel_1853/NB1 pixel_1853/VBIAS pixel_1853/NB2 pixel_1853/AMP_IN pixel_1853/SF_IB
+ pixel_1853/PIX_OUT pixel_1853/CSA_VREF pixel
Xpixel_1842 pixel_1842/gring pixel_1842/VDD pixel_1842/GND pixel_1842/VREF pixel_1842/ROW_SEL
+ pixel_1842/NB1 pixel_1842/VBIAS pixel_1842/NB2 pixel_1842/AMP_IN pixel_1842/SF_IB
+ pixel_1842/PIX_OUT pixel_1842/CSA_VREF pixel
Xpixel_1831 pixel_1831/gring pixel_1831/VDD pixel_1831/GND pixel_1831/VREF pixel_1831/ROW_SEL
+ pixel_1831/NB1 pixel_1831/VBIAS pixel_1831/NB2 pixel_1831/AMP_IN pixel_1831/SF_IB
+ pixel_1831/PIX_OUT pixel_1831/CSA_VREF pixel
Xpixel_1820 pixel_1820/gring pixel_1820/VDD pixel_1820/GND pixel_1820/VREF pixel_1820/ROW_SEL
+ pixel_1820/NB1 pixel_1820/VBIAS pixel_1820/NB2 pixel_1820/AMP_IN pixel_1820/SF_IB
+ pixel_1820/PIX_OUT pixel_1820/CSA_VREF pixel
Xpixel_2598 pixel_2598/gring pixel_2598/VDD pixel_2598/GND pixel_2598/VREF pixel_2598/ROW_SEL
+ pixel_2598/NB1 pixel_2598/VBIAS pixel_2598/NB2 pixel_2598/AMP_IN pixel_2598/SF_IB
+ pixel_2598/PIX_OUT pixel_2598/CSA_VREF pixel
Xpixel_2587 pixel_2587/gring pixel_2587/VDD pixel_2587/GND pixel_2587/VREF pixel_2587/ROW_SEL
+ pixel_2587/NB1 pixel_2587/VBIAS pixel_2587/NB2 pixel_2587/AMP_IN pixel_2587/SF_IB
+ pixel_2587/PIX_OUT pixel_2587/CSA_VREF pixel
Xpixel_2576 pixel_2576/gring pixel_2576/VDD pixel_2576/GND pixel_2576/VREF pixel_2576/ROW_SEL
+ pixel_2576/NB1 pixel_2576/VBIAS pixel_2576/NB2 pixel_2576/AMP_IN pixel_2576/SF_IB
+ pixel_2576/PIX_OUT pixel_2576/CSA_VREF pixel
Xpixel_2565 pixel_2565/gring pixel_2565/VDD pixel_2565/GND pixel_2565/VREF pixel_2565/ROW_SEL
+ pixel_2565/NB1 pixel_2565/VBIAS pixel_2565/NB2 pixel_2565/AMP_IN pixel_2565/SF_IB
+ pixel_2565/PIX_OUT pixel_2565/CSA_VREF pixel
Xpixel_1886 pixel_1886/gring pixel_1886/VDD pixel_1886/GND pixel_1886/VREF pixel_1886/ROW_SEL
+ pixel_1886/NB1 pixel_1886/VBIAS pixel_1886/NB2 pixel_1886/AMP_IN pixel_1886/SF_IB
+ pixel_1886/PIX_OUT pixel_1886/CSA_VREF pixel
Xpixel_1875 pixel_1875/gring pixel_1875/VDD pixel_1875/GND pixel_1875/VREF pixel_1875/ROW_SEL
+ pixel_1875/NB1 pixel_1875/VBIAS pixel_1875/NB2 pixel_1875/AMP_IN pixel_1875/SF_IB
+ pixel_1875/PIX_OUT pixel_1875/CSA_VREF pixel
Xpixel_1864 pixel_1864/gring pixel_1864/VDD pixel_1864/GND pixel_1864/VREF pixel_1864/ROW_SEL
+ pixel_1864/NB1 pixel_1864/VBIAS pixel_1864/NB2 pixel_1864/AMP_IN pixel_1864/SF_IB
+ pixel_1864/PIX_OUT pixel_1864/CSA_VREF pixel
Xpixel_1897 pixel_1897/gring pixel_1897/VDD pixel_1897/GND pixel_1897/VREF pixel_1897/ROW_SEL
+ pixel_1897/NB1 pixel_1897/VBIAS pixel_1897/NB2 pixel_1897/AMP_IN pixel_1897/SF_IB
+ pixel_1897/PIX_OUT pixel_1897/CSA_VREF pixel
Xpixel_5180 pixel_5180/gring pixel_5180/VDD pixel_5180/GND pixel_5180/VREF pixel_5180/ROW_SEL
+ pixel_5180/NB1 pixel_5180/VBIAS pixel_5180/NB2 pixel_5180/AMP_IN pixel_5180/SF_IB
+ pixel_5180/PIX_OUT pixel_5180/CSA_VREF pixel
Xpixel_5191 pixel_5191/gring pixel_5191/VDD pixel_5191/GND pixel_5191/VREF pixel_5191/ROW_SEL
+ pixel_5191/NB1 pixel_5191/VBIAS pixel_5191/NB2 pixel_5191/AMP_IN pixel_5191/SF_IB
+ pixel_5191/PIX_OUT pixel_5191/CSA_VREF pixel
Xpixel_4490 pixel_4490/gring pixel_4490/VDD pixel_4490/GND pixel_4490/VREF pixel_4490/ROW_SEL
+ pixel_4490/NB1 pixel_4490/VBIAS pixel_4490/NB2 pixel_4490/AMP_IN pixel_4490/SF_IB
+ pixel_4490/PIX_OUT pixel_4490/CSA_VREF pixel
Xpixel_6809 pixel_6809/gring pixel_6809/VDD pixel_6809/GND pixel_6809/VREF pixel_6809/ROW_SEL
+ pixel_6809/NB1 pixel_6809/VBIAS pixel_6809/NB2 pixel_6809/AMP_IN pixel_6809/SF_IB
+ pixel_6809/PIX_OUT pixel_6809/CSA_VREF pixel
Xpixel_1105 pixel_1105/gring pixel_1105/VDD pixel_1105/GND pixel_1105/VREF pixel_1105/ROW_SEL
+ pixel_1105/NB1 pixel_1105/VBIAS pixel_1105/NB2 pixel_1105/AMP_IN pixel_1105/SF_IB
+ pixel_1105/PIX_OUT pixel_1105/CSA_VREF pixel
Xpixel_1138 pixel_1138/gring pixel_1138/VDD pixel_1138/GND pixel_1138/VREF pixel_1138/ROW_SEL
+ pixel_1138/NB1 pixel_1138/VBIAS pixel_1138/NB2 pixel_1138/AMP_IN pixel_1138/SF_IB
+ pixel_1138/PIX_OUT pixel_1138/CSA_VREF pixel
Xpixel_1127 pixel_1127/gring pixel_1127/VDD pixel_1127/GND pixel_1127/VREF pixel_1127/ROW_SEL
+ pixel_1127/NB1 pixel_1127/VBIAS pixel_1127/NB2 pixel_1127/AMP_IN pixel_1127/SF_IB
+ pixel_1127/PIX_OUT pixel_1127/CSA_VREF pixel
Xpixel_1116 pixel_1116/gring pixel_1116/VDD pixel_1116/GND pixel_1116/VREF pixel_1116/ROW_SEL
+ pixel_1116/NB1 pixel_1116/VBIAS pixel_1116/NB2 pixel_1116/AMP_IN pixel_1116/SF_IB
+ pixel_1116/PIX_OUT pixel_1116/CSA_VREF pixel
Xpixel_1149 pixel_1149/gring pixel_1149/VDD pixel_1149/GND pixel_1149/VREF pixel_1149/ROW_SEL
+ pixel_1149/NB1 pixel_1149/VBIAS pixel_1149/NB2 pixel_1149/AMP_IN pixel_1149/SF_IB
+ pixel_1149/PIX_OUT pixel_1149/CSA_VREF pixel
Xpixel_9413 pixel_9413/gring pixel_9413/VDD pixel_9413/GND pixel_9413/VREF pixel_9413/ROW_SEL
+ pixel_9413/NB1 pixel_9413/VBIAS pixel_9413/NB2 pixel_9413/AMP_IN pixel_9413/SF_IB
+ pixel_9413/PIX_OUT pixel_9413/CSA_VREF pixel
Xpixel_9402 pixel_9402/gring pixel_9402/VDD pixel_9402/GND pixel_9402/VREF pixel_9402/ROW_SEL
+ pixel_9402/NB1 pixel_9402/VBIAS pixel_9402/NB2 pixel_9402/AMP_IN pixel_9402/SF_IB
+ pixel_9402/PIX_OUT pixel_9402/CSA_VREF pixel
Xpixel_8712 pixel_8712/gring pixel_8712/VDD pixel_8712/GND pixel_8712/VREF pixel_8712/ROW_SEL
+ pixel_8712/NB1 pixel_8712/VBIAS pixel_8712/NB2 pixel_8712/AMP_IN pixel_8712/SF_IB
+ pixel_8712/PIX_OUT pixel_8712/CSA_VREF pixel
Xpixel_8701 pixel_8701/gring pixel_8701/VDD pixel_8701/GND pixel_8701/VREF pixel_8701/ROW_SEL
+ pixel_8701/NB1 pixel_8701/VBIAS pixel_8701/NB2 pixel_8701/AMP_IN pixel_8701/SF_IB
+ pixel_8701/PIX_OUT pixel_8701/CSA_VREF pixel
Xpixel_9446 pixel_9446/gring pixel_9446/VDD pixel_9446/GND pixel_9446/VREF pixel_9446/ROW_SEL
+ pixel_9446/NB1 pixel_9446/VBIAS pixel_9446/NB2 pixel_9446/AMP_IN pixel_9446/SF_IB
+ pixel_9446/PIX_OUT pixel_9446/CSA_VREF pixel
Xpixel_9435 pixel_9435/gring pixel_9435/VDD pixel_9435/GND pixel_9435/VREF pixel_9435/ROW_SEL
+ pixel_9435/NB1 pixel_9435/VBIAS pixel_9435/NB2 pixel_9435/AMP_IN pixel_9435/SF_IB
+ pixel_9435/PIX_OUT pixel_9435/CSA_VREF pixel
Xpixel_9424 pixel_9424/gring pixel_9424/VDD pixel_9424/GND pixel_9424/VREF pixel_9424/ROW_SEL
+ pixel_9424/NB1 pixel_9424/VBIAS pixel_9424/NB2 pixel_9424/AMP_IN pixel_9424/SF_IB
+ pixel_9424/PIX_OUT pixel_9424/CSA_VREF pixel
Xpixel_8745 pixel_8745/gring pixel_8745/VDD pixel_8745/GND pixel_8745/VREF pixel_8745/ROW_SEL
+ pixel_8745/NB1 pixel_8745/VBIAS pixel_8745/NB2 pixel_8745/AMP_IN pixel_8745/SF_IB
+ pixel_8745/PIX_OUT pixel_8745/CSA_VREF pixel
Xpixel_8734 pixel_8734/gring pixel_8734/VDD pixel_8734/GND pixel_8734/VREF pixel_8734/ROW_SEL
+ pixel_8734/NB1 pixel_8734/VBIAS pixel_8734/NB2 pixel_8734/AMP_IN pixel_8734/SF_IB
+ pixel_8734/PIX_OUT pixel_8734/CSA_VREF pixel
Xpixel_8723 pixel_8723/gring pixel_8723/VDD pixel_8723/GND pixel_8723/VREF pixel_8723/ROW_SEL
+ pixel_8723/NB1 pixel_8723/VBIAS pixel_8723/NB2 pixel_8723/AMP_IN pixel_8723/SF_IB
+ pixel_8723/PIX_OUT pixel_8723/CSA_VREF pixel
Xpixel_9479 pixel_9479/gring pixel_9479/VDD pixel_9479/GND pixel_9479/VREF pixel_9479/ROW_SEL
+ pixel_9479/NB1 pixel_9479/VBIAS pixel_9479/NB2 pixel_9479/AMP_IN pixel_9479/SF_IB
+ pixel_9479/PIX_OUT pixel_9479/CSA_VREF pixel
Xpixel_9468 pixel_9468/gring pixel_9468/VDD pixel_9468/GND pixel_9468/VREF pixel_9468/ROW_SEL
+ pixel_9468/NB1 pixel_9468/VBIAS pixel_9468/NB2 pixel_9468/AMP_IN pixel_9468/SF_IB
+ pixel_9468/PIX_OUT pixel_9468/CSA_VREF pixel
Xpixel_9457 pixel_9457/gring pixel_9457/VDD pixel_9457/GND pixel_9457/VREF pixel_9457/ROW_SEL
+ pixel_9457/NB1 pixel_9457/VBIAS pixel_9457/NB2 pixel_9457/AMP_IN pixel_9457/SF_IB
+ pixel_9457/PIX_OUT pixel_9457/CSA_VREF pixel
Xpixel_8778 pixel_8778/gring pixel_8778/VDD pixel_8778/GND pixel_8778/VREF pixel_8778/ROW_SEL
+ pixel_8778/NB1 pixel_8778/VBIAS pixel_8778/NB2 pixel_8778/AMP_IN pixel_8778/SF_IB
+ pixel_8778/PIX_OUT pixel_8778/CSA_VREF pixel
Xpixel_8767 pixel_8767/gring pixel_8767/VDD pixel_8767/GND pixel_8767/VREF pixel_8767/ROW_SEL
+ pixel_8767/NB1 pixel_8767/VBIAS pixel_8767/NB2 pixel_8767/AMP_IN pixel_8767/SF_IB
+ pixel_8767/PIX_OUT pixel_8767/CSA_VREF pixel
Xpixel_8756 pixel_8756/gring pixel_8756/VDD pixel_8756/GND pixel_8756/VREF pixel_8756/ROW_SEL
+ pixel_8756/NB1 pixel_8756/VBIAS pixel_8756/NB2 pixel_8756/AMP_IN pixel_8756/SF_IB
+ pixel_8756/PIX_OUT pixel_8756/CSA_VREF pixel
Xpixel_8789 pixel_8789/gring pixel_8789/VDD pixel_8789/GND pixel_8789/VREF pixel_8789/ROW_SEL
+ pixel_8789/NB1 pixel_8789/VBIAS pixel_8789/NB2 pixel_8789/AMP_IN pixel_8789/SF_IB
+ pixel_8789/PIX_OUT pixel_8789/CSA_VREF pixel
Xpixel_3041 pixel_3041/gring pixel_3041/VDD pixel_3041/GND pixel_3041/VREF pixel_3041/ROW_SEL
+ pixel_3041/NB1 pixel_3041/VBIAS pixel_3041/NB2 pixel_3041/AMP_IN pixel_3041/SF_IB
+ pixel_3041/PIX_OUT pixel_3041/CSA_VREF pixel
Xpixel_3030 pixel_3030/gring pixel_3030/VDD pixel_3030/GND pixel_3030/VREF pixel_3030/ROW_SEL
+ pixel_3030/NB1 pixel_3030/VBIAS pixel_3030/NB2 pixel_3030/AMP_IN pixel_3030/SF_IB
+ pixel_3030/PIX_OUT pixel_3030/CSA_VREF pixel
Xpixel_3074 pixel_3074/gring pixel_3074/VDD pixel_3074/GND pixel_3074/VREF pixel_3074/ROW_SEL
+ pixel_3074/NB1 pixel_3074/VBIAS pixel_3074/NB2 pixel_3074/AMP_IN pixel_3074/SF_IB
+ pixel_3074/PIX_OUT pixel_3074/CSA_VREF pixel
Xpixel_3063 pixel_3063/gring pixel_3063/VDD pixel_3063/GND pixel_3063/VREF pixel_3063/ROW_SEL
+ pixel_3063/NB1 pixel_3063/VBIAS pixel_3063/NB2 pixel_3063/AMP_IN pixel_3063/SF_IB
+ pixel_3063/PIX_OUT pixel_3063/CSA_VREF pixel
Xpixel_3052 pixel_3052/gring pixel_3052/VDD pixel_3052/GND pixel_3052/VREF pixel_3052/ROW_SEL
+ pixel_3052/NB1 pixel_3052/VBIAS pixel_3052/NB2 pixel_3052/AMP_IN pixel_3052/SF_IB
+ pixel_3052/PIX_OUT pixel_3052/CSA_VREF pixel
Xpixel_2373 pixel_2373/gring pixel_2373/VDD pixel_2373/GND pixel_2373/VREF pixel_2373/ROW_SEL
+ pixel_2373/NB1 pixel_2373/VBIAS pixel_2373/NB2 pixel_2373/AMP_IN pixel_2373/SF_IB
+ pixel_2373/PIX_OUT pixel_2373/CSA_VREF pixel
Xpixel_2362 pixel_2362/gring pixel_2362/VDD pixel_2362/GND pixel_2362/VREF pixel_2362/ROW_SEL
+ pixel_2362/NB1 pixel_2362/VBIAS pixel_2362/NB2 pixel_2362/AMP_IN pixel_2362/SF_IB
+ pixel_2362/PIX_OUT pixel_2362/CSA_VREF pixel
Xpixel_2351 pixel_2351/gring pixel_2351/VDD pixel_2351/GND pixel_2351/VREF pixel_2351/ROW_SEL
+ pixel_2351/NB1 pixel_2351/VBIAS pixel_2351/NB2 pixel_2351/AMP_IN pixel_2351/SF_IB
+ pixel_2351/PIX_OUT pixel_2351/CSA_VREF pixel
Xpixel_2340 pixel_2340/gring pixel_2340/VDD pixel_2340/GND pixel_2340/VREF pixel_2340/ROW_SEL
+ pixel_2340/NB1 pixel_2340/VBIAS pixel_2340/NB2 pixel_2340/AMP_IN pixel_2340/SF_IB
+ pixel_2340/PIX_OUT pixel_2340/CSA_VREF pixel
Xpixel_3096 pixel_3096/gring pixel_3096/VDD pixel_3096/GND pixel_3096/VREF pixel_3096/ROW_SEL
+ pixel_3096/NB1 pixel_3096/VBIAS pixel_3096/NB2 pixel_3096/AMP_IN pixel_3096/SF_IB
+ pixel_3096/PIX_OUT pixel_3096/CSA_VREF pixel
Xpixel_3085 pixel_3085/gring pixel_3085/VDD pixel_3085/GND pixel_3085/VREF pixel_3085/ROW_SEL
+ pixel_3085/NB1 pixel_3085/VBIAS pixel_3085/NB2 pixel_3085/AMP_IN pixel_3085/SF_IB
+ pixel_3085/PIX_OUT pixel_3085/CSA_VREF pixel
Xpixel_1661 pixel_1661/gring pixel_1661/VDD pixel_1661/GND pixel_1661/VREF pixel_1661/ROW_SEL
+ pixel_1661/NB1 pixel_1661/VBIAS pixel_1661/NB2 pixel_1661/AMP_IN pixel_1661/SF_IB
+ pixel_1661/PIX_OUT pixel_1661/CSA_VREF pixel
Xpixel_1650 pixel_1650/gring pixel_1650/VDD pixel_1650/GND pixel_1650/VREF pixel_1650/ROW_SEL
+ pixel_1650/NB1 pixel_1650/VBIAS pixel_1650/NB2 pixel_1650/AMP_IN pixel_1650/SF_IB
+ pixel_1650/PIX_OUT pixel_1650/CSA_VREF pixel
Xpixel_2395 pixel_2395/gring pixel_2395/VDD pixel_2395/GND pixel_2395/VREF pixel_2395/ROW_SEL
+ pixel_2395/NB1 pixel_2395/VBIAS pixel_2395/NB2 pixel_2395/AMP_IN pixel_2395/SF_IB
+ pixel_2395/PIX_OUT pixel_2395/CSA_VREF pixel
Xpixel_2384 pixel_2384/gring pixel_2384/VDD pixel_2384/GND pixel_2384/VREF pixel_2384/ROW_SEL
+ pixel_2384/NB1 pixel_2384/VBIAS pixel_2384/NB2 pixel_2384/AMP_IN pixel_2384/SF_IB
+ pixel_2384/PIX_OUT pixel_2384/CSA_VREF pixel
Xpixel_1694 pixel_1694/gring pixel_1694/VDD pixel_1694/GND pixel_1694/VREF pixel_1694/ROW_SEL
+ pixel_1694/NB1 pixel_1694/VBIAS pixel_1694/NB2 pixel_1694/AMP_IN pixel_1694/SF_IB
+ pixel_1694/PIX_OUT pixel_1694/CSA_VREF pixel
Xpixel_1683 pixel_1683/gring pixel_1683/VDD pixel_1683/GND pixel_1683/VREF pixel_1683/ROW_SEL
+ pixel_1683/NB1 pixel_1683/VBIAS pixel_1683/NB2 pixel_1683/AMP_IN pixel_1683/SF_IB
+ pixel_1683/PIX_OUT pixel_1683/CSA_VREF pixel
Xpixel_1672 pixel_1672/gring pixel_1672/VDD pixel_1672/GND pixel_1672/VREF pixel_1672/ROW_SEL
+ pixel_1672/NB1 pixel_1672/VBIAS pixel_1672/NB2 pixel_1672/AMP_IN pixel_1672/SF_IB
+ pixel_1672/PIX_OUT pixel_1672/CSA_VREF pixel
Xpixel_9980 pixel_9980/gring pixel_9980/VDD pixel_9980/GND pixel_9980/VREF pixel_9980/ROW_SEL
+ pixel_9980/NB1 pixel_9980/VBIAS pixel_9980/NB2 pixel_9980/AMP_IN pixel_9980/SF_IB
+ pixel_9980/PIX_OUT pixel_9980/CSA_VREF pixel
Xpixel_9991 pixel_9991/gring pixel_9991/VDD pixel_9991/GND pixel_9991/VREF pixel_9991/ROW_SEL
+ pixel_9991/NB1 pixel_9991/VBIAS pixel_9991/NB2 pixel_9991/AMP_IN pixel_9991/SF_IB
+ pixel_9991/PIX_OUT pixel_9991/CSA_VREF pixel
Xpixel_709 pixel_709/gring pixel_709/VDD pixel_709/GND pixel_709/VREF pixel_709/ROW_SEL
+ pixel_709/NB1 pixel_709/VBIAS pixel_709/NB2 pixel_709/AMP_IN pixel_709/SF_IB pixel_709/PIX_OUT
+ pixel_709/CSA_VREF pixel
Xpixel_8008 pixel_8008/gring pixel_8008/VDD pixel_8008/GND pixel_8008/VREF pixel_8008/ROW_SEL
+ pixel_8008/NB1 pixel_8008/VBIAS pixel_8008/NB2 pixel_8008/AMP_IN pixel_8008/SF_IB
+ pixel_8008/PIX_OUT pixel_8008/CSA_VREF pixel
Xpixel_8019 pixel_8019/gring pixel_8019/VDD pixel_8019/GND pixel_8019/VREF pixel_8019/ROW_SEL
+ pixel_8019/NB1 pixel_8019/VBIAS pixel_8019/NB2 pixel_8019/AMP_IN pixel_8019/SF_IB
+ pixel_8019/PIX_OUT pixel_8019/CSA_VREF pixel
Xpixel_7307 pixel_7307/gring pixel_7307/VDD pixel_7307/GND pixel_7307/VREF pixel_7307/ROW_SEL
+ pixel_7307/NB1 pixel_7307/VBIAS pixel_7307/NB2 pixel_7307/AMP_IN pixel_7307/SF_IB
+ pixel_7307/PIX_OUT pixel_7307/CSA_VREF pixel
Xpixel_7318 pixel_7318/gring pixel_7318/VDD pixel_7318/GND pixel_7318/VREF pixel_7318/ROW_SEL
+ pixel_7318/NB1 pixel_7318/VBIAS pixel_7318/NB2 pixel_7318/AMP_IN pixel_7318/SF_IB
+ pixel_7318/PIX_OUT pixel_7318/CSA_VREF pixel
Xpixel_7329 pixel_7329/gring pixel_7329/VDD pixel_7329/GND pixel_7329/VREF pixel_7329/ROW_SEL
+ pixel_7329/NB1 pixel_7329/VBIAS pixel_7329/NB2 pixel_7329/AMP_IN pixel_7329/SF_IB
+ pixel_7329/PIX_OUT pixel_7329/CSA_VREF pixel
Xpixel_6606 pixel_6606/gring pixel_6606/VDD pixel_6606/GND pixel_6606/VREF pixel_6606/ROW_SEL
+ pixel_6606/NB1 pixel_6606/VBIAS pixel_6606/NB2 pixel_6606/AMP_IN pixel_6606/SF_IB
+ pixel_6606/PIX_OUT pixel_6606/CSA_VREF pixel
Xpixel_6617 pixel_6617/gring pixel_6617/VDD pixel_6617/GND pixel_6617/VREF pixel_6617/ROW_SEL
+ pixel_6617/NB1 pixel_6617/VBIAS pixel_6617/NB2 pixel_6617/AMP_IN pixel_6617/SF_IB
+ pixel_6617/PIX_OUT pixel_6617/CSA_VREF pixel
Xpixel_6628 pixel_6628/gring pixel_6628/VDD pixel_6628/GND pixel_6628/VREF pixel_6628/ROW_SEL
+ pixel_6628/NB1 pixel_6628/VBIAS pixel_6628/NB2 pixel_6628/AMP_IN pixel_6628/SF_IB
+ pixel_6628/PIX_OUT pixel_6628/CSA_VREF pixel
Xpixel_6639 pixel_6639/gring pixel_6639/VDD pixel_6639/GND pixel_6639/VREF pixel_6639/ROW_SEL
+ pixel_6639/NB1 pixel_6639/VBIAS pixel_6639/NB2 pixel_6639/AMP_IN pixel_6639/SF_IB
+ pixel_6639/PIX_OUT pixel_6639/CSA_VREF pixel
Xpixel_5905 pixel_5905/gring pixel_5905/VDD pixel_5905/GND pixel_5905/VREF pixel_5905/ROW_SEL
+ pixel_5905/NB1 pixel_5905/VBIAS pixel_5905/NB2 pixel_5905/AMP_IN pixel_5905/SF_IB
+ pixel_5905/PIX_OUT pixel_5905/CSA_VREF pixel
Xpixel_5916 pixel_5916/gring pixel_5916/VDD pixel_5916/GND pixel_5916/VREF pixel_5916/ROW_SEL
+ pixel_5916/NB1 pixel_5916/VBIAS pixel_5916/NB2 pixel_5916/AMP_IN pixel_5916/SF_IB
+ pixel_5916/PIX_OUT pixel_5916/CSA_VREF pixel
Xpixel_5927 pixel_5927/gring pixel_5927/VDD pixel_5927/GND pixel_5927/VREF pixel_5927/ROW_SEL
+ pixel_5927/NB1 pixel_5927/VBIAS pixel_5927/NB2 pixel_5927/AMP_IN pixel_5927/SF_IB
+ pixel_5927/PIX_OUT pixel_5927/CSA_VREF pixel
Xpixel_5938 pixel_5938/gring pixel_5938/VDD pixel_5938/GND pixel_5938/VREF pixel_5938/ROW_SEL
+ pixel_5938/NB1 pixel_5938/VBIAS pixel_5938/NB2 pixel_5938/AMP_IN pixel_5938/SF_IB
+ pixel_5938/PIX_OUT pixel_5938/CSA_VREF pixel
Xpixel_5949 pixel_5949/gring pixel_5949/VDD pixel_5949/GND pixel_5949/VREF pixel_5949/ROW_SEL
+ pixel_5949/NB1 pixel_5949/VBIAS pixel_5949/NB2 pixel_5949/AMP_IN pixel_5949/SF_IB
+ pixel_5949/PIX_OUT pixel_5949/CSA_VREF pixel
Xpixel_9221 pixel_9221/gring pixel_9221/VDD pixel_9221/GND pixel_9221/VREF pixel_9221/ROW_SEL
+ pixel_9221/NB1 pixel_9221/VBIAS pixel_9221/NB2 pixel_9221/AMP_IN pixel_9221/SF_IB
+ pixel_9221/PIX_OUT pixel_9221/CSA_VREF pixel
Xpixel_9210 pixel_9210/gring pixel_9210/VDD pixel_9210/GND pixel_9210/VREF pixel_9210/ROW_SEL
+ pixel_9210/NB1 pixel_9210/VBIAS pixel_9210/NB2 pixel_9210/AMP_IN pixel_9210/SF_IB
+ pixel_9210/PIX_OUT pixel_9210/CSA_VREF pixel
Xpixel_8520 pixel_8520/gring pixel_8520/VDD pixel_8520/GND pixel_8520/VREF pixel_8520/ROW_SEL
+ pixel_8520/NB1 pixel_8520/VBIAS pixel_8520/NB2 pixel_8520/AMP_IN pixel_8520/SF_IB
+ pixel_8520/PIX_OUT pixel_8520/CSA_VREF pixel
Xpixel_9265 pixel_9265/gring pixel_9265/VDD pixel_9265/GND pixel_9265/VREF pixel_9265/ROW_SEL
+ pixel_9265/NB1 pixel_9265/VBIAS pixel_9265/NB2 pixel_9265/AMP_IN pixel_9265/SF_IB
+ pixel_9265/PIX_OUT pixel_9265/CSA_VREF pixel
Xpixel_9254 pixel_9254/gring pixel_9254/VDD pixel_9254/GND pixel_9254/VREF pixel_9254/ROW_SEL
+ pixel_9254/NB1 pixel_9254/VBIAS pixel_9254/NB2 pixel_9254/AMP_IN pixel_9254/SF_IB
+ pixel_9254/PIX_OUT pixel_9254/CSA_VREF pixel
Xpixel_9243 pixel_9243/gring pixel_9243/VDD pixel_9243/GND pixel_9243/VREF pixel_9243/ROW_SEL
+ pixel_9243/NB1 pixel_9243/VBIAS pixel_9243/NB2 pixel_9243/AMP_IN pixel_9243/SF_IB
+ pixel_9243/PIX_OUT pixel_9243/CSA_VREF pixel
Xpixel_9232 pixel_9232/gring pixel_9232/VDD pixel_9232/GND pixel_9232/VREF pixel_9232/ROW_SEL
+ pixel_9232/NB1 pixel_9232/VBIAS pixel_9232/NB2 pixel_9232/AMP_IN pixel_9232/SF_IB
+ pixel_9232/PIX_OUT pixel_9232/CSA_VREF pixel
Xpixel_8553 pixel_8553/gring pixel_8553/VDD pixel_8553/GND pixel_8553/VREF pixel_8553/ROW_SEL
+ pixel_8553/NB1 pixel_8553/VBIAS pixel_8553/NB2 pixel_8553/AMP_IN pixel_8553/SF_IB
+ pixel_8553/PIX_OUT pixel_8553/CSA_VREF pixel
Xpixel_8542 pixel_8542/gring pixel_8542/VDD pixel_8542/GND pixel_8542/VREF pixel_8542/ROW_SEL
+ pixel_8542/NB1 pixel_8542/VBIAS pixel_8542/NB2 pixel_8542/AMP_IN pixel_8542/SF_IB
+ pixel_8542/PIX_OUT pixel_8542/CSA_VREF pixel
Xpixel_8531 pixel_8531/gring pixel_8531/VDD pixel_8531/GND pixel_8531/VREF pixel_8531/ROW_SEL
+ pixel_8531/NB1 pixel_8531/VBIAS pixel_8531/NB2 pixel_8531/AMP_IN pixel_8531/SF_IB
+ pixel_8531/PIX_OUT pixel_8531/CSA_VREF pixel
Xpixel_9298 pixel_9298/gring pixel_9298/VDD pixel_9298/GND pixel_9298/VREF pixel_9298/ROW_SEL
+ pixel_9298/NB1 pixel_9298/VBIAS pixel_9298/NB2 pixel_9298/AMP_IN pixel_9298/SF_IB
+ pixel_9298/PIX_OUT pixel_9298/CSA_VREF pixel
Xpixel_9287 pixel_9287/gring pixel_9287/VDD pixel_9287/GND pixel_9287/VREF pixel_9287/ROW_SEL
+ pixel_9287/NB1 pixel_9287/VBIAS pixel_9287/NB2 pixel_9287/AMP_IN pixel_9287/SF_IB
+ pixel_9287/PIX_OUT pixel_9287/CSA_VREF pixel
Xpixel_9276 pixel_9276/gring pixel_9276/VDD pixel_9276/GND pixel_9276/VREF pixel_9276/ROW_SEL
+ pixel_9276/NB1 pixel_9276/VBIAS pixel_9276/NB2 pixel_9276/AMP_IN pixel_9276/SF_IB
+ pixel_9276/PIX_OUT pixel_9276/CSA_VREF pixel
Xpixel_8586 pixel_8586/gring pixel_8586/VDD pixel_8586/GND pixel_8586/VREF pixel_8586/ROW_SEL
+ pixel_8586/NB1 pixel_8586/VBIAS pixel_8586/NB2 pixel_8586/AMP_IN pixel_8586/SF_IB
+ pixel_8586/PIX_OUT pixel_8586/CSA_VREF pixel
Xpixel_8575 pixel_8575/gring pixel_8575/VDD pixel_8575/GND pixel_8575/VREF pixel_8575/ROW_SEL
+ pixel_8575/NB1 pixel_8575/VBIAS pixel_8575/NB2 pixel_8575/AMP_IN pixel_8575/SF_IB
+ pixel_8575/PIX_OUT pixel_8575/CSA_VREF pixel
Xpixel_8564 pixel_8564/gring pixel_8564/VDD pixel_8564/GND pixel_8564/VREF pixel_8564/ROW_SEL
+ pixel_8564/NB1 pixel_8564/VBIAS pixel_8564/NB2 pixel_8564/AMP_IN pixel_8564/SF_IB
+ pixel_8564/PIX_OUT pixel_8564/CSA_VREF pixel
Xpixel_7830 pixel_7830/gring pixel_7830/VDD pixel_7830/GND pixel_7830/VREF pixel_7830/ROW_SEL
+ pixel_7830/NB1 pixel_7830/VBIAS pixel_7830/NB2 pixel_7830/AMP_IN pixel_7830/SF_IB
+ pixel_7830/PIX_OUT pixel_7830/CSA_VREF pixel
Xpixel_7841 pixel_7841/gring pixel_7841/VDD pixel_7841/GND pixel_7841/VREF pixel_7841/ROW_SEL
+ pixel_7841/NB1 pixel_7841/VBIAS pixel_7841/NB2 pixel_7841/AMP_IN pixel_7841/SF_IB
+ pixel_7841/PIX_OUT pixel_7841/CSA_VREF pixel
Xpixel_7852 pixel_7852/gring pixel_7852/VDD pixel_7852/GND pixel_7852/VREF pixel_7852/ROW_SEL
+ pixel_7852/NB1 pixel_7852/VBIAS pixel_7852/NB2 pixel_7852/AMP_IN pixel_7852/SF_IB
+ pixel_7852/PIX_OUT pixel_7852/CSA_VREF pixel
Xpixel_8597 pixel_8597/gring pixel_8597/VDD pixel_8597/GND pixel_8597/VREF pixel_8597/ROW_SEL
+ pixel_8597/NB1 pixel_8597/VBIAS pixel_8597/NB2 pixel_8597/AMP_IN pixel_8597/SF_IB
+ pixel_8597/PIX_OUT pixel_8597/CSA_VREF pixel
Xpixel_7863 pixel_7863/gring pixel_7863/VDD pixel_7863/GND pixel_7863/VREF pixel_7863/ROW_SEL
+ pixel_7863/NB1 pixel_7863/VBIAS pixel_7863/NB2 pixel_7863/AMP_IN pixel_7863/SF_IB
+ pixel_7863/PIX_OUT pixel_7863/CSA_VREF pixel
Xpixel_7874 pixel_7874/gring pixel_7874/VDD pixel_7874/GND pixel_7874/VREF pixel_7874/ROW_SEL
+ pixel_7874/NB1 pixel_7874/VBIAS pixel_7874/NB2 pixel_7874/AMP_IN pixel_7874/SF_IB
+ pixel_7874/PIX_OUT pixel_7874/CSA_VREF pixel
Xpixel_7885 pixel_7885/gring pixel_7885/VDD pixel_7885/GND pixel_7885/VREF pixel_7885/ROW_SEL
+ pixel_7885/NB1 pixel_7885/VBIAS pixel_7885/NB2 pixel_7885/AMP_IN pixel_7885/SF_IB
+ pixel_7885/PIX_OUT pixel_7885/CSA_VREF pixel
Xpixel_7896 pixel_7896/gring pixel_7896/VDD pixel_7896/GND pixel_7896/VREF pixel_7896/ROW_SEL
+ pixel_7896/NB1 pixel_7896/VBIAS pixel_7896/NB2 pixel_7896/AMP_IN pixel_7896/SF_IB
+ pixel_7896/PIX_OUT pixel_7896/CSA_VREF pixel
Xpixel_2181 pixel_2181/gring pixel_2181/VDD pixel_2181/GND pixel_2181/VREF pixel_2181/ROW_SEL
+ pixel_2181/NB1 pixel_2181/VBIAS pixel_2181/NB2 pixel_2181/AMP_IN pixel_2181/SF_IB
+ pixel_2181/PIX_OUT pixel_2181/CSA_VREF pixel
Xpixel_2170 pixel_2170/gring pixel_2170/VDD pixel_2170/GND pixel_2170/VREF pixel_2170/ROW_SEL
+ pixel_2170/NB1 pixel_2170/VBIAS pixel_2170/NB2 pixel_2170/AMP_IN pixel_2170/SF_IB
+ pixel_2170/PIX_OUT pixel_2170/CSA_VREF pixel
Xpixel_2192 pixel_2192/gring pixel_2192/VDD pixel_2192/GND pixel_2192/VREF pixel_2192/ROW_SEL
+ pixel_2192/NB1 pixel_2192/VBIAS pixel_2192/NB2 pixel_2192/AMP_IN pixel_2192/SF_IB
+ pixel_2192/PIX_OUT pixel_2192/CSA_VREF pixel
Xpixel_1491 pixel_1491/gring pixel_1491/VDD pixel_1491/GND pixel_1491/VREF pixel_1491/ROW_SEL
+ pixel_1491/NB1 pixel_1491/VBIAS pixel_1491/NB2 pixel_1491/AMP_IN pixel_1491/SF_IB
+ pixel_1491/PIX_OUT pixel_1491/CSA_VREF pixel
Xpixel_1480 pixel_1480/gring pixel_1480/VDD pixel_1480/GND pixel_1480/VREF pixel_1480/ROW_SEL
+ pixel_1480/NB1 pixel_1480/VBIAS pixel_1480/NB2 pixel_1480/AMP_IN pixel_1480/SF_IB
+ pixel_1480/PIX_OUT pixel_1480/CSA_VREF pixel
Xpixel_539 pixel_539/gring pixel_539/VDD pixel_539/GND pixel_539/VREF pixel_539/ROW_SEL
+ pixel_539/NB1 pixel_539/VBIAS pixel_539/NB2 pixel_539/AMP_IN pixel_539/SF_IB pixel_539/PIX_OUT
+ pixel_539/CSA_VREF pixel
Xpixel_528 pixel_528/gring pixel_528/VDD pixel_528/GND pixel_528/VREF pixel_528/ROW_SEL
+ pixel_528/NB1 pixel_528/VBIAS pixel_528/NB2 pixel_528/AMP_IN pixel_528/SF_IB pixel_528/PIX_OUT
+ pixel_528/CSA_VREF pixel
Xpixel_517 pixel_517/gring pixel_517/VDD pixel_517/GND pixel_517/VREF pixel_517/ROW_SEL
+ pixel_517/NB1 pixel_517/VBIAS pixel_517/NB2 pixel_517/AMP_IN pixel_517/SF_IB pixel_517/PIX_OUT
+ pixel_517/CSA_VREF pixel
Xpixel_506 pixel_506/gring pixel_506/VDD pixel_506/GND pixel_506/VREF pixel_506/ROW_SEL
+ pixel_506/NB1 pixel_506/VBIAS pixel_506/NB2 pixel_506/AMP_IN pixel_506/SF_IB pixel_506/PIX_OUT
+ pixel_506/CSA_VREF pixel
Xpixel_7104 pixel_7104/gring pixel_7104/VDD pixel_7104/GND pixel_7104/VREF pixel_7104/ROW_SEL
+ pixel_7104/NB1 pixel_7104/VBIAS pixel_7104/NB2 pixel_7104/AMP_IN pixel_7104/SF_IB
+ pixel_7104/PIX_OUT pixel_7104/CSA_VREF pixel
Xpixel_7115 pixel_7115/gring pixel_7115/VDD pixel_7115/GND pixel_7115/VREF pixel_7115/ROW_SEL
+ pixel_7115/NB1 pixel_7115/VBIAS pixel_7115/NB2 pixel_7115/AMP_IN pixel_7115/SF_IB
+ pixel_7115/PIX_OUT pixel_7115/CSA_VREF pixel
Xpixel_7126 pixel_7126/gring pixel_7126/VDD pixel_7126/GND pixel_7126/VREF pixel_7126/ROW_SEL
+ pixel_7126/NB1 pixel_7126/VBIAS pixel_7126/NB2 pixel_7126/AMP_IN pixel_7126/SF_IB
+ pixel_7126/PIX_OUT pixel_7126/CSA_VREF pixel
Xpixel_7137 pixel_7137/gring pixel_7137/VDD pixel_7137/GND pixel_7137/VREF pixel_7137/ROW_SEL
+ pixel_7137/NB1 pixel_7137/VBIAS pixel_7137/NB2 pixel_7137/AMP_IN pixel_7137/SF_IB
+ pixel_7137/PIX_OUT pixel_7137/CSA_VREF pixel
Xpixel_7148 pixel_7148/gring pixel_7148/VDD pixel_7148/GND pixel_7148/VREF pixel_7148/ROW_SEL
+ pixel_7148/NB1 pixel_7148/VBIAS pixel_7148/NB2 pixel_7148/AMP_IN pixel_7148/SF_IB
+ pixel_7148/PIX_OUT pixel_7148/CSA_VREF pixel
Xpixel_7159 pixel_7159/gring pixel_7159/VDD pixel_7159/GND pixel_7159/VREF pixel_7159/ROW_SEL
+ pixel_7159/NB1 pixel_7159/VBIAS pixel_7159/NB2 pixel_7159/AMP_IN pixel_7159/SF_IB
+ pixel_7159/PIX_OUT pixel_7159/CSA_VREF pixel
Xpixel_6403 pixel_6403/gring pixel_6403/VDD pixel_6403/GND pixel_6403/VREF pixel_6403/ROW_SEL
+ pixel_6403/NB1 pixel_6403/VBIAS pixel_6403/NB2 pixel_6403/AMP_IN pixel_6403/SF_IB
+ pixel_6403/PIX_OUT pixel_6403/CSA_VREF pixel
Xpixel_6414 pixel_6414/gring pixel_6414/VDD pixel_6414/GND pixel_6414/VREF pixel_6414/ROW_SEL
+ pixel_6414/NB1 pixel_6414/VBIAS pixel_6414/NB2 pixel_6414/AMP_IN pixel_6414/SF_IB
+ pixel_6414/PIX_OUT pixel_6414/CSA_VREF pixel
Xpixel_6425 pixel_6425/gring pixel_6425/VDD pixel_6425/GND pixel_6425/VREF pixel_6425/ROW_SEL
+ pixel_6425/NB1 pixel_6425/VBIAS pixel_6425/NB2 pixel_6425/AMP_IN pixel_6425/SF_IB
+ pixel_6425/PIX_OUT pixel_6425/CSA_VREF pixel
Xpixel_6436 pixel_6436/gring pixel_6436/VDD pixel_6436/GND pixel_6436/VREF pixel_6436/ROW_SEL
+ pixel_6436/NB1 pixel_6436/VBIAS pixel_6436/NB2 pixel_6436/AMP_IN pixel_6436/SF_IB
+ pixel_6436/PIX_OUT pixel_6436/CSA_VREF pixel
Xpixel_6447 pixel_6447/gring pixel_6447/VDD pixel_6447/GND pixel_6447/VREF pixel_6447/ROW_SEL
+ pixel_6447/NB1 pixel_6447/VBIAS pixel_6447/NB2 pixel_6447/AMP_IN pixel_6447/SF_IB
+ pixel_6447/PIX_OUT pixel_6447/CSA_VREF pixel
Xpixel_6458 pixel_6458/gring pixel_6458/VDD pixel_6458/GND pixel_6458/VREF pixel_6458/ROW_SEL
+ pixel_6458/NB1 pixel_6458/VBIAS pixel_6458/NB2 pixel_6458/AMP_IN pixel_6458/SF_IB
+ pixel_6458/PIX_OUT pixel_6458/CSA_VREF pixel
Xpixel_6469 pixel_6469/gring pixel_6469/VDD pixel_6469/GND pixel_6469/VREF pixel_6469/ROW_SEL
+ pixel_6469/NB1 pixel_6469/VBIAS pixel_6469/NB2 pixel_6469/AMP_IN pixel_6469/SF_IB
+ pixel_6469/PIX_OUT pixel_6469/CSA_VREF pixel
Xpixel_5702 pixel_5702/gring pixel_5702/VDD pixel_5702/GND pixel_5702/VREF pixel_5702/ROW_SEL
+ pixel_5702/NB1 pixel_5702/VBIAS pixel_5702/NB2 pixel_5702/AMP_IN pixel_5702/SF_IB
+ pixel_5702/PIX_OUT pixel_5702/CSA_VREF pixel
Xpixel_5713 pixel_5713/gring pixel_5713/VDD pixel_5713/GND pixel_5713/VREF pixel_5713/ROW_SEL
+ pixel_5713/NB1 pixel_5713/VBIAS pixel_5713/NB2 pixel_5713/AMP_IN pixel_5713/SF_IB
+ pixel_5713/PIX_OUT pixel_5713/CSA_VREF pixel
Xpixel_5724 pixel_5724/gring pixel_5724/VDD pixel_5724/GND pixel_5724/VREF pixel_5724/ROW_SEL
+ pixel_5724/NB1 pixel_5724/VBIAS pixel_5724/NB2 pixel_5724/AMP_IN pixel_5724/SF_IB
+ pixel_5724/PIX_OUT pixel_5724/CSA_VREF pixel
Xpixel_5735 pixel_5735/gring pixel_5735/VDD pixel_5735/GND pixel_5735/VREF pixel_5735/ROW_SEL
+ pixel_5735/NB1 pixel_5735/VBIAS pixel_5735/NB2 pixel_5735/AMP_IN pixel_5735/SF_IB
+ pixel_5735/PIX_OUT pixel_5735/CSA_VREF pixel
Xpixel_5746 pixel_5746/gring pixel_5746/VDD pixel_5746/GND pixel_5746/VREF pixel_5746/ROW_SEL
+ pixel_5746/NB1 pixel_5746/VBIAS pixel_5746/NB2 pixel_5746/AMP_IN pixel_5746/SF_IB
+ pixel_5746/PIX_OUT pixel_5746/CSA_VREF pixel
Xpixel_5757 pixel_5757/gring pixel_5757/VDD pixel_5757/GND pixel_5757/VREF pixel_5757/ROW_SEL
+ pixel_5757/NB1 pixel_5757/VBIAS pixel_5757/NB2 pixel_5757/AMP_IN pixel_5757/SF_IB
+ pixel_5757/PIX_OUT pixel_5757/CSA_VREF pixel
Xpixel_5768 pixel_5768/gring pixel_5768/VDD pixel_5768/GND pixel_5768/VREF pixel_5768/ROW_SEL
+ pixel_5768/NB1 pixel_5768/VBIAS pixel_5768/NB2 pixel_5768/AMP_IN pixel_5768/SF_IB
+ pixel_5768/PIX_OUT pixel_5768/CSA_VREF pixel
Xpixel_5779 pixel_5779/gring pixel_5779/VDD pixel_5779/GND pixel_5779/VREF pixel_5779/ROW_SEL
+ pixel_5779/NB1 pixel_5779/VBIAS pixel_5779/NB2 pixel_5779/AMP_IN pixel_5779/SF_IB
+ pixel_5779/PIX_OUT pixel_5779/CSA_VREF pixel
Xpixel_9040 pixel_9040/gring pixel_9040/VDD pixel_9040/GND pixel_9040/VREF pixel_9040/ROW_SEL
+ pixel_9040/NB1 pixel_9040/VBIAS pixel_9040/NB2 pixel_9040/AMP_IN pixel_9040/SF_IB
+ pixel_9040/PIX_OUT pixel_9040/CSA_VREF pixel
Xpixel_9073 pixel_9073/gring pixel_9073/VDD pixel_9073/GND pixel_9073/VREF pixel_9073/ROW_SEL
+ pixel_9073/NB1 pixel_9073/VBIAS pixel_9073/NB2 pixel_9073/AMP_IN pixel_9073/SF_IB
+ pixel_9073/PIX_OUT pixel_9073/CSA_VREF pixel
Xpixel_9062 pixel_9062/gring pixel_9062/VDD pixel_9062/GND pixel_9062/VREF pixel_9062/ROW_SEL
+ pixel_9062/NB1 pixel_9062/VBIAS pixel_9062/NB2 pixel_9062/AMP_IN pixel_9062/SF_IB
+ pixel_9062/PIX_OUT pixel_9062/CSA_VREF pixel
Xpixel_9051 pixel_9051/gring pixel_9051/VDD pixel_9051/GND pixel_9051/VREF pixel_9051/ROW_SEL
+ pixel_9051/NB1 pixel_9051/VBIAS pixel_9051/NB2 pixel_9051/AMP_IN pixel_9051/SF_IB
+ pixel_9051/PIX_OUT pixel_9051/CSA_VREF pixel
Xpixel_9095 pixel_9095/gring pixel_9095/VDD pixel_9095/GND pixel_9095/VREF pixel_9095/ROW_SEL
+ pixel_9095/NB1 pixel_9095/VBIAS pixel_9095/NB2 pixel_9095/AMP_IN pixel_9095/SF_IB
+ pixel_9095/PIX_OUT pixel_9095/CSA_VREF pixel
Xpixel_9084 pixel_9084/gring pixel_9084/VDD pixel_9084/GND pixel_9084/VREF pixel_9084/ROW_SEL
+ pixel_9084/NB1 pixel_9084/VBIAS pixel_9084/NB2 pixel_9084/AMP_IN pixel_9084/SF_IB
+ pixel_9084/PIX_OUT pixel_9084/CSA_VREF pixel
Xpixel_8350 pixel_8350/gring pixel_8350/VDD pixel_8350/GND pixel_8350/VREF pixel_8350/ROW_SEL
+ pixel_8350/NB1 pixel_8350/VBIAS pixel_8350/NB2 pixel_8350/AMP_IN pixel_8350/SF_IB
+ pixel_8350/PIX_OUT pixel_8350/CSA_VREF pixel
Xpixel_8361 pixel_8361/gring pixel_8361/VDD pixel_8361/GND pixel_8361/VREF pixel_8361/ROW_SEL
+ pixel_8361/NB1 pixel_8361/VBIAS pixel_8361/NB2 pixel_8361/AMP_IN pixel_8361/SF_IB
+ pixel_8361/PIX_OUT pixel_8361/CSA_VREF pixel
Xpixel_8372 pixel_8372/gring pixel_8372/VDD pixel_8372/GND pixel_8372/VREF pixel_8372/ROW_SEL
+ pixel_8372/NB1 pixel_8372/VBIAS pixel_8372/NB2 pixel_8372/AMP_IN pixel_8372/SF_IB
+ pixel_8372/PIX_OUT pixel_8372/CSA_VREF pixel
Xpixel_8383 pixel_8383/gring pixel_8383/VDD pixel_8383/GND pixel_8383/VREF pixel_8383/ROW_SEL
+ pixel_8383/NB1 pixel_8383/VBIAS pixel_8383/NB2 pixel_8383/AMP_IN pixel_8383/SF_IB
+ pixel_8383/PIX_OUT pixel_8383/CSA_VREF pixel
Xpixel_8394 pixel_8394/gring pixel_8394/VDD pixel_8394/GND pixel_8394/VREF pixel_8394/ROW_SEL
+ pixel_8394/NB1 pixel_8394/VBIAS pixel_8394/NB2 pixel_8394/AMP_IN pixel_8394/SF_IB
+ pixel_8394/PIX_OUT pixel_8394/CSA_VREF pixel
Xpixel_7660 pixel_7660/gring pixel_7660/VDD pixel_7660/GND pixel_7660/VREF pixel_7660/ROW_SEL
+ pixel_7660/NB1 pixel_7660/VBIAS pixel_7660/NB2 pixel_7660/AMP_IN pixel_7660/SF_IB
+ pixel_7660/PIX_OUT pixel_7660/CSA_VREF pixel
Xpixel_7671 pixel_7671/gring pixel_7671/VDD pixel_7671/GND pixel_7671/VREF pixel_7671/ROW_SEL
+ pixel_7671/NB1 pixel_7671/VBIAS pixel_7671/NB2 pixel_7671/AMP_IN pixel_7671/SF_IB
+ pixel_7671/PIX_OUT pixel_7671/CSA_VREF pixel
Xpixel_7682 pixel_7682/gring pixel_7682/VDD pixel_7682/GND pixel_7682/VREF pixel_7682/ROW_SEL
+ pixel_7682/NB1 pixel_7682/VBIAS pixel_7682/NB2 pixel_7682/AMP_IN pixel_7682/SF_IB
+ pixel_7682/PIX_OUT pixel_7682/CSA_VREF pixel
Xpixel_7693 pixel_7693/gring pixel_7693/VDD pixel_7693/GND pixel_7693/VREF pixel_7693/ROW_SEL
+ pixel_7693/NB1 pixel_7693/VBIAS pixel_7693/NB2 pixel_7693/AMP_IN pixel_7693/SF_IB
+ pixel_7693/PIX_OUT pixel_7693/CSA_VREF pixel
Xpixel_6970 pixel_6970/gring pixel_6970/VDD pixel_6970/GND pixel_6970/VREF pixel_6970/ROW_SEL
+ pixel_6970/NB1 pixel_6970/VBIAS pixel_6970/NB2 pixel_6970/AMP_IN pixel_6970/SF_IB
+ pixel_6970/PIX_OUT pixel_6970/CSA_VREF pixel
Xpixel_6981 pixel_6981/gring pixel_6981/VDD pixel_6981/GND pixel_6981/VREF pixel_6981/ROW_SEL
+ pixel_6981/NB1 pixel_6981/VBIAS pixel_6981/NB2 pixel_6981/AMP_IN pixel_6981/SF_IB
+ pixel_6981/PIX_OUT pixel_6981/CSA_VREF pixel
Xpixel_73 pixel_73/gring pixel_73/VDD pixel_73/GND pixel_73/VREF pixel_73/ROW_SEL
+ pixel_73/NB1 pixel_73/VBIAS pixel_73/NB2 pixel_73/AMP_IN pixel_73/SF_IB pixel_73/PIX_OUT
+ pixel_73/CSA_VREF pixel
Xpixel_62 pixel_62/gring pixel_62/VDD pixel_62/GND pixel_62/VREF pixel_62/ROW_SEL
+ pixel_62/NB1 pixel_62/VBIAS pixel_62/NB2 pixel_62/AMP_IN pixel_62/SF_IB pixel_62/PIX_OUT
+ pixel_62/CSA_VREF pixel
Xpixel_51 pixel_51/gring pixel_51/VDD pixel_51/GND pixel_51/VREF pixel_51/ROW_SEL
+ pixel_51/NB1 pixel_51/VBIAS pixel_51/NB2 pixel_51/AMP_IN pixel_51/SF_IB pixel_51/PIX_OUT
+ pixel_51/CSA_VREF pixel
Xpixel_40 pixel_40/gring pixel_40/VDD pixel_40/GND pixel_40/VREF pixel_40/ROW_SEL
+ pixel_40/NB1 pixel_40/VBIAS pixel_40/NB2 pixel_40/AMP_IN pixel_40/SF_IB pixel_40/PIX_OUT
+ pixel_40/CSA_VREF pixel
Xpixel_6992 pixel_6992/gring pixel_6992/VDD pixel_6992/GND pixel_6992/VREF pixel_6992/ROW_SEL
+ pixel_6992/NB1 pixel_6992/VBIAS pixel_6992/NB2 pixel_6992/AMP_IN pixel_6992/SF_IB
+ pixel_6992/PIX_OUT pixel_6992/CSA_VREF pixel
Xpixel_95 pixel_95/gring pixel_95/VDD pixel_95/GND pixel_95/VREF pixel_95/ROW_SEL
+ pixel_95/NB1 pixel_95/VBIAS pixel_95/NB2 pixel_95/AMP_IN pixel_95/SF_IB pixel_95/PIX_OUT
+ pixel_95/CSA_VREF pixel
Xpixel_84 pixel_84/gring pixel_84/VDD pixel_84/GND pixel_84/VREF pixel_84/ROW_SEL
+ pixel_84/NB1 pixel_84/VBIAS pixel_84/NB2 pixel_84/AMP_IN pixel_84/SF_IB pixel_84/PIX_OUT
+ pixel_84/CSA_VREF pixel
Xpixel_5009 pixel_5009/gring pixel_5009/VDD pixel_5009/GND pixel_5009/VREF pixel_5009/ROW_SEL
+ pixel_5009/NB1 pixel_5009/VBIAS pixel_5009/NB2 pixel_5009/AMP_IN pixel_5009/SF_IB
+ pixel_5009/PIX_OUT pixel_5009/CSA_VREF pixel
Xpixel_303 pixel_303/gring pixel_303/VDD pixel_303/GND pixel_303/VREF pixel_303/ROW_SEL
+ pixel_303/NB1 pixel_303/VBIAS pixel_303/NB2 pixel_303/AMP_IN pixel_303/SF_IB pixel_303/PIX_OUT
+ pixel_303/CSA_VREF pixel
Xpixel_4308 pixel_4308/gring pixel_4308/VDD pixel_4308/GND pixel_4308/VREF pixel_4308/ROW_SEL
+ pixel_4308/NB1 pixel_4308/VBIAS pixel_4308/NB2 pixel_4308/AMP_IN pixel_4308/SF_IB
+ pixel_4308/PIX_OUT pixel_4308/CSA_VREF pixel
Xpixel_347 pixel_347/gring pixel_347/VDD pixel_347/GND pixel_347/VREF pixel_347/ROW_SEL
+ pixel_347/NB1 pixel_347/VBIAS pixel_347/NB2 pixel_347/AMP_IN pixel_347/SF_IB pixel_347/PIX_OUT
+ pixel_347/CSA_VREF pixel
Xpixel_336 pixel_336/gring pixel_336/VDD pixel_336/GND pixel_336/VREF pixel_336/ROW_SEL
+ pixel_336/NB1 pixel_336/VBIAS pixel_336/NB2 pixel_336/AMP_IN pixel_336/SF_IB pixel_336/PIX_OUT
+ pixel_336/CSA_VREF pixel
Xpixel_325 pixel_325/gring pixel_325/VDD pixel_325/GND pixel_325/VREF pixel_325/ROW_SEL
+ pixel_325/NB1 pixel_325/VBIAS pixel_325/NB2 pixel_325/AMP_IN pixel_325/SF_IB pixel_325/PIX_OUT
+ pixel_325/CSA_VREF pixel
Xpixel_314 pixel_314/gring pixel_314/VDD pixel_314/GND pixel_314/VREF pixel_314/ROW_SEL
+ pixel_314/NB1 pixel_314/VBIAS pixel_314/NB2 pixel_314/AMP_IN pixel_314/SF_IB pixel_314/PIX_OUT
+ pixel_314/CSA_VREF pixel
Xpixel_3607 pixel_3607/gring pixel_3607/VDD pixel_3607/GND pixel_3607/VREF pixel_3607/ROW_SEL
+ pixel_3607/NB1 pixel_3607/VBIAS pixel_3607/NB2 pixel_3607/AMP_IN pixel_3607/SF_IB
+ pixel_3607/PIX_OUT pixel_3607/CSA_VREF pixel
Xpixel_4319 pixel_4319/gring pixel_4319/VDD pixel_4319/GND pixel_4319/VREF pixel_4319/ROW_SEL
+ pixel_4319/NB1 pixel_4319/VBIAS pixel_4319/NB2 pixel_4319/AMP_IN pixel_4319/SF_IB
+ pixel_4319/PIX_OUT pixel_4319/CSA_VREF pixel
Xpixel_369 pixel_369/gring pixel_369/VDD pixel_369/GND pixel_369/VREF pixel_369/ROW_SEL
+ pixel_369/NB1 pixel_369/VBIAS pixel_369/NB2 pixel_369/AMP_IN pixel_369/SF_IB pixel_369/PIX_OUT
+ pixel_369/CSA_VREF pixel
Xpixel_358 pixel_358/gring pixel_358/VDD pixel_358/GND pixel_358/VREF pixel_358/ROW_SEL
+ pixel_358/NB1 pixel_358/VBIAS pixel_358/NB2 pixel_358/AMP_IN pixel_358/SF_IB pixel_358/PIX_OUT
+ pixel_358/CSA_VREF pixel
Xpixel_3629 pixel_3629/gring pixel_3629/VDD pixel_3629/GND pixel_3629/VREF pixel_3629/ROW_SEL
+ pixel_3629/NB1 pixel_3629/VBIAS pixel_3629/NB2 pixel_3629/AMP_IN pixel_3629/SF_IB
+ pixel_3629/PIX_OUT pixel_3629/CSA_VREF pixel
Xpixel_3618 pixel_3618/gring pixel_3618/VDD pixel_3618/GND pixel_3618/VREF pixel_3618/ROW_SEL
+ pixel_3618/NB1 pixel_3618/VBIAS pixel_3618/NB2 pixel_3618/AMP_IN pixel_3618/SF_IB
+ pixel_3618/PIX_OUT pixel_3618/CSA_VREF pixel
Xpixel_2928 pixel_2928/gring pixel_2928/VDD pixel_2928/GND pixel_2928/VREF pixel_2928/ROW_SEL
+ pixel_2928/NB1 pixel_2928/VBIAS pixel_2928/NB2 pixel_2928/AMP_IN pixel_2928/SF_IB
+ pixel_2928/PIX_OUT pixel_2928/CSA_VREF pixel
Xpixel_2917 pixel_2917/gring pixel_2917/VDD pixel_2917/GND pixel_2917/VREF pixel_2917/ROW_SEL
+ pixel_2917/NB1 pixel_2917/VBIAS pixel_2917/NB2 pixel_2917/AMP_IN pixel_2917/SF_IB
+ pixel_2917/PIX_OUT pixel_2917/CSA_VREF pixel
Xpixel_2906 pixel_2906/gring pixel_2906/VDD pixel_2906/GND pixel_2906/VREF pixel_2906/ROW_SEL
+ pixel_2906/NB1 pixel_2906/VBIAS pixel_2906/NB2 pixel_2906/AMP_IN pixel_2906/SF_IB
+ pixel_2906/PIX_OUT pixel_2906/CSA_VREF pixel
Xpixel_2939 pixel_2939/gring pixel_2939/VDD pixel_2939/GND pixel_2939/VREF pixel_2939/ROW_SEL
+ pixel_2939/NB1 pixel_2939/VBIAS pixel_2939/NB2 pixel_2939/AMP_IN pixel_2939/SF_IB
+ pixel_2939/PIX_OUT pixel_2939/CSA_VREF pixel
Xpixel_6200 pixel_6200/gring pixel_6200/VDD pixel_6200/GND pixel_6200/VREF pixel_6200/ROW_SEL
+ pixel_6200/NB1 pixel_6200/VBIAS pixel_6200/NB2 pixel_6200/AMP_IN pixel_6200/SF_IB
+ pixel_6200/PIX_OUT pixel_6200/CSA_VREF pixel
Xpixel_6211 pixel_6211/gring pixel_6211/VDD pixel_6211/GND pixel_6211/VREF pixel_6211/ROW_SEL
+ pixel_6211/NB1 pixel_6211/VBIAS pixel_6211/NB2 pixel_6211/AMP_IN pixel_6211/SF_IB
+ pixel_6211/PIX_OUT pixel_6211/CSA_VREF pixel
Xpixel_6222 pixel_6222/gring pixel_6222/VDD pixel_6222/GND pixel_6222/VREF pixel_6222/ROW_SEL
+ pixel_6222/NB1 pixel_6222/VBIAS pixel_6222/NB2 pixel_6222/AMP_IN pixel_6222/SF_IB
+ pixel_6222/PIX_OUT pixel_6222/CSA_VREF pixel
Xpixel_6233 pixel_6233/gring pixel_6233/VDD pixel_6233/GND pixel_6233/VREF pixel_6233/ROW_SEL
+ pixel_6233/NB1 pixel_6233/VBIAS pixel_6233/NB2 pixel_6233/AMP_IN pixel_6233/SF_IB
+ pixel_6233/PIX_OUT pixel_6233/CSA_VREF pixel
Xpixel_6244 pixel_6244/gring pixel_6244/VDD pixel_6244/GND pixel_6244/VREF pixel_6244/ROW_SEL
+ pixel_6244/NB1 pixel_6244/VBIAS pixel_6244/NB2 pixel_6244/AMP_IN pixel_6244/SF_IB
+ pixel_6244/PIX_OUT pixel_6244/CSA_VREF pixel
Xpixel_6255 pixel_6255/gring pixel_6255/VDD pixel_6255/GND pixel_6255/VREF pixel_6255/ROW_SEL
+ pixel_6255/NB1 pixel_6255/VBIAS pixel_6255/NB2 pixel_6255/AMP_IN pixel_6255/SF_IB
+ pixel_6255/PIX_OUT pixel_6255/CSA_VREF pixel
Xpixel_6266 pixel_6266/gring pixel_6266/VDD pixel_6266/GND pixel_6266/VREF pixel_6266/ROW_SEL
+ pixel_6266/NB1 pixel_6266/VBIAS pixel_6266/NB2 pixel_6266/AMP_IN pixel_6266/SF_IB
+ pixel_6266/PIX_OUT pixel_6266/CSA_VREF pixel
Xpixel_6277 pixel_6277/gring pixel_6277/VDD pixel_6277/GND pixel_6277/VREF pixel_6277/ROW_SEL
+ pixel_6277/NB1 pixel_6277/VBIAS pixel_6277/NB2 pixel_6277/AMP_IN pixel_6277/SF_IB
+ pixel_6277/PIX_OUT pixel_6277/CSA_VREF pixel
Xpixel_5510 pixel_5510/gring pixel_5510/VDD pixel_5510/GND pixel_5510/VREF pixel_5510/ROW_SEL
+ pixel_5510/NB1 pixel_5510/VBIAS pixel_5510/NB2 pixel_5510/AMP_IN pixel_5510/SF_IB
+ pixel_5510/PIX_OUT pixel_5510/CSA_VREF pixel
Xpixel_5521 pixel_5521/gring pixel_5521/VDD pixel_5521/GND pixel_5521/VREF pixel_5521/ROW_SEL
+ pixel_5521/NB1 pixel_5521/VBIAS pixel_5521/NB2 pixel_5521/AMP_IN pixel_5521/SF_IB
+ pixel_5521/PIX_OUT pixel_5521/CSA_VREF pixel
Xpixel_5532 pixel_5532/gring pixel_5532/VDD pixel_5532/GND pixel_5532/VREF pixel_5532/ROW_SEL
+ pixel_5532/NB1 pixel_5532/VBIAS pixel_5532/NB2 pixel_5532/AMP_IN pixel_5532/SF_IB
+ pixel_5532/PIX_OUT pixel_5532/CSA_VREF pixel
Xpixel_6288 pixel_6288/gring pixel_6288/VDD pixel_6288/GND pixel_6288/VREF pixel_6288/ROW_SEL
+ pixel_6288/NB1 pixel_6288/VBIAS pixel_6288/NB2 pixel_6288/AMP_IN pixel_6288/SF_IB
+ pixel_6288/PIX_OUT pixel_6288/CSA_VREF pixel
Xpixel_6299 pixel_6299/gring pixel_6299/VDD pixel_6299/GND pixel_6299/VREF pixel_6299/ROW_SEL
+ pixel_6299/NB1 pixel_6299/VBIAS pixel_6299/NB2 pixel_6299/AMP_IN pixel_6299/SF_IB
+ pixel_6299/PIX_OUT pixel_6299/CSA_VREF pixel
Xpixel_5543 pixel_5543/gring pixel_5543/VDD pixel_5543/GND pixel_5543/VREF pixel_5543/ROW_SEL
+ pixel_5543/NB1 pixel_5543/VBIAS pixel_5543/NB2 pixel_5543/AMP_IN pixel_5543/SF_IB
+ pixel_5543/PIX_OUT pixel_5543/CSA_VREF pixel
Xpixel_5554 pixel_5554/gring pixel_5554/VDD pixel_5554/GND pixel_5554/VREF pixel_5554/ROW_SEL
+ pixel_5554/NB1 pixel_5554/VBIAS pixel_5554/NB2 pixel_5554/AMP_IN pixel_5554/SF_IB
+ pixel_5554/PIX_OUT pixel_5554/CSA_VREF pixel
Xpixel_5565 pixel_5565/gring pixel_5565/VDD pixel_5565/GND pixel_5565/VREF pixel_5565/ROW_SEL
+ pixel_5565/NB1 pixel_5565/VBIAS pixel_5565/NB2 pixel_5565/AMP_IN pixel_5565/SF_IB
+ pixel_5565/PIX_OUT pixel_5565/CSA_VREF pixel
Xpixel_5576 pixel_5576/gring pixel_5576/VDD pixel_5576/GND pixel_5576/VREF pixel_5576/ROW_SEL
+ pixel_5576/NB1 pixel_5576/VBIAS pixel_5576/NB2 pixel_5576/AMP_IN pixel_5576/SF_IB
+ pixel_5576/PIX_OUT pixel_5576/CSA_VREF pixel
Xpixel_4820 pixel_4820/gring pixel_4820/VDD pixel_4820/GND pixel_4820/VREF pixel_4820/ROW_SEL
+ pixel_4820/NB1 pixel_4820/VBIAS pixel_4820/NB2 pixel_4820/AMP_IN pixel_4820/SF_IB
+ pixel_4820/PIX_OUT pixel_4820/CSA_VREF pixel
Xpixel_4831 pixel_4831/gring pixel_4831/VDD pixel_4831/GND pixel_4831/VREF pixel_4831/ROW_SEL
+ pixel_4831/NB1 pixel_4831/VBIAS pixel_4831/NB2 pixel_4831/AMP_IN pixel_4831/SF_IB
+ pixel_4831/PIX_OUT pixel_4831/CSA_VREF pixel
Xpixel_5587 pixel_5587/gring pixel_5587/VDD pixel_5587/GND pixel_5587/VREF pixel_5587/ROW_SEL
+ pixel_5587/NB1 pixel_5587/VBIAS pixel_5587/NB2 pixel_5587/AMP_IN pixel_5587/SF_IB
+ pixel_5587/PIX_OUT pixel_5587/CSA_VREF pixel
Xpixel_5598 pixel_5598/gring pixel_5598/VDD pixel_5598/GND pixel_5598/VREF pixel_5598/ROW_SEL
+ pixel_5598/NB1 pixel_5598/VBIAS pixel_5598/NB2 pixel_5598/AMP_IN pixel_5598/SF_IB
+ pixel_5598/PIX_OUT pixel_5598/CSA_VREF pixel
Xpixel_4842 pixel_4842/gring pixel_4842/VDD pixel_4842/GND pixel_4842/VREF pixel_4842/ROW_SEL
+ pixel_4842/NB1 pixel_4842/VBIAS pixel_4842/NB2 pixel_4842/AMP_IN pixel_4842/SF_IB
+ pixel_4842/PIX_OUT pixel_4842/CSA_VREF pixel
Xpixel_4853 pixel_4853/gring pixel_4853/VDD pixel_4853/GND pixel_4853/VREF pixel_4853/ROW_SEL
+ pixel_4853/NB1 pixel_4853/VBIAS pixel_4853/NB2 pixel_4853/AMP_IN pixel_4853/SF_IB
+ pixel_4853/PIX_OUT pixel_4853/CSA_VREF pixel
Xpixel_4864 pixel_4864/gring pixel_4864/VDD pixel_4864/GND pixel_4864/VREF pixel_4864/ROW_SEL
+ pixel_4864/NB1 pixel_4864/VBIAS pixel_4864/NB2 pixel_4864/AMP_IN pixel_4864/SF_IB
+ pixel_4864/PIX_OUT pixel_4864/CSA_VREF pixel
Xpixel_892 pixel_892/gring pixel_892/VDD pixel_892/GND pixel_892/VREF pixel_892/ROW_SEL
+ pixel_892/NB1 pixel_892/VBIAS pixel_892/NB2 pixel_892/AMP_IN pixel_892/SF_IB pixel_892/PIX_OUT
+ pixel_892/CSA_VREF pixel
Xpixel_881 pixel_881/gring pixel_881/VDD pixel_881/GND pixel_881/VREF pixel_881/ROW_SEL
+ pixel_881/NB1 pixel_881/VBIAS pixel_881/NB2 pixel_881/AMP_IN pixel_881/SF_IB pixel_881/PIX_OUT
+ pixel_881/CSA_VREF pixel
Xpixel_870 pixel_870/gring pixel_870/VDD pixel_870/GND pixel_870/VREF pixel_870/ROW_SEL
+ pixel_870/NB1 pixel_870/VBIAS pixel_870/NB2 pixel_870/AMP_IN pixel_870/SF_IB pixel_870/PIX_OUT
+ pixel_870/CSA_VREF pixel
Xpixel_4875 pixel_4875/gring pixel_4875/VDD pixel_4875/GND pixel_4875/VREF pixel_4875/ROW_SEL
+ pixel_4875/NB1 pixel_4875/VBIAS pixel_4875/NB2 pixel_4875/AMP_IN pixel_4875/SF_IB
+ pixel_4875/PIX_OUT pixel_4875/CSA_VREF pixel
Xpixel_4886 pixel_4886/gring pixel_4886/VDD pixel_4886/GND pixel_4886/VREF pixel_4886/ROW_SEL
+ pixel_4886/NB1 pixel_4886/VBIAS pixel_4886/NB2 pixel_4886/AMP_IN pixel_4886/SF_IB
+ pixel_4886/PIX_OUT pixel_4886/CSA_VREF pixel
Xpixel_4897 pixel_4897/gring pixel_4897/VDD pixel_4897/GND pixel_4897/VREF pixel_4897/ROW_SEL
+ pixel_4897/NB1 pixel_4897/VBIAS pixel_4897/NB2 pixel_4897/AMP_IN pixel_4897/SF_IB
+ pixel_4897/PIX_OUT pixel_4897/CSA_VREF pixel
Xpixel_8180 pixel_8180/gring pixel_8180/VDD pixel_8180/GND pixel_8180/VREF pixel_8180/ROW_SEL
+ pixel_8180/NB1 pixel_8180/VBIAS pixel_8180/NB2 pixel_8180/AMP_IN pixel_8180/SF_IB
+ pixel_8180/PIX_OUT pixel_8180/CSA_VREF pixel
Xpixel_8191 pixel_8191/gring pixel_8191/VDD pixel_8191/GND pixel_8191/VREF pixel_8191/ROW_SEL
+ pixel_8191/NB1 pixel_8191/VBIAS pixel_8191/NB2 pixel_8191/AMP_IN pixel_8191/SF_IB
+ pixel_8191/PIX_OUT pixel_8191/CSA_VREF pixel
Xpixel_7490 pixel_7490/gring pixel_7490/VDD pixel_7490/GND pixel_7490/VREF pixel_7490/ROW_SEL
+ pixel_7490/NB1 pixel_7490/VBIAS pixel_7490/NB2 pixel_7490/AMP_IN pixel_7490/SF_IB
+ pixel_7490/PIX_OUT pixel_7490/CSA_VREF pixel
Xpixel_9809 pixel_9809/gring pixel_9809/VDD pixel_9809/GND pixel_9809/VREF pixel_9809/ROW_SEL
+ pixel_9809/NB1 pixel_9809/VBIAS pixel_9809/NB2 pixel_9809/AMP_IN pixel_9809/SF_IB
+ pixel_9809/PIX_OUT pixel_9809/CSA_VREF pixel
Xpixel_122 pixel_122/gring pixel_122/VDD pixel_122/GND pixel_122/VREF pixel_122/ROW_SEL
+ pixel_122/NB1 pixel_122/VBIAS pixel_122/NB2 pixel_122/AMP_IN pixel_122/SF_IB pixel_122/PIX_OUT
+ pixel_122/CSA_VREF pixel
Xpixel_111 pixel_111/gring pixel_111/VDD pixel_111/GND pixel_111/VREF pixel_111/ROW_SEL
+ pixel_111/NB1 pixel_111/VBIAS pixel_111/NB2 pixel_111/AMP_IN pixel_111/SF_IB pixel_111/PIX_OUT
+ pixel_111/CSA_VREF pixel
Xpixel_100 pixel_100/gring pixel_100/VDD pixel_100/GND pixel_100/VREF pixel_100/ROW_SEL
+ pixel_100/NB1 pixel_100/VBIAS pixel_100/NB2 pixel_100/AMP_IN pixel_100/SF_IB pixel_100/PIX_OUT
+ pixel_100/CSA_VREF pixel
Xpixel_4105 pixel_4105/gring pixel_4105/VDD pixel_4105/GND pixel_4105/VREF pixel_4105/ROW_SEL
+ pixel_4105/NB1 pixel_4105/VBIAS pixel_4105/NB2 pixel_4105/AMP_IN pixel_4105/SF_IB
+ pixel_4105/PIX_OUT pixel_4105/CSA_VREF pixel
Xpixel_4116 pixel_4116/gring pixel_4116/VDD pixel_4116/GND pixel_4116/VREF pixel_4116/ROW_SEL
+ pixel_4116/NB1 pixel_4116/VBIAS pixel_4116/NB2 pixel_4116/AMP_IN pixel_4116/SF_IB
+ pixel_4116/PIX_OUT pixel_4116/CSA_VREF pixel
Xpixel_155 pixel_155/gring pixel_155/VDD pixel_155/GND pixel_155/VREF pixel_155/ROW_SEL
+ pixel_155/NB1 pixel_155/VBIAS pixel_155/NB2 pixel_155/AMP_IN pixel_155/SF_IB pixel_155/PIX_OUT
+ pixel_155/CSA_VREF pixel
Xpixel_144 pixel_144/gring pixel_144/VDD pixel_144/GND pixel_144/VREF pixel_144/ROW_SEL
+ pixel_144/NB1 pixel_144/VBIAS pixel_144/NB2 pixel_144/AMP_IN pixel_144/SF_IB pixel_144/PIX_OUT
+ pixel_144/CSA_VREF pixel
Xpixel_133 pixel_133/gring pixel_133/VDD pixel_133/GND pixel_133/VREF pixel_133/ROW_SEL
+ pixel_133/NB1 pixel_133/VBIAS pixel_133/NB2 pixel_133/AMP_IN pixel_133/SF_IB pixel_133/PIX_OUT
+ pixel_133/CSA_VREF pixel
Xpixel_3415 pixel_3415/gring pixel_3415/VDD pixel_3415/GND pixel_3415/VREF pixel_3415/ROW_SEL
+ pixel_3415/NB1 pixel_3415/VBIAS pixel_3415/NB2 pixel_3415/AMP_IN pixel_3415/SF_IB
+ pixel_3415/PIX_OUT pixel_3415/CSA_VREF pixel
Xpixel_3404 pixel_3404/gring pixel_3404/VDD pixel_3404/GND pixel_3404/VREF pixel_3404/ROW_SEL
+ pixel_3404/NB1 pixel_3404/VBIAS pixel_3404/NB2 pixel_3404/AMP_IN pixel_3404/SF_IB
+ pixel_3404/PIX_OUT pixel_3404/CSA_VREF pixel
Xpixel_4127 pixel_4127/gring pixel_4127/VDD pixel_4127/GND pixel_4127/VREF pixel_4127/ROW_SEL
+ pixel_4127/NB1 pixel_4127/VBIAS pixel_4127/NB2 pixel_4127/AMP_IN pixel_4127/SF_IB
+ pixel_4127/PIX_OUT pixel_4127/CSA_VREF pixel
Xpixel_4138 pixel_4138/gring pixel_4138/VDD pixel_4138/GND pixel_4138/VREF pixel_4138/ROW_SEL
+ pixel_4138/NB1 pixel_4138/VBIAS pixel_4138/NB2 pixel_4138/AMP_IN pixel_4138/SF_IB
+ pixel_4138/PIX_OUT pixel_4138/CSA_VREF pixel
Xpixel_4149 pixel_4149/gring pixel_4149/VDD pixel_4149/GND pixel_4149/VREF pixel_4149/ROW_SEL
+ pixel_4149/NB1 pixel_4149/VBIAS pixel_4149/NB2 pixel_4149/AMP_IN pixel_4149/SF_IB
+ pixel_4149/PIX_OUT pixel_4149/CSA_VREF pixel
Xpixel_188 pixel_188/gring pixel_188/VDD pixel_188/GND pixel_188/VREF pixel_188/ROW_SEL
+ pixel_188/NB1 pixel_188/VBIAS pixel_188/NB2 pixel_188/AMP_IN pixel_188/SF_IB pixel_188/PIX_OUT
+ pixel_188/CSA_VREF pixel
Xpixel_177 pixel_177/gring pixel_177/VDD pixel_177/GND pixel_177/VREF pixel_177/ROW_SEL
+ pixel_177/NB1 pixel_177/VBIAS pixel_177/NB2 pixel_177/AMP_IN pixel_177/SF_IB pixel_177/PIX_OUT
+ pixel_177/CSA_VREF pixel
Xpixel_166 pixel_166/gring pixel_166/VDD pixel_166/GND pixel_166/VREF pixel_166/ROW_SEL
+ pixel_166/NB1 pixel_166/VBIAS pixel_166/NB2 pixel_166/AMP_IN pixel_166/SF_IB pixel_166/PIX_OUT
+ pixel_166/CSA_VREF pixel
Xpixel_2703 pixel_2703/gring pixel_2703/VDD pixel_2703/GND pixel_2703/VREF pixel_2703/ROW_SEL
+ pixel_2703/NB1 pixel_2703/VBIAS pixel_2703/NB2 pixel_2703/AMP_IN pixel_2703/SF_IB
+ pixel_2703/PIX_OUT pixel_2703/CSA_VREF pixel
Xpixel_3448 pixel_3448/gring pixel_3448/VDD pixel_3448/GND pixel_3448/VREF pixel_3448/ROW_SEL
+ pixel_3448/NB1 pixel_3448/VBIAS pixel_3448/NB2 pixel_3448/AMP_IN pixel_3448/SF_IB
+ pixel_3448/PIX_OUT pixel_3448/CSA_VREF pixel
Xpixel_3437 pixel_3437/gring pixel_3437/VDD pixel_3437/GND pixel_3437/VREF pixel_3437/ROW_SEL
+ pixel_3437/NB1 pixel_3437/VBIAS pixel_3437/NB2 pixel_3437/AMP_IN pixel_3437/SF_IB
+ pixel_3437/PIX_OUT pixel_3437/CSA_VREF pixel
Xpixel_3426 pixel_3426/gring pixel_3426/VDD pixel_3426/GND pixel_3426/VREF pixel_3426/ROW_SEL
+ pixel_3426/NB1 pixel_3426/VBIAS pixel_3426/NB2 pixel_3426/AMP_IN pixel_3426/SF_IB
+ pixel_3426/PIX_OUT pixel_3426/CSA_VREF pixel
Xpixel_199 pixel_199/gring pixel_199/VDD pixel_199/GND pixel_199/VREF pixel_199/ROW_SEL
+ pixel_199/NB1 pixel_199/VBIAS pixel_199/NB2 pixel_199/AMP_IN pixel_199/SF_IB pixel_199/PIX_OUT
+ pixel_199/CSA_VREF pixel
Xpixel_2747 pixel_2747/gring pixel_2747/VDD pixel_2747/GND pixel_2747/VREF pixel_2747/ROW_SEL
+ pixel_2747/NB1 pixel_2747/VBIAS pixel_2747/NB2 pixel_2747/AMP_IN pixel_2747/SF_IB
+ pixel_2747/PIX_OUT pixel_2747/CSA_VREF pixel
Xpixel_2736 pixel_2736/gring pixel_2736/VDD pixel_2736/GND pixel_2736/VREF pixel_2736/ROW_SEL
+ pixel_2736/NB1 pixel_2736/VBIAS pixel_2736/NB2 pixel_2736/AMP_IN pixel_2736/SF_IB
+ pixel_2736/PIX_OUT pixel_2736/CSA_VREF pixel
Xpixel_2725 pixel_2725/gring pixel_2725/VDD pixel_2725/GND pixel_2725/VREF pixel_2725/ROW_SEL
+ pixel_2725/NB1 pixel_2725/VBIAS pixel_2725/NB2 pixel_2725/AMP_IN pixel_2725/SF_IB
+ pixel_2725/PIX_OUT pixel_2725/CSA_VREF pixel
Xpixel_2714 pixel_2714/gring pixel_2714/VDD pixel_2714/GND pixel_2714/VREF pixel_2714/ROW_SEL
+ pixel_2714/NB1 pixel_2714/VBIAS pixel_2714/NB2 pixel_2714/AMP_IN pixel_2714/SF_IB
+ pixel_2714/PIX_OUT pixel_2714/CSA_VREF pixel
Xpixel_3459 pixel_3459/gring pixel_3459/VDD pixel_3459/GND pixel_3459/VREF pixel_3459/ROW_SEL
+ pixel_3459/NB1 pixel_3459/VBIAS pixel_3459/NB2 pixel_3459/AMP_IN pixel_3459/SF_IB
+ pixel_3459/PIX_OUT pixel_3459/CSA_VREF pixel
Xpixel_2769 pixel_2769/gring pixel_2769/VDD pixel_2769/GND pixel_2769/VREF pixel_2769/ROW_SEL
+ pixel_2769/NB1 pixel_2769/VBIAS pixel_2769/NB2 pixel_2769/AMP_IN pixel_2769/SF_IB
+ pixel_2769/PIX_OUT pixel_2769/CSA_VREF pixel
Xpixel_2758 pixel_2758/gring pixel_2758/VDD pixel_2758/GND pixel_2758/VREF pixel_2758/ROW_SEL
+ pixel_2758/NB1 pixel_2758/VBIAS pixel_2758/NB2 pixel_2758/AMP_IN pixel_2758/SF_IB
+ pixel_2758/PIX_OUT pixel_2758/CSA_VREF pixel
Xpixel_6030 pixel_6030/gring pixel_6030/VDD pixel_6030/GND pixel_6030/VREF pixel_6030/ROW_SEL
+ pixel_6030/NB1 pixel_6030/VBIAS pixel_6030/NB2 pixel_6030/AMP_IN pixel_6030/SF_IB
+ pixel_6030/PIX_OUT pixel_6030/CSA_VREF pixel
Xpixel_6041 pixel_6041/gring pixel_6041/VDD pixel_6041/GND pixel_6041/VREF pixel_6041/ROW_SEL
+ pixel_6041/NB1 pixel_6041/VBIAS pixel_6041/NB2 pixel_6041/AMP_IN pixel_6041/SF_IB
+ pixel_6041/PIX_OUT pixel_6041/CSA_VREF pixel
Xpixel_6052 pixel_6052/gring pixel_6052/VDD pixel_6052/GND pixel_6052/VREF pixel_6052/ROW_SEL
+ pixel_6052/NB1 pixel_6052/VBIAS pixel_6052/NB2 pixel_6052/AMP_IN pixel_6052/SF_IB
+ pixel_6052/PIX_OUT pixel_6052/CSA_VREF pixel
Xpixel_6063 pixel_6063/gring pixel_6063/VDD pixel_6063/GND pixel_6063/VREF pixel_6063/ROW_SEL
+ pixel_6063/NB1 pixel_6063/VBIAS pixel_6063/NB2 pixel_6063/AMP_IN pixel_6063/SF_IB
+ pixel_6063/PIX_OUT pixel_6063/CSA_VREF pixel
Xpixel_6074 pixel_6074/gring pixel_6074/VDD pixel_6074/GND pixel_6074/VREF pixel_6074/ROW_SEL
+ pixel_6074/NB1 pixel_6074/VBIAS pixel_6074/NB2 pixel_6074/AMP_IN pixel_6074/SF_IB
+ pixel_6074/PIX_OUT pixel_6074/CSA_VREF pixel
Xpixel_6085 pixel_6085/gring pixel_6085/VDD pixel_6085/GND pixel_6085/VREF pixel_6085/ROW_SEL
+ pixel_6085/NB1 pixel_6085/VBIAS pixel_6085/NB2 pixel_6085/AMP_IN pixel_6085/SF_IB
+ pixel_6085/PIX_OUT pixel_6085/CSA_VREF pixel
Xpixel_5340 pixel_5340/gring pixel_5340/VDD pixel_5340/GND pixel_5340/VREF pixel_5340/ROW_SEL
+ pixel_5340/NB1 pixel_5340/VBIAS pixel_5340/NB2 pixel_5340/AMP_IN pixel_5340/SF_IB
+ pixel_5340/PIX_OUT pixel_5340/CSA_VREF pixel
Xpixel_5351 pixel_5351/gring pixel_5351/VDD pixel_5351/GND pixel_5351/VREF pixel_5351/ROW_SEL
+ pixel_5351/NB1 pixel_5351/VBIAS pixel_5351/NB2 pixel_5351/AMP_IN pixel_5351/SF_IB
+ pixel_5351/PIX_OUT pixel_5351/CSA_VREF pixel
Xpixel_6096 pixel_6096/gring pixel_6096/VDD pixel_6096/GND pixel_6096/VREF pixel_6096/ROW_SEL
+ pixel_6096/NB1 pixel_6096/VBIAS pixel_6096/NB2 pixel_6096/AMP_IN pixel_6096/SF_IB
+ pixel_6096/PIX_OUT pixel_6096/CSA_VREF pixel
Xpixel_5362 pixel_5362/gring pixel_5362/VDD pixel_5362/GND pixel_5362/VREF pixel_5362/ROW_SEL
+ pixel_5362/NB1 pixel_5362/VBIAS pixel_5362/NB2 pixel_5362/AMP_IN pixel_5362/SF_IB
+ pixel_5362/PIX_OUT pixel_5362/CSA_VREF pixel
Xpixel_5373 pixel_5373/gring pixel_5373/VDD pixel_5373/GND pixel_5373/VREF pixel_5373/ROW_SEL
+ pixel_5373/NB1 pixel_5373/VBIAS pixel_5373/NB2 pixel_5373/AMP_IN pixel_5373/SF_IB
+ pixel_5373/PIX_OUT pixel_5373/CSA_VREF pixel
Xpixel_5384 pixel_5384/gring pixel_5384/VDD pixel_5384/GND pixel_5384/VREF pixel_5384/ROW_SEL
+ pixel_5384/NB1 pixel_5384/VBIAS pixel_5384/NB2 pixel_5384/AMP_IN pixel_5384/SF_IB
+ pixel_5384/PIX_OUT pixel_5384/CSA_VREF pixel
Xpixel_5395 pixel_5395/gring pixel_5395/VDD pixel_5395/GND pixel_5395/VREF pixel_5395/ROW_SEL
+ pixel_5395/NB1 pixel_5395/VBIAS pixel_5395/NB2 pixel_5395/AMP_IN pixel_5395/SF_IB
+ pixel_5395/PIX_OUT pixel_5395/CSA_VREF pixel
Xpixel_4650 pixel_4650/gring pixel_4650/VDD pixel_4650/GND pixel_4650/VREF pixel_4650/ROW_SEL
+ pixel_4650/NB1 pixel_4650/VBIAS pixel_4650/NB2 pixel_4650/AMP_IN pixel_4650/SF_IB
+ pixel_4650/PIX_OUT pixel_4650/CSA_VREF pixel
Xpixel_4661 pixel_4661/gring pixel_4661/VDD pixel_4661/GND pixel_4661/VREF pixel_4661/ROW_SEL
+ pixel_4661/NB1 pixel_4661/VBIAS pixel_4661/NB2 pixel_4661/AMP_IN pixel_4661/SF_IB
+ pixel_4661/PIX_OUT pixel_4661/CSA_VREF pixel
Xpixel_4672 pixel_4672/gring pixel_4672/VDD pixel_4672/GND pixel_4672/VREF pixel_4672/ROW_SEL
+ pixel_4672/NB1 pixel_4672/VBIAS pixel_4672/NB2 pixel_4672/AMP_IN pixel_4672/SF_IB
+ pixel_4672/PIX_OUT pixel_4672/CSA_VREF pixel
Xpixel_4683 pixel_4683/gring pixel_4683/VDD pixel_4683/GND pixel_4683/VREF pixel_4683/ROW_SEL
+ pixel_4683/NB1 pixel_4683/VBIAS pixel_4683/NB2 pixel_4683/AMP_IN pixel_4683/SF_IB
+ pixel_4683/PIX_OUT pixel_4683/CSA_VREF pixel
Xpixel_4694 pixel_4694/gring pixel_4694/VDD pixel_4694/GND pixel_4694/VREF pixel_4694/ROW_SEL
+ pixel_4694/NB1 pixel_4694/VBIAS pixel_4694/NB2 pixel_4694/AMP_IN pixel_4694/SF_IB
+ pixel_4694/PIX_OUT pixel_4694/CSA_VREF pixel
Xpixel_3960 pixel_3960/gring pixel_3960/VDD pixel_3960/GND pixel_3960/VREF pixel_3960/ROW_SEL
+ pixel_3960/NB1 pixel_3960/VBIAS pixel_3960/NB2 pixel_3960/AMP_IN pixel_3960/SF_IB
+ pixel_3960/PIX_OUT pixel_3960/CSA_VREF pixel
Xpixel_3971 pixel_3971/gring pixel_3971/VDD pixel_3971/GND pixel_3971/VREF pixel_3971/ROW_SEL
+ pixel_3971/NB1 pixel_3971/VBIAS pixel_3971/NB2 pixel_3971/AMP_IN pixel_3971/SF_IB
+ pixel_3971/PIX_OUT pixel_3971/CSA_VREF pixel
Xpixel_3982 pixel_3982/gring pixel_3982/VDD pixel_3982/GND pixel_3982/VREF pixel_3982/ROW_SEL
+ pixel_3982/NB1 pixel_3982/VBIAS pixel_3982/NB2 pixel_3982/AMP_IN pixel_3982/SF_IB
+ pixel_3982/PIX_OUT pixel_3982/CSA_VREF pixel
Xpixel_3993 pixel_3993/gring pixel_3993/VDD pixel_3993/GND pixel_3993/VREF pixel_3993/ROW_SEL
+ pixel_3993/NB1 pixel_3993/VBIAS pixel_3993/NB2 pixel_3993/AMP_IN pixel_3993/SF_IB
+ pixel_3993/PIX_OUT pixel_3993/CSA_VREF pixel
Xpixel_3 pixel_3/gring pixel_3/VDD pixel_3/GND pixel_3/VREF pixel_3/ROW_SEL pixel_3/NB1
+ pixel_3/VBIAS pixel_3/NB2 pixel_3/AMP_IN pixel_3/SF_IB pixel_3/PIX_OUT pixel_3/CSA_VREF
+ pixel
Xpixel_1309 pixel_1309/gring pixel_1309/VDD pixel_1309/GND pixel_1309/VREF pixel_1309/ROW_SEL
+ pixel_1309/NB1 pixel_1309/VBIAS pixel_1309/NB2 pixel_1309/AMP_IN pixel_1309/SF_IB
+ pixel_1309/PIX_OUT pixel_1309/CSA_VREF pixel
Xpixel_9606 pixel_9606/gring pixel_9606/VDD pixel_9606/GND pixel_9606/VREF pixel_9606/ROW_SEL
+ pixel_9606/NB1 pixel_9606/VBIAS pixel_9606/NB2 pixel_9606/AMP_IN pixel_9606/SF_IB
+ pixel_9606/PIX_OUT pixel_9606/CSA_VREF pixel
Xpixel_9617 pixel_9617/gring pixel_9617/VDD pixel_9617/GND pixel_9617/VREF pixel_9617/ROW_SEL
+ pixel_9617/NB1 pixel_9617/VBIAS pixel_9617/NB2 pixel_9617/AMP_IN pixel_9617/SF_IB
+ pixel_9617/PIX_OUT pixel_9617/CSA_VREF pixel
Xpixel_9628 pixel_9628/gring pixel_9628/VDD pixel_9628/GND pixel_9628/VREF pixel_9628/ROW_SEL
+ pixel_9628/NB1 pixel_9628/VBIAS pixel_9628/NB2 pixel_9628/AMP_IN pixel_9628/SF_IB
+ pixel_9628/PIX_OUT pixel_9628/CSA_VREF pixel
Xpixel_9639 pixel_9639/gring pixel_9639/VDD pixel_9639/GND pixel_9639/VREF pixel_9639/ROW_SEL
+ pixel_9639/NB1 pixel_9639/VBIAS pixel_9639/NB2 pixel_9639/AMP_IN pixel_9639/SF_IB
+ pixel_9639/PIX_OUT pixel_9639/CSA_VREF pixel
Xpixel_8927 pixel_8927/gring pixel_8927/VDD pixel_8927/GND pixel_8927/VREF pixel_8927/ROW_SEL
+ pixel_8927/NB1 pixel_8927/VBIAS pixel_8927/NB2 pixel_8927/AMP_IN pixel_8927/SF_IB
+ pixel_8927/PIX_OUT pixel_8927/CSA_VREF pixel
Xpixel_8916 pixel_8916/gring pixel_8916/VDD pixel_8916/GND pixel_8916/VREF pixel_8916/ROW_SEL
+ pixel_8916/NB1 pixel_8916/VBIAS pixel_8916/NB2 pixel_8916/AMP_IN pixel_8916/SF_IB
+ pixel_8916/PIX_OUT pixel_8916/CSA_VREF pixel
Xpixel_8905 pixel_8905/gring pixel_8905/VDD pixel_8905/GND pixel_8905/VREF pixel_8905/ROW_SEL
+ pixel_8905/NB1 pixel_8905/VBIAS pixel_8905/NB2 pixel_8905/AMP_IN pixel_8905/SF_IB
+ pixel_8905/PIX_OUT pixel_8905/CSA_VREF pixel
Xpixel_8949 pixel_8949/gring pixel_8949/VDD pixel_8949/GND pixel_8949/VREF pixel_8949/ROW_SEL
+ pixel_8949/NB1 pixel_8949/VBIAS pixel_8949/NB2 pixel_8949/AMP_IN pixel_8949/SF_IB
+ pixel_8949/PIX_OUT pixel_8949/CSA_VREF pixel
Xpixel_8938 pixel_8938/gring pixel_8938/VDD pixel_8938/GND pixel_8938/VREF pixel_8938/ROW_SEL
+ pixel_8938/NB1 pixel_8938/VBIAS pixel_8938/NB2 pixel_8938/AMP_IN pixel_8938/SF_IB
+ pixel_8938/PIX_OUT pixel_8938/CSA_VREF pixel
Xpixel_3223 pixel_3223/gring pixel_3223/VDD pixel_3223/GND pixel_3223/VREF pixel_3223/ROW_SEL
+ pixel_3223/NB1 pixel_3223/VBIAS pixel_3223/NB2 pixel_3223/AMP_IN pixel_3223/SF_IB
+ pixel_3223/PIX_OUT pixel_3223/CSA_VREF pixel
Xpixel_3212 pixel_3212/gring pixel_3212/VDD pixel_3212/GND pixel_3212/VREF pixel_3212/ROW_SEL
+ pixel_3212/NB1 pixel_3212/VBIAS pixel_3212/NB2 pixel_3212/AMP_IN pixel_3212/SF_IB
+ pixel_3212/PIX_OUT pixel_3212/CSA_VREF pixel
Xpixel_3201 pixel_3201/gring pixel_3201/VDD pixel_3201/GND pixel_3201/VREF pixel_3201/ROW_SEL
+ pixel_3201/NB1 pixel_3201/VBIAS pixel_3201/NB2 pixel_3201/AMP_IN pixel_3201/SF_IB
+ pixel_3201/PIX_OUT pixel_3201/CSA_VREF pixel
Xpixel_2522 pixel_2522/gring pixel_2522/VDD pixel_2522/GND pixel_2522/VREF pixel_2522/ROW_SEL
+ pixel_2522/NB1 pixel_2522/VBIAS pixel_2522/NB2 pixel_2522/AMP_IN pixel_2522/SF_IB
+ pixel_2522/PIX_OUT pixel_2522/CSA_VREF pixel
Xpixel_2511 pixel_2511/gring pixel_2511/VDD pixel_2511/GND pixel_2511/VREF pixel_2511/ROW_SEL
+ pixel_2511/NB1 pixel_2511/VBIAS pixel_2511/NB2 pixel_2511/AMP_IN pixel_2511/SF_IB
+ pixel_2511/PIX_OUT pixel_2511/CSA_VREF pixel
Xpixel_2500 pixel_2500/gring pixel_2500/VDD pixel_2500/GND pixel_2500/VREF pixel_2500/ROW_SEL
+ pixel_2500/NB1 pixel_2500/VBIAS pixel_2500/NB2 pixel_2500/AMP_IN pixel_2500/SF_IB
+ pixel_2500/PIX_OUT pixel_2500/CSA_VREF pixel
Xpixel_3256 pixel_3256/gring pixel_3256/VDD pixel_3256/GND pixel_3256/VREF pixel_3256/ROW_SEL
+ pixel_3256/NB1 pixel_3256/VBIAS pixel_3256/NB2 pixel_3256/AMP_IN pixel_3256/SF_IB
+ pixel_3256/PIX_OUT pixel_3256/CSA_VREF pixel
Xpixel_3245 pixel_3245/gring pixel_3245/VDD pixel_3245/GND pixel_3245/VREF pixel_3245/ROW_SEL
+ pixel_3245/NB1 pixel_3245/VBIAS pixel_3245/NB2 pixel_3245/AMP_IN pixel_3245/SF_IB
+ pixel_3245/PIX_OUT pixel_3245/CSA_VREF pixel
Xpixel_3234 pixel_3234/gring pixel_3234/VDD pixel_3234/GND pixel_3234/VREF pixel_3234/ROW_SEL
+ pixel_3234/NB1 pixel_3234/VBIAS pixel_3234/NB2 pixel_3234/AMP_IN pixel_3234/SF_IB
+ pixel_3234/PIX_OUT pixel_3234/CSA_VREF pixel
Xpixel_1810 pixel_1810/gring pixel_1810/VDD pixel_1810/GND pixel_1810/VREF pixel_1810/ROW_SEL
+ pixel_1810/NB1 pixel_1810/VBIAS pixel_1810/NB2 pixel_1810/AMP_IN pixel_1810/SF_IB
+ pixel_1810/PIX_OUT pixel_1810/CSA_VREF pixel
Xpixel_2555 pixel_2555/gring pixel_2555/VDD pixel_2555/GND pixel_2555/VREF pixel_2555/ROW_SEL
+ pixel_2555/NB1 pixel_2555/VBIAS pixel_2555/NB2 pixel_2555/AMP_IN pixel_2555/SF_IB
+ pixel_2555/PIX_OUT pixel_2555/CSA_VREF pixel
Xpixel_2544 pixel_2544/gring pixel_2544/VDD pixel_2544/GND pixel_2544/VREF pixel_2544/ROW_SEL
+ pixel_2544/NB1 pixel_2544/VBIAS pixel_2544/NB2 pixel_2544/AMP_IN pixel_2544/SF_IB
+ pixel_2544/PIX_OUT pixel_2544/CSA_VREF pixel
Xpixel_2533 pixel_2533/gring pixel_2533/VDD pixel_2533/GND pixel_2533/VREF pixel_2533/ROW_SEL
+ pixel_2533/NB1 pixel_2533/VBIAS pixel_2533/NB2 pixel_2533/AMP_IN pixel_2533/SF_IB
+ pixel_2533/PIX_OUT pixel_2533/CSA_VREF pixel
Xpixel_3289 pixel_3289/gring pixel_3289/VDD pixel_3289/GND pixel_3289/VREF pixel_3289/ROW_SEL
+ pixel_3289/NB1 pixel_3289/VBIAS pixel_3289/NB2 pixel_3289/AMP_IN pixel_3289/SF_IB
+ pixel_3289/PIX_OUT pixel_3289/CSA_VREF pixel
Xpixel_3278 pixel_3278/gring pixel_3278/VDD pixel_3278/GND pixel_3278/VREF pixel_3278/ROW_SEL
+ pixel_3278/NB1 pixel_3278/VBIAS pixel_3278/NB2 pixel_3278/AMP_IN pixel_3278/SF_IB
+ pixel_3278/PIX_OUT pixel_3278/CSA_VREF pixel
Xpixel_3267 pixel_3267/gring pixel_3267/VDD pixel_3267/GND pixel_3267/VREF pixel_3267/ROW_SEL
+ pixel_3267/NB1 pixel_3267/VBIAS pixel_3267/NB2 pixel_3267/AMP_IN pixel_3267/SF_IB
+ pixel_3267/PIX_OUT pixel_3267/CSA_VREF pixel
Xpixel_1843 pixel_1843/gring pixel_1843/VDD pixel_1843/GND pixel_1843/VREF pixel_1843/ROW_SEL
+ pixel_1843/NB1 pixel_1843/VBIAS pixel_1843/NB2 pixel_1843/AMP_IN pixel_1843/SF_IB
+ pixel_1843/PIX_OUT pixel_1843/CSA_VREF pixel
Xpixel_1832 pixel_1832/gring pixel_1832/VDD pixel_1832/GND pixel_1832/VREF pixel_1832/ROW_SEL
+ pixel_1832/NB1 pixel_1832/VBIAS pixel_1832/NB2 pixel_1832/AMP_IN pixel_1832/SF_IB
+ pixel_1832/PIX_OUT pixel_1832/CSA_VREF pixel
Xpixel_1821 pixel_1821/gring pixel_1821/VDD pixel_1821/GND pixel_1821/VREF pixel_1821/ROW_SEL
+ pixel_1821/NB1 pixel_1821/VBIAS pixel_1821/NB2 pixel_1821/AMP_IN pixel_1821/SF_IB
+ pixel_1821/PIX_OUT pixel_1821/CSA_VREF pixel
Xpixel_2588 pixel_2588/gring pixel_2588/VDD pixel_2588/GND pixel_2588/VREF pixel_2588/ROW_SEL
+ pixel_2588/NB1 pixel_2588/VBIAS pixel_2588/NB2 pixel_2588/AMP_IN pixel_2588/SF_IB
+ pixel_2588/PIX_OUT pixel_2588/CSA_VREF pixel
Xpixel_2577 pixel_2577/gring pixel_2577/VDD pixel_2577/GND pixel_2577/VREF pixel_2577/ROW_SEL
+ pixel_2577/NB1 pixel_2577/VBIAS pixel_2577/NB2 pixel_2577/AMP_IN pixel_2577/SF_IB
+ pixel_2577/PIX_OUT pixel_2577/CSA_VREF pixel
Xpixel_2566 pixel_2566/gring pixel_2566/VDD pixel_2566/GND pixel_2566/VREF pixel_2566/ROW_SEL
+ pixel_2566/NB1 pixel_2566/VBIAS pixel_2566/NB2 pixel_2566/AMP_IN pixel_2566/SF_IB
+ pixel_2566/PIX_OUT pixel_2566/CSA_VREF pixel
Xpixel_1887 pixel_1887/gring pixel_1887/VDD pixel_1887/GND pixel_1887/VREF pixel_1887/ROW_SEL
+ pixel_1887/NB1 pixel_1887/VBIAS pixel_1887/NB2 pixel_1887/AMP_IN pixel_1887/SF_IB
+ pixel_1887/PIX_OUT pixel_1887/CSA_VREF pixel
Xpixel_1876 pixel_1876/gring pixel_1876/VDD pixel_1876/GND pixel_1876/VREF pixel_1876/ROW_SEL
+ pixel_1876/NB1 pixel_1876/VBIAS pixel_1876/NB2 pixel_1876/AMP_IN pixel_1876/SF_IB
+ pixel_1876/PIX_OUT pixel_1876/CSA_VREF pixel
Xpixel_1865 pixel_1865/gring pixel_1865/VDD pixel_1865/GND pixel_1865/VREF pixel_1865/ROW_SEL
+ pixel_1865/NB1 pixel_1865/VBIAS pixel_1865/NB2 pixel_1865/AMP_IN pixel_1865/SF_IB
+ pixel_1865/PIX_OUT pixel_1865/CSA_VREF pixel
Xpixel_1854 pixel_1854/gring pixel_1854/VDD pixel_1854/GND pixel_1854/VREF pixel_1854/ROW_SEL
+ pixel_1854/NB1 pixel_1854/VBIAS pixel_1854/NB2 pixel_1854/AMP_IN pixel_1854/SF_IB
+ pixel_1854/PIX_OUT pixel_1854/CSA_VREF pixel
Xpixel_2599 pixel_2599/gring pixel_2599/VDD pixel_2599/GND pixel_2599/VREF pixel_2599/ROW_SEL
+ pixel_2599/NB1 pixel_2599/VBIAS pixel_2599/NB2 pixel_2599/AMP_IN pixel_2599/SF_IB
+ pixel_2599/PIX_OUT pixel_2599/CSA_VREF pixel
Xpixel_1898 pixel_1898/gring pixel_1898/VDD pixel_1898/GND pixel_1898/VREF pixel_1898/ROW_SEL
+ pixel_1898/NB1 pixel_1898/VBIAS pixel_1898/NB2 pixel_1898/AMP_IN pixel_1898/SF_IB
+ pixel_1898/PIX_OUT pixel_1898/CSA_VREF pixel
Xpixel_5170 pixel_5170/gring pixel_5170/VDD pixel_5170/GND pixel_5170/VREF pixel_5170/ROW_SEL
+ pixel_5170/NB1 pixel_5170/VBIAS pixel_5170/NB2 pixel_5170/AMP_IN pixel_5170/SF_IB
+ pixel_5170/PIX_OUT pixel_5170/CSA_VREF pixel
Xpixel_5181 pixel_5181/gring pixel_5181/VDD pixel_5181/GND pixel_5181/VREF pixel_5181/ROW_SEL
+ pixel_5181/NB1 pixel_5181/VBIAS pixel_5181/NB2 pixel_5181/AMP_IN pixel_5181/SF_IB
+ pixel_5181/PIX_OUT pixel_5181/CSA_VREF pixel
Xpixel_5192 pixel_5192/gring pixel_5192/VDD pixel_5192/GND pixel_5192/VREF pixel_5192/ROW_SEL
+ pixel_5192/NB1 pixel_5192/VBIAS pixel_5192/NB2 pixel_5192/AMP_IN pixel_5192/SF_IB
+ pixel_5192/PIX_OUT pixel_5192/CSA_VREF pixel
Xpixel_4480 pixel_4480/gring pixel_4480/VDD pixel_4480/GND pixel_4480/VREF pixel_4480/ROW_SEL
+ pixel_4480/NB1 pixel_4480/VBIAS pixel_4480/NB2 pixel_4480/AMP_IN pixel_4480/SF_IB
+ pixel_4480/PIX_OUT pixel_4480/CSA_VREF pixel
Xpixel_4491 pixel_4491/gring pixel_4491/VDD pixel_4491/GND pixel_4491/VREF pixel_4491/ROW_SEL
+ pixel_4491/NB1 pixel_4491/VBIAS pixel_4491/NB2 pixel_4491/AMP_IN pixel_4491/SF_IB
+ pixel_4491/PIX_OUT pixel_4491/CSA_VREF pixel
Xpixel_3790 pixel_3790/gring pixel_3790/VDD pixel_3790/GND pixel_3790/VREF pixel_3790/ROW_SEL
+ pixel_3790/NB1 pixel_3790/VBIAS pixel_3790/NB2 pixel_3790/AMP_IN pixel_3790/SF_IB
+ pixel_3790/PIX_OUT pixel_3790/CSA_VREF pixel
Xpixel_1106 pixel_1106/gring pixel_1106/VDD pixel_1106/GND pixel_1106/VREF pixel_1106/ROW_SEL
+ pixel_1106/NB1 pixel_1106/VBIAS pixel_1106/NB2 pixel_1106/AMP_IN pixel_1106/SF_IB
+ pixel_1106/PIX_OUT pixel_1106/CSA_VREF pixel
Xpixel_1139 pixel_1139/gring pixel_1139/VDD pixel_1139/GND pixel_1139/VREF pixel_1139/ROW_SEL
+ pixel_1139/NB1 pixel_1139/VBIAS pixel_1139/NB2 pixel_1139/AMP_IN pixel_1139/SF_IB
+ pixel_1139/PIX_OUT pixel_1139/CSA_VREF pixel
Xpixel_1128 pixel_1128/gring pixel_1128/VDD pixel_1128/GND pixel_1128/VREF pixel_1128/ROW_SEL
+ pixel_1128/NB1 pixel_1128/VBIAS pixel_1128/NB2 pixel_1128/AMP_IN pixel_1128/SF_IB
+ pixel_1128/PIX_OUT pixel_1128/CSA_VREF pixel
Xpixel_1117 pixel_1117/gring pixel_1117/VDD pixel_1117/GND pixel_1117/VREF pixel_1117/ROW_SEL
+ pixel_1117/NB1 pixel_1117/VBIAS pixel_1117/NB2 pixel_1117/AMP_IN pixel_1117/SF_IB
+ pixel_1117/PIX_OUT pixel_1117/CSA_VREF pixel
Xpixel_9414 pixel_9414/gring pixel_9414/VDD pixel_9414/GND pixel_9414/VREF pixel_9414/ROW_SEL
+ pixel_9414/NB1 pixel_9414/VBIAS pixel_9414/NB2 pixel_9414/AMP_IN pixel_9414/SF_IB
+ pixel_9414/PIX_OUT pixel_9414/CSA_VREF pixel
Xpixel_9403 pixel_9403/gring pixel_9403/VDD pixel_9403/GND pixel_9403/VREF pixel_9403/ROW_SEL
+ pixel_9403/NB1 pixel_9403/VBIAS pixel_9403/NB2 pixel_9403/AMP_IN pixel_9403/SF_IB
+ pixel_9403/PIX_OUT pixel_9403/CSA_VREF pixel
Xpixel_8702 pixel_8702/gring pixel_8702/VDD pixel_8702/GND pixel_8702/VREF pixel_8702/ROW_SEL
+ pixel_8702/NB1 pixel_8702/VBIAS pixel_8702/NB2 pixel_8702/AMP_IN pixel_8702/SF_IB
+ pixel_8702/PIX_OUT pixel_8702/CSA_VREF pixel
Xpixel_9447 pixel_9447/gring pixel_9447/VDD pixel_9447/GND pixel_9447/VREF pixel_9447/ROW_SEL
+ pixel_9447/NB1 pixel_9447/VBIAS pixel_9447/NB2 pixel_9447/AMP_IN pixel_9447/SF_IB
+ pixel_9447/PIX_OUT pixel_9447/CSA_VREF pixel
Xpixel_9436 pixel_9436/gring pixel_9436/VDD pixel_9436/GND pixel_9436/VREF pixel_9436/ROW_SEL
+ pixel_9436/NB1 pixel_9436/VBIAS pixel_9436/NB2 pixel_9436/AMP_IN pixel_9436/SF_IB
+ pixel_9436/PIX_OUT pixel_9436/CSA_VREF pixel
Xpixel_9425 pixel_9425/gring pixel_9425/VDD pixel_9425/GND pixel_9425/VREF pixel_9425/ROW_SEL
+ pixel_9425/NB1 pixel_9425/VBIAS pixel_9425/NB2 pixel_9425/AMP_IN pixel_9425/SF_IB
+ pixel_9425/PIX_OUT pixel_9425/CSA_VREF pixel
Xpixel_8735 pixel_8735/gring pixel_8735/VDD pixel_8735/GND pixel_8735/VREF pixel_8735/ROW_SEL
+ pixel_8735/NB1 pixel_8735/VBIAS pixel_8735/NB2 pixel_8735/AMP_IN pixel_8735/SF_IB
+ pixel_8735/PIX_OUT pixel_8735/CSA_VREF pixel
Xpixel_8724 pixel_8724/gring pixel_8724/VDD pixel_8724/GND pixel_8724/VREF pixel_8724/ROW_SEL
+ pixel_8724/NB1 pixel_8724/VBIAS pixel_8724/NB2 pixel_8724/AMP_IN pixel_8724/SF_IB
+ pixel_8724/PIX_OUT pixel_8724/CSA_VREF pixel
Xpixel_8713 pixel_8713/gring pixel_8713/VDD pixel_8713/GND pixel_8713/VREF pixel_8713/ROW_SEL
+ pixel_8713/NB1 pixel_8713/VBIAS pixel_8713/NB2 pixel_8713/AMP_IN pixel_8713/SF_IB
+ pixel_8713/PIX_OUT pixel_8713/CSA_VREF pixel
Xpixel_9469 pixel_9469/gring pixel_9469/VDD pixel_9469/GND pixel_9469/VREF pixel_9469/ROW_SEL
+ pixel_9469/NB1 pixel_9469/VBIAS pixel_9469/NB2 pixel_9469/AMP_IN pixel_9469/SF_IB
+ pixel_9469/PIX_OUT pixel_9469/CSA_VREF pixel
Xpixel_9458 pixel_9458/gring pixel_9458/VDD pixel_9458/GND pixel_9458/VREF pixel_9458/ROW_SEL
+ pixel_9458/NB1 pixel_9458/VBIAS pixel_9458/NB2 pixel_9458/AMP_IN pixel_9458/SF_IB
+ pixel_9458/PIX_OUT pixel_9458/CSA_VREF pixel
Xpixel_8779 pixel_8779/gring pixel_8779/VDD pixel_8779/GND pixel_8779/VREF pixel_8779/ROW_SEL
+ pixel_8779/NB1 pixel_8779/VBIAS pixel_8779/NB2 pixel_8779/AMP_IN pixel_8779/SF_IB
+ pixel_8779/PIX_OUT pixel_8779/CSA_VREF pixel
Xpixel_8768 pixel_8768/gring pixel_8768/VDD pixel_8768/GND pixel_8768/VREF pixel_8768/ROW_SEL
+ pixel_8768/NB1 pixel_8768/VBIAS pixel_8768/NB2 pixel_8768/AMP_IN pixel_8768/SF_IB
+ pixel_8768/PIX_OUT pixel_8768/CSA_VREF pixel
Xpixel_8757 pixel_8757/gring pixel_8757/VDD pixel_8757/GND pixel_8757/VREF pixel_8757/ROW_SEL
+ pixel_8757/NB1 pixel_8757/VBIAS pixel_8757/NB2 pixel_8757/AMP_IN pixel_8757/SF_IB
+ pixel_8757/PIX_OUT pixel_8757/CSA_VREF pixel
Xpixel_8746 pixel_8746/gring pixel_8746/VDD pixel_8746/GND pixel_8746/VREF pixel_8746/ROW_SEL
+ pixel_8746/NB1 pixel_8746/VBIAS pixel_8746/NB2 pixel_8746/AMP_IN pixel_8746/SF_IB
+ pixel_8746/PIX_OUT pixel_8746/CSA_VREF pixel
Xpixel_3031 pixel_3031/gring pixel_3031/VDD pixel_3031/GND pixel_3031/VREF pixel_3031/ROW_SEL
+ pixel_3031/NB1 pixel_3031/VBIAS pixel_3031/NB2 pixel_3031/AMP_IN pixel_3031/SF_IB
+ pixel_3031/PIX_OUT pixel_3031/CSA_VREF pixel
Xpixel_3020 pixel_3020/gring pixel_3020/VDD pixel_3020/GND pixel_3020/VREF pixel_3020/ROW_SEL
+ pixel_3020/NB1 pixel_3020/VBIAS pixel_3020/NB2 pixel_3020/AMP_IN pixel_3020/SF_IB
+ pixel_3020/PIX_OUT pixel_3020/CSA_VREF pixel
Xpixel_2330 pixel_2330/gring pixel_2330/VDD pixel_2330/GND pixel_2330/VREF pixel_2330/ROW_SEL
+ pixel_2330/NB1 pixel_2330/VBIAS pixel_2330/NB2 pixel_2330/AMP_IN pixel_2330/SF_IB
+ pixel_2330/PIX_OUT pixel_2330/CSA_VREF pixel
Xpixel_3075 pixel_3075/gring pixel_3075/VDD pixel_3075/GND pixel_3075/VREF pixel_3075/ROW_SEL
+ pixel_3075/NB1 pixel_3075/VBIAS pixel_3075/NB2 pixel_3075/AMP_IN pixel_3075/SF_IB
+ pixel_3075/PIX_OUT pixel_3075/CSA_VREF pixel
Xpixel_3064 pixel_3064/gring pixel_3064/VDD pixel_3064/GND pixel_3064/VREF pixel_3064/ROW_SEL
+ pixel_3064/NB1 pixel_3064/VBIAS pixel_3064/NB2 pixel_3064/AMP_IN pixel_3064/SF_IB
+ pixel_3064/PIX_OUT pixel_3064/CSA_VREF pixel
Xpixel_3053 pixel_3053/gring pixel_3053/VDD pixel_3053/GND pixel_3053/VREF pixel_3053/ROW_SEL
+ pixel_3053/NB1 pixel_3053/VBIAS pixel_3053/NB2 pixel_3053/AMP_IN pixel_3053/SF_IB
+ pixel_3053/PIX_OUT pixel_3053/CSA_VREF pixel
Xpixel_3042 pixel_3042/gring pixel_3042/VDD pixel_3042/GND pixel_3042/VREF pixel_3042/ROW_SEL
+ pixel_3042/NB1 pixel_3042/VBIAS pixel_3042/NB2 pixel_3042/AMP_IN pixel_3042/SF_IB
+ pixel_3042/PIX_OUT pixel_3042/CSA_VREF pixel
Xpixel_2363 pixel_2363/gring pixel_2363/VDD pixel_2363/GND pixel_2363/VREF pixel_2363/ROW_SEL
+ pixel_2363/NB1 pixel_2363/VBIAS pixel_2363/NB2 pixel_2363/AMP_IN pixel_2363/SF_IB
+ pixel_2363/PIX_OUT pixel_2363/CSA_VREF pixel
Xpixel_2352 pixel_2352/gring pixel_2352/VDD pixel_2352/GND pixel_2352/VREF pixel_2352/ROW_SEL
+ pixel_2352/NB1 pixel_2352/VBIAS pixel_2352/NB2 pixel_2352/AMP_IN pixel_2352/SF_IB
+ pixel_2352/PIX_OUT pixel_2352/CSA_VREF pixel
Xpixel_2341 pixel_2341/gring pixel_2341/VDD pixel_2341/GND pixel_2341/VREF pixel_2341/ROW_SEL
+ pixel_2341/NB1 pixel_2341/VBIAS pixel_2341/NB2 pixel_2341/AMP_IN pixel_2341/SF_IB
+ pixel_2341/PIX_OUT pixel_2341/CSA_VREF pixel
Xpixel_3097 pixel_3097/gring pixel_3097/VDD pixel_3097/GND pixel_3097/VREF pixel_3097/ROW_SEL
+ pixel_3097/NB1 pixel_3097/VBIAS pixel_3097/NB2 pixel_3097/AMP_IN pixel_3097/SF_IB
+ pixel_3097/PIX_OUT pixel_3097/CSA_VREF pixel
Xpixel_3086 pixel_3086/gring pixel_3086/VDD pixel_3086/GND pixel_3086/VREF pixel_3086/ROW_SEL
+ pixel_3086/NB1 pixel_3086/VBIAS pixel_3086/NB2 pixel_3086/AMP_IN pixel_3086/SF_IB
+ pixel_3086/PIX_OUT pixel_3086/CSA_VREF pixel
Xpixel_1651 pixel_1651/gring pixel_1651/VDD pixel_1651/GND pixel_1651/VREF pixel_1651/ROW_SEL
+ pixel_1651/NB1 pixel_1651/VBIAS pixel_1651/NB2 pixel_1651/AMP_IN pixel_1651/SF_IB
+ pixel_1651/PIX_OUT pixel_1651/CSA_VREF pixel
Xpixel_1640 pixel_1640/gring pixel_1640/VDD pixel_1640/GND pixel_1640/VREF pixel_1640/ROW_SEL
+ pixel_1640/NB1 pixel_1640/VBIAS pixel_1640/NB2 pixel_1640/AMP_IN pixel_1640/SF_IB
+ pixel_1640/PIX_OUT pixel_1640/CSA_VREF pixel
Xpixel_2396 pixel_2396/gring pixel_2396/VDD pixel_2396/GND pixel_2396/VREF pixel_2396/ROW_SEL
+ pixel_2396/NB1 pixel_2396/VBIAS pixel_2396/NB2 pixel_2396/AMP_IN pixel_2396/SF_IB
+ pixel_2396/PIX_OUT pixel_2396/CSA_VREF pixel
Xpixel_2385 pixel_2385/gring pixel_2385/VDD pixel_2385/GND pixel_2385/VREF pixel_2385/ROW_SEL
+ pixel_2385/NB1 pixel_2385/VBIAS pixel_2385/NB2 pixel_2385/AMP_IN pixel_2385/SF_IB
+ pixel_2385/PIX_OUT pixel_2385/CSA_VREF pixel
Xpixel_2374 pixel_2374/gring pixel_2374/VDD pixel_2374/GND pixel_2374/VREF pixel_2374/ROW_SEL
+ pixel_2374/NB1 pixel_2374/VBIAS pixel_2374/NB2 pixel_2374/AMP_IN pixel_2374/SF_IB
+ pixel_2374/PIX_OUT pixel_2374/CSA_VREF pixel
Xpixel_1695 pixel_1695/gring pixel_1695/VDD pixel_1695/GND pixel_1695/VREF pixel_1695/ROW_SEL
+ pixel_1695/NB1 pixel_1695/VBIAS pixel_1695/NB2 pixel_1695/AMP_IN pixel_1695/SF_IB
+ pixel_1695/PIX_OUT pixel_1695/CSA_VREF pixel
Xpixel_1684 pixel_1684/gring pixel_1684/VDD pixel_1684/GND pixel_1684/VREF pixel_1684/ROW_SEL
+ pixel_1684/NB1 pixel_1684/VBIAS pixel_1684/NB2 pixel_1684/AMP_IN pixel_1684/SF_IB
+ pixel_1684/PIX_OUT pixel_1684/CSA_VREF pixel
Xpixel_1673 pixel_1673/gring pixel_1673/VDD pixel_1673/GND pixel_1673/VREF pixel_1673/ROW_SEL
+ pixel_1673/NB1 pixel_1673/VBIAS pixel_1673/NB2 pixel_1673/AMP_IN pixel_1673/SF_IB
+ pixel_1673/PIX_OUT pixel_1673/CSA_VREF pixel
Xpixel_1662 pixel_1662/gring pixel_1662/VDD pixel_1662/GND pixel_1662/VREF pixel_1662/ROW_SEL
+ pixel_1662/NB1 pixel_1662/VBIAS pixel_1662/NB2 pixel_1662/AMP_IN pixel_1662/SF_IB
+ pixel_1662/PIX_OUT pixel_1662/CSA_VREF pixel
Xpixel_9970 pixel_9970/gring pixel_9970/VDD pixel_9970/GND pixel_9970/VREF pixel_9970/ROW_SEL
+ pixel_9970/NB1 pixel_9970/VBIAS pixel_9970/NB2 pixel_9970/AMP_IN pixel_9970/SF_IB
+ pixel_9970/PIX_OUT pixel_9970/CSA_VREF pixel
Xpixel_9981 pixel_9981/gring pixel_9981/VDD pixel_9981/GND pixel_9981/VREF pixel_9981/ROW_SEL
+ pixel_9981/NB1 pixel_9981/VBIAS pixel_9981/NB2 pixel_9981/AMP_IN pixel_9981/SF_IB
+ pixel_9981/PIX_OUT pixel_9981/CSA_VREF pixel
Xpixel_9992 pixel_9992/gring pixel_9992/VDD pixel_9992/GND pixel_9992/VREF pixel_9992/ROW_SEL
+ pixel_9992/NB1 pixel_9992/VBIAS pixel_9992/NB2 pixel_9992/AMP_IN pixel_9992/SF_IB
+ pixel_9992/PIX_OUT pixel_9992/CSA_VREF pixel
Xpixel_8009 pixel_8009/gring pixel_8009/VDD pixel_8009/GND pixel_8009/VREF pixel_8009/ROW_SEL
+ pixel_8009/NB1 pixel_8009/VBIAS pixel_8009/NB2 pixel_8009/AMP_IN pixel_8009/SF_IB
+ pixel_8009/PIX_OUT pixel_8009/CSA_VREF pixel
Xpixel_7308 pixel_7308/gring pixel_7308/VDD pixel_7308/GND pixel_7308/VREF pixel_7308/ROW_SEL
+ pixel_7308/NB1 pixel_7308/VBIAS pixel_7308/NB2 pixel_7308/AMP_IN pixel_7308/SF_IB
+ pixel_7308/PIX_OUT pixel_7308/CSA_VREF pixel
Xpixel_7319 pixel_7319/gring pixel_7319/VDD pixel_7319/GND pixel_7319/VREF pixel_7319/ROW_SEL
+ pixel_7319/NB1 pixel_7319/VBIAS pixel_7319/NB2 pixel_7319/AMP_IN pixel_7319/SF_IB
+ pixel_7319/PIX_OUT pixel_7319/CSA_VREF pixel
Xpixel_6607 pixel_6607/gring pixel_6607/VDD pixel_6607/GND pixel_6607/VREF pixel_6607/ROW_SEL
+ pixel_6607/NB1 pixel_6607/VBIAS pixel_6607/NB2 pixel_6607/AMP_IN pixel_6607/SF_IB
+ pixel_6607/PIX_OUT pixel_6607/CSA_VREF pixel
Xpixel_6618 pixel_6618/gring pixel_6618/VDD pixel_6618/GND pixel_6618/VREF pixel_6618/ROW_SEL
+ pixel_6618/NB1 pixel_6618/VBIAS pixel_6618/NB2 pixel_6618/AMP_IN pixel_6618/SF_IB
+ pixel_6618/PIX_OUT pixel_6618/CSA_VREF pixel
Xpixel_6629 pixel_6629/gring pixel_6629/VDD pixel_6629/GND pixel_6629/VREF pixel_6629/ROW_SEL
+ pixel_6629/NB1 pixel_6629/VBIAS pixel_6629/NB2 pixel_6629/AMP_IN pixel_6629/SF_IB
+ pixel_6629/PIX_OUT pixel_6629/CSA_VREF pixel
Xpixel_5906 pixel_5906/gring pixel_5906/VDD pixel_5906/GND pixel_5906/VREF pixel_5906/ROW_SEL
+ pixel_5906/NB1 pixel_5906/VBIAS pixel_5906/NB2 pixel_5906/AMP_IN pixel_5906/SF_IB
+ pixel_5906/PIX_OUT pixel_5906/CSA_VREF pixel
Xpixel_5917 pixel_5917/gring pixel_5917/VDD pixel_5917/GND pixel_5917/VREF pixel_5917/ROW_SEL
+ pixel_5917/NB1 pixel_5917/VBIAS pixel_5917/NB2 pixel_5917/AMP_IN pixel_5917/SF_IB
+ pixel_5917/PIX_OUT pixel_5917/CSA_VREF pixel
Xpixel_5928 pixel_5928/gring pixel_5928/VDD pixel_5928/GND pixel_5928/VREF pixel_5928/ROW_SEL
+ pixel_5928/NB1 pixel_5928/VBIAS pixel_5928/NB2 pixel_5928/AMP_IN pixel_5928/SF_IB
+ pixel_5928/PIX_OUT pixel_5928/CSA_VREF pixel
Xpixel_5939 pixel_5939/gring pixel_5939/VDD pixel_5939/GND pixel_5939/VREF pixel_5939/ROW_SEL
+ pixel_5939/NB1 pixel_5939/VBIAS pixel_5939/NB2 pixel_5939/AMP_IN pixel_5939/SF_IB
+ pixel_5939/PIX_OUT pixel_5939/CSA_VREF pixel
Xpixel_9222 pixel_9222/gring pixel_9222/VDD pixel_9222/GND pixel_9222/VREF pixel_9222/ROW_SEL
+ pixel_9222/NB1 pixel_9222/VBIAS pixel_9222/NB2 pixel_9222/AMP_IN pixel_9222/SF_IB
+ pixel_9222/PIX_OUT pixel_9222/CSA_VREF pixel
Xpixel_9211 pixel_9211/gring pixel_9211/VDD pixel_9211/GND pixel_9211/VREF pixel_9211/ROW_SEL
+ pixel_9211/NB1 pixel_9211/VBIAS pixel_9211/NB2 pixel_9211/AMP_IN pixel_9211/SF_IB
+ pixel_9211/PIX_OUT pixel_9211/CSA_VREF pixel
Xpixel_9200 pixel_9200/gring pixel_9200/VDD pixel_9200/GND pixel_9200/VREF pixel_9200/ROW_SEL
+ pixel_9200/NB1 pixel_9200/VBIAS pixel_9200/NB2 pixel_9200/AMP_IN pixel_9200/SF_IB
+ pixel_9200/PIX_OUT pixel_9200/CSA_VREF pixel
Xpixel_8510 pixel_8510/gring pixel_8510/VDD pixel_8510/GND pixel_8510/VREF pixel_8510/ROW_SEL
+ pixel_8510/NB1 pixel_8510/VBIAS pixel_8510/NB2 pixel_8510/AMP_IN pixel_8510/SF_IB
+ pixel_8510/PIX_OUT pixel_8510/CSA_VREF pixel
Xpixel_9255 pixel_9255/gring pixel_9255/VDD pixel_9255/GND pixel_9255/VREF pixel_9255/ROW_SEL
+ pixel_9255/NB1 pixel_9255/VBIAS pixel_9255/NB2 pixel_9255/AMP_IN pixel_9255/SF_IB
+ pixel_9255/PIX_OUT pixel_9255/CSA_VREF pixel
Xpixel_9244 pixel_9244/gring pixel_9244/VDD pixel_9244/GND pixel_9244/VREF pixel_9244/ROW_SEL
+ pixel_9244/NB1 pixel_9244/VBIAS pixel_9244/NB2 pixel_9244/AMP_IN pixel_9244/SF_IB
+ pixel_9244/PIX_OUT pixel_9244/CSA_VREF pixel
Xpixel_9233 pixel_9233/gring pixel_9233/VDD pixel_9233/GND pixel_9233/VREF pixel_9233/ROW_SEL
+ pixel_9233/NB1 pixel_9233/VBIAS pixel_9233/NB2 pixel_9233/AMP_IN pixel_9233/SF_IB
+ pixel_9233/PIX_OUT pixel_9233/CSA_VREF pixel
Xpixel_8554 pixel_8554/gring pixel_8554/VDD pixel_8554/GND pixel_8554/VREF pixel_8554/ROW_SEL
+ pixel_8554/NB1 pixel_8554/VBIAS pixel_8554/NB2 pixel_8554/AMP_IN pixel_8554/SF_IB
+ pixel_8554/PIX_OUT pixel_8554/CSA_VREF pixel
Xpixel_8543 pixel_8543/gring pixel_8543/VDD pixel_8543/GND pixel_8543/VREF pixel_8543/ROW_SEL
+ pixel_8543/NB1 pixel_8543/VBIAS pixel_8543/NB2 pixel_8543/AMP_IN pixel_8543/SF_IB
+ pixel_8543/PIX_OUT pixel_8543/CSA_VREF pixel
Xpixel_8532 pixel_8532/gring pixel_8532/VDD pixel_8532/GND pixel_8532/VREF pixel_8532/ROW_SEL
+ pixel_8532/NB1 pixel_8532/VBIAS pixel_8532/NB2 pixel_8532/AMP_IN pixel_8532/SF_IB
+ pixel_8532/PIX_OUT pixel_8532/CSA_VREF pixel
Xpixel_8521 pixel_8521/gring pixel_8521/VDD pixel_8521/GND pixel_8521/VREF pixel_8521/ROW_SEL
+ pixel_8521/NB1 pixel_8521/VBIAS pixel_8521/NB2 pixel_8521/AMP_IN pixel_8521/SF_IB
+ pixel_8521/PIX_OUT pixel_8521/CSA_VREF pixel
Xpixel_9288 pixel_9288/gring pixel_9288/VDD pixel_9288/GND pixel_9288/VREF pixel_9288/ROW_SEL
+ pixel_9288/NB1 pixel_9288/VBIAS pixel_9288/NB2 pixel_9288/AMP_IN pixel_9288/SF_IB
+ pixel_9288/PIX_OUT pixel_9288/CSA_VREF pixel
Xpixel_9277 pixel_9277/gring pixel_9277/VDD pixel_9277/GND pixel_9277/VREF pixel_9277/ROW_SEL
+ pixel_9277/NB1 pixel_9277/VBIAS pixel_9277/NB2 pixel_9277/AMP_IN pixel_9277/SF_IB
+ pixel_9277/PIX_OUT pixel_9277/CSA_VREF pixel
Xpixel_9266 pixel_9266/gring pixel_9266/VDD pixel_9266/GND pixel_9266/VREF pixel_9266/ROW_SEL
+ pixel_9266/NB1 pixel_9266/VBIAS pixel_9266/NB2 pixel_9266/AMP_IN pixel_9266/SF_IB
+ pixel_9266/PIX_OUT pixel_9266/CSA_VREF pixel
Xpixel_8587 pixel_8587/gring pixel_8587/VDD pixel_8587/GND pixel_8587/VREF pixel_8587/ROW_SEL
+ pixel_8587/NB1 pixel_8587/VBIAS pixel_8587/NB2 pixel_8587/AMP_IN pixel_8587/SF_IB
+ pixel_8587/PIX_OUT pixel_8587/CSA_VREF pixel
Xpixel_8576 pixel_8576/gring pixel_8576/VDD pixel_8576/GND pixel_8576/VREF pixel_8576/ROW_SEL
+ pixel_8576/NB1 pixel_8576/VBIAS pixel_8576/NB2 pixel_8576/AMP_IN pixel_8576/SF_IB
+ pixel_8576/PIX_OUT pixel_8576/CSA_VREF pixel
Xpixel_8565 pixel_8565/gring pixel_8565/VDD pixel_8565/GND pixel_8565/VREF pixel_8565/ROW_SEL
+ pixel_8565/NB1 pixel_8565/VBIAS pixel_8565/NB2 pixel_8565/AMP_IN pixel_8565/SF_IB
+ pixel_8565/PIX_OUT pixel_8565/CSA_VREF pixel
Xpixel_9299 pixel_9299/gring pixel_9299/VDD pixel_9299/GND pixel_9299/VREF pixel_9299/ROW_SEL
+ pixel_9299/NB1 pixel_9299/VBIAS pixel_9299/NB2 pixel_9299/AMP_IN pixel_9299/SF_IB
+ pixel_9299/PIX_OUT pixel_9299/CSA_VREF pixel
Xpixel_7820 pixel_7820/gring pixel_7820/VDD pixel_7820/GND pixel_7820/VREF pixel_7820/ROW_SEL
+ pixel_7820/NB1 pixel_7820/VBIAS pixel_7820/NB2 pixel_7820/AMP_IN pixel_7820/SF_IB
+ pixel_7820/PIX_OUT pixel_7820/CSA_VREF pixel
Xpixel_7831 pixel_7831/gring pixel_7831/VDD pixel_7831/GND pixel_7831/VREF pixel_7831/ROW_SEL
+ pixel_7831/NB1 pixel_7831/VBIAS pixel_7831/NB2 pixel_7831/AMP_IN pixel_7831/SF_IB
+ pixel_7831/PIX_OUT pixel_7831/CSA_VREF pixel
Xpixel_7842 pixel_7842/gring pixel_7842/VDD pixel_7842/GND pixel_7842/VREF pixel_7842/ROW_SEL
+ pixel_7842/NB1 pixel_7842/VBIAS pixel_7842/NB2 pixel_7842/AMP_IN pixel_7842/SF_IB
+ pixel_7842/PIX_OUT pixel_7842/CSA_VREF pixel
Xpixel_8598 pixel_8598/gring pixel_8598/VDD pixel_8598/GND pixel_8598/VREF pixel_8598/ROW_SEL
+ pixel_8598/NB1 pixel_8598/VBIAS pixel_8598/NB2 pixel_8598/AMP_IN pixel_8598/SF_IB
+ pixel_8598/PIX_OUT pixel_8598/CSA_VREF pixel
Xpixel_7853 pixel_7853/gring pixel_7853/VDD pixel_7853/GND pixel_7853/VREF pixel_7853/ROW_SEL
+ pixel_7853/NB1 pixel_7853/VBIAS pixel_7853/NB2 pixel_7853/AMP_IN pixel_7853/SF_IB
+ pixel_7853/PIX_OUT pixel_7853/CSA_VREF pixel
Xpixel_7864 pixel_7864/gring pixel_7864/VDD pixel_7864/GND pixel_7864/VREF pixel_7864/ROW_SEL
+ pixel_7864/NB1 pixel_7864/VBIAS pixel_7864/NB2 pixel_7864/AMP_IN pixel_7864/SF_IB
+ pixel_7864/PIX_OUT pixel_7864/CSA_VREF pixel
Xpixel_7875 pixel_7875/gring pixel_7875/VDD pixel_7875/GND pixel_7875/VREF pixel_7875/ROW_SEL
+ pixel_7875/NB1 pixel_7875/VBIAS pixel_7875/NB2 pixel_7875/AMP_IN pixel_7875/SF_IB
+ pixel_7875/PIX_OUT pixel_7875/CSA_VREF pixel
Xpixel_7886 pixel_7886/gring pixel_7886/VDD pixel_7886/GND pixel_7886/VREF pixel_7886/ROW_SEL
+ pixel_7886/NB1 pixel_7886/VBIAS pixel_7886/NB2 pixel_7886/AMP_IN pixel_7886/SF_IB
+ pixel_7886/PIX_OUT pixel_7886/CSA_VREF pixel
Xpixel_7897 pixel_7897/gring pixel_7897/VDD pixel_7897/GND pixel_7897/VREF pixel_7897/ROW_SEL
+ pixel_7897/NB1 pixel_7897/VBIAS pixel_7897/NB2 pixel_7897/AMP_IN pixel_7897/SF_IB
+ pixel_7897/PIX_OUT pixel_7897/CSA_VREF pixel
Xpixel_2171 pixel_2171/gring pixel_2171/VDD pixel_2171/GND pixel_2171/VREF pixel_2171/ROW_SEL
+ pixel_2171/NB1 pixel_2171/VBIAS pixel_2171/NB2 pixel_2171/AMP_IN pixel_2171/SF_IB
+ pixel_2171/PIX_OUT pixel_2171/CSA_VREF pixel
Xpixel_2160 pixel_2160/gring pixel_2160/VDD pixel_2160/GND pixel_2160/VREF pixel_2160/ROW_SEL
+ pixel_2160/NB1 pixel_2160/VBIAS pixel_2160/NB2 pixel_2160/AMP_IN pixel_2160/SF_IB
+ pixel_2160/PIX_OUT pixel_2160/CSA_VREF pixel
Xpixel_1470 pixel_1470/gring pixel_1470/VDD pixel_1470/GND pixel_1470/VREF pixel_1470/ROW_SEL
+ pixel_1470/NB1 pixel_1470/VBIAS pixel_1470/NB2 pixel_1470/AMP_IN pixel_1470/SF_IB
+ pixel_1470/PIX_OUT pixel_1470/CSA_VREF pixel
Xpixel_2193 pixel_2193/gring pixel_2193/VDD pixel_2193/GND pixel_2193/VREF pixel_2193/ROW_SEL
+ pixel_2193/NB1 pixel_2193/VBIAS pixel_2193/NB2 pixel_2193/AMP_IN pixel_2193/SF_IB
+ pixel_2193/PIX_OUT pixel_2193/CSA_VREF pixel
Xpixel_2182 pixel_2182/gring pixel_2182/VDD pixel_2182/GND pixel_2182/VREF pixel_2182/ROW_SEL
+ pixel_2182/NB1 pixel_2182/VBIAS pixel_2182/NB2 pixel_2182/AMP_IN pixel_2182/SF_IB
+ pixel_2182/PIX_OUT pixel_2182/CSA_VREF pixel
Xpixel_1492 pixel_1492/gring pixel_1492/VDD pixel_1492/GND pixel_1492/VREF pixel_1492/ROW_SEL
+ pixel_1492/NB1 pixel_1492/VBIAS pixel_1492/NB2 pixel_1492/AMP_IN pixel_1492/SF_IB
+ pixel_1492/PIX_OUT pixel_1492/CSA_VREF pixel
Xpixel_1481 pixel_1481/gring pixel_1481/VDD pixel_1481/GND pixel_1481/VREF pixel_1481/ROW_SEL
+ pixel_1481/NB1 pixel_1481/VBIAS pixel_1481/NB2 pixel_1481/AMP_IN pixel_1481/SF_IB
+ pixel_1481/PIX_OUT pixel_1481/CSA_VREF pixel
Xpixel_529 pixel_529/gring pixel_529/VDD pixel_529/GND pixel_529/VREF pixel_529/ROW_SEL
+ pixel_529/NB1 pixel_529/VBIAS pixel_529/NB2 pixel_529/AMP_IN pixel_529/SF_IB pixel_529/PIX_OUT
+ pixel_529/CSA_VREF pixel
Xpixel_518 pixel_518/gring pixel_518/VDD pixel_518/GND pixel_518/VREF pixel_518/ROW_SEL
+ pixel_518/NB1 pixel_518/VBIAS pixel_518/NB2 pixel_518/AMP_IN pixel_518/SF_IB pixel_518/PIX_OUT
+ pixel_518/CSA_VREF pixel
Xpixel_507 pixel_507/gring pixel_507/VDD pixel_507/GND pixel_507/VREF pixel_507/ROW_SEL
+ pixel_507/NB1 pixel_507/VBIAS pixel_507/NB2 pixel_507/AMP_IN pixel_507/SF_IB pixel_507/PIX_OUT
+ pixel_507/CSA_VREF pixel
Xpixel_7105 pixel_7105/gring pixel_7105/VDD pixel_7105/GND pixel_7105/VREF pixel_7105/ROW_SEL
+ pixel_7105/NB1 pixel_7105/VBIAS pixel_7105/NB2 pixel_7105/AMP_IN pixel_7105/SF_IB
+ pixel_7105/PIX_OUT pixel_7105/CSA_VREF pixel
Xpixel_7116 pixel_7116/gring pixel_7116/VDD pixel_7116/GND pixel_7116/VREF pixel_7116/ROW_SEL
+ pixel_7116/NB1 pixel_7116/VBIAS pixel_7116/NB2 pixel_7116/AMP_IN pixel_7116/SF_IB
+ pixel_7116/PIX_OUT pixel_7116/CSA_VREF pixel
Xpixel_7127 pixel_7127/gring pixel_7127/VDD pixel_7127/GND pixel_7127/VREF pixel_7127/ROW_SEL
+ pixel_7127/NB1 pixel_7127/VBIAS pixel_7127/NB2 pixel_7127/AMP_IN pixel_7127/SF_IB
+ pixel_7127/PIX_OUT pixel_7127/CSA_VREF pixel
Xpixel_7138 pixel_7138/gring pixel_7138/VDD pixel_7138/GND pixel_7138/VREF pixel_7138/ROW_SEL
+ pixel_7138/NB1 pixel_7138/VBIAS pixel_7138/NB2 pixel_7138/AMP_IN pixel_7138/SF_IB
+ pixel_7138/PIX_OUT pixel_7138/CSA_VREF pixel
Xpixel_7149 pixel_7149/gring pixel_7149/VDD pixel_7149/GND pixel_7149/VREF pixel_7149/ROW_SEL
+ pixel_7149/NB1 pixel_7149/VBIAS pixel_7149/NB2 pixel_7149/AMP_IN pixel_7149/SF_IB
+ pixel_7149/PIX_OUT pixel_7149/CSA_VREF pixel
Xpixel_6404 pixel_6404/gring pixel_6404/VDD pixel_6404/GND pixel_6404/VREF pixel_6404/ROW_SEL
+ pixel_6404/NB1 pixel_6404/VBIAS pixel_6404/NB2 pixel_6404/AMP_IN pixel_6404/SF_IB
+ pixel_6404/PIX_OUT pixel_6404/CSA_VREF pixel
Xpixel_6415 pixel_6415/gring pixel_6415/VDD pixel_6415/GND pixel_6415/VREF pixel_6415/ROW_SEL
+ pixel_6415/NB1 pixel_6415/VBIAS pixel_6415/NB2 pixel_6415/AMP_IN pixel_6415/SF_IB
+ pixel_6415/PIX_OUT pixel_6415/CSA_VREF pixel
Xpixel_6426 pixel_6426/gring pixel_6426/VDD pixel_6426/GND pixel_6426/VREF pixel_6426/ROW_SEL
+ pixel_6426/NB1 pixel_6426/VBIAS pixel_6426/NB2 pixel_6426/AMP_IN pixel_6426/SF_IB
+ pixel_6426/PIX_OUT pixel_6426/CSA_VREF pixel
Xpixel_6437 pixel_6437/gring pixel_6437/VDD pixel_6437/GND pixel_6437/VREF pixel_6437/ROW_SEL
+ pixel_6437/NB1 pixel_6437/VBIAS pixel_6437/NB2 pixel_6437/AMP_IN pixel_6437/SF_IB
+ pixel_6437/PIX_OUT pixel_6437/CSA_VREF pixel
Xpixel_6448 pixel_6448/gring pixel_6448/VDD pixel_6448/GND pixel_6448/VREF pixel_6448/ROW_SEL
+ pixel_6448/NB1 pixel_6448/VBIAS pixel_6448/NB2 pixel_6448/AMP_IN pixel_6448/SF_IB
+ pixel_6448/PIX_OUT pixel_6448/CSA_VREF pixel
Xpixel_6459 pixel_6459/gring pixel_6459/VDD pixel_6459/GND pixel_6459/VREF pixel_6459/ROW_SEL
+ pixel_6459/NB1 pixel_6459/VBIAS pixel_6459/NB2 pixel_6459/AMP_IN pixel_6459/SF_IB
+ pixel_6459/PIX_OUT pixel_6459/CSA_VREF pixel
Xpixel_5703 pixel_5703/gring pixel_5703/VDD pixel_5703/GND pixel_5703/VREF pixel_5703/ROW_SEL
+ pixel_5703/NB1 pixel_5703/VBIAS pixel_5703/NB2 pixel_5703/AMP_IN pixel_5703/SF_IB
+ pixel_5703/PIX_OUT pixel_5703/CSA_VREF pixel
Xpixel_5714 pixel_5714/gring pixel_5714/VDD pixel_5714/GND pixel_5714/VREF pixel_5714/ROW_SEL
+ pixel_5714/NB1 pixel_5714/VBIAS pixel_5714/NB2 pixel_5714/AMP_IN pixel_5714/SF_IB
+ pixel_5714/PIX_OUT pixel_5714/CSA_VREF pixel
Xpixel_5725 pixel_5725/gring pixel_5725/VDD pixel_5725/GND pixel_5725/VREF pixel_5725/ROW_SEL
+ pixel_5725/NB1 pixel_5725/VBIAS pixel_5725/NB2 pixel_5725/AMP_IN pixel_5725/SF_IB
+ pixel_5725/PIX_OUT pixel_5725/CSA_VREF pixel
Xpixel_5736 pixel_5736/gring pixel_5736/VDD pixel_5736/GND pixel_5736/VREF pixel_5736/ROW_SEL
+ pixel_5736/NB1 pixel_5736/VBIAS pixel_5736/NB2 pixel_5736/AMP_IN pixel_5736/SF_IB
+ pixel_5736/PIX_OUT pixel_5736/CSA_VREF pixel
Xpixel_5747 pixel_5747/gring pixel_5747/VDD pixel_5747/GND pixel_5747/VREF pixel_5747/ROW_SEL
+ pixel_5747/NB1 pixel_5747/VBIAS pixel_5747/NB2 pixel_5747/AMP_IN pixel_5747/SF_IB
+ pixel_5747/PIX_OUT pixel_5747/CSA_VREF pixel
Xpixel_5758 pixel_5758/gring pixel_5758/VDD pixel_5758/GND pixel_5758/VREF pixel_5758/ROW_SEL
+ pixel_5758/NB1 pixel_5758/VBIAS pixel_5758/NB2 pixel_5758/AMP_IN pixel_5758/SF_IB
+ pixel_5758/PIX_OUT pixel_5758/CSA_VREF pixel
Xpixel_5769 pixel_5769/gring pixel_5769/VDD pixel_5769/GND pixel_5769/VREF pixel_5769/ROW_SEL
+ pixel_5769/NB1 pixel_5769/VBIAS pixel_5769/NB2 pixel_5769/AMP_IN pixel_5769/SF_IB
+ pixel_5769/PIX_OUT pixel_5769/CSA_VREF pixel
Xpixel_9030 pixel_9030/gring pixel_9030/VDD pixel_9030/GND pixel_9030/VREF pixel_9030/ROW_SEL
+ pixel_9030/NB1 pixel_9030/VBIAS pixel_9030/NB2 pixel_9030/AMP_IN pixel_9030/SF_IB
+ pixel_9030/PIX_OUT pixel_9030/CSA_VREF pixel
Xpixel_9063 pixel_9063/gring pixel_9063/VDD pixel_9063/GND pixel_9063/VREF pixel_9063/ROW_SEL
+ pixel_9063/NB1 pixel_9063/VBIAS pixel_9063/NB2 pixel_9063/AMP_IN pixel_9063/SF_IB
+ pixel_9063/PIX_OUT pixel_9063/CSA_VREF pixel
Xpixel_9052 pixel_9052/gring pixel_9052/VDD pixel_9052/GND pixel_9052/VREF pixel_9052/ROW_SEL
+ pixel_9052/NB1 pixel_9052/VBIAS pixel_9052/NB2 pixel_9052/AMP_IN pixel_9052/SF_IB
+ pixel_9052/PIX_OUT pixel_9052/CSA_VREF pixel
Xpixel_9041 pixel_9041/gring pixel_9041/VDD pixel_9041/GND pixel_9041/VREF pixel_9041/ROW_SEL
+ pixel_9041/NB1 pixel_9041/VBIAS pixel_9041/NB2 pixel_9041/AMP_IN pixel_9041/SF_IB
+ pixel_9041/PIX_OUT pixel_9041/CSA_VREF pixel
Xpixel_9096 pixel_9096/gring pixel_9096/VDD pixel_9096/GND pixel_9096/VREF pixel_9096/ROW_SEL
+ pixel_9096/NB1 pixel_9096/VBIAS pixel_9096/NB2 pixel_9096/AMP_IN pixel_9096/SF_IB
+ pixel_9096/PIX_OUT pixel_9096/CSA_VREF pixel
Xpixel_9085 pixel_9085/gring pixel_9085/VDD pixel_9085/GND pixel_9085/VREF pixel_9085/ROW_SEL
+ pixel_9085/NB1 pixel_9085/VBIAS pixel_9085/NB2 pixel_9085/AMP_IN pixel_9085/SF_IB
+ pixel_9085/PIX_OUT pixel_9085/CSA_VREF pixel
Xpixel_9074 pixel_9074/gring pixel_9074/VDD pixel_9074/GND pixel_9074/VREF pixel_9074/ROW_SEL
+ pixel_9074/NB1 pixel_9074/VBIAS pixel_9074/NB2 pixel_9074/AMP_IN pixel_9074/SF_IB
+ pixel_9074/PIX_OUT pixel_9074/CSA_VREF pixel
Xpixel_8340 pixel_8340/gring pixel_8340/VDD pixel_8340/GND pixel_8340/VREF pixel_8340/ROW_SEL
+ pixel_8340/NB1 pixel_8340/VBIAS pixel_8340/NB2 pixel_8340/AMP_IN pixel_8340/SF_IB
+ pixel_8340/PIX_OUT pixel_8340/CSA_VREF pixel
Xpixel_8351 pixel_8351/gring pixel_8351/VDD pixel_8351/GND pixel_8351/VREF pixel_8351/ROW_SEL
+ pixel_8351/NB1 pixel_8351/VBIAS pixel_8351/NB2 pixel_8351/AMP_IN pixel_8351/SF_IB
+ pixel_8351/PIX_OUT pixel_8351/CSA_VREF pixel
Xpixel_8362 pixel_8362/gring pixel_8362/VDD pixel_8362/GND pixel_8362/VREF pixel_8362/ROW_SEL
+ pixel_8362/NB1 pixel_8362/VBIAS pixel_8362/NB2 pixel_8362/AMP_IN pixel_8362/SF_IB
+ pixel_8362/PIX_OUT pixel_8362/CSA_VREF pixel
Xpixel_8373 pixel_8373/gring pixel_8373/VDD pixel_8373/GND pixel_8373/VREF pixel_8373/ROW_SEL
+ pixel_8373/NB1 pixel_8373/VBIAS pixel_8373/NB2 pixel_8373/AMP_IN pixel_8373/SF_IB
+ pixel_8373/PIX_OUT pixel_8373/CSA_VREF pixel
Xpixel_8384 pixel_8384/gring pixel_8384/VDD pixel_8384/GND pixel_8384/VREF pixel_8384/ROW_SEL
+ pixel_8384/NB1 pixel_8384/VBIAS pixel_8384/NB2 pixel_8384/AMP_IN pixel_8384/SF_IB
+ pixel_8384/PIX_OUT pixel_8384/CSA_VREF pixel
Xpixel_8395 pixel_8395/gring pixel_8395/VDD pixel_8395/GND pixel_8395/VREF pixel_8395/ROW_SEL
+ pixel_8395/NB1 pixel_8395/VBIAS pixel_8395/NB2 pixel_8395/AMP_IN pixel_8395/SF_IB
+ pixel_8395/PIX_OUT pixel_8395/CSA_VREF pixel
Xpixel_7650 pixel_7650/gring pixel_7650/VDD pixel_7650/GND pixel_7650/VREF pixel_7650/ROW_SEL
+ pixel_7650/NB1 pixel_7650/VBIAS pixel_7650/NB2 pixel_7650/AMP_IN pixel_7650/SF_IB
+ pixel_7650/PIX_OUT pixel_7650/CSA_VREF pixel
Xpixel_7661 pixel_7661/gring pixel_7661/VDD pixel_7661/GND pixel_7661/VREF pixel_7661/ROW_SEL
+ pixel_7661/NB1 pixel_7661/VBIAS pixel_7661/NB2 pixel_7661/AMP_IN pixel_7661/SF_IB
+ pixel_7661/PIX_OUT pixel_7661/CSA_VREF pixel
Xpixel_7672 pixel_7672/gring pixel_7672/VDD pixel_7672/GND pixel_7672/VREF pixel_7672/ROW_SEL
+ pixel_7672/NB1 pixel_7672/VBIAS pixel_7672/NB2 pixel_7672/AMP_IN pixel_7672/SF_IB
+ pixel_7672/PIX_OUT pixel_7672/CSA_VREF pixel
Xpixel_7683 pixel_7683/gring pixel_7683/VDD pixel_7683/GND pixel_7683/VREF pixel_7683/ROW_SEL
+ pixel_7683/NB1 pixel_7683/VBIAS pixel_7683/NB2 pixel_7683/AMP_IN pixel_7683/SF_IB
+ pixel_7683/PIX_OUT pixel_7683/CSA_VREF pixel
Xpixel_7694 pixel_7694/gring pixel_7694/VDD pixel_7694/GND pixel_7694/VREF pixel_7694/ROW_SEL
+ pixel_7694/NB1 pixel_7694/VBIAS pixel_7694/NB2 pixel_7694/AMP_IN pixel_7694/SF_IB
+ pixel_7694/PIX_OUT pixel_7694/CSA_VREF pixel
Xpixel_30 pixel_30/gring pixel_30/VDD pixel_30/GND pixel_30/VREF pixel_30/ROW_SEL
+ pixel_30/NB1 pixel_30/VBIAS pixel_30/NB2 pixel_30/AMP_IN pixel_30/SF_IB pixel_30/PIX_OUT
+ pixel_30/CSA_VREF pixel
Xpixel_6960 pixel_6960/gring pixel_6960/VDD pixel_6960/GND pixel_6960/VREF pixel_6960/ROW_SEL
+ pixel_6960/NB1 pixel_6960/VBIAS pixel_6960/NB2 pixel_6960/AMP_IN pixel_6960/SF_IB
+ pixel_6960/PIX_OUT pixel_6960/CSA_VREF pixel
Xpixel_6971 pixel_6971/gring pixel_6971/VDD pixel_6971/GND pixel_6971/VREF pixel_6971/ROW_SEL
+ pixel_6971/NB1 pixel_6971/VBIAS pixel_6971/NB2 pixel_6971/AMP_IN pixel_6971/SF_IB
+ pixel_6971/PIX_OUT pixel_6971/CSA_VREF pixel
Xpixel_6982 pixel_6982/gring pixel_6982/VDD pixel_6982/GND pixel_6982/VREF pixel_6982/ROW_SEL
+ pixel_6982/NB1 pixel_6982/VBIAS pixel_6982/NB2 pixel_6982/AMP_IN pixel_6982/SF_IB
+ pixel_6982/PIX_OUT pixel_6982/CSA_VREF pixel
Xpixel_63 pixel_63/gring pixel_63/VDD pixel_63/GND pixel_63/VREF pixel_63/ROW_SEL
+ pixel_63/NB1 pixel_63/VBIAS pixel_63/NB2 pixel_63/AMP_IN pixel_63/SF_IB pixel_63/PIX_OUT
+ pixel_63/CSA_VREF pixel
Xpixel_52 pixel_52/gring pixel_52/VDD pixel_52/GND pixel_52/VREF pixel_52/ROW_SEL
+ pixel_52/NB1 pixel_52/VBIAS pixel_52/NB2 pixel_52/AMP_IN pixel_52/SF_IB pixel_52/PIX_OUT
+ pixel_52/CSA_VREF pixel
Xpixel_41 pixel_41/gring pixel_41/VDD pixel_41/GND pixel_41/VREF pixel_41/ROW_SEL
+ pixel_41/NB1 pixel_41/VBIAS pixel_41/NB2 pixel_41/AMP_IN pixel_41/SF_IB pixel_41/PIX_OUT
+ pixel_41/CSA_VREF pixel
Xpixel_6993 pixel_6993/gring pixel_6993/VDD pixel_6993/GND pixel_6993/VREF pixel_6993/ROW_SEL
+ pixel_6993/NB1 pixel_6993/VBIAS pixel_6993/NB2 pixel_6993/AMP_IN pixel_6993/SF_IB
+ pixel_6993/PIX_OUT pixel_6993/CSA_VREF pixel
Xpixel_96 pixel_96/gring pixel_96/VDD pixel_96/GND pixel_96/VREF pixel_96/ROW_SEL
+ pixel_96/NB1 pixel_96/VBIAS pixel_96/NB2 pixel_96/AMP_IN pixel_96/SF_IB pixel_96/PIX_OUT
+ pixel_96/CSA_VREF pixel
Xpixel_85 pixel_85/gring pixel_85/VDD pixel_85/GND pixel_85/VREF pixel_85/ROW_SEL
+ pixel_85/NB1 pixel_85/VBIAS pixel_85/NB2 pixel_85/AMP_IN pixel_85/SF_IB pixel_85/PIX_OUT
+ pixel_85/CSA_VREF pixel
Xpixel_74 pixel_74/gring pixel_74/VDD pixel_74/GND pixel_74/VREF pixel_74/ROW_SEL
+ pixel_74/NB1 pixel_74/VBIAS pixel_74/NB2 pixel_74/AMP_IN pixel_74/SF_IB pixel_74/PIX_OUT
+ pixel_74/CSA_VREF pixel
Xpixel_304 pixel_304/gring pixel_304/VDD pixel_304/GND pixel_304/VREF pixel_304/ROW_SEL
+ pixel_304/NB1 pixel_304/VBIAS pixel_304/NB2 pixel_304/AMP_IN pixel_304/SF_IB pixel_304/PIX_OUT
+ pixel_304/CSA_VREF pixel
Xpixel_4309 pixel_4309/gring pixel_4309/VDD pixel_4309/GND pixel_4309/VREF pixel_4309/ROW_SEL
+ pixel_4309/NB1 pixel_4309/VBIAS pixel_4309/NB2 pixel_4309/AMP_IN pixel_4309/SF_IB
+ pixel_4309/PIX_OUT pixel_4309/CSA_VREF pixel
Xpixel_337 pixel_337/gring pixel_337/VDD pixel_337/GND pixel_337/VREF pixel_337/ROW_SEL
+ pixel_337/NB1 pixel_337/VBIAS pixel_337/NB2 pixel_337/AMP_IN pixel_337/SF_IB pixel_337/PIX_OUT
+ pixel_337/CSA_VREF pixel
Xpixel_326 pixel_326/gring pixel_326/VDD pixel_326/GND pixel_326/VREF pixel_326/ROW_SEL
+ pixel_326/NB1 pixel_326/VBIAS pixel_326/NB2 pixel_326/AMP_IN pixel_326/SF_IB pixel_326/PIX_OUT
+ pixel_326/CSA_VREF pixel
Xpixel_315 pixel_315/gring pixel_315/VDD pixel_315/GND pixel_315/VREF pixel_315/ROW_SEL
+ pixel_315/NB1 pixel_315/VBIAS pixel_315/NB2 pixel_315/AMP_IN pixel_315/SF_IB pixel_315/PIX_OUT
+ pixel_315/CSA_VREF pixel
Xpixel_359 pixel_359/gring pixel_359/VDD pixel_359/GND pixel_359/VREF pixel_359/ROW_SEL
+ pixel_359/NB1 pixel_359/VBIAS pixel_359/NB2 pixel_359/AMP_IN pixel_359/SF_IB pixel_359/PIX_OUT
+ pixel_359/CSA_VREF pixel
Xpixel_348 pixel_348/gring pixel_348/VDD pixel_348/GND pixel_348/VREF pixel_348/ROW_SEL
+ pixel_348/NB1 pixel_348/VBIAS pixel_348/NB2 pixel_348/AMP_IN pixel_348/SF_IB pixel_348/PIX_OUT
+ pixel_348/CSA_VREF pixel
Xpixel_3619 pixel_3619/gring pixel_3619/VDD pixel_3619/GND pixel_3619/VREF pixel_3619/ROW_SEL
+ pixel_3619/NB1 pixel_3619/VBIAS pixel_3619/NB2 pixel_3619/AMP_IN pixel_3619/SF_IB
+ pixel_3619/PIX_OUT pixel_3619/CSA_VREF pixel
Xpixel_3608 pixel_3608/gring pixel_3608/VDD pixel_3608/GND pixel_3608/VREF pixel_3608/ROW_SEL
+ pixel_3608/NB1 pixel_3608/VBIAS pixel_3608/NB2 pixel_3608/AMP_IN pixel_3608/SF_IB
+ pixel_3608/PIX_OUT pixel_3608/CSA_VREF pixel
Xpixel_2929 pixel_2929/gring pixel_2929/VDD pixel_2929/GND pixel_2929/VREF pixel_2929/ROW_SEL
+ pixel_2929/NB1 pixel_2929/VBIAS pixel_2929/NB2 pixel_2929/AMP_IN pixel_2929/SF_IB
+ pixel_2929/PIX_OUT pixel_2929/CSA_VREF pixel
Xpixel_2918 pixel_2918/gring pixel_2918/VDD pixel_2918/GND pixel_2918/VREF pixel_2918/ROW_SEL
+ pixel_2918/NB1 pixel_2918/VBIAS pixel_2918/NB2 pixel_2918/AMP_IN pixel_2918/SF_IB
+ pixel_2918/PIX_OUT pixel_2918/CSA_VREF pixel
Xpixel_2907 pixel_2907/gring pixel_2907/VDD pixel_2907/GND pixel_2907/VREF pixel_2907/ROW_SEL
+ pixel_2907/NB1 pixel_2907/VBIAS pixel_2907/NB2 pixel_2907/AMP_IN pixel_2907/SF_IB
+ pixel_2907/PIX_OUT pixel_2907/CSA_VREF pixel
Xpixel_6201 pixel_6201/gring pixel_6201/VDD pixel_6201/GND pixel_6201/VREF pixel_6201/ROW_SEL
+ pixel_6201/NB1 pixel_6201/VBIAS pixel_6201/NB2 pixel_6201/AMP_IN pixel_6201/SF_IB
+ pixel_6201/PIX_OUT pixel_6201/CSA_VREF pixel
Xpixel_6212 pixel_6212/gring pixel_6212/VDD pixel_6212/GND pixel_6212/VREF pixel_6212/ROW_SEL
+ pixel_6212/NB1 pixel_6212/VBIAS pixel_6212/NB2 pixel_6212/AMP_IN pixel_6212/SF_IB
+ pixel_6212/PIX_OUT pixel_6212/CSA_VREF pixel
Xpixel_6223 pixel_6223/gring pixel_6223/VDD pixel_6223/GND pixel_6223/VREF pixel_6223/ROW_SEL
+ pixel_6223/NB1 pixel_6223/VBIAS pixel_6223/NB2 pixel_6223/AMP_IN pixel_6223/SF_IB
+ pixel_6223/PIX_OUT pixel_6223/CSA_VREF pixel
Xpixel_6234 pixel_6234/gring pixel_6234/VDD pixel_6234/GND pixel_6234/VREF pixel_6234/ROW_SEL
+ pixel_6234/NB1 pixel_6234/VBIAS pixel_6234/NB2 pixel_6234/AMP_IN pixel_6234/SF_IB
+ pixel_6234/PIX_OUT pixel_6234/CSA_VREF pixel
Xpixel_6245 pixel_6245/gring pixel_6245/VDD pixel_6245/GND pixel_6245/VREF pixel_6245/ROW_SEL
+ pixel_6245/NB1 pixel_6245/VBIAS pixel_6245/NB2 pixel_6245/AMP_IN pixel_6245/SF_IB
+ pixel_6245/PIX_OUT pixel_6245/CSA_VREF pixel
Xpixel_6256 pixel_6256/gring pixel_6256/VDD pixel_6256/GND pixel_6256/VREF pixel_6256/ROW_SEL
+ pixel_6256/NB1 pixel_6256/VBIAS pixel_6256/NB2 pixel_6256/AMP_IN pixel_6256/SF_IB
+ pixel_6256/PIX_OUT pixel_6256/CSA_VREF pixel
Xpixel_6267 pixel_6267/gring pixel_6267/VDD pixel_6267/GND pixel_6267/VREF pixel_6267/ROW_SEL
+ pixel_6267/NB1 pixel_6267/VBIAS pixel_6267/NB2 pixel_6267/AMP_IN pixel_6267/SF_IB
+ pixel_6267/PIX_OUT pixel_6267/CSA_VREF pixel
Xpixel_6278 pixel_6278/gring pixel_6278/VDD pixel_6278/GND pixel_6278/VREF pixel_6278/ROW_SEL
+ pixel_6278/NB1 pixel_6278/VBIAS pixel_6278/NB2 pixel_6278/AMP_IN pixel_6278/SF_IB
+ pixel_6278/PIX_OUT pixel_6278/CSA_VREF pixel
Xpixel_5500 pixel_5500/gring pixel_5500/VDD pixel_5500/GND pixel_5500/VREF pixel_5500/ROW_SEL
+ pixel_5500/NB1 pixel_5500/VBIAS pixel_5500/NB2 pixel_5500/AMP_IN pixel_5500/SF_IB
+ pixel_5500/PIX_OUT pixel_5500/CSA_VREF pixel
Xpixel_5511 pixel_5511/gring pixel_5511/VDD pixel_5511/GND pixel_5511/VREF pixel_5511/ROW_SEL
+ pixel_5511/NB1 pixel_5511/VBIAS pixel_5511/NB2 pixel_5511/AMP_IN pixel_5511/SF_IB
+ pixel_5511/PIX_OUT pixel_5511/CSA_VREF pixel
Xpixel_5522 pixel_5522/gring pixel_5522/VDD pixel_5522/GND pixel_5522/VREF pixel_5522/ROW_SEL
+ pixel_5522/NB1 pixel_5522/VBIAS pixel_5522/NB2 pixel_5522/AMP_IN pixel_5522/SF_IB
+ pixel_5522/PIX_OUT pixel_5522/CSA_VREF pixel
Xpixel_5533 pixel_5533/gring pixel_5533/VDD pixel_5533/GND pixel_5533/VREF pixel_5533/ROW_SEL
+ pixel_5533/NB1 pixel_5533/VBIAS pixel_5533/NB2 pixel_5533/AMP_IN pixel_5533/SF_IB
+ pixel_5533/PIX_OUT pixel_5533/CSA_VREF pixel
Xpixel_6289 pixel_6289/gring pixel_6289/VDD pixel_6289/GND pixel_6289/VREF pixel_6289/ROW_SEL
+ pixel_6289/NB1 pixel_6289/VBIAS pixel_6289/NB2 pixel_6289/AMP_IN pixel_6289/SF_IB
+ pixel_6289/PIX_OUT pixel_6289/CSA_VREF pixel
Xpixel_5544 pixel_5544/gring pixel_5544/VDD pixel_5544/GND pixel_5544/VREF pixel_5544/ROW_SEL
+ pixel_5544/NB1 pixel_5544/VBIAS pixel_5544/NB2 pixel_5544/AMP_IN pixel_5544/SF_IB
+ pixel_5544/PIX_OUT pixel_5544/CSA_VREF pixel
Xpixel_5555 pixel_5555/gring pixel_5555/VDD pixel_5555/GND pixel_5555/VREF pixel_5555/ROW_SEL
+ pixel_5555/NB1 pixel_5555/VBIAS pixel_5555/NB2 pixel_5555/AMP_IN pixel_5555/SF_IB
+ pixel_5555/PIX_OUT pixel_5555/CSA_VREF pixel
Xpixel_5566 pixel_5566/gring pixel_5566/VDD pixel_5566/GND pixel_5566/VREF pixel_5566/ROW_SEL
+ pixel_5566/NB1 pixel_5566/VBIAS pixel_5566/NB2 pixel_5566/AMP_IN pixel_5566/SF_IB
+ pixel_5566/PIX_OUT pixel_5566/CSA_VREF pixel
Xpixel_4810 pixel_4810/gring pixel_4810/VDD pixel_4810/GND pixel_4810/VREF pixel_4810/ROW_SEL
+ pixel_4810/NB1 pixel_4810/VBIAS pixel_4810/NB2 pixel_4810/AMP_IN pixel_4810/SF_IB
+ pixel_4810/PIX_OUT pixel_4810/CSA_VREF pixel
Xpixel_4821 pixel_4821/gring pixel_4821/VDD pixel_4821/GND pixel_4821/VREF pixel_4821/ROW_SEL
+ pixel_4821/NB1 pixel_4821/VBIAS pixel_4821/NB2 pixel_4821/AMP_IN pixel_4821/SF_IB
+ pixel_4821/PIX_OUT pixel_4821/CSA_VREF pixel
Xpixel_860 pixel_860/gring pixel_860/VDD pixel_860/GND pixel_860/VREF pixel_860/ROW_SEL
+ pixel_860/NB1 pixel_860/VBIAS pixel_860/NB2 pixel_860/AMP_IN pixel_860/SF_IB pixel_860/PIX_OUT
+ pixel_860/CSA_VREF pixel
Xpixel_5577 pixel_5577/gring pixel_5577/VDD pixel_5577/GND pixel_5577/VREF pixel_5577/ROW_SEL
+ pixel_5577/NB1 pixel_5577/VBIAS pixel_5577/NB2 pixel_5577/AMP_IN pixel_5577/SF_IB
+ pixel_5577/PIX_OUT pixel_5577/CSA_VREF pixel
Xpixel_5588 pixel_5588/gring pixel_5588/VDD pixel_5588/GND pixel_5588/VREF pixel_5588/ROW_SEL
+ pixel_5588/NB1 pixel_5588/VBIAS pixel_5588/NB2 pixel_5588/AMP_IN pixel_5588/SF_IB
+ pixel_5588/PIX_OUT pixel_5588/CSA_VREF pixel
Xpixel_5599 pixel_5599/gring pixel_5599/VDD pixel_5599/GND pixel_5599/VREF pixel_5599/ROW_SEL
+ pixel_5599/NB1 pixel_5599/VBIAS pixel_5599/NB2 pixel_5599/AMP_IN pixel_5599/SF_IB
+ pixel_5599/PIX_OUT pixel_5599/CSA_VREF pixel
Xpixel_4832 pixel_4832/gring pixel_4832/VDD pixel_4832/GND pixel_4832/VREF pixel_4832/ROW_SEL
+ pixel_4832/NB1 pixel_4832/VBIAS pixel_4832/NB2 pixel_4832/AMP_IN pixel_4832/SF_IB
+ pixel_4832/PIX_OUT pixel_4832/CSA_VREF pixel
Xpixel_4843 pixel_4843/gring pixel_4843/VDD pixel_4843/GND pixel_4843/VREF pixel_4843/ROW_SEL
+ pixel_4843/NB1 pixel_4843/VBIAS pixel_4843/NB2 pixel_4843/AMP_IN pixel_4843/SF_IB
+ pixel_4843/PIX_OUT pixel_4843/CSA_VREF pixel
Xpixel_4854 pixel_4854/gring pixel_4854/VDD pixel_4854/GND pixel_4854/VREF pixel_4854/ROW_SEL
+ pixel_4854/NB1 pixel_4854/VBIAS pixel_4854/NB2 pixel_4854/AMP_IN pixel_4854/SF_IB
+ pixel_4854/PIX_OUT pixel_4854/CSA_VREF pixel
Xpixel_4865 pixel_4865/gring pixel_4865/VDD pixel_4865/GND pixel_4865/VREF pixel_4865/ROW_SEL
+ pixel_4865/NB1 pixel_4865/VBIAS pixel_4865/NB2 pixel_4865/AMP_IN pixel_4865/SF_IB
+ pixel_4865/PIX_OUT pixel_4865/CSA_VREF pixel
Xpixel_893 pixel_893/gring pixel_893/VDD pixel_893/GND pixel_893/VREF pixel_893/ROW_SEL
+ pixel_893/NB1 pixel_893/VBIAS pixel_893/NB2 pixel_893/AMP_IN pixel_893/SF_IB pixel_893/PIX_OUT
+ pixel_893/CSA_VREF pixel
Xpixel_882 pixel_882/gring pixel_882/VDD pixel_882/GND pixel_882/VREF pixel_882/ROW_SEL
+ pixel_882/NB1 pixel_882/VBIAS pixel_882/NB2 pixel_882/AMP_IN pixel_882/SF_IB pixel_882/PIX_OUT
+ pixel_882/CSA_VREF pixel
Xpixel_871 pixel_871/gring pixel_871/VDD pixel_871/GND pixel_871/VREF pixel_871/ROW_SEL
+ pixel_871/NB1 pixel_871/VBIAS pixel_871/NB2 pixel_871/AMP_IN pixel_871/SF_IB pixel_871/PIX_OUT
+ pixel_871/CSA_VREF pixel
Xpixel_4876 pixel_4876/gring pixel_4876/VDD pixel_4876/GND pixel_4876/VREF pixel_4876/ROW_SEL
+ pixel_4876/NB1 pixel_4876/VBIAS pixel_4876/NB2 pixel_4876/AMP_IN pixel_4876/SF_IB
+ pixel_4876/PIX_OUT pixel_4876/CSA_VREF pixel
Xpixel_4887 pixel_4887/gring pixel_4887/VDD pixel_4887/GND pixel_4887/VREF pixel_4887/ROW_SEL
+ pixel_4887/NB1 pixel_4887/VBIAS pixel_4887/NB2 pixel_4887/AMP_IN pixel_4887/SF_IB
+ pixel_4887/PIX_OUT pixel_4887/CSA_VREF pixel
Xpixel_4898 pixel_4898/gring pixel_4898/VDD pixel_4898/GND pixel_4898/VREF pixel_4898/ROW_SEL
+ pixel_4898/NB1 pixel_4898/VBIAS pixel_4898/NB2 pixel_4898/AMP_IN pixel_4898/SF_IB
+ pixel_4898/PIX_OUT pixel_4898/CSA_VREF pixel
Xpixel_8170 pixel_8170/gring pixel_8170/VDD pixel_8170/GND pixel_8170/VREF pixel_8170/ROW_SEL
+ pixel_8170/NB1 pixel_8170/VBIAS pixel_8170/NB2 pixel_8170/AMP_IN pixel_8170/SF_IB
+ pixel_8170/PIX_OUT pixel_8170/CSA_VREF pixel
Xpixel_8181 pixel_8181/gring pixel_8181/VDD pixel_8181/GND pixel_8181/VREF pixel_8181/ROW_SEL
+ pixel_8181/NB1 pixel_8181/VBIAS pixel_8181/NB2 pixel_8181/AMP_IN pixel_8181/SF_IB
+ pixel_8181/PIX_OUT pixel_8181/CSA_VREF pixel
Xpixel_8192 pixel_8192/gring pixel_8192/VDD pixel_8192/GND pixel_8192/VREF pixel_8192/ROW_SEL
+ pixel_8192/NB1 pixel_8192/VBIAS pixel_8192/NB2 pixel_8192/AMP_IN pixel_8192/SF_IB
+ pixel_8192/PIX_OUT pixel_8192/CSA_VREF pixel
Xpixel_7480 pixel_7480/gring pixel_7480/VDD pixel_7480/GND pixel_7480/VREF pixel_7480/ROW_SEL
+ pixel_7480/NB1 pixel_7480/VBIAS pixel_7480/NB2 pixel_7480/AMP_IN pixel_7480/SF_IB
+ pixel_7480/PIX_OUT pixel_7480/CSA_VREF pixel
Xpixel_7491 pixel_7491/gring pixel_7491/VDD pixel_7491/GND pixel_7491/VREF pixel_7491/ROW_SEL
+ pixel_7491/NB1 pixel_7491/VBIAS pixel_7491/NB2 pixel_7491/AMP_IN pixel_7491/SF_IB
+ pixel_7491/PIX_OUT pixel_7491/CSA_VREF pixel
Xpixel_6790 pixel_6790/gring pixel_6790/VDD pixel_6790/GND pixel_6790/VREF pixel_6790/ROW_SEL
+ pixel_6790/NB1 pixel_6790/VBIAS pixel_6790/NB2 pixel_6790/AMP_IN pixel_6790/SF_IB
+ pixel_6790/PIX_OUT pixel_6790/CSA_VREF pixel
Xpixel_112 pixel_112/gring pixel_112/VDD pixel_112/GND pixel_112/VREF pixel_112/ROW_SEL
+ pixel_112/NB1 pixel_112/VBIAS pixel_112/NB2 pixel_112/AMP_IN pixel_112/SF_IB pixel_112/PIX_OUT
+ pixel_112/CSA_VREF pixel
Xpixel_101 pixel_101/gring pixel_101/VDD pixel_101/GND pixel_101/VREF pixel_101/ROW_SEL
+ pixel_101/NB1 pixel_101/VBIAS pixel_101/NB2 pixel_101/AMP_IN pixel_101/SF_IB pixel_101/PIX_OUT
+ pixel_101/CSA_VREF pixel
Xpixel_4106 pixel_4106/gring pixel_4106/VDD pixel_4106/GND pixel_4106/VREF pixel_4106/ROW_SEL
+ pixel_4106/NB1 pixel_4106/VBIAS pixel_4106/NB2 pixel_4106/AMP_IN pixel_4106/SF_IB
+ pixel_4106/PIX_OUT pixel_4106/CSA_VREF pixel
Xpixel_4117 pixel_4117/gring pixel_4117/VDD pixel_4117/GND pixel_4117/VREF pixel_4117/ROW_SEL
+ pixel_4117/NB1 pixel_4117/VBIAS pixel_4117/NB2 pixel_4117/AMP_IN pixel_4117/SF_IB
+ pixel_4117/PIX_OUT pixel_4117/CSA_VREF pixel
Xpixel_145 pixel_145/gring pixel_145/VDD pixel_145/GND pixel_145/VREF pixel_145/ROW_SEL
+ pixel_145/NB1 pixel_145/VBIAS pixel_145/NB2 pixel_145/AMP_IN pixel_145/SF_IB pixel_145/PIX_OUT
+ pixel_145/CSA_VREF pixel
Xpixel_134 pixel_134/gring pixel_134/VDD pixel_134/GND pixel_134/VREF pixel_134/ROW_SEL
+ pixel_134/NB1 pixel_134/VBIAS pixel_134/NB2 pixel_134/AMP_IN pixel_134/SF_IB pixel_134/PIX_OUT
+ pixel_134/CSA_VREF pixel
Xpixel_123 pixel_123/gring pixel_123/VDD pixel_123/GND pixel_123/VREF pixel_123/ROW_SEL
+ pixel_123/NB1 pixel_123/VBIAS pixel_123/NB2 pixel_123/AMP_IN pixel_123/SF_IB pixel_123/PIX_OUT
+ pixel_123/CSA_VREF pixel
Xpixel_3405 pixel_3405/gring pixel_3405/VDD pixel_3405/GND pixel_3405/VREF pixel_3405/ROW_SEL
+ pixel_3405/NB1 pixel_3405/VBIAS pixel_3405/NB2 pixel_3405/AMP_IN pixel_3405/SF_IB
+ pixel_3405/PIX_OUT pixel_3405/CSA_VREF pixel
Xpixel_4128 pixel_4128/gring pixel_4128/VDD pixel_4128/GND pixel_4128/VREF pixel_4128/ROW_SEL
+ pixel_4128/NB1 pixel_4128/VBIAS pixel_4128/NB2 pixel_4128/AMP_IN pixel_4128/SF_IB
+ pixel_4128/PIX_OUT pixel_4128/CSA_VREF pixel
Xpixel_4139 pixel_4139/gring pixel_4139/VDD pixel_4139/GND pixel_4139/VREF pixel_4139/ROW_SEL
+ pixel_4139/NB1 pixel_4139/VBIAS pixel_4139/NB2 pixel_4139/AMP_IN pixel_4139/SF_IB
+ pixel_4139/PIX_OUT pixel_4139/CSA_VREF pixel
Xpixel_189 pixel_189/gring pixel_189/VDD pixel_189/GND pixel_189/VREF pixel_189/ROW_SEL
+ pixel_189/NB1 pixel_189/VBIAS pixel_189/NB2 pixel_189/AMP_IN pixel_189/SF_IB pixel_189/PIX_OUT
+ pixel_189/CSA_VREF pixel
Xpixel_178 pixel_178/gring pixel_178/VDD pixel_178/GND pixel_178/VREF pixel_178/ROW_SEL
+ pixel_178/NB1 pixel_178/VBIAS pixel_178/NB2 pixel_178/AMP_IN pixel_178/SF_IB pixel_178/PIX_OUT
+ pixel_178/CSA_VREF pixel
Xpixel_167 pixel_167/gring pixel_167/VDD pixel_167/GND pixel_167/VREF pixel_167/ROW_SEL
+ pixel_167/NB1 pixel_167/VBIAS pixel_167/NB2 pixel_167/AMP_IN pixel_167/SF_IB pixel_167/PIX_OUT
+ pixel_167/CSA_VREF pixel
Xpixel_156 pixel_156/gring pixel_156/VDD pixel_156/GND pixel_156/VREF pixel_156/ROW_SEL
+ pixel_156/NB1 pixel_156/VBIAS pixel_156/NB2 pixel_156/AMP_IN pixel_156/SF_IB pixel_156/PIX_OUT
+ pixel_156/CSA_VREF pixel
Xpixel_2704 pixel_2704/gring pixel_2704/VDD pixel_2704/GND pixel_2704/VREF pixel_2704/ROW_SEL
+ pixel_2704/NB1 pixel_2704/VBIAS pixel_2704/NB2 pixel_2704/AMP_IN pixel_2704/SF_IB
+ pixel_2704/PIX_OUT pixel_2704/CSA_VREF pixel
Xpixel_3449 pixel_3449/gring pixel_3449/VDD pixel_3449/GND pixel_3449/VREF pixel_3449/ROW_SEL
+ pixel_3449/NB1 pixel_3449/VBIAS pixel_3449/NB2 pixel_3449/AMP_IN pixel_3449/SF_IB
+ pixel_3449/PIX_OUT pixel_3449/CSA_VREF pixel
Xpixel_3438 pixel_3438/gring pixel_3438/VDD pixel_3438/GND pixel_3438/VREF pixel_3438/ROW_SEL
+ pixel_3438/NB1 pixel_3438/VBIAS pixel_3438/NB2 pixel_3438/AMP_IN pixel_3438/SF_IB
+ pixel_3438/PIX_OUT pixel_3438/CSA_VREF pixel
Xpixel_3427 pixel_3427/gring pixel_3427/VDD pixel_3427/GND pixel_3427/VREF pixel_3427/ROW_SEL
+ pixel_3427/NB1 pixel_3427/VBIAS pixel_3427/NB2 pixel_3427/AMP_IN pixel_3427/SF_IB
+ pixel_3427/PIX_OUT pixel_3427/CSA_VREF pixel
Xpixel_3416 pixel_3416/gring pixel_3416/VDD pixel_3416/GND pixel_3416/VREF pixel_3416/ROW_SEL
+ pixel_3416/NB1 pixel_3416/VBIAS pixel_3416/NB2 pixel_3416/AMP_IN pixel_3416/SF_IB
+ pixel_3416/PIX_OUT pixel_3416/CSA_VREF pixel
Xpixel_2737 pixel_2737/gring pixel_2737/VDD pixel_2737/GND pixel_2737/VREF pixel_2737/ROW_SEL
+ pixel_2737/NB1 pixel_2737/VBIAS pixel_2737/NB2 pixel_2737/AMP_IN pixel_2737/SF_IB
+ pixel_2737/PIX_OUT pixel_2737/CSA_VREF pixel
Xpixel_2726 pixel_2726/gring pixel_2726/VDD pixel_2726/GND pixel_2726/VREF pixel_2726/ROW_SEL
+ pixel_2726/NB1 pixel_2726/VBIAS pixel_2726/NB2 pixel_2726/AMP_IN pixel_2726/SF_IB
+ pixel_2726/PIX_OUT pixel_2726/CSA_VREF pixel
Xpixel_2715 pixel_2715/gring pixel_2715/VDD pixel_2715/GND pixel_2715/VREF pixel_2715/ROW_SEL
+ pixel_2715/NB1 pixel_2715/VBIAS pixel_2715/NB2 pixel_2715/AMP_IN pixel_2715/SF_IB
+ pixel_2715/PIX_OUT pixel_2715/CSA_VREF pixel
Xpixel_2759 pixel_2759/gring pixel_2759/VDD pixel_2759/GND pixel_2759/VREF pixel_2759/ROW_SEL
+ pixel_2759/NB1 pixel_2759/VBIAS pixel_2759/NB2 pixel_2759/AMP_IN pixel_2759/SF_IB
+ pixel_2759/PIX_OUT pixel_2759/CSA_VREF pixel
Xpixel_2748 pixel_2748/gring pixel_2748/VDD pixel_2748/GND pixel_2748/VREF pixel_2748/ROW_SEL
+ pixel_2748/NB1 pixel_2748/VBIAS pixel_2748/NB2 pixel_2748/AMP_IN pixel_2748/SF_IB
+ pixel_2748/PIX_OUT pixel_2748/CSA_VREF pixel
Xpixel_6020 pixel_6020/gring pixel_6020/VDD pixel_6020/GND pixel_6020/VREF pixel_6020/ROW_SEL
+ pixel_6020/NB1 pixel_6020/VBIAS pixel_6020/NB2 pixel_6020/AMP_IN pixel_6020/SF_IB
+ pixel_6020/PIX_OUT pixel_6020/CSA_VREF pixel
Xpixel_6031 pixel_6031/gring pixel_6031/VDD pixel_6031/GND pixel_6031/VREF pixel_6031/ROW_SEL
+ pixel_6031/NB1 pixel_6031/VBIAS pixel_6031/NB2 pixel_6031/AMP_IN pixel_6031/SF_IB
+ pixel_6031/PIX_OUT pixel_6031/CSA_VREF pixel
Xpixel_6042 pixel_6042/gring pixel_6042/VDD pixel_6042/GND pixel_6042/VREF pixel_6042/ROW_SEL
+ pixel_6042/NB1 pixel_6042/VBIAS pixel_6042/NB2 pixel_6042/AMP_IN pixel_6042/SF_IB
+ pixel_6042/PIX_OUT pixel_6042/CSA_VREF pixel
Xpixel_6053 pixel_6053/gring pixel_6053/VDD pixel_6053/GND pixel_6053/VREF pixel_6053/ROW_SEL
+ pixel_6053/NB1 pixel_6053/VBIAS pixel_6053/NB2 pixel_6053/AMP_IN pixel_6053/SF_IB
+ pixel_6053/PIX_OUT pixel_6053/CSA_VREF pixel
Xpixel_6064 pixel_6064/gring pixel_6064/VDD pixel_6064/GND pixel_6064/VREF pixel_6064/ROW_SEL
+ pixel_6064/NB1 pixel_6064/VBIAS pixel_6064/NB2 pixel_6064/AMP_IN pixel_6064/SF_IB
+ pixel_6064/PIX_OUT pixel_6064/CSA_VREF pixel
Xpixel_6075 pixel_6075/gring pixel_6075/VDD pixel_6075/GND pixel_6075/VREF pixel_6075/ROW_SEL
+ pixel_6075/NB1 pixel_6075/VBIAS pixel_6075/NB2 pixel_6075/AMP_IN pixel_6075/SF_IB
+ pixel_6075/PIX_OUT pixel_6075/CSA_VREF pixel
Xpixel_6086 pixel_6086/gring pixel_6086/VDD pixel_6086/GND pixel_6086/VREF pixel_6086/ROW_SEL
+ pixel_6086/NB1 pixel_6086/VBIAS pixel_6086/NB2 pixel_6086/AMP_IN pixel_6086/SF_IB
+ pixel_6086/PIX_OUT pixel_6086/CSA_VREF pixel
Xpixel_5330 pixel_5330/gring pixel_5330/VDD pixel_5330/GND pixel_5330/VREF pixel_5330/ROW_SEL
+ pixel_5330/NB1 pixel_5330/VBIAS pixel_5330/NB2 pixel_5330/AMP_IN pixel_5330/SF_IB
+ pixel_5330/PIX_OUT pixel_5330/CSA_VREF pixel
Xpixel_5341 pixel_5341/gring pixel_5341/VDD pixel_5341/GND pixel_5341/VREF pixel_5341/ROW_SEL
+ pixel_5341/NB1 pixel_5341/VBIAS pixel_5341/NB2 pixel_5341/AMP_IN pixel_5341/SF_IB
+ pixel_5341/PIX_OUT pixel_5341/CSA_VREF pixel
Xpixel_6097 pixel_6097/gring pixel_6097/VDD pixel_6097/GND pixel_6097/VREF pixel_6097/ROW_SEL
+ pixel_6097/NB1 pixel_6097/VBIAS pixel_6097/NB2 pixel_6097/AMP_IN pixel_6097/SF_IB
+ pixel_6097/PIX_OUT pixel_6097/CSA_VREF pixel
Xpixel_5352 pixel_5352/gring pixel_5352/VDD pixel_5352/GND pixel_5352/VREF pixel_5352/ROW_SEL
+ pixel_5352/NB1 pixel_5352/VBIAS pixel_5352/NB2 pixel_5352/AMP_IN pixel_5352/SF_IB
+ pixel_5352/PIX_OUT pixel_5352/CSA_VREF pixel
Xpixel_5363 pixel_5363/gring pixel_5363/VDD pixel_5363/GND pixel_5363/VREF pixel_5363/ROW_SEL
+ pixel_5363/NB1 pixel_5363/VBIAS pixel_5363/NB2 pixel_5363/AMP_IN pixel_5363/SF_IB
+ pixel_5363/PIX_OUT pixel_5363/CSA_VREF pixel
Xpixel_5374 pixel_5374/gring pixel_5374/VDD pixel_5374/GND pixel_5374/VREF pixel_5374/ROW_SEL
+ pixel_5374/NB1 pixel_5374/VBIAS pixel_5374/NB2 pixel_5374/AMP_IN pixel_5374/SF_IB
+ pixel_5374/PIX_OUT pixel_5374/CSA_VREF pixel
Xpixel_5385 pixel_5385/gring pixel_5385/VDD pixel_5385/GND pixel_5385/VREF pixel_5385/ROW_SEL
+ pixel_5385/NB1 pixel_5385/VBIAS pixel_5385/NB2 pixel_5385/AMP_IN pixel_5385/SF_IB
+ pixel_5385/PIX_OUT pixel_5385/CSA_VREF pixel
Xpixel_5396 pixel_5396/gring pixel_5396/VDD pixel_5396/GND pixel_5396/VREF pixel_5396/ROW_SEL
+ pixel_5396/NB1 pixel_5396/VBIAS pixel_5396/NB2 pixel_5396/AMP_IN pixel_5396/SF_IB
+ pixel_5396/PIX_OUT pixel_5396/CSA_VREF pixel
Xpixel_4640 pixel_4640/gring pixel_4640/VDD pixel_4640/GND pixel_4640/VREF pixel_4640/ROW_SEL
+ pixel_4640/NB1 pixel_4640/VBIAS pixel_4640/NB2 pixel_4640/AMP_IN pixel_4640/SF_IB
+ pixel_4640/PIX_OUT pixel_4640/CSA_VREF pixel
Xpixel_4651 pixel_4651/gring pixel_4651/VDD pixel_4651/GND pixel_4651/VREF pixel_4651/ROW_SEL
+ pixel_4651/NB1 pixel_4651/VBIAS pixel_4651/NB2 pixel_4651/AMP_IN pixel_4651/SF_IB
+ pixel_4651/PIX_OUT pixel_4651/CSA_VREF pixel
Xpixel_4662 pixel_4662/gring pixel_4662/VDD pixel_4662/GND pixel_4662/VREF pixel_4662/ROW_SEL
+ pixel_4662/NB1 pixel_4662/VBIAS pixel_4662/NB2 pixel_4662/AMP_IN pixel_4662/SF_IB
+ pixel_4662/PIX_OUT pixel_4662/CSA_VREF pixel
Xpixel_4673 pixel_4673/gring pixel_4673/VDD pixel_4673/GND pixel_4673/VREF pixel_4673/ROW_SEL
+ pixel_4673/NB1 pixel_4673/VBIAS pixel_4673/NB2 pixel_4673/AMP_IN pixel_4673/SF_IB
+ pixel_4673/PIX_OUT pixel_4673/CSA_VREF pixel
Xpixel_690 pixel_690/gring pixel_690/VDD pixel_690/GND pixel_690/VREF pixel_690/ROW_SEL
+ pixel_690/NB1 pixel_690/VBIAS pixel_690/NB2 pixel_690/AMP_IN pixel_690/SF_IB pixel_690/PIX_OUT
+ pixel_690/CSA_VREF pixel
Xpixel_4684 pixel_4684/gring pixel_4684/VDD pixel_4684/GND pixel_4684/VREF pixel_4684/ROW_SEL
+ pixel_4684/NB1 pixel_4684/VBIAS pixel_4684/NB2 pixel_4684/AMP_IN pixel_4684/SF_IB
+ pixel_4684/PIX_OUT pixel_4684/CSA_VREF pixel
Xpixel_4695 pixel_4695/gring pixel_4695/VDD pixel_4695/GND pixel_4695/VREF pixel_4695/ROW_SEL
+ pixel_4695/NB1 pixel_4695/VBIAS pixel_4695/NB2 pixel_4695/AMP_IN pixel_4695/SF_IB
+ pixel_4695/PIX_OUT pixel_4695/CSA_VREF pixel
Xpixel_3950 pixel_3950/gring pixel_3950/VDD pixel_3950/GND pixel_3950/VREF pixel_3950/ROW_SEL
+ pixel_3950/NB1 pixel_3950/VBIAS pixel_3950/NB2 pixel_3950/AMP_IN pixel_3950/SF_IB
+ pixel_3950/PIX_OUT pixel_3950/CSA_VREF pixel
Xpixel_3961 pixel_3961/gring pixel_3961/VDD pixel_3961/GND pixel_3961/VREF pixel_3961/ROW_SEL
+ pixel_3961/NB1 pixel_3961/VBIAS pixel_3961/NB2 pixel_3961/AMP_IN pixel_3961/SF_IB
+ pixel_3961/PIX_OUT pixel_3961/CSA_VREF pixel
Xpixel_3972 pixel_3972/gring pixel_3972/VDD pixel_3972/GND pixel_3972/VREF pixel_3972/ROW_SEL
+ pixel_3972/NB1 pixel_3972/VBIAS pixel_3972/NB2 pixel_3972/AMP_IN pixel_3972/SF_IB
+ pixel_3972/PIX_OUT pixel_3972/CSA_VREF pixel
Xpixel_3983 pixel_3983/gring pixel_3983/VDD pixel_3983/GND pixel_3983/VREF pixel_3983/ROW_SEL
+ pixel_3983/NB1 pixel_3983/VBIAS pixel_3983/NB2 pixel_3983/AMP_IN pixel_3983/SF_IB
+ pixel_3983/PIX_OUT pixel_3983/CSA_VREF pixel
Xpixel_3994 pixel_3994/gring pixel_3994/VDD pixel_3994/GND pixel_3994/VREF pixel_3994/ROW_SEL
+ pixel_3994/NB1 pixel_3994/VBIAS pixel_3994/NB2 pixel_3994/AMP_IN pixel_3994/SF_IB
+ pixel_3994/PIX_OUT pixel_3994/CSA_VREF pixel
Xpixel_4 pixel_4/gring pixel_4/VDD pixel_4/GND pixel_4/VREF pixel_4/ROW_SEL pixel_4/NB1
+ pixel_4/VBIAS pixel_4/NB2 pixel_4/AMP_IN pixel_4/SF_IB pixel_4/PIX_OUT pixel_4/CSA_VREF
+ pixel
Xpixel_9607 pixel_9607/gring pixel_9607/VDD pixel_9607/GND pixel_9607/VREF pixel_9607/ROW_SEL
+ pixel_9607/NB1 pixel_9607/VBIAS pixel_9607/NB2 pixel_9607/AMP_IN pixel_9607/SF_IB
+ pixel_9607/PIX_OUT pixel_9607/CSA_VREF pixel
Xpixel_9618 pixel_9618/gring pixel_9618/VDD pixel_9618/GND pixel_9618/VREF pixel_9618/ROW_SEL
+ pixel_9618/NB1 pixel_9618/VBIAS pixel_9618/NB2 pixel_9618/AMP_IN pixel_9618/SF_IB
+ pixel_9618/PIX_OUT pixel_9618/CSA_VREF pixel
Xpixel_9629 pixel_9629/gring pixel_9629/VDD pixel_9629/GND pixel_9629/VREF pixel_9629/ROW_SEL
+ pixel_9629/NB1 pixel_9629/VBIAS pixel_9629/NB2 pixel_9629/AMP_IN pixel_9629/SF_IB
+ pixel_9629/PIX_OUT pixel_9629/CSA_VREF pixel
Xpixel_8928 pixel_8928/gring pixel_8928/VDD pixel_8928/GND pixel_8928/VREF pixel_8928/ROW_SEL
+ pixel_8928/NB1 pixel_8928/VBIAS pixel_8928/NB2 pixel_8928/AMP_IN pixel_8928/SF_IB
+ pixel_8928/PIX_OUT pixel_8928/CSA_VREF pixel
Xpixel_8917 pixel_8917/gring pixel_8917/VDD pixel_8917/GND pixel_8917/VREF pixel_8917/ROW_SEL
+ pixel_8917/NB1 pixel_8917/VBIAS pixel_8917/NB2 pixel_8917/AMP_IN pixel_8917/SF_IB
+ pixel_8917/PIX_OUT pixel_8917/CSA_VREF pixel
Xpixel_8906 pixel_8906/gring pixel_8906/VDD pixel_8906/GND pixel_8906/VREF pixel_8906/ROW_SEL
+ pixel_8906/NB1 pixel_8906/VBIAS pixel_8906/NB2 pixel_8906/AMP_IN pixel_8906/SF_IB
+ pixel_8906/PIX_OUT pixel_8906/CSA_VREF pixel
Xpixel_8939 pixel_8939/gring pixel_8939/VDD pixel_8939/GND pixel_8939/VREF pixel_8939/ROW_SEL
+ pixel_8939/NB1 pixel_8939/VBIAS pixel_8939/NB2 pixel_8939/AMP_IN pixel_8939/SF_IB
+ pixel_8939/PIX_OUT pixel_8939/CSA_VREF pixel
Xpixel_3224 pixel_3224/gring pixel_3224/VDD pixel_3224/GND pixel_3224/VREF pixel_3224/ROW_SEL
+ pixel_3224/NB1 pixel_3224/VBIAS pixel_3224/NB2 pixel_3224/AMP_IN pixel_3224/SF_IB
+ pixel_3224/PIX_OUT pixel_3224/CSA_VREF pixel
Xpixel_3213 pixel_3213/gring pixel_3213/VDD pixel_3213/GND pixel_3213/VREF pixel_3213/ROW_SEL
+ pixel_3213/NB1 pixel_3213/VBIAS pixel_3213/NB2 pixel_3213/AMP_IN pixel_3213/SF_IB
+ pixel_3213/PIX_OUT pixel_3213/CSA_VREF pixel
Xpixel_3202 pixel_3202/gring pixel_3202/VDD pixel_3202/GND pixel_3202/VREF pixel_3202/ROW_SEL
+ pixel_3202/NB1 pixel_3202/VBIAS pixel_3202/NB2 pixel_3202/AMP_IN pixel_3202/SF_IB
+ pixel_3202/PIX_OUT pixel_3202/CSA_VREF pixel
Xpixel_2512 pixel_2512/gring pixel_2512/VDD pixel_2512/GND pixel_2512/VREF pixel_2512/ROW_SEL
+ pixel_2512/NB1 pixel_2512/VBIAS pixel_2512/NB2 pixel_2512/AMP_IN pixel_2512/SF_IB
+ pixel_2512/PIX_OUT pixel_2512/CSA_VREF pixel
Xpixel_2501 pixel_2501/gring pixel_2501/VDD pixel_2501/GND pixel_2501/VREF pixel_2501/ROW_SEL
+ pixel_2501/NB1 pixel_2501/VBIAS pixel_2501/NB2 pixel_2501/AMP_IN pixel_2501/SF_IB
+ pixel_2501/PIX_OUT pixel_2501/CSA_VREF pixel
Xpixel_3257 pixel_3257/gring pixel_3257/VDD pixel_3257/GND pixel_3257/VREF pixel_3257/ROW_SEL
+ pixel_3257/NB1 pixel_3257/VBIAS pixel_3257/NB2 pixel_3257/AMP_IN pixel_3257/SF_IB
+ pixel_3257/PIX_OUT pixel_3257/CSA_VREF pixel
Xpixel_3246 pixel_3246/gring pixel_3246/VDD pixel_3246/GND pixel_3246/VREF pixel_3246/ROW_SEL
+ pixel_3246/NB1 pixel_3246/VBIAS pixel_3246/NB2 pixel_3246/AMP_IN pixel_3246/SF_IB
+ pixel_3246/PIX_OUT pixel_3246/CSA_VREF pixel
Xpixel_3235 pixel_3235/gring pixel_3235/VDD pixel_3235/GND pixel_3235/VREF pixel_3235/ROW_SEL
+ pixel_3235/NB1 pixel_3235/VBIAS pixel_3235/NB2 pixel_3235/AMP_IN pixel_3235/SF_IB
+ pixel_3235/PIX_OUT pixel_3235/CSA_VREF pixel
Xpixel_1800 pixel_1800/gring pixel_1800/VDD pixel_1800/GND pixel_1800/VREF pixel_1800/ROW_SEL
+ pixel_1800/NB1 pixel_1800/VBIAS pixel_1800/NB2 pixel_1800/AMP_IN pixel_1800/SF_IB
+ pixel_1800/PIX_OUT pixel_1800/CSA_VREF pixel
Xpixel_2545 pixel_2545/gring pixel_2545/VDD pixel_2545/GND pixel_2545/VREF pixel_2545/ROW_SEL
+ pixel_2545/NB1 pixel_2545/VBIAS pixel_2545/NB2 pixel_2545/AMP_IN pixel_2545/SF_IB
+ pixel_2545/PIX_OUT pixel_2545/CSA_VREF pixel
Xpixel_2534 pixel_2534/gring pixel_2534/VDD pixel_2534/GND pixel_2534/VREF pixel_2534/ROW_SEL
+ pixel_2534/NB1 pixel_2534/VBIAS pixel_2534/NB2 pixel_2534/AMP_IN pixel_2534/SF_IB
+ pixel_2534/PIX_OUT pixel_2534/CSA_VREF pixel
Xpixel_2523 pixel_2523/gring pixel_2523/VDD pixel_2523/GND pixel_2523/VREF pixel_2523/ROW_SEL
+ pixel_2523/NB1 pixel_2523/VBIAS pixel_2523/NB2 pixel_2523/AMP_IN pixel_2523/SF_IB
+ pixel_2523/PIX_OUT pixel_2523/CSA_VREF pixel
Xpixel_3279 pixel_3279/gring pixel_3279/VDD pixel_3279/GND pixel_3279/VREF pixel_3279/ROW_SEL
+ pixel_3279/NB1 pixel_3279/VBIAS pixel_3279/NB2 pixel_3279/AMP_IN pixel_3279/SF_IB
+ pixel_3279/PIX_OUT pixel_3279/CSA_VREF pixel
Xpixel_3268 pixel_3268/gring pixel_3268/VDD pixel_3268/GND pixel_3268/VREF pixel_3268/ROW_SEL
+ pixel_3268/NB1 pixel_3268/VBIAS pixel_3268/NB2 pixel_3268/AMP_IN pixel_3268/SF_IB
+ pixel_3268/PIX_OUT pixel_3268/CSA_VREF pixel
Xpixel_1844 pixel_1844/gring pixel_1844/VDD pixel_1844/GND pixel_1844/VREF pixel_1844/ROW_SEL
+ pixel_1844/NB1 pixel_1844/VBIAS pixel_1844/NB2 pixel_1844/AMP_IN pixel_1844/SF_IB
+ pixel_1844/PIX_OUT pixel_1844/CSA_VREF pixel
Xpixel_1833 pixel_1833/gring pixel_1833/VDD pixel_1833/GND pixel_1833/VREF pixel_1833/ROW_SEL
+ pixel_1833/NB1 pixel_1833/VBIAS pixel_1833/NB2 pixel_1833/AMP_IN pixel_1833/SF_IB
+ pixel_1833/PIX_OUT pixel_1833/CSA_VREF pixel
Xpixel_1822 pixel_1822/gring pixel_1822/VDD pixel_1822/GND pixel_1822/VREF pixel_1822/ROW_SEL
+ pixel_1822/NB1 pixel_1822/VBIAS pixel_1822/NB2 pixel_1822/AMP_IN pixel_1822/SF_IB
+ pixel_1822/PIX_OUT pixel_1822/CSA_VREF pixel
Xpixel_1811 pixel_1811/gring pixel_1811/VDD pixel_1811/GND pixel_1811/VREF pixel_1811/ROW_SEL
+ pixel_1811/NB1 pixel_1811/VBIAS pixel_1811/NB2 pixel_1811/AMP_IN pixel_1811/SF_IB
+ pixel_1811/PIX_OUT pixel_1811/CSA_VREF pixel
Xpixel_2589 pixel_2589/gring pixel_2589/VDD pixel_2589/GND pixel_2589/VREF pixel_2589/ROW_SEL
+ pixel_2589/NB1 pixel_2589/VBIAS pixel_2589/NB2 pixel_2589/AMP_IN pixel_2589/SF_IB
+ pixel_2589/PIX_OUT pixel_2589/CSA_VREF pixel
Xpixel_2578 pixel_2578/gring pixel_2578/VDD pixel_2578/GND pixel_2578/VREF pixel_2578/ROW_SEL
+ pixel_2578/NB1 pixel_2578/VBIAS pixel_2578/NB2 pixel_2578/AMP_IN pixel_2578/SF_IB
+ pixel_2578/PIX_OUT pixel_2578/CSA_VREF pixel
Xpixel_2567 pixel_2567/gring pixel_2567/VDD pixel_2567/GND pixel_2567/VREF pixel_2567/ROW_SEL
+ pixel_2567/NB1 pixel_2567/VBIAS pixel_2567/NB2 pixel_2567/AMP_IN pixel_2567/SF_IB
+ pixel_2567/PIX_OUT pixel_2567/CSA_VREF pixel
Xpixel_2556 pixel_2556/gring pixel_2556/VDD pixel_2556/GND pixel_2556/VREF pixel_2556/ROW_SEL
+ pixel_2556/NB1 pixel_2556/VBIAS pixel_2556/NB2 pixel_2556/AMP_IN pixel_2556/SF_IB
+ pixel_2556/PIX_OUT pixel_2556/CSA_VREF pixel
Xpixel_1877 pixel_1877/gring pixel_1877/VDD pixel_1877/GND pixel_1877/VREF pixel_1877/ROW_SEL
+ pixel_1877/NB1 pixel_1877/VBIAS pixel_1877/NB2 pixel_1877/AMP_IN pixel_1877/SF_IB
+ pixel_1877/PIX_OUT pixel_1877/CSA_VREF pixel
Xpixel_1866 pixel_1866/gring pixel_1866/VDD pixel_1866/GND pixel_1866/VREF pixel_1866/ROW_SEL
+ pixel_1866/NB1 pixel_1866/VBIAS pixel_1866/NB2 pixel_1866/AMP_IN pixel_1866/SF_IB
+ pixel_1866/PIX_OUT pixel_1866/CSA_VREF pixel
Xpixel_1855 pixel_1855/gring pixel_1855/VDD pixel_1855/GND pixel_1855/VREF pixel_1855/ROW_SEL
+ pixel_1855/NB1 pixel_1855/VBIAS pixel_1855/NB2 pixel_1855/AMP_IN pixel_1855/SF_IB
+ pixel_1855/PIX_OUT pixel_1855/CSA_VREF pixel
Xpixel_1899 pixel_1899/gring pixel_1899/VDD pixel_1899/GND pixel_1899/VREF pixel_1899/ROW_SEL
+ pixel_1899/NB1 pixel_1899/VBIAS pixel_1899/NB2 pixel_1899/AMP_IN pixel_1899/SF_IB
+ pixel_1899/PIX_OUT pixel_1899/CSA_VREF pixel
Xpixel_1888 pixel_1888/gring pixel_1888/VDD pixel_1888/GND pixel_1888/VREF pixel_1888/ROW_SEL
+ pixel_1888/NB1 pixel_1888/VBIAS pixel_1888/NB2 pixel_1888/AMP_IN pixel_1888/SF_IB
+ pixel_1888/PIX_OUT pixel_1888/CSA_VREF pixel
Xpixel_5160 pixel_5160/gring pixel_5160/VDD pixel_5160/GND pixel_5160/VREF pixel_5160/ROW_SEL
+ pixel_5160/NB1 pixel_5160/VBIAS pixel_5160/NB2 pixel_5160/AMP_IN pixel_5160/SF_IB
+ pixel_5160/PIX_OUT pixel_5160/CSA_VREF pixel
Xpixel_5171 pixel_5171/gring pixel_5171/VDD pixel_5171/GND pixel_5171/VREF pixel_5171/ROW_SEL
+ pixel_5171/NB1 pixel_5171/VBIAS pixel_5171/NB2 pixel_5171/AMP_IN pixel_5171/SF_IB
+ pixel_5171/PIX_OUT pixel_5171/CSA_VREF pixel
Xpixel_5182 pixel_5182/gring pixel_5182/VDD pixel_5182/GND pixel_5182/VREF pixel_5182/ROW_SEL
+ pixel_5182/NB1 pixel_5182/VBIAS pixel_5182/NB2 pixel_5182/AMP_IN pixel_5182/SF_IB
+ pixel_5182/PIX_OUT pixel_5182/CSA_VREF pixel
Xpixel_5193 pixel_5193/gring pixel_5193/VDD pixel_5193/GND pixel_5193/VREF pixel_5193/ROW_SEL
+ pixel_5193/NB1 pixel_5193/VBIAS pixel_5193/NB2 pixel_5193/AMP_IN pixel_5193/SF_IB
+ pixel_5193/PIX_OUT pixel_5193/CSA_VREF pixel
Xpixel_4470 pixel_4470/gring pixel_4470/VDD pixel_4470/GND pixel_4470/VREF pixel_4470/ROW_SEL
+ pixel_4470/NB1 pixel_4470/VBIAS pixel_4470/NB2 pixel_4470/AMP_IN pixel_4470/SF_IB
+ pixel_4470/PIX_OUT pixel_4470/CSA_VREF pixel
Xpixel_4481 pixel_4481/gring pixel_4481/VDD pixel_4481/GND pixel_4481/VREF pixel_4481/ROW_SEL
+ pixel_4481/NB1 pixel_4481/VBIAS pixel_4481/NB2 pixel_4481/AMP_IN pixel_4481/SF_IB
+ pixel_4481/PIX_OUT pixel_4481/CSA_VREF pixel
Xpixel_4492 pixel_4492/gring pixel_4492/VDD pixel_4492/GND pixel_4492/VREF pixel_4492/ROW_SEL
+ pixel_4492/NB1 pixel_4492/VBIAS pixel_4492/NB2 pixel_4492/AMP_IN pixel_4492/SF_IB
+ pixel_4492/PIX_OUT pixel_4492/CSA_VREF pixel
Xpixel_3791 pixel_3791/gring pixel_3791/VDD pixel_3791/GND pixel_3791/VREF pixel_3791/ROW_SEL
+ pixel_3791/NB1 pixel_3791/VBIAS pixel_3791/NB2 pixel_3791/AMP_IN pixel_3791/SF_IB
+ pixel_3791/PIX_OUT pixel_3791/CSA_VREF pixel
Xpixel_3780 pixel_3780/gring pixel_3780/VDD pixel_3780/GND pixel_3780/VREF pixel_3780/ROW_SEL
+ pixel_3780/NB1 pixel_3780/VBIAS pixel_3780/NB2 pixel_3780/AMP_IN pixel_3780/SF_IB
+ pixel_3780/PIX_OUT pixel_3780/CSA_VREF pixel
Xpixel_1129 pixel_1129/gring pixel_1129/VDD pixel_1129/GND pixel_1129/VREF pixel_1129/ROW_SEL
+ pixel_1129/NB1 pixel_1129/VBIAS pixel_1129/NB2 pixel_1129/AMP_IN pixel_1129/SF_IB
+ pixel_1129/PIX_OUT pixel_1129/CSA_VREF pixel
Xpixel_1118 pixel_1118/gring pixel_1118/VDD pixel_1118/GND pixel_1118/VREF pixel_1118/ROW_SEL
+ pixel_1118/NB1 pixel_1118/VBIAS pixel_1118/NB2 pixel_1118/AMP_IN pixel_1118/SF_IB
+ pixel_1118/PIX_OUT pixel_1118/CSA_VREF pixel
Xpixel_1107 pixel_1107/gring pixel_1107/VDD pixel_1107/GND pixel_1107/VREF pixel_1107/ROW_SEL
+ pixel_1107/NB1 pixel_1107/VBIAS pixel_1107/NB2 pixel_1107/AMP_IN pixel_1107/SF_IB
+ pixel_1107/PIX_OUT pixel_1107/CSA_VREF pixel
Xpixel_9404 pixel_9404/gring pixel_9404/VDD pixel_9404/GND pixel_9404/VREF pixel_9404/ROW_SEL
+ pixel_9404/NB1 pixel_9404/VBIAS pixel_9404/NB2 pixel_9404/AMP_IN pixel_9404/SF_IB
+ pixel_9404/PIX_OUT pixel_9404/CSA_VREF pixel
Xpixel_8703 pixel_8703/gring pixel_8703/VDD pixel_8703/GND pixel_8703/VREF pixel_8703/ROW_SEL
+ pixel_8703/NB1 pixel_8703/VBIAS pixel_8703/NB2 pixel_8703/AMP_IN pixel_8703/SF_IB
+ pixel_8703/PIX_OUT pixel_8703/CSA_VREF pixel
Xpixel_9437 pixel_9437/gring pixel_9437/VDD pixel_9437/GND pixel_9437/VREF pixel_9437/ROW_SEL
+ pixel_9437/NB1 pixel_9437/VBIAS pixel_9437/NB2 pixel_9437/AMP_IN pixel_9437/SF_IB
+ pixel_9437/PIX_OUT pixel_9437/CSA_VREF pixel
Xpixel_9426 pixel_9426/gring pixel_9426/VDD pixel_9426/GND pixel_9426/VREF pixel_9426/ROW_SEL
+ pixel_9426/NB1 pixel_9426/VBIAS pixel_9426/NB2 pixel_9426/AMP_IN pixel_9426/SF_IB
+ pixel_9426/PIX_OUT pixel_9426/CSA_VREF pixel
Xpixel_9415 pixel_9415/gring pixel_9415/VDD pixel_9415/GND pixel_9415/VREF pixel_9415/ROW_SEL
+ pixel_9415/NB1 pixel_9415/VBIAS pixel_9415/NB2 pixel_9415/AMP_IN pixel_9415/SF_IB
+ pixel_9415/PIX_OUT pixel_9415/CSA_VREF pixel
Xpixel_8736 pixel_8736/gring pixel_8736/VDD pixel_8736/GND pixel_8736/VREF pixel_8736/ROW_SEL
+ pixel_8736/NB1 pixel_8736/VBIAS pixel_8736/NB2 pixel_8736/AMP_IN pixel_8736/SF_IB
+ pixel_8736/PIX_OUT pixel_8736/CSA_VREF pixel
Xpixel_8725 pixel_8725/gring pixel_8725/VDD pixel_8725/GND pixel_8725/VREF pixel_8725/ROW_SEL
+ pixel_8725/NB1 pixel_8725/VBIAS pixel_8725/NB2 pixel_8725/AMP_IN pixel_8725/SF_IB
+ pixel_8725/PIX_OUT pixel_8725/CSA_VREF pixel
Xpixel_8714 pixel_8714/gring pixel_8714/VDD pixel_8714/GND pixel_8714/VREF pixel_8714/ROW_SEL
+ pixel_8714/NB1 pixel_8714/VBIAS pixel_8714/NB2 pixel_8714/AMP_IN pixel_8714/SF_IB
+ pixel_8714/PIX_OUT pixel_8714/CSA_VREF pixel
Xpixel_9459 pixel_9459/gring pixel_9459/VDD pixel_9459/GND pixel_9459/VREF pixel_9459/ROW_SEL
+ pixel_9459/NB1 pixel_9459/VBIAS pixel_9459/NB2 pixel_9459/AMP_IN pixel_9459/SF_IB
+ pixel_9459/PIX_OUT pixel_9459/CSA_VREF pixel
Xpixel_9448 pixel_9448/gring pixel_9448/VDD pixel_9448/GND pixel_9448/VREF pixel_9448/ROW_SEL
+ pixel_9448/NB1 pixel_9448/VBIAS pixel_9448/NB2 pixel_9448/AMP_IN pixel_9448/SF_IB
+ pixel_9448/PIX_OUT pixel_9448/CSA_VREF pixel
Xpixel_8769 pixel_8769/gring pixel_8769/VDD pixel_8769/GND pixel_8769/VREF pixel_8769/ROW_SEL
+ pixel_8769/NB1 pixel_8769/VBIAS pixel_8769/NB2 pixel_8769/AMP_IN pixel_8769/SF_IB
+ pixel_8769/PIX_OUT pixel_8769/CSA_VREF pixel
Xpixel_8758 pixel_8758/gring pixel_8758/VDD pixel_8758/GND pixel_8758/VREF pixel_8758/ROW_SEL
+ pixel_8758/NB1 pixel_8758/VBIAS pixel_8758/NB2 pixel_8758/AMP_IN pixel_8758/SF_IB
+ pixel_8758/PIX_OUT pixel_8758/CSA_VREF pixel
Xpixel_8747 pixel_8747/gring pixel_8747/VDD pixel_8747/GND pixel_8747/VREF pixel_8747/ROW_SEL
+ pixel_8747/NB1 pixel_8747/VBIAS pixel_8747/NB2 pixel_8747/AMP_IN pixel_8747/SF_IB
+ pixel_8747/PIX_OUT pixel_8747/CSA_VREF pixel
Xpixel_3032 pixel_3032/gring pixel_3032/VDD pixel_3032/GND pixel_3032/VREF pixel_3032/ROW_SEL
+ pixel_3032/NB1 pixel_3032/VBIAS pixel_3032/NB2 pixel_3032/AMP_IN pixel_3032/SF_IB
+ pixel_3032/PIX_OUT pixel_3032/CSA_VREF pixel
Xpixel_3021 pixel_3021/gring pixel_3021/VDD pixel_3021/GND pixel_3021/VREF pixel_3021/ROW_SEL
+ pixel_3021/NB1 pixel_3021/VBIAS pixel_3021/NB2 pixel_3021/AMP_IN pixel_3021/SF_IB
+ pixel_3021/PIX_OUT pixel_3021/CSA_VREF pixel
Xpixel_3010 pixel_3010/gring pixel_3010/VDD pixel_3010/GND pixel_3010/VREF pixel_3010/ROW_SEL
+ pixel_3010/NB1 pixel_3010/VBIAS pixel_3010/NB2 pixel_3010/AMP_IN pixel_3010/SF_IB
+ pixel_3010/PIX_OUT pixel_3010/CSA_VREF pixel
Xpixel_2320 pixel_2320/gring pixel_2320/VDD pixel_2320/GND pixel_2320/VREF pixel_2320/ROW_SEL
+ pixel_2320/NB1 pixel_2320/VBIAS pixel_2320/NB2 pixel_2320/AMP_IN pixel_2320/SF_IB
+ pixel_2320/PIX_OUT pixel_2320/CSA_VREF pixel
Xpixel_3065 pixel_3065/gring pixel_3065/VDD pixel_3065/GND pixel_3065/VREF pixel_3065/ROW_SEL
+ pixel_3065/NB1 pixel_3065/VBIAS pixel_3065/NB2 pixel_3065/AMP_IN pixel_3065/SF_IB
+ pixel_3065/PIX_OUT pixel_3065/CSA_VREF pixel
Xpixel_3054 pixel_3054/gring pixel_3054/VDD pixel_3054/GND pixel_3054/VREF pixel_3054/ROW_SEL
+ pixel_3054/NB1 pixel_3054/VBIAS pixel_3054/NB2 pixel_3054/AMP_IN pixel_3054/SF_IB
+ pixel_3054/PIX_OUT pixel_3054/CSA_VREF pixel
Xpixel_3043 pixel_3043/gring pixel_3043/VDD pixel_3043/GND pixel_3043/VREF pixel_3043/ROW_SEL
+ pixel_3043/NB1 pixel_3043/VBIAS pixel_3043/NB2 pixel_3043/AMP_IN pixel_3043/SF_IB
+ pixel_3043/PIX_OUT pixel_3043/CSA_VREF pixel
Xpixel_2364 pixel_2364/gring pixel_2364/VDD pixel_2364/GND pixel_2364/VREF pixel_2364/ROW_SEL
+ pixel_2364/NB1 pixel_2364/VBIAS pixel_2364/NB2 pixel_2364/AMP_IN pixel_2364/SF_IB
+ pixel_2364/PIX_OUT pixel_2364/CSA_VREF pixel
Xpixel_2353 pixel_2353/gring pixel_2353/VDD pixel_2353/GND pixel_2353/VREF pixel_2353/ROW_SEL
+ pixel_2353/NB1 pixel_2353/VBIAS pixel_2353/NB2 pixel_2353/AMP_IN pixel_2353/SF_IB
+ pixel_2353/PIX_OUT pixel_2353/CSA_VREF pixel
Xpixel_2342 pixel_2342/gring pixel_2342/VDD pixel_2342/GND pixel_2342/VREF pixel_2342/ROW_SEL
+ pixel_2342/NB1 pixel_2342/VBIAS pixel_2342/NB2 pixel_2342/AMP_IN pixel_2342/SF_IB
+ pixel_2342/PIX_OUT pixel_2342/CSA_VREF pixel
Xpixel_2331 pixel_2331/gring pixel_2331/VDD pixel_2331/GND pixel_2331/VREF pixel_2331/ROW_SEL
+ pixel_2331/NB1 pixel_2331/VBIAS pixel_2331/NB2 pixel_2331/AMP_IN pixel_2331/SF_IB
+ pixel_2331/PIX_OUT pixel_2331/CSA_VREF pixel
Xpixel_3098 pixel_3098/gring pixel_3098/VDD pixel_3098/GND pixel_3098/VREF pixel_3098/ROW_SEL
+ pixel_3098/NB1 pixel_3098/VBIAS pixel_3098/NB2 pixel_3098/AMP_IN pixel_3098/SF_IB
+ pixel_3098/PIX_OUT pixel_3098/CSA_VREF pixel
Xpixel_3087 pixel_3087/gring pixel_3087/VDD pixel_3087/GND pixel_3087/VREF pixel_3087/ROW_SEL
+ pixel_3087/NB1 pixel_3087/VBIAS pixel_3087/NB2 pixel_3087/AMP_IN pixel_3087/SF_IB
+ pixel_3087/PIX_OUT pixel_3087/CSA_VREF pixel
Xpixel_3076 pixel_3076/gring pixel_3076/VDD pixel_3076/GND pixel_3076/VREF pixel_3076/ROW_SEL
+ pixel_3076/NB1 pixel_3076/VBIAS pixel_3076/NB2 pixel_3076/AMP_IN pixel_3076/SF_IB
+ pixel_3076/PIX_OUT pixel_3076/CSA_VREF pixel
Xpixel_1652 pixel_1652/gring pixel_1652/VDD pixel_1652/GND pixel_1652/VREF pixel_1652/ROW_SEL
+ pixel_1652/NB1 pixel_1652/VBIAS pixel_1652/NB2 pixel_1652/AMP_IN pixel_1652/SF_IB
+ pixel_1652/PIX_OUT pixel_1652/CSA_VREF pixel
Xpixel_1641 pixel_1641/gring pixel_1641/VDD pixel_1641/GND pixel_1641/VREF pixel_1641/ROW_SEL
+ pixel_1641/NB1 pixel_1641/VBIAS pixel_1641/NB2 pixel_1641/AMP_IN pixel_1641/SF_IB
+ pixel_1641/PIX_OUT pixel_1641/CSA_VREF pixel
Xpixel_1630 pixel_1630/gring pixel_1630/VDD pixel_1630/GND pixel_1630/VREF pixel_1630/ROW_SEL
+ pixel_1630/NB1 pixel_1630/VBIAS pixel_1630/NB2 pixel_1630/AMP_IN pixel_1630/SF_IB
+ pixel_1630/PIX_OUT pixel_1630/CSA_VREF pixel
Xpixel_2397 pixel_2397/gring pixel_2397/VDD pixel_2397/GND pixel_2397/VREF pixel_2397/ROW_SEL
+ pixel_2397/NB1 pixel_2397/VBIAS pixel_2397/NB2 pixel_2397/AMP_IN pixel_2397/SF_IB
+ pixel_2397/PIX_OUT pixel_2397/CSA_VREF pixel
Xpixel_2386 pixel_2386/gring pixel_2386/VDD pixel_2386/GND pixel_2386/VREF pixel_2386/ROW_SEL
+ pixel_2386/NB1 pixel_2386/VBIAS pixel_2386/NB2 pixel_2386/AMP_IN pixel_2386/SF_IB
+ pixel_2386/PIX_OUT pixel_2386/CSA_VREF pixel
Xpixel_2375 pixel_2375/gring pixel_2375/VDD pixel_2375/GND pixel_2375/VREF pixel_2375/ROW_SEL
+ pixel_2375/NB1 pixel_2375/VBIAS pixel_2375/NB2 pixel_2375/AMP_IN pixel_2375/SF_IB
+ pixel_2375/PIX_OUT pixel_2375/CSA_VREF pixel
Xpixel_1685 pixel_1685/gring pixel_1685/VDD pixel_1685/GND pixel_1685/VREF pixel_1685/ROW_SEL
+ pixel_1685/NB1 pixel_1685/VBIAS pixel_1685/NB2 pixel_1685/AMP_IN pixel_1685/SF_IB
+ pixel_1685/PIX_OUT pixel_1685/CSA_VREF pixel
Xpixel_1674 pixel_1674/gring pixel_1674/VDD pixel_1674/GND pixel_1674/VREF pixel_1674/ROW_SEL
+ pixel_1674/NB1 pixel_1674/VBIAS pixel_1674/NB2 pixel_1674/AMP_IN pixel_1674/SF_IB
+ pixel_1674/PIX_OUT pixel_1674/CSA_VREF pixel
Xpixel_1663 pixel_1663/gring pixel_1663/VDD pixel_1663/GND pixel_1663/VREF pixel_1663/ROW_SEL
+ pixel_1663/NB1 pixel_1663/VBIAS pixel_1663/NB2 pixel_1663/AMP_IN pixel_1663/SF_IB
+ pixel_1663/PIX_OUT pixel_1663/CSA_VREF pixel
Xpixel_1696 pixel_1696/gring pixel_1696/VDD pixel_1696/GND pixel_1696/VREF pixel_1696/ROW_SEL
+ pixel_1696/NB1 pixel_1696/VBIAS pixel_1696/NB2 pixel_1696/AMP_IN pixel_1696/SF_IB
+ pixel_1696/PIX_OUT pixel_1696/CSA_VREF pixel
Xpixel_9960 pixel_9960/gring pixel_9960/VDD pixel_9960/GND pixel_9960/VREF pixel_9960/ROW_SEL
+ pixel_9960/NB1 pixel_9960/VBIAS pixel_9960/NB2 pixel_9960/AMP_IN pixel_9960/SF_IB
+ pixel_9960/PIX_OUT pixel_9960/CSA_VREF pixel
Xpixel_9971 pixel_9971/gring pixel_9971/VDD pixel_9971/GND pixel_9971/VREF pixel_9971/ROW_SEL
+ pixel_9971/NB1 pixel_9971/VBIAS pixel_9971/NB2 pixel_9971/AMP_IN pixel_9971/SF_IB
+ pixel_9971/PIX_OUT pixel_9971/CSA_VREF pixel
Xpixel_9982 pixel_9982/gring pixel_9982/VDD pixel_9982/GND pixel_9982/VREF pixel_9982/ROW_SEL
+ pixel_9982/NB1 pixel_9982/VBIAS pixel_9982/NB2 pixel_9982/AMP_IN pixel_9982/SF_IB
+ pixel_9982/PIX_OUT pixel_9982/CSA_VREF pixel
Xpixel_9993 pixel_9993/gring pixel_9993/VDD pixel_9993/GND pixel_9993/VREF pixel_9993/ROW_SEL
+ pixel_9993/NB1 pixel_9993/VBIAS pixel_9993/NB2 pixel_9993/AMP_IN pixel_9993/SF_IB
+ pixel_9993/PIX_OUT pixel_9993/CSA_VREF pixel
Xpixel_7309 pixel_7309/gring pixel_7309/VDD pixel_7309/GND pixel_7309/VREF pixel_7309/ROW_SEL
+ pixel_7309/NB1 pixel_7309/VBIAS pixel_7309/NB2 pixel_7309/AMP_IN pixel_7309/SF_IB
+ pixel_7309/PIX_OUT pixel_7309/CSA_VREF pixel
Xpixel_6608 pixel_6608/gring pixel_6608/VDD pixel_6608/GND pixel_6608/VREF pixel_6608/ROW_SEL
+ pixel_6608/NB1 pixel_6608/VBIAS pixel_6608/NB2 pixel_6608/AMP_IN pixel_6608/SF_IB
+ pixel_6608/PIX_OUT pixel_6608/CSA_VREF pixel
Xpixel_6619 pixel_6619/gring pixel_6619/VDD pixel_6619/GND pixel_6619/VREF pixel_6619/ROW_SEL
+ pixel_6619/NB1 pixel_6619/VBIAS pixel_6619/NB2 pixel_6619/AMP_IN pixel_6619/SF_IB
+ pixel_6619/PIX_OUT pixel_6619/CSA_VREF pixel
Xpixel_5907 pixel_5907/gring pixel_5907/VDD pixel_5907/GND pixel_5907/VREF pixel_5907/ROW_SEL
+ pixel_5907/NB1 pixel_5907/VBIAS pixel_5907/NB2 pixel_5907/AMP_IN pixel_5907/SF_IB
+ pixel_5907/PIX_OUT pixel_5907/CSA_VREF pixel
Xpixel_5918 pixel_5918/gring pixel_5918/VDD pixel_5918/GND pixel_5918/VREF pixel_5918/ROW_SEL
+ pixel_5918/NB1 pixel_5918/VBIAS pixel_5918/NB2 pixel_5918/AMP_IN pixel_5918/SF_IB
+ pixel_5918/PIX_OUT pixel_5918/CSA_VREF pixel
Xpixel_5929 pixel_5929/gring pixel_5929/VDD pixel_5929/GND pixel_5929/VREF pixel_5929/ROW_SEL
+ pixel_5929/NB1 pixel_5929/VBIAS pixel_5929/NB2 pixel_5929/AMP_IN pixel_5929/SF_IB
+ pixel_5929/PIX_OUT pixel_5929/CSA_VREF pixel
Xpixel_9212 pixel_9212/gring pixel_9212/VDD pixel_9212/GND pixel_9212/VREF pixel_9212/ROW_SEL
+ pixel_9212/NB1 pixel_9212/VBIAS pixel_9212/NB2 pixel_9212/AMP_IN pixel_9212/SF_IB
+ pixel_9212/PIX_OUT pixel_9212/CSA_VREF pixel
Xpixel_9201 pixel_9201/gring pixel_9201/VDD pixel_9201/GND pixel_9201/VREF pixel_9201/ROW_SEL
+ pixel_9201/NB1 pixel_9201/VBIAS pixel_9201/NB2 pixel_9201/AMP_IN pixel_9201/SF_IB
+ pixel_9201/PIX_OUT pixel_9201/CSA_VREF pixel
Xpixel_8511 pixel_8511/gring pixel_8511/VDD pixel_8511/GND pixel_8511/VREF pixel_8511/ROW_SEL
+ pixel_8511/NB1 pixel_8511/VBIAS pixel_8511/NB2 pixel_8511/AMP_IN pixel_8511/SF_IB
+ pixel_8511/PIX_OUT pixel_8511/CSA_VREF pixel
Xpixel_8500 pixel_8500/gring pixel_8500/VDD pixel_8500/GND pixel_8500/VREF pixel_8500/ROW_SEL
+ pixel_8500/NB1 pixel_8500/VBIAS pixel_8500/NB2 pixel_8500/AMP_IN pixel_8500/SF_IB
+ pixel_8500/PIX_OUT pixel_8500/CSA_VREF pixel
Xpixel_9256 pixel_9256/gring pixel_9256/VDD pixel_9256/GND pixel_9256/VREF pixel_9256/ROW_SEL
+ pixel_9256/NB1 pixel_9256/VBIAS pixel_9256/NB2 pixel_9256/AMP_IN pixel_9256/SF_IB
+ pixel_9256/PIX_OUT pixel_9256/CSA_VREF pixel
Xpixel_9245 pixel_9245/gring pixel_9245/VDD pixel_9245/GND pixel_9245/VREF pixel_9245/ROW_SEL
+ pixel_9245/NB1 pixel_9245/VBIAS pixel_9245/NB2 pixel_9245/AMP_IN pixel_9245/SF_IB
+ pixel_9245/PIX_OUT pixel_9245/CSA_VREF pixel
Xpixel_9234 pixel_9234/gring pixel_9234/VDD pixel_9234/GND pixel_9234/VREF pixel_9234/ROW_SEL
+ pixel_9234/NB1 pixel_9234/VBIAS pixel_9234/NB2 pixel_9234/AMP_IN pixel_9234/SF_IB
+ pixel_9234/PIX_OUT pixel_9234/CSA_VREF pixel
Xpixel_9223 pixel_9223/gring pixel_9223/VDD pixel_9223/GND pixel_9223/VREF pixel_9223/ROW_SEL
+ pixel_9223/NB1 pixel_9223/VBIAS pixel_9223/NB2 pixel_9223/AMP_IN pixel_9223/SF_IB
+ pixel_9223/PIX_OUT pixel_9223/CSA_VREF pixel
Xpixel_8544 pixel_8544/gring pixel_8544/VDD pixel_8544/GND pixel_8544/VREF pixel_8544/ROW_SEL
+ pixel_8544/NB1 pixel_8544/VBIAS pixel_8544/NB2 pixel_8544/AMP_IN pixel_8544/SF_IB
+ pixel_8544/PIX_OUT pixel_8544/CSA_VREF pixel
Xpixel_8533 pixel_8533/gring pixel_8533/VDD pixel_8533/GND pixel_8533/VREF pixel_8533/ROW_SEL
+ pixel_8533/NB1 pixel_8533/VBIAS pixel_8533/NB2 pixel_8533/AMP_IN pixel_8533/SF_IB
+ pixel_8533/PIX_OUT pixel_8533/CSA_VREF pixel
Xpixel_8522 pixel_8522/gring pixel_8522/VDD pixel_8522/GND pixel_8522/VREF pixel_8522/ROW_SEL
+ pixel_8522/NB1 pixel_8522/VBIAS pixel_8522/NB2 pixel_8522/AMP_IN pixel_8522/SF_IB
+ pixel_8522/PIX_OUT pixel_8522/CSA_VREF pixel
Xpixel_9289 pixel_9289/gring pixel_9289/VDD pixel_9289/GND pixel_9289/VREF pixel_9289/ROW_SEL
+ pixel_9289/NB1 pixel_9289/VBIAS pixel_9289/NB2 pixel_9289/AMP_IN pixel_9289/SF_IB
+ pixel_9289/PIX_OUT pixel_9289/CSA_VREF pixel
Xpixel_9278 pixel_9278/gring pixel_9278/VDD pixel_9278/GND pixel_9278/VREF pixel_9278/ROW_SEL
+ pixel_9278/NB1 pixel_9278/VBIAS pixel_9278/NB2 pixel_9278/AMP_IN pixel_9278/SF_IB
+ pixel_9278/PIX_OUT pixel_9278/CSA_VREF pixel
Xpixel_9267 pixel_9267/gring pixel_9267/VDD pixel_9267/GND pixel_9267/VREF pixel_9267/ROW_SEL
+ pixel_9267/NB1 pixel_9267/VBIAS pixel_9267/NB2 pixel_9267/AMP_IN pixel_9267/SF_IB
+ pixel_9267/PIX_OUT pixel_9267/CSA_VREF pixel
Xpixel_8577 pixel_8577/gring pixel_8577/VDD pixel_8577/GND pixel_8577/VREF pixel_8577/ROW_SEL
+ pixel_8577/NB1 pixel_8577/VBIAS pixel_8577/NB2 pixel_8577/AMP_IN pixel_8577/SF_IB
+ pixel_8577/PIX_OUT pixel_8577/CSA_VREF pixel
Xpixel_8566 pixel_8566/gring pixel_8566/VDD pixel_8566/GND pixel_8566/VREF pixel_8566/ROW_SEL
+ pixel_8566/NB1 pixel_8566/VBIAS pixel_8566/NB2 pixel_8566/AMP_IN pixel_8566/SF_IB
+ pixel_8566/PIX_OUT pixel_8566/CSA_VREF pixel
Xpixel_8555 pixel_8555/gring pixel_8555/VDD pixel_8555/GND pixel_8555/VREF pixel_8555/ROW_SEL
+ pixel_8555/NB1 pixel_8555/VBIAS pixel_8555/NB2 pixel_8555/AMP_IN pixel_8555/SF_IB
+ pixel_8555/PIX_OUT pixel_8555/CSA_VREF pixel
Xpixel_7810 pixel_7810/gring pixel_7810/VDD pixel_7810/GND pixel_7810/VREF pixel_7810/ROW_SEL
+ pixel_7810/NB1 pixel_7810/VBIAS pixel_7810/NB2 pixel_7810/AMP_IN pixel_7810/SF_IB
+ pixel_7810/PIX_OUT pixel_7810/CSA_VREF pixel
Xpixel_7821 pixel_7821/gring pixel_7821/VDD pixel_7821/GND pixel_7821/VREF pixel_7821/ROW_SEL
+ pixel_7821/NB1 pixel_7821/VBIAS pixel_7821/NB2 pixel_7821/AMP_IN pixel_7821/SF_IB
+ pixel_7821/PIX_OUT pixel_7821/CSA_VREF pixel
Xpixel_7832 pixel_7832/gring pixel_7832/VDD pixel_7832/GND pixel_7832/VREF pixel_7832/ROW_SEL
+ pixel_7832/NB1 pixel_7832/VBIAS pixel_7832/NB2 pixel_7832/AMP_IN pixel_7832/SF_IB
+ pixel_7832/PIX_OUT pixel_7832/CSA_VREF pixel
Xpixel_7843 pixel_7843/gring pixel_7843/VDD pixel_7843/GND pixel_7843/VREF pixel_7843/ROW_SEL
+ pixel_7843/NB1 pixel_7843/VBIAS pixel_7843/NB2 pixel_7843/AMP_IN pixel_7843/SF_IB
+ pixel_7843/PIX_OUT pixel_7843/CSA_VREF pixel
Xpixel_8599 pixel_8599/gring pixel_8599/VDD pixel_8599/GND pixel_8599/VREF pixel_8599/ROW_SEL
+ pixel_8599/NB1 pixel_8599/VBIAS pixel_8599/NB2 pixel_8599/AMP_IN pixel_8599/SF_IB
+ pixel_8599/PIX_OUT pixel_8599/CSA_VREF pixel
Xpixel_8588 pixel_8588/gring pixel_8588/VDD pixel_8588/GND pixel_8588/VREF pixel_8588/ROW_SEL
+ pixel_8588/NB1 pixel_8588/VBIAS pixel_8588/NB2 pixel_8588/AMP_IN pixel_8588/SF_IB
+ pixel_8588/PIX_OUT pixel_8588/CSA_VREF pixel
Xpixel_7854 pixel_7854/gring pixel_7854/VDD pixel_7854/GND pixel_7854/VREF pixel_7854/ROW_SEL
+ pixel_7854/NB1 pixel_7854/VBIAS pixel_7854/NB2 pixel_7854/AMP_IN pixel_7854/SF_IB
+ pixel_7854/PIX_OUT pixel_7854/CSA_VREF pixel
Xpixel_7865 pixel_7865/gring pixel_7865/VDD pixel_7865/GND pixel_7865/VREF pixel_7865/ROW_SEL
+ pixel_7865/NB1 pixel_7865/VBIAS pixel_7865/NB2 pixel_7865/AMP_IN pixel_7865/SF_IB
+ pixel_7865/PIX_OUT pixel_7865/CSA_VREF pixel
Xpixel_7876 pixel_7876/gring pixel_7876/VDD pixel_7876/GND pixel_7876/VREF pixel_7876/ROW_SEL
+ pixel_7876/NB1 pixel_7876/VBIAS pixel_7876/NB2 pixel_7876/AMP_IN pixel_7876/SF_IB
+ pixel_7876/PIX_OUT pixel_7876/CSA_VREF pixel
Xpixel_7887 pixel_7887/gring pixel_7887/VDD pixel_7887/GND pixel_7887/VREF pixel_7887/ROW_SEL
+ pixel_7887/NB1 pixel_7887/VBIAS pixel_7887/NB2 pixel_7887/AMP_IN pixel_7887/SF_IB
+ pixel_7887/PIX_OUT pixel_7887/CSA_VREF pixel
Xpixel_7898 pixel_7898/gring pixel_7898/VDD pixel_7898/GND pixel_7898/VREF pixel_7898/ROW_SEL
+ pixel_7898/NB1 pixel_7898/VBIAS pixel_7898/NB2 pixel_7898/AMP_IN pixel_7898/SF_IB
+ pixel_7898/PIX_OUT pixel_7898/CSA_VREF pixel
Xpixel_2172 pixel_2172/gring pixel_2172/VDD pixel_2172/GND pixel_2172/VREF pixel_2172/ROW_SEL
+ pixel_2172/NB1 pixel_2172/VBIAS pixel_2172/NB2 pixel_2172/AMP_IN pixel_2172/SF_IB
+ pixel_2172/PIX_OUT pixel_2172/CSA_VREF pixel
Xpixel_2161 pixel_2161/gring pixel_2161/VDD pixel_2161/GND pixel_2161/VREF pixel_2161/ROW_SEL
+ pixel_2161/NB1 pixel_2161/VBIAS pixel_2161/NB2 pixel_2161/AMP_IN pixel_2161/SF_IB
+ pixel_2161/PIX_OUT pixel_2161/CSA_VREF pixel
Xpixel_2150 pixel_2150/gring pixel_2150/VDD pixel_2150/GND pixel_2150/VREF pixel_2150/ROW_SEL
+ pixel_2150/NB1 pixel_2150/VBIAS pixel_2150/NB2 pixel_2150/AMP_IN pixel_2150/SF_IB
+ pixel_2150/PIX_OUT pixel_2150/CSA_VREF pixel
Xpixel_1460 pixel_1460/gring pixel_1460/VDD pixel_1460/GND pixel_1460/VREF pixel_1460/ROW_SEL
+ pixel_1460/NB1 pixel_1460/VBIAS pixel_1460/NB2 pixel_1460/AMP_IN pixel_1460/SF_IB
+ pixel_1460/PIX_OUT pixel_1460/CSA_VREF pixel
Xpixel_2194 pixel_2194/gring pixel_2194/VDD pixel_2194/GND pixel_2194/VREF pixel_2194/ROW_SEL
+ pixel_2194/NB1 pixel_2194/VBIAS pixel_2194/NB2 pixel_2194/AMP_IN pixel_2194/SF_IB
+ pixel_2194/PIX_OUT pixel_2194/CSA_VREF pixel
Xpixel_2183 pixel_2183/gring pixel_2183/VDD pixel_2183/GND pixel_2183/VREF pixel_2183/ROW_SEL
+ pixel_2183/NB1 pixel_2183/VBIAS pixel_2183/NB2 pixel_2183/AMP_IN pixel_2183/SF_IB
+ pixel_2183/PIX_OUT pixel_2183/CSA_VREF pixel
Xpixel_1493 pixel_1493/gring pixel_1493/VDD pixel_1493/GND pixel_1493/VREF pixel_1493/ROW_SEL
+ pixel_1493/NB1 pixel_1493/VBIAS pixel_1493/NB2 pixel_1493/AMP_IN pixel_1493/SF_IB
+ pixel_1493/PIX_OUT pixel_1493/CSA_VREF pixel
Xpixel_1482 pixel_1482/gring pixel_1482/VDD pixel_1482/GND pixel_1482/VREF pixel_1482/ROW_SEL
+ pixel_1482/NB1 pixel_1482/VBIAS pixel_1482/NB2 pixel_1482/AMP_IN pixel_1482/SF_IB
+ pixel_1482/PIX_OUT pixel_1482/CSA_VREF pixel
Xpixel_1471 pixel_1471/gring pixel_1471/VDD pixel_1471/GND pixel_1471/VREF pixel_1471/ROW_SEL
+ pixel_1471/NB1 pixel_1471/VBIAS pixel_1471/NB2 pixel_1471/AMP_IN pixel_1471/SF_IB
+ pixel_1471/PIX_OUT pixel_1471/CSA_VREF pixel
Xpixel_9790 pixel_9790/gring pixel_9790/VDD pixel_9790/GND pixel_9790/VREF pixel_9790/ROW_SEL
+ pixel_9790/NB1 pixel_9790/VBIAS pixel_9790/NB2 pixel_9790/AMP_IN pixel_9790/SF_IB
+ pixel_9790/PIX_OUT pixel_9790/CSA_VREF pixel
Xpixel_519 pixel_519/gring pixel_519/VDD pixel_519/GND pixel_519/VREF pixel_519/ROW_SEL
+ pixel_519/NB1 pixel_519/VBIAS pixel_519/NB2 pixel_519/AMP_IN pixel_519/SF_IB pixel_519/PIX_OUT
+ pixel_519/CSA_VREF pixel
Xpixel_508 pixel_508/gring pixel_508/VDD pixel_508/GND pixel_508/VREF pixel_508/ROW_SEL
+ pixel_508/NB1 pixel_508/VBIAS pixel_508/NB2 pixel_508/AMP_IN pixel_508/SF_IB pixel_508/PIX_OUT
+ pixel_508/CSA_VREF pixel
Xpixel_7106 pixel_7106/gring pixel_7106/VDD pixel_7106/GND pixel_7106/VREF pixel_7106/ROW_SEL
+ pixel_7106/NB1 pixel_7106/VBIAS pixel_7106/NB2 pixel_7106/AMP_IN pixel_7106/SF_IB
+ pixel_7106/PIX_OUT pixel_7106/CSA_VREF pixel
Xpixel_7117 pixel_7117/gring pixel_7117/VDD pixel_7117/GND pixel_7117/VREF pixel_7117/ROW_SEL
+ pixel_7117/NB1 pixel_7117/VBIAS pixel_7117/NB2 pixel_7117/AMP_IN pixel_7117/SF_IB
+ pixel_7117/PIX_OUT pixel_7117/CSA_VREF pixel
Xpixel_7128 pixel_7128/gring pixel_7128/VDD pixel_7128/GND pixel_7128/VREF pixel_7128/ROW_SEL
+ pixel_7128/NB1 pixel_7128/VBIAS pixel_7128/NB2 pixel_7128/AMP_IN pixel_7128/SF_IB
+ pixel_7128/PIX_OUT pixel_7128/CSA_VREF pixel
Xpixel_7139 pixel_7139/gring pixel_7139/VDD pixel_7139/GND pixel_7139/VREF pixel_7139/ROW_SEL
+ pixel_7139/NB1 pixel_7139/VBIAS pixel_7139/NB2 pixel_7139/AMP_IN pixel_7139/SF_IB
+ pixel_7139/PIX_OUT pixel_7139/CSA_VREF pixel
Xpixel_6405 pixel_6405/gring pixel_6405/VDD pixel_6405/GND pixel_6405/VREF pixel_6405/ROW_SEL
+ pixel_6405/NB1 pixel_6405/VBIAS pixel_6405/NB2 pixel_6405/AMP_IN pixel_6405/SF_IB
+ pixel_6405/PIX_OUT pixel_6405/CSA_VREF pixel
Xpixel_6416 pixel_6416/gring pixel_6416/VDD pixel_6416/GND pixel_6416/VREF pixel_6416/ROW_SEL
+ pixel_6416/NB1 pixel_6416/VBIAS pixel_6416/NB2 pixel_6416/AMP_IN pixel_6416/SF_IB
+ pixel_6416/PIX_OUT pixel_6416/CSA_VREF pixel
Xpixel_6427 pixel_6427/gring pixel_6427/VDD pixel_6427/GND pixel_6427/VREF pixel_6427/ROW_SEL
+ pixel_6427/NB1 pixel_6427/VBIAS pixel_6427/NB2 pixel_6427/AMP_IN pixel_6427/SF_IB
+ pixel_6427/PIX_OUT pixel_6427/CSA_VREF pixel
Xpixel_6438 pixel_6438/gring pixel_6438/VDD pixel_6438/GND pixel_6438/VREF pixel_6438/ROW_SEL
+ pixel_6438/NB1 pixel_6438/VBIAS pixel_6438/NB2 pixel_6438/AMP_IN pixel_6438/SF_IB
+ pixel_6438/PIX_OUT pixel_6438/CSA_VREF pixel
Xpixel_6449 pixel_6449/gring pixel_6449/VDD pixel_6449/GND pixel_6449/VREF pixel_6449/ROW_SEL
+ pixel_6449/NB1 pixel_6449/VBIAS pixel_6449/NB2 pixel_6449/AMP_IN pixel_6449/SF_IB
+ pixel_6449/PIX_OUT pixel_6449/CSA_VREF pixel
Xpixel_5704 pixel_5704/gring pixel_5704/VDD pixel_5704/GND pixel_5704/VREF pixel_5704/ROW_SEL
+ pixel_5704/NB1 pixel_5704/VBIAS pixel_5704/NB2 pixel_5704/AMP_IN pixel_5704/SF_IB
+ pixel_5704/PIX_OUT pixel_5704/CSA_VREF pixel
Xpixel_5715 pixel_5715/gring pixel_5715/VDD pixel_5715/GND pixel_5715/VREF pixel_5715/ROW_SEL
+ pixel_5715/NB1 pixel_5715/VBIAS pixel_5715/NB2 pixel_5715/AMP_IN pixel_5715/SF_IB
+ pixel_5715/PIX_OUT pixel_5715/CSA_VREF pixel
Xpixel_5726 pixel_5726/gring pixel_5726/VDD pixel_5726/GND pixel_5726/VREF pixel_5726/ROW_SEL
+ pixel_5726/NB1 pixel_5726/VBIAS pixel_5726/NB2 pixel_5726/AMP_IN pixel_5726/SF_IB
+ pixel_5726/PIX_OUT pixel_5726/CSA_VREF pixel
Xpixel_5737 pixel_5737/gring pixel_5737/VDD pixel_5737/GND pixel_5737/VREF pixel_5737/ROW_SEL
+ pixel_5737/NB1 pixel_5737/VBIAS pixel_5737/NB2 pixel_5737/AMP_IN pixel_5737/SF_IB
+ pixel_5737/PIX_OUT pixel_5737/CSA_VREF pixel
Xpixel_5748 pixel_5748/gring pixel_5748/VDD pixel_5748/GND pixel_5748/VREF pixel_5748/ROW_SEL
+ pixel_5748/NB1 pixel_5748/VBIAS pixel_5748/NB2 pixel_5748/AMP_IN pixel_5748/SF_IB
+ pixel_5748/PIX_OUT pixel_5748/CSA_VREF pixel
Xpixel_5759 pixel_5759/gring pixel_5759/VDD pixel_5759/GND pixel_5759/VREF pixel_5759/ROW_SEL
+ pixel_5759/NB1 pixel_5759/VBIAS pixel_5759/NB2 pixel_5759/AMP_IN pixel_5759/SF_IB
+ pixel_5759/PIX_OUT pixel_5759/CSA_VREF pixel
Xpixel_9031 pixel_9031/gring pixel_9031/VDD pixel_9031/GND pixel_9031/VREF pixel_9031/ROW_SEL
+ pixel_9031/NB1 pixel_9031/VBIAS pixel_9031/NB2 pixel_9031/AMP_IN pixel_9031/SF_IB
+ pixel_9031/PIX_OUT pixel_9031/CSA_VREF pixel
Xpixel_9020 pixel_9020/gring pixel_9020/VDD pixel_9020/GND pixel_9020/VREF pixel_9020/ROW_SEL
+ pixel_9020/NB1 pixel_9020/VBIAS pixel_9020/NB2 pixel_9020/AMP_IN pixel_9020/SF_IB
+ pixel_9020/PIX_OUT pixel_9020/CSA_VREF pixel
Xpixel_9064 pixel_9064/gring pixel_9064/VDD pixel_9064/GND pixel_9064/VREF pixel_9064/ROW_SEL
+ pixel_9064/NB1 pixel_9064/VBIAS pixel_9064/NB2 pixel_9064/AMP_IN pixel_9064/SF_IB
+ pixel_9064/PIX_OUT pixel_9064/CSA_VREF pixel
Xpixel_9053 pixel_9053/gring pixel_9053/VDD pixel_9053/GND pixel_9053/VREF pixel_9053/ROW_SEL
+ pixel_9053/NB1 pixel_9053/VBIAS pixel_9053/NB2 pixel_9053/AMP_IN pixel_9053/SF_IB
+ pixel_9053/PIX_OUT pixel_9053/CSA_VREF pixel
Xpixel_9042 pixel_9042/gring pixel_9042/VDD pixel_9042/GND pixel_9042/VREF pixel_9042/ROW_SEL
+ pixel_9042/NB1 pixel_9042/VBIAS pixel_9042/NB2 pixel_9042/AMP_IN pixel_9042/SF_IB
+ pixel_9042/PIX_OUT pixel_9042/CSA_VREF pixel
Xpixel_9097 pixel_9097/gring pixel_9097/VDD pixel_9097/GND pixel_9097/VREF pixel_9097/ROW_SEL
+ pixel_9097/NB1 pixel_9097/VBIAS pixel_9097/NB2 pixel_9097/AMP_IN pixel_9097/SF_IB
+ pixel_9097/PIX_OUT pixel_9097/CSA_VREF pixel
Xpixel_9086 pixel_9086/gring pixel_9086/VDD pixel_9086/GND pixel_9086/VREF pixel_9086/ROW_SEL
+ pixel_9086/NB1 pixel_9086/VBIAS pixel_9086/NB2 pixel_9086/AMP_IN pixel_9086/SF_IB
+ pixel_9086/PIX_OUT pixel_9086/CSA_VREF pixel
Xpixel_9075 pixel_9075/gring pixel_9075/VDD pixel_9075/GND pixel_9075/VREF pixel_9075/ROW_SEL
+ pixel_9075/NB1 pixel_9075/VBIAS pixel_9075/NB2 pixel_9075/AMP_IN pixel_9075/SF_IB
+ pixel_9075/PIX_OUT pixel_9075/CSA_VREF pixel
Xpixel_8330 pixel_8330/gring pixel_8330/VDD pixel_8330/GND pixel_8330/VREF pixel_8330/ROW_SEL
+ pixel_8330/NB1 pixel_8330/VBIAS pixel_8330/NB2 pixel_8330/AMP_IN pixel_8330/SF_IB
+ pixel_8330/PIX_OUT pixel_8330/CSA_VREF pixel
Xpixel_8341 pixel_8341/gring pixel_8341/VDD pixel_8341/GND pixel_8341/VREF pixel_8341/ROW_SEL
+ pixel_8341/NB1 pixel_8341/VBIAS pixel_8341/NB2 pixel_8341/AMP_IN pixel_8341/SF_IB
+ pixel_8341/PIX_OUT pixel_8341/CSA_VREF pixel
Xpixel_8352 pixel_8352/gring pixel_8352/VDD pixel_8352/GND pixel_8352/VREF pixel_8352/ROW_SEL
+ pixel_8352/NB1 pixel_8352/VBIAS pixel_8352/NB2 pixel_8352/AMP_IN pixel_8352/SF_IB
+ pixel_8352/PIX_OUT pixel_8352/CSA_VREF pixel
Xpixel_8363 pixel_8363/gring pixel_8363/VDD pixel_8363/GND pixel_8363/VREF pixel_8363/ROW_SEL
+ pixel_8363/NB1 pixel_8363/VBIAS pixel_8363/NB2 pixel_8363/AMP_IN pixel_8363/SF_IB
+ pixel_8363/PIX_OUT pixel_8363/CSA_VREF pixel
Xpixel_8374 pixel_8374/gring pixel_8374/VDD pixel_8374/GND pixel_8374/VREF pixel_8374/ROW_SEL
+ pixel_8374/NB1 pixel_8374/VBIAS pixel_8374/NB2 pixel_8374/AMP_IN pixel_8374/SF_IB
+ pixel_8374/PIX_OUT pixel_8374/CSA_VREF pixel
Xpixel_8385 pixel_8385/gring pixel_8385/VDD pixel_8385/GND pixel_8385/VREF pixel_8385/ROW_SEL
+ pixel_8385/NB1 pixel_8385/VBIAS pixel_8385/NB2 pixel_8385/AMP_IN pixel_8385/SF_IB
+ pixel_8385/PIX_OUT pixel_8385/CSA_VREF pixel
Xpixel_8396 pixel_8396/gring pixel_8396/VDD pixel_8396/GND pixel_8396/VREF pixel_8396/ROW_SEL
+ pixel_8396/NB1 pixel_8396/VBIAS pixel_8396/NB2 pixel_8396/AMP_IN pixel_8396/SF_IB
+ pixel_8396/PIX_OUT pixel_8396/CSA_VREF pixel
Xpixel_7640 pixel_7640/gring pixel_7640/VDD pixel_7640/GND pixel_7640/VREF pixel_7640/ROW_SEL
+ pixel_7640/NB1 pixel_7640/VBIAS pixel_7640/NB2 pixel_7640/AMP_IN pixel_7640/SF_IB
+ pixel_7640/PIX_OUT pixel_7640/CSA_VREF pixel
Xpixel_7651 pixel_7651/gring pixel_7651/VDD pixel_7651/GND pixel_7651/VREF pixel_7651/ROW_SEL
+ pixel_7651/NB1 pixel_7651/VBIAS pixel_7651/NB2 pixel_7651/AMP_IN pixel_7651/SF_IB
+ pixel_7651/PIX_OUT pixel_7651/CSA_VREF pixel
Xpixel_7662 pixel_7662/gring pixel_7662/VDD pixel_7662/GND pixel_7662/VREF pixel_7662/ROW_SEL
+ pixel_7662/NB1 pixel_7662/VBIAS pixel_7662/NB2 pixel_7662/AMP_IN pixel_7662/SF_IB
+ pixel_7662/PIX_OUT pixel_7662/CSA_VREF pixel
Xpixel_7673 pixel_7673/gring pixel_7673/VDD pixel_7673/GND pixel_7673/VREF pixel_7673/ROW_SEL
+ pixel_7673/NB1 pixel_7673/VBIAS pixel_7673/NB2 pixel_7673/AMP_IN pixel_7673/SF_IB
+ pixel_7673/PIX_OUT pixel_7673/CSA_VREF pixel
Xpixel_7684 pixel_7684/gring pixel_7684/VDD pixel_7684/GND pixel_7684/VREF pixel_7684/ROW_SEL
+ pixel_7684/NB1 pixel_7684/VBIAS pixel_7684/NB2 pixel_7684/AMP_IN pixel_7684/SF_IB
+ pixel_7684/PIX_OUT pixel_7684/CSA_VREF pixel
Xpixel_20 pixel_20/gring pixel_20/VDD pixel_20/GND pixel_20/VREF pixel_20/ROW_SEL
+ pixel_20/NB1 pixel_20/VBIAS pixel_20/NB2 pixel_20/AMP_IN pixel_20/SF_IB pixel_20/PIX_OUT
+ pixel_20/CSA_VREF pixel
Xpixel_7695 pixel_7695/gring pixel_7695/VDD pixel_7695/GND pixel_7695/VREF pixel_7695/ROW_SEL
+ pixel_7695/NB1 pixel_7695/VBIAS pixel_7695/NB2 pixel_7695/AMP_IN pixel_7695/SF_IB
+ pixel_7695/PIX_OUT pixel_7695/CSA_VREF pixel
Xpixel_6950 pixel_6950/gring pixel_6950/VDD pixel_6950/GND pixel_6950/VREF pixel_6950/ROW_SEL
+ pixel_6950/NB1 pixel_6950/VBIAS pixel_6950/NB2 pixel_6950/AMP_IN pixel_6950/SF_IB
+ pixel_6950/PIX_OUT pixel_6950/CSA_VREF pixel
Xpixel_6961 pixel_6961/gring pixel_6961/VDD pixel_6961/GND pixel_6961/VREF pixel_6961/ROW_SEL
+ pixel_6961/NB1 pixel_6961/VBIAS pixel_6961/NB2 pixel_6961/AMP_IN pixel_6961/SF_IB
+ pixel_6961/PIX_OUT pixel_6961/CSA_VREF pixel
Xpixel_6972 pixel_6972/gring pixel_6972/VDD pixel_6972/GND pixel_6972/VREF pixel_6972/ROW_SEL
+ pixel_6972/NB1 pixel_6972/VBIAS pixel_6972/NB2 pixel_6972/AMP_IN pixel_6972/SF_IB
+ pixel_6972/PIX_OUT pixel_6972/CSA_VREF pixel
Xpixel_64 pixel_64/gring pixel_64/VDD pixel_64/GND pixel_64/VREF pixel_64/ROW_SEL
+ pixel_64/NB1 pixel_64/VBIAS pixel_64/NB2 pixel_64/AMP_IN pixel_64/SF_IB pixel_64/PIX_OUT
+ pixel_64/CSA_VREF pixel
Xpixel_53 pixel_53/gring pixel_53/VDD pixel_53/GND pixel_53/VREF pixel_53/ROW_SEL
+ pixel_53/NB1 pixel_53/VBIAS pixel_53/NB2 pixel_53/AMP_IN pixel_53/SF_IB pixel_53/PIX_OUT
+ pixel_53/CSA_VREF pixel
Xpixel_42 pixel_42/gring pixel_42/VDD pixel_42/GND pixel_42/VREF pixel_42/ROW_SEL
+ pixel_42/NB1 pixel_42/VBIAS pixel_42/NB2 pixel_42/AMP_IN pixel_42/SF_IB pixel_42/PIX_OUT
+ pixel_42/CSA_VREF pixel
Xpixel_31 pixel_31/gring pixel_31/VDD pixel_31/GND pixel_31/VREF pixel_31/ROW_SEL
+ pixel_31/NB1 pixel_31/VBIAS pixel_31/NB2 pixel_31/AMP_IN pixel_31/SF_IB pixel_31/PIX_OUT
+ pixel_31/CSA_VREF pixel
Xpixel_6983 pixel_6983/gring pixel_6983/VDD pixel_6983/GND pixel_6983/VREF pixel_6983/ROW_SEL
+ pixel_6983/NB1 pixel_6983/VBIAS pixel_6983/NB2 pixel_6983/AMP_IN pixel_6983/SF_IB
+ pixel_6983/PIX_OUT pixel_6983/CSA_VREF pixel
Xpixel_6994 pixel_6994/gring pixel_6994/VDD pixel_6994/GND pixel_6994/VREF pixel_6994/ROW_SEL
+ pixel_6994/NB1 pixel_6994/VBIAS pixel_6994/NB2 pixel_6994/AMP_IN pixel_6994/SF_IB
+ pixel_6994/PIX_OUT pixel_6994/CSA_VREF pixel
Xpixel_97 pixel_97/gring pixel_97/VDD pixel_97/GND pixel_97/VREF pixel_97/ROW_SEL
+ pixel_97/NB1 pixel_97/VBIAS pixel_97/NB2 pixel_97/AMP_IN pixel_97/SF_IB pixel_97/PIX_OUT
+ pixel_97/CSA_VREF pixel
Xpixel_86 pixel_86/gring pixel_86/VDD pixel_86/GND pixel_86/VREF pixel_86/ROW_SEL
+ pixel_86/NB1 pixel_86/VBIAS pixel_86/NB2 pixel_86/AMP_IN pixel_86/SF_IB pixel_86/PIX_OUT
+ pixel_86/CSA_VREF pixel
Xpixel_75 pixel_75/gring pixel_75/VDD pixel_75/GND pixel_75/VREF pixel_75/ROW_SEL
+ pixel_75/NB1 pixel_75/VBIAS pixel_75/NB2 pixel_75/AMP_IN pixel_75/SF_IB pixel_75/PIX_OUT
+ pixel_75/CSA_VREF pixel
Xpixel_1290 pixel_1290/gring pixel_1290/VDD pixel_1290/GND pixel_1290/VREF pixel_1290/ROW_SEL
+ pixel_1290/NB1 pixel_1290/VBIAS pixel_1290/NB2 pixel_1290/AMP_IN pixel_1290/SF_IB
+ pixel_1290/PIX_OUT pixel_1290/CSA_VREF pixel
Xpixel_338 pixel_338/gring pixel_338/VDD pixel_338/GND pixel_338/VREF pixel_338/ROW_SEL
+ pixel_338/NB1 pixel_338/VBIAS pixel_338/NB2 pixel_338/AMP_IN pixel_338/SF_IB pixel_338/PIX_OUT
+ pixel_338/CSA_VREF pixel
Xpixel_327 pixel_327/gring pixel_327/VDD pixel_327/GND pixel_327/VREF pixel_327/ROW_SEL
+ pixel_327/NB1 pixel_327/VBIAS pixel_327/NB2 pixel_327/AMP_IN pixel_327/SF_IB pixel_327/PIX_OUT
+ pixel_327/CSA_VREF pixel
Xpixel_316 pixel_316/gring pixel_316/VDD pixel_316/GND pixel_316/VREF pixel_316/ROW_SEL
+ pixel_316/NB1 pixel_316/VBIAS pixel_316/NB2 pixel_316/AMP_IN pixel_316/SF_IB pixel_316/PIX_OUT
+ pixel_316/CSA_VREF pixel
Xpixel_305 pixel_305/gring pixel_305/VDD pixel_305/GND pixel_305/VREF pixel_305/ROW_SEL
+ pixel_305/NB1 pixel_305/VBIAS pixel_305/NB2 pixel_305/AMP_IN pixel_305/SF_IB pixel_305/PIX_OUT
+ pixel_305/CSA_VREF pixel
Xpixel_349 pixel_349/gring pixel_349/VDD pixel_349/GND pixel_349/VREF pixel_349/ROW_SEL
+ pixel_349/NB1 pixel_349/VBIAS pixel_349/NB2 pixel_349/AMP_IN pixel_349/SF_IB pixel_349/PIX_OUT
+ pixel_349/CSA_VREF pixel
Xpixel_3609 pixel_3609/gring pixel_3609/VDD pixel_3609/GND pixel_3609/VREF pixel_3609/ROW_SEL
+ pixel_3609/NB1 pixel_3609/VBIAS pixel_3609/NB2 pixel_3609/AMP_IN pixel_3609/SF_IB
+ pixel_3609/PIX_OUT pixel_3609/CSA_VREF pixel
Xpixel_2919 pixel_2919/gring pixel_2919/VDD pixel_2919/GND pixel_2919/VREF pixel_2919/ROW_SEL
+ pixel_2919/NB1 pixel_2919/VBIAS pixel_2919/NB2 pixel_2919/AMP_IN pixel_2919/SF_IB
+ pixel_2919/PIX_OUT pixel_2919/CSA_VREF pixel
Xpixel_2908 pixel_2908/gring pixel_2908/VDD pixel_2908/GND pixel_2908/VREF pixel_2908/ROW_SEL
+ pixel_2908/NB1 pixel_2908/VBIAS pixel_2908/NB2 pixel_2908/AMP_IN pixel_2908/SF_IB
+ pixel_2908/PIX_OUT pixel_2908/CSA_VREF pixel
Xpixel_6202 pixel_6202/gring pixel_6202/VDD pixel_6202/GND pixel_6202/VREF pixel_6202/ROW_SEL
+ pixel_6202/NB1 pixel_6202/VBIAS pixel_6202/NB2 pixel_6202/AMP_IN pixel_6202/SF_IB
+ pixel_6202/PIX_OUT pixel_6202/CSA_VREF pixel
Xpixel_6213 pixel_6213/gring pixel_6213/VDD pixel_6213/GND pixel_6213/VREF pixel_6213/ROW_SEL
+ pixel_6213/NB1 pixel_6213/VBIAS pixel_6213/NB2 pixel_6213/AMP_IN pixel_6213/SF_IB
+ pixel_6213/PIX_OUT pixel_6213/CSA_VREF pixel
Xpixel_6224 pixel_6224/gring pixel_6224/VDD pixel_6224/GND pixel_6224/VREF pixel_6224/ROW_SEL
+ pixel_6224/NB1 pixel_6224/VBIAS pixel_6224/NB2 pixel_6224/AMP_IN pixel_6224/SF_IB
+ pixel_6224/PIX_OUT pixel_6224/CSA_VREF pixel
Xpixel_6235 pixel_6235/gring pixel_6235/VDD pixel_6235/GND pixel_6235/VREF pixel_6235/ROW_SEL
+ pixel_6235/NB1 pixel_6235/VBIAS pixel_6235/NB2 pixel_6235/AMP_IN pixel_6235/SF_IB
+ pixel_6235/PIX_OUT pixel_6235/CSA_VREF pixel
Xpixel_6246 pixel_6246/gring pixel_6246/VDD pixel_6246/GND pixel_6246/VREF pixel_6246/ROW_SEL
+ pixel_6246/NB1 pixel_6246/VBIAS pixel_6246/NB2 pixel_6246/AMP_IN pixel_6246/SF_IB
+ pixel_6246/PIX_OUT pixel_6246/CSA_VREF pixel
Xpixel_6257 pixel_6257/gring pixel_6257/VDD pixel_6257/GND pixel_6257/VREF pixel_6257/ROW_SEL
+ pixel_6257/NB1 pixel_6257/VBIAS pixel_6257/NB2 pixel_6257/AMP_IN pixel_6257/SF_IB
+ pixel_6257/PIX_OUT pixel_6257/CSA_VREF pixel
Xpixel_6268 pixel_6268/gring pixel_6268/VDD pixel_6268/GND pixel_6268/VREF pixel_6268/ROW_SEL
+ pixel_6268/NB1 pixel_6268/VBIAS pixel_6268/NB2 pixel_6268/AMP_IN pixel_6268/SF_IB
+ pixel_6268/PIX_OUT pixel_6268/CSA_VREF pixel
Xpixel_5501 pixel_5501/gring pixel_5501/VDD pixel_5501/GND pixel_5501/VREF pixel_5501/ROW_SEL
+ pixel_5501/NB1 pixel_5501/VBIAS pixel_5501/NB2 pixel_5501/AMP_IN pixel_5501/SF_IB
+ pixel_5501/PIX_OUT pixel_5501/CSA_VREF pixel
Xpixel_5512 pixel_5512/gring pixel_5512/VDD pixel_5512/GND pixel_5512/VREF pixel_5512/ROW_SEL
+ pixel_5512/NB1 pixel_5512/VBIAS pixel_5512/NB2 pixel_5512/AMP_IN pixel_5512/SF_IB
+ pixel_5512/PIX_OUT pixel_5512/CSA_VREF pixel
Xpixel_5523 pixel_5523/gring pixel_5523/VDD pixel_5523/GND pixel_5523/VREF pixel_5523/ROW_SEL
+ pixel_5523/NB1 pixel_5523/VBIAS pixel_5523/NB2 pixel_5523/AMP_IN pixel_5523/SF_IB
+ pixel_5523/PIX_OUT pixel_5523/CSA_VREF pixel
Xpixel_6279 pixel_6279/gring pixel_6279/VDD pixel_6279/GND pixel_6279/VREF pixel_6279/ROW_SEL
+ pixel_6279/NB1 pixel_6279/VBIAS pixel_6279/NB2 pixel_6279/AMP_IN pixel_6279/SF_IB
+ pixel_6279/PIX_OUT pixel_6279/CSA_VREF pixel
Xpixel_5534 pixel_5534/gring pixel_5534/VDD pixel_5534/GND pixel_5534/VREF pixel_5534/ROW_SEL
+ pixel_5534/NB1 pixel_5534/VBIAS pixel_5534/NB2 pixel_5534/AMP_IN pixel_5534/SF_IB
+ pixel_5534/PIX_OUT pixel_5534/CSA_VREF pixel
Xpixel_5545 pixel_5545/gring pixel_5545/VDD pixel_5545/GND pixel_5545/VREF pixel_5545/ROW_SEL
+ pixel_5545/NB1 pixel_5545/VBIAS pixel_5545/NB2 pixel_5545/AMP_IN pixel_5545/SF_IB
+ pixel_5545/PIX_OUT pixel_5545/CSA_VREF pixel
Xpixel_5556 pixel_5556/gring pixel_5556/VDD pixel_5556/GND pixel_5556/VREF pixel_5556/ROW_SEL
+ pixel_5556/NB1 pixel_5556/VBIAS pixel_5556/NB2 pixel_5556/AMP_IN pixel_5556/SF_IB
+ pixel_5556/PIX_OUT pixel_5556/CSA_VREF pixel
Xpixel_5567 pixel_5567/gring pixel_5567/VDD pixel_5567/GND pixel_5567/VREF pixel_5567/ROW_SEL
+ pixel_5567/NB1 pixel_5567/VBIAS pixel_5567/NB2 pixel_5567/AMP_IN pixel_5567/SF_IB
+ pixel_5567/PIX_OUT pixel_5567/CSA_VREF pixel
Xpixel_4800 pixel_4800/gring pixel_4800/VDD pixel_4800/GND pixel_4800/VREF pixel_4800/ROW_SEL
+ pixel_4800/NB1 pixel_4800/VBIAS pixel_4800/NB2 pixel_4800/AMP_IN pixel_4800/SF_IB
+ pixel_4800/PIX_OUT pixel_4800/CSA_VREF pixel
Xpixel_4811 pixel_4811/gring pixel_4811/VDD pixel_4811/GND pixel_4811/VREF pixel_4811/ROW_SEL
+ pixel_4811/NB1 pixel_4811/VBIAS pixel_4811/NB2 pixel_4811/AMP_IN pixel_4811/SF_IB
+ pixel_4811/PIX_OUT pixel_4811/CSA_VREF pixel
Xpixel_4822 pixel_4822/gring pixel_4822/VDD pixel_4822/GND pixel_4822/VREF pixel_4822/ROW_SEL
+ pixel_4822/NB1 pixel_4822/VBIAS pixel_4822/NB2 pixel_4822/AMP_IN pixel_4822/SF_IB
+ pixel_4822/PIX_OUT pixel_4822/CSA_VREF pixel
Xpixel_850 pixel_850/gring pixel_850/VDD pixel_850/GND pixel_850/VREF pixel_850/ROW_SEL
+ pixel_850/NB1 pixel_850/VBIAS pixel_850/NB2 pixel_850/AMP_IN pixel_850/SF_IB pixel_850/PIX_OUT
+ pixel_850/CSA_VREF pixel
Xpixel_5578 pixel_5578/gring pixel_5578/VDD pixel_5578/GND pixel_5578/VREF pixel_5578/ROW_SEL
+ pixel_5578/NB1 pixel_5578/VBIAS pixel_5578/NB2 pixel_5578/AMP_IN pixel_5578/SF_IB
+ pixel_5578/PIX_OUT pixel_5578/CSA_VREF pixel
Xpixel_5589 pixel_5589/gring pixel_5589/VDD pixel_5589/GND pixel_5589/VREF pixel_5589/ROW_SEL
+ pixel_5589/NB1 pixel_5589/VBIAS pixel_5589/NB2 pixel_5589/AMP_IN pixel_5589/SF_IB
+ pixel_5589/PIX_OUT pixel_5589/CSA_VREF pixel
Xpixel_4833 pixel_4833/gring pixel_4833/VDD pixel_4833/GND pixel_4833/VREF pixel_4833/ROW_SEL
+ pixel_4833/NB1 pixel_4833/VBIAS pixel_4833/NB2 pixel_4833/AMP_IN pixel_4833/SF_IB
+ pixel_4833/PIX_OUT pixel_4833/CSA_VREF pixel
Xpixel_4844 pixel_4844/gring pixel_4844/VDD pixel_4844/GND pixel_4844/VREF pixel_4844/ROW_SEL
+ pixel_4844/NB1 pixel_4844/VBIAS pixel_4844/NB2 pixel_4844/AMP_IN pixel_4844/SF_IB
+ pixel_4844/PIX_OUT pixel_4844/CSA_VREF pixel
Xpixel_4855 pixel_4855/gring pixel_4855/VDD pixel_4855/GND pixel_4855/VREF pixel_4855/ROW_SEL
+ pixel_4855/NB1 pixel_4855/VBIAS pixel_4855/NB2 pixel_4855/AMP_IN pixel_4855/SF_IB
+ pixel_4855/PIX_OUT pixel_4855/CSA_VREF pixel
Xpixel_894 pixel_894/gring pixel_894/VDD pixel_894/GND pixel_894/VREF pixel_894/ROW_SEL
+ pixel_894/NB1 pixel_894/VBIAS pixel_894/NB2 pixel_894/AMP_IN pixel_894/SF_IB pixel_894/PIX_OUT
+ pixel_894/CSA_VREF pixel
Xpixel_883 pixel_883/gring pixel_883/VDD pixel_883/GND pixel_883/VREF pixel_883/ROW_SEL
+ pixel_883/NB1 pixel_883/VBIAS pixel_883/NB2 pixel_883/AMP_IN pixel_883/SF_IB pixel_883/PIX_OUT
+ pixel_883/CSA_VREF pixel
Xpixel_872 pixel_872/gring pixel_872/VDD pixel_872/GND pixel_872/VREF pixel_872/ROW_SEL
+ pixel_872/NB1 pixel_872/VBIAS pixel_872/NB2 pixel_872/AMP_IN pixel_872/SF_IB pixel_872/PIX_OUT
+ pixel_872/CSA_VREF pixel
Xpixel_861 pixel_861/gring pixel_861/VDD pixel_861/GND pixel_861/VREF pixel_861/ROW_SEL
+ pixel_861/NB1 pixel_861/VBIAS pixel_861/NB2 pixel_861/AMP_IN pixel_861/SF_IB pixel_861/PIX_OUT
+ pixel_861/CSA_VREF pixel
Xpixel_4866 pixel_4866/gring pixel_4866/VDD pixel_4866/GND pixel_4866/VREF pixel_4866/ROW_SEL
+ pixel_4866/NB1 pixel_4866/VBIAS pixel_4866/NB2 pixel_4866/AMP_IN pixel_4866/SF_IB
+ pixel_4866/PIX_OUT pixel_4866/CSA_VREF pixel
Xpixel_4877 pixel_4877/gring pixel_4877/VDD pixel_4877/GND pixel_4877/VREF pixel_4877/ROW_SEL
+ pixel_4877/NB1 pixel_4877/VBIAS pixel_4877/NB2 pixel_4877/AMP_IN pixel_4877/SF_IB
+ pixel_4877/PIX_OUT pixel_4877/CSA_VREF pixel
Xpixel_4888 pixel_4888/gring pixel_4888/VDD pixel_4888/GND pixel_4888/VREF pixel_4888/ROW_SEL
+ pixel_4888/NB1 pixel_4888/VBIAS pixel_4888/NB2 pixel_4888/AMP_IN pixel_4888/SF_IB
+ pixel_4888/PIX_OUT pixel_4888/CSA_VREF pixel
Xpixel_4899 pixel_4899/gring pixel_4899/VDD pixel_4899/GND pixel_4899/VREF pixel_4899/ROW_SEL
+ pixel_4899/NB1 pixel_4899/VBIAS pixel_4899/NB2 pixel_4899/AMP_IN pixel_4899/SF_IB
+ pixel_4899/PIX_OUT pixel_4899/CSA_VREF pixel
Xpixel_8160 pixel_8160/gring pixel_8160/VDD pixel_8160/GND pixel_8160/VREF pixel_8160/ROW_SEL
+ pixel_8160/NB1 pixel_8160/VBIAS pixel_8160/NB2 pixel_8160/AMP_IN pixel_8160/SF_IB
+ pixel_8160/PIX_OUT pixel_8160/CSA_VREF pixel
Xpixel_8171 pixel_8171/gring pixel_8171/VDD pixel_8171/GND pixel_8171/VREF pixel_8171/ROW_SEL
+ pixel_8171/NB1 pixel_8171/VBIAS pixel_8171/NB2 pixel_8171/AMP_IN pixel_8171/SF_IB
+ pixel_8171/PIX_OUT pixel_8171/CSA_VREF pixel
Xpixel_8182 pixel_8182/gring pixel_8182/VDD pixel_8182/GND pixel_8182/VREF pixel_8182/ROW_SEL
+ pixel_8182/NB1 pixel_8182/VBIAS pixel_8182/NB2 pixel_8182/AMP_IN pixel_8182/SF_IB
+ pixel_8182/PIX_OUT pixel_8182/CSA_VREF pixel
Xpixel_8193 pixel_8193/gring pixel_8193/VDD pixel_8193/GND pixel_8193/VREF pixel_8193/ROW_SEL
+ pixel_8193/NB1 pixel_8193/VBIAS pixel_8193/NB2 pixel_8193/AMP_IN pixel_8193/SF_IB
+ pixel_8193/PIX_OUT pixel_8193/CSA_VREF pixel
Xpixel_7470 pixel_7470/gring pixel_7470/VDD pixel_7470/GND pixel_7470/VREF pixel_7470/ROW_SEL
+ pixel_7470/NB1 pixel_7470/VBIAS pixel_7470/NB2 pixel_7470/AMP_IN pixel_7470/SF_IB
+ pixel_7470/PIX_OUT pixel_7470/CSA_VREF pixel
Xpixel_7481 pixel_7481/gring pixel_7481/VDD pixel_7481/GND pixel_7481/VREF pixel_7481/ROW_SEL
+ pixel_7481/NB1 pixel_7481/VBIAS pixel_7481/NB2 pixel_7481/AMP_IN pixel_7481/SF_IB
+ pixel_7481/PIX_OUT pixel_7481/CSA_VREF pixel
Xpixel_7492 pixel_7492/gring pixel_7492/VDD pixel_7492/GND pixel_7492/VREF pixel_7492/ROW_SEL
+ pixel_7492/NB1 pixel_7492/VBIAS pixel_7492/NB2 pixel_7492/AMP_IN pixel_7492/SF_IB
+ pixel_7492/PIX_OUT pixel_7492/CSA_VREF pixel
Xpixel_6780 pixel_6780/gring pixel_6780/VDD pixel_6780/GND pixel_6780/VREF pixel_6780/ROW_SEL
+ pixel_6780/NB1 pixel_6780/VBIAS pixel_6780/NB2 pixel_6780/AMP_IN pixel_6780/SF_IB
+ pixel_6780/PIX_OUT pixel_6780/CSA_VREF pixel
Xpixel_6791 pixel_6791/gring pixel_6791/VDD pixel_6791/GND pixel_6791/VREF pixel_6791/ROW_SEL
+ pixel_6791/NB1 pixel_6791/VBIAS pixel_6791/NB2 pixel_6791/AMP_IN pixel_6791/SF_IB
+ pixel_6791/PIX_OUT pixel_6791/CSA_VREF pixel
Xpixel_113 pixel_113/gring pixel_113/VDD pixel_113/GND pixel_113/VREF pixel_113/ROW_SEL
+ pixel_113/NB1 pixel_113/VBIAS pixel_113/NB2 pixel_113/AMP_IN pixel_113/SF_IB pixel_113/PIX_OUT
+ pixel_113/CSA_VREF pixel
Xpixel_102 pixel_102/gring pixel_102/VDD pixel_102/GND pixel_102/VREF pixel_102/ROW_SEL
+ pixel_102/NB1 pixel_102/VBIAS pixel_102/NB2 pixel_102/AMP_IN pixel_102/SF_IB pixel_102/PIX_OUT
+ pixel_102/CSA_VREF pixel
Xpixel_4107 pixel_4107/gring pixel_4107/VDD pixel_4107/GND pixel_4107/VREF pixel_4107/ROW_SEL
+ pixel_4107/NB1 pixel_4107/VBIAS pixel_4107/NB2 pixel_4107/AMP_IN pixel_4107/SF_IB
+ pixel_4107/PIX_OUT pixel_4107/CSA_VREF pixel
Xpixel_146 pixel_146/gring pixel_146/VDD pixel_146/GND pixel_146/VREF pixel_146/ROW_SEL
+ pixel_146/NB1 pixel_146/VBIAS pixel_146/NB2 pixel_146/AMP_IN pixel_146/SF_IB pixel_146/PIX_OUT
+ pixel_146/CSA_VREF pixel
Xpixel_135 pixel_135/gring pixel_135/VDD pixel_135/GND pixel_135/VREF pixel_135/ROW_SEL
+ pixel_135/NB1 pixel_135/VBIAS pixel_135/NB2 pixel_135/AMP_IN pixel_135/SF_IB pixel_135/PIX_OUT
+ pixel_135/CSA_VREF pixel
Xpixel_124 pixel_124/gring pixel_124/VDD pixel_124/GND pixel_124/VREF pixel_124/ROW_SEL
+ pixel_124/NB1 pixel_124/VBIAS pixel_124/NB2 pixel_124/AMP_IN pixel_124/SF_IB pixel_124/PIX_OUT
+ pixel_124/CSA_VREF pixel
Xpixel_3406 pixel_3406/gring pixel_3406/VDD pixel_3406/GND pixel_3406/VREF pixel_3406/ROW_SEL
+ pixel_3406/NB1 pixel_3406/VBIAS pixel_3406/NB2 pixel_3406/AMP_IN pixel_3406/SF_IB
+ pixel_3406/PIX_OUT pixel_3406/CSA_VREF pixel
Xpixel_4118 pixel_4118/gring pixel_4118/VDD pixel_4118/GND pixel_4118/VREF pixel_4118/ROW_SEL
+ pixel_4118/NB1 pixel_4118/VBIAS pixel_4118/NB2 pixel_4118/AMP_IN pixel_4118/SF_IB
+ pixel_4118/PIX_OUT pixel_4118/CSA_VREF pixel
Xpixel_4129 pixel_4129/gring pixel_4129/VDD pixel_4129/GND pixel_4129/VREF pixel_4129/ROW_SEL
+ pixel_4129/NB1 pixel_4129/VBIAS pixel_4129/NB2 pixel_4129/AMP_IN pixel_4129/SF_IB
+ pixel_4129/PIX_OUT pixel_4129/CSA_VREF pixel
Xpixel_179 pixel_179/gring pixel_179/VDD pixel_179/GND pixel_179/VREF pixel_179/ROW_SEL
+ pixel_179/NB1 pixel_179/VBIAS pixel_179/NB2 pixel_179/AMP_IN pixel_179/SF_IB pixel_179/PIX_OUT
+ pixel_179/CSA_VREF pixel
Xpixel_168 pixel_168/gring pixel_168/VDD pixel_168/GND pixel_168/VREF pixel_168/ROW_SEL
+ pixel_168/NB1 pixel_168/VBIAS pixel_168/NB2 pixel_168/AMP_IN pixel_168/SF_IB pixel_168/PIX_OUT
+ pixel_168/CSA_VREF pixel
Xpixel_157 pixel_157/gring pixel_157/VDD pixel_157/GND pixel_157/VREF pixel_157/ROW_SEL
+ pixel_157/NB1 pixel_157/VBIAS pixel_157/NB2 pixel_157/AMP_IN pixel_157/SF_IB pixel_157/PIX_OUT
+ pixel_157/CSA_VREF pixel
Xpixel_3439 pixel_3439/gring pixel_3439/VDD pixel_3439/GND pixel_3439/VREF pixel_3439/ROW_SEL
+ pixel_3439/NB1 pixel_3439/VBIAS pixel_3439/NB2 pixel_3439/AMP_IN pixel_3439/SF_IB
+ pixel_3439/PIX_OUT pixel_3439/CSA_VREF pixel
Xpixel_3428 pixel_3428/gring pixel_3428/VDD pixel_3428/GND pixel_3428/VREF pixel_3428/ROW_SEL
+ pixel_3428/NB1 pixel_3428/VBIAS pixel_3428/NB2 pixel_3428/AMP_IN pixel_3428/SF_IB
+ pixel_3428/PIX_OUT pixel_3428/CSA_VREF pixel
Xpixel_3417 pixel_3417/gring pixel_3417/VDD pixel_3417/GND pixel_3417/VREF pixel_3417/ROW_SEL
+ pixel_3417/NB1 pixel_3417/VBIAS pixel_3417/NB2 pixel_3417/AMP_IN pixel_3417/SF_IB
+ pixel_3417/PIX_OUT pixel_3417/CSA_VREF pixel
Xpixel_2738 pixel_2738/gring pixel_2738/VDD pixel_2738/GND pixel_2738/VREF pixel_2738/ROW_SEL
+ pixel_2738/NB1 pixel_2738/VBIAS pixel_2738/NB2 pixel_2738/AMP_IN pixel_2738/SF_IB
+ pixel_2738/PIX_OUT pixel_2738/CSA_VREF pixel
Xpixel_2727 pixel_2727/gring pixel_2727/VDD pixel_2727/GND pixel_2727/VREF pixel_2727/ROW_SEL
+ pixel_2727/NB1 pixel_2727/VBIAS pixel_2727/NB2 pixel_2727/AMP_IN pixel_2727/SF_IB
+ pixel_2727/PIX_OUT pixel_2727/CSA_VREF pixel
Xpixel_2716 pixel_2716/gring pixel_2716/VDD pixel_2716/GND pixel_2716/VREF pixel_2716/ROW_SEL
+ pixel_2716/NB1 pixel_2716/VBIAS pixel_2716/NB2 pixel_2716/AMP_IN pixel_2716/SF_IB
+ pixel_2716/PIX_OUT pixel_2716/CSA_VREF pixel
Xpixel_2705 pixel_2705/gring pixel_2705/VDD pixel_2705/GND pixel_2705/VREF pixel_2705/ROW_SEL
+ pixel_2705/NB1 pixel_2705/VBIAS pixel_2705/NB2 pixel_2705/AMP_IN pixel_2705/SF_IB
+ pixel_2705/PIX_OUT pixel_2705/CSA_VREF pixel
Xpixel_2749 pixel_2749/gring pixel_2749/VDD pixel_2749/GND pixel_2749/VREF pixel_2749/ROW_SEL
+ pixel_2749/NB1 pixel_2749/VBIAS pixel_2749/NB2 pixel_2749/AMP_IN pixel_2749/SF_IB
+ pixel_2749/PIX_OUT pixel_2749/CSA_VREF pixel
Xpixel_6010 pixel_6010/gring pixel_6010/VDD pixel_6010/GND pixel_6010/VREF pixel_6010/ROW_SEL
+ pixel_6010/NB1 pixel_6010/VBIAS pixel_6010/NB2 pixel_6010/AMP_IN pixel_6010/SF_IB
+ pixel_6010/PIX_OUT pixel_6010/CSA_VREF pixel
Xpixel_6021 pixel_6021/gring pixel_6021/VDD pixel_6021/GND pixel_6021/VREF pixel_6021/ROW_SEL
+ pixel_6021/NB1 pixel_6021/VBIAS pixel_6021/NB2 pixel_6021/AMP_IN pixel_6021/SF_IB
+ pixel_6021/PIX_OUT pixel_6021/CSA_VREF pixel
Xpixel_6032 pixel_6032/gring pixel_6032/VDD pixel_6032/GND pixel_6032/VREF pixel_6032/ROW_SEL
+ pixel_6032/NB1 pixel_6032/VBIAS pixel_6032/NB2 pixel_6032/AMP_IN pixel_6032/SF_IB
+ pixel_6032/PIX_OUT pixel_6032/CSA_VREF pixel
Xpixel_6043 pixel_6043/gring pixel_6043/VDD pixel_6043/GND pixel_6043/VREF pixel_6043/ROW_SEL
+ pixel_6043/NB1 pixel_6043/VBIAS pixel_6043/NB2 pixel_6043/AMP_IN pixel_6043/SF_IB
+ pixel_6043/PIX_OUT pixel_6043/CSA_VREF pixel
Xpixel_6054 pixel_6054/gring pixel_6054/VDD pixel_6054/GND pixel_6054/VREF pixel_6054/ROW_SEL
+ pixel_6054/NB1 pixel_6054/VBIAS pixel_6054/NB2 pixel_6054/AMP_IN pixel_6054/SF_IB
+ pixel_6054/PIX_OUT pixel_6054/CSA_VREF pixel
Xpixel_6065 pixel_6065/gring pixel_6065/VDD pixel_6065/GND pixel_6065/VREF pixel_6065/ROW_SEL
+ pixel_6065/NB1 pixel_6065/VBIAS pixel_6065/NB2 pixel_6065/AMP_IN pixel_6065/SF_IB
+ pixel_6065/PIX_OUT pixel_6065/CSA_VREF pixel
Xpixel_6076 pixel_6076/gring pixel_6076/VDD pixel_6076/GND pixel_6076/VREF pixel_6076/ROW_SEL
+ pixel_6076/NB1 pixel_6076/VBIAS pixel_6076/NB2 pixel_6076/AMP_IN pixel_6076/SF_IB
+ pixel_6076/PIX_OUT pixel_6076/CSA_VREF pixel
Xpixel_5320 pixel_5320/gring pixel_5320/VDD pixel_5320/GND pixel_5320/VREF pixel_5320/ROW_SEL
+ pixel_5320/NB1 pixel_5320/VBIAS pixel_5320/NB2 pixel_5320/AMP_IN pixel_5320/SF_IB
+ pixel_5320/PIX_OUT pixel_5320/CSA_VREF pixel
Xpixel_5331 pixel_5331/gring pixel_5331/VDD pixel_5331/GND pixel_5331/VREF pixel_5331/ROW_SEL
+ pixel_5331/NB1 pixel_5331/VBIAS pixel_5331/NB2 pixel_5331/AMP_IN pixel_5331/SF_IB
+ pixel_5331/PIX_OUT pixel_5331/CSA_VREF pixel
Xpixel_6087 pixel_6087/gring pixel_6087/VDD pixel_6087/GND pixel_6087/VREF pixel_6087/ROW_SEL
+ pixel_6087/NB1 pixel_6087/VBIAS pixel_6087/NB2 pixel_6087/AMP_IN pixel_6087/SF_IB
+ pixel_6087/PIX_OUT pixel_6087/CSA_VREF pixel
Xpixel_6098 pixel_6098/gring pixel_6098/VDD pixel_6098/GND pixel_6098/VREF pixel_6098/ROW_SEL
+ pixel_6098/NB1 pixel_6098/VBIAS pixel_6098/NB2 pixel_6098/AMP_IN pixel_6098/SF_IB
+ pixel_6098/PIX_OUT pixel_6098/CSA_VREF pixel
Xpixel_5342 pixel_5342/gring pixel_5342/VDD pixel_5342/GND pixel_5342/VREF pixel_5342/ROW_SEL
+ pixel_5342/NB1 pixel_5342/VBIAS pixel_5342/NB2 pixel_5342/AMP_IN pixel_5342/SF_IB
+ pixel_5342/PIX_OUT pixel_5342/CSA_VREF pixel
Xpixel_5353 pixel_5353/gring pixel_5353/VDD pixel_5353/GND pixel_5353/VREF pixel_5353/ROW_SEL
+ pixel_5353/NB1 pixel_5353/VBIAS pixel_5353/NB2 pixel_5353/AMP_IN pixel_5353/SF_IB
+ pixel_5353/PIX_OUT pixel_5353/CSA_VREF pixel
Xpixel_5364 pixel_5364/gring pixel_5364/VDD pixel_5364/GND pixel_5364/VREF pixel_5364/ROW_SEL
+ pixel_5364/NB1 pixel_5364/VBIAS pixel_5364/NB2 pixel_5364/AMP_IN pixel_5364/SF_IB
+ pixel_5364/PIX_OUT pixel_5364/CSA_VREF pixel
Xpixel_5375 pixel_5375/gring pixel_5375/VDD pixel_5375/GND pixel_5375/VREF pixel_5375/ROW_SEL
+ pixel_5375/NB1 pixel_5375/VBIAS pixel_5375/NB2 pixel_5375/AMP_IN pixel_5375/SF_IB
+ pixel_5375/PIX_OUT pixel_5375/CSA_VREF pixel
Xpixel_4630 pixel_4630/gring pixel_4630/VDD pixel_4630/GND pixel_4630/VREF pixel_4630/ROW_SEL
+ pixel_4630/NB1 pixel_4630/VBIAS pixel_4630/NB2 pixel_4630/AMP_IN pixel_4630/SF_IB
+ pixel_4630/PIX_OUT pixel_4630/CSA_VREF pixel
Xpixel_5386 pixel_5386/gring pixel_5386/VDD pixel_5386/GND pixel_5386/VREF pixel_5386/ROW_SEL
+ pixel_5386/NB1 pixel_5386/VBIAS pixel_5386/NB2 pixel_5386/AMP_IN pixel_5386/SF_IB
+ pixel_5386/PIX_OUT pixel_5386/CSA_VREF pixel
Xpixel_5397 pixel_5397/gring pixel_5397/VDD pixel_5397/GND pixel_5397/VREF pixel_5397/ROW_SEL
+ pixel_5397/NB1 pixel_5397/VBIAS pixel_5397/NB2 pixel_5397/AMP_IN pixel_5397/SF_IB
+ pixel_5397/PIX_OUT pixel_5397/CSA_VREF pixel
Xpixel_4641 pixel_4641/gring pixel_4641/VDD pixel_4641/GND pixel_4641/VREF pixel_4641/ROW_SEL
+ pixel_4641/NB1 pixel_4641/VBIAS pixel_4641/NB2 pixel_4641/AMP_IN pixel_4641/SF_IB
+ pixel_4641/PIX_OUT pixel_4641/CSA_VREF pixel
Xpixel_4652 pixel_4652/gring pixel_4652/VDD pixel_4652/GND pixel_4652/VREF pixel_4652/ROW_SEL
+ pixel_4652/NB1 pixel_4652/VBIAS pixel_4652/NB2 pixel_4652/AMP_IN pixel_4652/SF_IB
+ pixel_4652/PIX_OUT pixel_4652/CSA_VREF pixel
Xpixel_4663 pixel_4663/gring pixel_4663/VDD pixel_4663/GND pixel_4663/VREF pixel_4663/ROW_SEL
+ pixel_4663/NB1 pixel_4663/VBIAS pixel_4663/NB2 pixel_4663/AMP_IN pixel_4663/SF_IB
+ pixel_4663/PIX_OUT pixel_4663/CSA_VREF pixel
Xpixel_691 pixel_691/gring pixel_691/VDD pixel_691/GND pixel_691/VREF pixel_691/ROW_SEL
+ pixel_691/NB1 pixel_691/VBIAS pixel_691/NB2 pixel_691/AMP_IN pixel_691/SF_IB pixel_691/PIX_OUT
+ pixel_691/CSA_VREF pixel
Xpixel_680 pixel_680/gring pixel_680/VDD pixel_680/GND pixel_680/VREF pixel_680/ROW_SEL
+ pixel_680/NB1 pixel_680/VBIAS pixel_680/NB2 pixel_680/AMP_IN pixel_680/SF_IB pixel_680/PIX_OUT
+ pixel_680/CSA_VREF pixel
Xpixel_4674 pixel_4674/gring pixel_4674/VDD pixel_4674/GND pixel_4674/VREF pixel_4674/ROW_SEL
+ pixel_4674/NB1 pixel_4674/VBIAS pixel_4674/NB2 pixel_4674/AMP_IN pixel_4674/SF_IB
+ pixel_4674/PIX_OUT pixel_4674/CSA_VREF pixel
Xpixel_4685 pixel_4685/gring pixel_4685/VDD pixel_4685/GND pixel_4685/VREF pixel_4685/ROW_SEL
+ pixel_4685/NB1 pixel_4685/VBIAS pixel_4685/NB2 pixel_4685/AMP_IN pixel_4685/SF_IB
+ pixel_4685/PIX_OUT pixel_4685/CSA_VREF pixel
Xpixel_4696 pixel_4696/gring pixel_4696/VDD pixel_4696/GND pixel_4696/VREF pixel_4696/ROW_SEL
+ pixel_4696/NB1 pixel_4696/VBIAS pixel_4696/NB2 pixel_4696/AMP_IN pixel_4696/SF_IB
+ pixel_4696/PIX_OUT pixel_4696/CSA_VREF pixel
Xpixel_3940 pixel_3940/gring pixel_3940/VDD pixel_3940/GND pixel_3940/VREF pixel_3940/ROW_SEL
+ pixel_3940/NB1 pixel_3940/VBIAS pixel_3940/NB2 pixel_3940/AMP_IN pixel_3940/SF_IB
+ pixel_3940/PIX_OUT pixel_3940/CSA_VREF pixel
Xpixel_3951 pixel_3951/gring pixel_3951/VDD pixel_3951/GND pixel_3951/VREF pixel_3951/ROW_SEL
+ pixel_3951/NB1 pixel_3951/VBIAS pixel_3951/NB2 pixel_3951/AMP_IN pixel_3951/SF_IB
+ pixel_3951/PIX_OUT pixel_3951/CSA_VREF pixel
Xpixel_3962 pixel_3962/gring pixel_3962/VDD pixel_3962/GND pixel_3962/VREF pixel_3962/ROW_SEL
+ pixel_3962/NB1 pixel_3962/VBIAS pixel_3962/NB2 pixel_3962/AMP_IN pixel_3962/SF_IB
+ pixel_3962/PIX_OUT pixel_3962/CSA_VREF pixel
Xpixel_3973 pixel_3973/gring pixel_3973/VDD pixel_3973/GND pixel_3973/VREF pixel_3973/ROW_SEL
+ pixel_3973/NB1 pixel_3973/VBIAS pixel_3973/NB2 pixel_3973/AMP_IN pixel_3973/SF_IB
+ pixel_3973/PIX_OUT pixel_3973/CSA_VREF pixel
Xpixel_3984 pixel_3984/gring pixel_3984/VDD pixel_3984/GND pixel_3984/VREF pixel_3984/ROW_SEL
+ pixel_3984/NB1 pixel_3984/VBIAS pixel_3984/NB2 pixel_3984/AMP_IN pixel_3984/SF_IB
+ pixel_3984/PIX_OUT pixel_3984/CSA_VREF pixel
Xpixel_3995 pixel_3995/gring pixel_3995/VDD pixel_3995/GND pixel_3995/VREF pixel_3995/ROW_SEL
+ pixel_3995/NB1 pixel_3995/VBIAS pixel_3995/NB2 pixel_3995/AMP_IN pixel_3995/SF_IB
+ pixel_3995/PIX_OUT pixel_3995/CSA_VREF pixel
Xpixel_5 pixel_5/gring pixel_5/VDD pixel_5/GND pixel_5/VREF pixel_5/ROW_SEL pixel_5/NB1
+ pixel_5/VBIAS pixel_5/NB2 pixel_5/AMP_IN pixel_5/SF_IB pixel_5/PIX_OUT pixel_5/CSA_VREF
+ pixel
Xpixel_9608 pixel_9608/gring pixel_9608/VDD pixel_9608/GND pixel_9608/VREF pixel_9608/ROW_SEL
+ pixel_9608/NB1 pixel_9608/VBIAS pixel_9608/NB2 pixel_9608/AMP_IN pixel_9608/SF_IB
+ pixel_9608/PIX_OUT pixel_9608/CSA_VREF pixel
Xpixel_9619 pixel_9619/gring pixel_9619/VDD pixel_9619/GND pixel_9619/VREF pixel_9619/ROW_SEL
+ pixel_9619/NB1 pixel_9619/VBIAS pixel_9619/NB2 pixel_9619/AMP_IN pixel_9619/SF_IB
+ pixel_9619/PIX_OUT pixel_9619/CSA_VREF pixel
Xpixel_8918 pixel_8918/gring pixel_8918/VDD pixel_8918/GND pixel_8918/VREF pixel_8918/ROW_SEL
+ pixel_8918/NB1 pixel_8918/VBIAS pixel_8918/NB2 pixel_8918/AMP_IN pixel_8918/SF_IB
+ pixel_8918/PIX_OUT pixel_8918/CSA_VREF pixel
Xpixel_8907 pixel_8907/gring pixel_8907/VDD pixel_8907/GND pixel_8907/VREF pixel_8907/ROW_SEL
+ pixel_8907/NB1 pixel_8907/VBIAS pixel_8907/NB2 pixel_8907/AMP_IN pixel_8907/SF_IB
+ pixel_8907/PIX_OUT pixel_8907/CSA_VREF pixel
Xpixel_8929 pixel_8929/gring pixel_8929/VDD pixel_8929/GND pixel_8929/VREF pixel_8929/ROW_SEL
+ pixel_8929/NB1 pixel_8929/VBIAS pixel_8929/NB2 pixel_8929/AMP_IN pixel_8929/SF_IB
+ pixel_8929/PIX_OUT pixel_8929/CSA_VREF pixel
Xpixel_3214 pixel_3214/gring pixel_3214/VDD pixel_3214/GND pixel_3214/VREF pixel_3214/ROW_SEL
+ pixel_3214/NB1 pixel_3214/VBIAS pixel_3214/NB2 pixel_3214/AMP_IN pixel_3214/SF_IB
+ pixel_3214/PIX_OUT pixel_3214/CSA_VREF pixel
Xpixel_3203 pixel_3203/gring pixel_3203/VDD pixel_3203/GND pixel_3203/VREF pixel_3203/ROW_SEL
+ pixel_3203/NB1 pixel_3203/VBIAS pixel_3203/NB2 pixel_3203/AMP_IN pixel_3203/SF_IB
+ pixel_3203/PIX_OUT pixel_3203/CSA_VREF pixel
Xpixel_2513 pixel_2513/gring pixel_2513/VDD pixel_2513/GND pixel_2513/VREF pixel_2513/ROW_SEL
+ pixel_2513/NB1 pixel_2513/VBIAS pixel_2513/NB2 pixel_2513/AMP_IN pixel_2513/SF_IB
+ pixel_2513/PIX_OUT pixel_2513/CSA_VREF pixel
Xpixel_2502 pixel_2502/gring pixel_2502/VDD pixel_2502/GND pixel_2502/VREF pixel_2502/ROW_SEL
+ pixel_2502/NB1 pixel_2502/VBIAS pixel_2502/NB2 pixel_2502/AMP_IN pixel_2502/SF_IB
+ pixel_2502/PIX_OUT pixel_2502/CSA_VREF pixel
Xpixel_3247 pixel_3247/gring pixel_3247/VDD pixel_3247/GND pixel_3247/VREF pixel_3247/ROW_SEL
+ pixel_3247/NB1 pixel_3247/VBIAS pixel_3247/NB2 pixel_3247/AMP_IN pixel_3247/SF_IB
+ pixel_3247/PIX_OUT pixel_3247/CSA_VREF pixel
Xpixel_3236 pixel_3236/gring pixel_3236/VDD pixel_3236/GND pixel_3236/VREF pixel_3236/ROW_SEL
+ pixel_3236/NB1 pixel_3236/VBIAS pixel_3236/NB2 pixel_3236/AMP_IN pixel_3236/SF_IB
+ pixel_3236/PIX_OUT pixel_3236/CSA_VREF pixel
Xpixel_3225 pixel_3225/gring pixel_3225/VDD pixel_3225/GND pixel_3225/VREF pixel_3225/ROW_SEL
+ pixel_3225/NB1 pixel_3225/VBIAS pixel_3225/NB2 pixel_3225/AMP_IN pixel_3225/SF_IB
+ pixel_3225/PIX_OUT pixel_3225/CSA_VREF pixel
Xpixel_1801 pixel_1801/gring pixel_1801/VDD pixel_1801/GND pixel_1801/VREF pixel_1801/ROW_SEL
+ pixel_1801/NB1 pixel_1801/VBIAS pixel_1801/NB2 pixel_1801/AMP_IN pixel_1801/SF_IB
+ pixel_1801/PIX_OUT pixel_1801/CSA_VREF pixel
Xpixel_2546 pixel_2546/gring pixel_2546/VDD pixel_2546/GND pixel_2546/VREF pixel_2546/ROW_SEL
+ pixel_2546/NB1 pixel_2546/VBIAS pixel_2546/NB2 pixel_2546/AMP_IN pixel_2546/SF_IB
+ pixel_2546/PIX_OUT pixel_2546/CSA_VREF pixel
Xpixel_2535 pixel_2535/gring pixel_2535/VDD pixel_2535/GND pixel_2535/VREF pixel_2535/ROW_SEL
+ pixel_2535/NB1 pixel_2535/VBIAS pixel_2535/NB2 pixel_2535/AMP_IN pixel_2535/SF_IB
+ pixel_2535/PIX_OUT pixel_2535/CSA_VREF pixel
Xpixel_2524 pixel_2524/gring pixel_2524/VDD pixel_2524/GND pixel_2524/VREF pixel_2524/ROW_SEL
+ pixel_2524/NB1 pixel_2524/VBIAS pixel_2524/NB2 pixel_2524/AMP_IN pixel_2524/SF_IB
+ pixel_2524/PIX_OUT pixel_2524/CSA_VREF pixel
Xpixel_3269 pixel_3269/gring pixel_3269/VDD pixel_3269/GND pixel_3269/VREF pixel_3269/ROW_SEL
+ pixel_3269/NB1 pixel_3269/VBIAS pixel_3269/NB2 pixel_3269/AMP_IN pixel_3269/SF_IB
+ pixel_3269/PIX_OUT pixel_3269/CSA_VREF pixel
Xpixel_3258 pixel_3258/gring pixel_3258/VDD pixel_3258/GND pixel_3258/VREF pixel_3258/ROW_SEL
+ pixel_3258/NB1 pixel_3258/VBIAS pixel_3258/NB2 pixel_3258/AMP_IN pixel_3258/SF_IB
+ pixel_3258/PIX_OUT pixel_3258/CSA_VREF pixel
Xpixel_1834 pixel_1834/gring pixel_1834/VDD pixel_1834/GND pixel_1834/VREF pixel_1834/ROW_SEL
+ pixel_1834/NB1 pixel_1834/VBIAS pixel_1834/NB2 pixel_1834/AMP_IN pixel_1834/SF_IB
+ pixel_1834/PIX_OUT pixel_1834/CSA_VREF pixel
Xpixel_1823 pixel_1823/gring pixel_1823/VDD pixel_1823/GND pixel_1823/VREF pixel_1823/ROW_SEL
+ pixel_1823/NB1 pixel_1823/VBIAS pixel_1823/NB2 pixel_1823/AMP_IN pixel_1823/SF_IB
+ pixel_1823/PIX_OUT pixel_1823/CSA_VREF pixel
Xpixel_1812 pixel_1812/gring pixel_1812/VDD pixel_1812/GND pixel_1812/VREF pixel_1812/ROW_SEL
+ pixel_1812/NB1 pixel_1812/VBIAS pixel_1812/NB2 pixel_1812/AMP_IN pixel_1812/SF_IB
+ pixel_1812/PIX_OUT pixel_1812/CSA_VREF pixel
Xpixel_2579 pixel_2579/gring pixel_2579/VDD pixel_2579/GND pixel_2579/VREF pixel_2579/ROW_SEL
+ pixel_2579/NB1 pixel_2579/VBIAS pixel_2579/NB2 pixel_2579/AMP_IN pixel_2579/SF_IB
+ pixel_2579/PIX_OUT pixel_2579/CSA_VREF pixel
Xpixel_2568 pixel_2568/gring pixel_2568/VDD pixel_2568/GND pixel_2568/VREF pixel_2568/ROW_SEL
+ pixel_2568/NB1 pixel_2568/VBIAS pixel_2568/NB2 pixel_2568/AMP_IN pixel_2568/SF_IB
+ pixel_2568/PIX_OUT pixel_2568/CSA_VREF pixel
Xpixel_2557 pixel_2557/gring pixel_2557/VDD pixel_2557/GND pixel_2557/VREF pixel_2557/ROW_SEL
+ pixel_2557/NB1 pixel_2557/VBIAS pixel_2557/NB2 pixel_2557/AMP_IN pixel_2557/SF_IB
+ pixel_2557/PIX_OUT pixel_2557/CSA_VREF pixel
Xpixel_1878 pixel_1878/gring pixel_1878/VDD pixel_1878/GND pixel_1878/VREF pixel_1878/ROW_SEL
+ pixel_1878/NB1 pixel_1878/VBIAS pixel_1878/NB2 pixel_1878/AMP_IN pixel_1878/SF_IB
+ pixel_1878/PIX_OUT pixel_1878/CSA_VREF pixel
Xpixel_1867 pixel_1867/gring pixel_1867/VDD pixel_1867/GND pixel_1867/VREF pixel_1867/ROW_SEL
+ pixel_1867/NB1 pixel_1867/VBIAS pixel_1867/NB2 pixel_1867/AMP_IN pixel_1867/SF_IB
+ pixel_1867/PIX_OUT pixel_1867/CSA_VREF pixel
Xpixel_1856 pixel_1856/gring pixel_1856/VDD pixel_1856/GND pixel_1856/VREF pixel_1856/ROW_SEL
+ pixel_1856/NB1 pixel_1856/VBIAS pixel_1856/NB2 pixel_1856/AMP_IN pixel_1856/SF_IB
+ pixel_1856/PIX_OUT pixel_1856/CSA_VREF pixel
Xpixel_1845 pixel_1845/gring pixel_1845/VDD pixel_1845/GND pixel_1845/VREF pixel_1845/ROW_SEL
+ pixel_1845/NB1 pixel_1845/VBIAS pixel_1845/NB2 pixel_1845/AMP_IN pixel_1845/SF_IB
+ pixel_1845/PIX_OUT pixel_1845/CSA_VREF pixel
Xpixel_1889 pixel_1889/gring pixel_1889/VDD pixel_1889/GND pixel_1889/VREF pixel_1889/ROW_SEL
+ pixel_1889/NB1 pixel_1889/VBIAS pixel_1889/NB2 pixel_1889/AMP_IN pixel_1889/SF_IB
+ pixel_1889/PIX_OUT pixel_1889/CSA_VREF pixel
Xpixel_5150 pixel_5150/gring pixel_5150/VDD pixel_5150/GND pixel_5150/VREF pixel_5150/ROW_SEL
+ pixel_5150/NB1 pixel_5150/VBIAS pixel_5150/NB2 pixel_5150/AMP_IN pixel_5150/SF_IB
+ pixel_5150/PIX_OUT pixel_5150/CSA_VREF pixel
Xpixel_5161 pixel_5161/gring pixel_5161/VDD pixel_5161/GND pixel_5161/VREF pixel_5161/ROW_SEL
+ pixel_5161/NB1 pixel_5161/VBIAS pixel_5161/NB2 pixel_5161/AMP_IN pixel_5161/SF_IB
+ pixel_5161/PIX_OUT pixel_5161/CSA_VREF pixel
Xpixel_5172 pixel_5172/gring pixel_5172/VDD pixel_5172/GND pixel_5172/VREF pixel_5172/ROW_SEL
+ pixel_5172/NB1 pixel_5172/VBIAS pixel_5172/NB2 pixel_5172/AMP_IN pixel_5172/SF_IB
+ pixel_5172/PIX_OUT pixel_5172/CSA_VREF pixel
Xpixel_5183 pixel_5183/gring pixel_5183/VDD pixel_5183/GND pixel_5183/VREF pixel_5183/ROW_SEL
+ pixel_5183/NB1 pixel_5183/VBIAS pixel_5183/NB2 pixel_5183/AMP_IN pixel_5183/SF_IB
+ pixel_5183/PIX_OUT pixel_5183/CSA_VREF pixel
Xpixel_5194 pixel_5194/gring pixel_5194/VDD pixel_5194/GND pixel_5194/VREF pixel_5194/ROW_SEL
+ pixel_5194/NB1 pixel_5194/VBIAS pixel_5194/NB2 pixel_5194/AMP_IN pixel_5194/SF_IB
+ pixel_5194/PIX_OUT pixel_5194/CSA_VREF pixel
Xpixel_4460 pixel_4460/gring pixel_4460/VDD pixel_4460/GND pixel_4460/VREF pixel_4460/ROW_SEL
+ pixel_4460/NB1 pixel_4460/VBIAS pixel_4460/NB2 pixel_4460/AMP_IN pixel_4460/SF_IB
+ pixel_4460/PIX_OUT pixel_4460/CSA_VREF pixel
Xpixel_4471 pixel_4471/gring pixel_4471/VDD pixel_4471/GND pixel_4471/VREF pixel_4471/ROW_SEL
+ pixel_4471/NB1 pixel_4471/VBIAS pixel_4471/NB2 pixel_4471/AMP_IN pixel_4471/SF_IB
+ pixel_4471/PIX_OUT pixel_4471/CSA_VREF pixel
Xpixel_3770 pixel_3770/gring pixel_3770/VDD pixel_3770/GND pixel_3770/VREF pixel_3770/ROW_SEL
+ pixel_3770/NB1 pixel_3770/VBIAS pixel_3770/NB2 pixel_3770/AMP_IN pixel_3770/SF_IB
+ pixel_3770/PIX_OUT pixel_3770/CSA_VREF pixel
Xpixel_4482 pixel_4482/gring pixel_4482/VDD pixel_4482/GND pixel_4482/VREF pixel_4482/ROW_SEL
+ pixel_4482/NB1 pixel_4482/VBIAS pixel_4482/NB2 pixel_4482/AMP_IN pixel_4482/SF_IB
+ pixel_4482/PIX_OUT pixel_4482/CSA_VREF pixel
Xpixel_4493 pixel_4493/gring pixel_4493/VDD pixel_4493/GND pixel_4493/VREF pixel_4493/ROW_SEL
+ pixel_4493/NB1 pixel_4493/VBIAS pixel_4493/NB2 pixel_4493/AMP_IN pixel_4493/SF_IB
+ pixel_4493/PIX_OUT pixel_4493/CSA_VREF pixel
Xpixel_3792 pixel_3792/gring pixel_3792/VDD pixel_3792/GND pixel_3792/VREF pixel_3792/ROW_SEL
+ pixel_3792/NB1 pixel_3792/VBIAS pixel_3792/NB2 pixel_3792/AMP_IN pixel_3792/SF_IB
+ pixel_3792/PIX_OUT pixel_3792/CSA_VREF pixel
Xpixel_3781 pixel_3781/gring pixel_3781/VDD pixel_3781/GND pixel_3781/VREF pixel_3781/ROW_SEL
+ pixel_3781/NB1 pixel_3781/VBIAS pixel_3781/NB2 pixel_3781/AMP_IN pixel_3781/SF_IB
+ pixel_3781/PIX_OUT pixel_3781/CSA_VREF pixel
Xpixel_1119 pixel_1119/gring pixel_1119/VDD pixel_1119/GND pixel_1119/VREF pixel_1119/ROW_SEL
+ pixel_1119/NB1 pixel_1119/VBIAS pixel_1119/NB2 pixel_1119/AMP_IN pixel_1119/SF_IB
+ pixel_1119/PIX_OUT pixel_1119/CSA_VREF pixel
Xpixel_1108 pixel_1108/gring pixel_1108/VDD pixel_1108/GND pixel_1108/VREF pixel_1108/ROW_SEL
+ pixel_1108/NB1 pixel_1108/VBIAS pixel_1108/NB2 pixel_1108/AMP_IN pixel_1108/SF_IB
+ pixel_1108/PIX_OUT pixel_1108/CSA_VREF pixel
Xpixel_9405 pixel_9405/gring pixel_9405/VDD pixel_9405/GND pixel_9405/VREF pixel_9405/ROW_SEL
+ pixel_9405/NB1 pixel_9405/VBIAS pixel_9405/NB2 pixel_9405/AMP_IN pixel_9405/SF_IB
+ pixel_9405/PIX_OUT pixel_9405/CSA_VREF pixel
Xpixel_9438 pixel_9438/gring pixel_9438/VDD pixel_9438/GND pixel_9438/VREF pixel_9438/ROW_SEL
+ pixel_9438/NB1 pixel_9438/VBIAS pixel_9438/NB2 pixel_9438/AMP_IN pixel_9438/SF_IB
+ pixel_9438/PIX_OUT pixel_9438/CSA_VREF pixel
Xpixel_9427 pixel_9427/gring pixel_9427/VDD pixel_9427/GND pixel_9427/VREF pixel_9427/ROW_SEL
+ pixel_9427/NB1 pixel_9427/VBIAS pixel_9427/NB2 pixel_9427/AMP_IN pixel_9427/SF_IB
+ pixel_9427/PIX_OUT pixel_9427/CSA_VREF pixel
Xpixel_9416 pixel_9416/gring pixel_9416/VDD pixel_9416/GND pixel_9416/VREF pixel_9416/ROW_SEL
+ pixel_9416/NB1 pixel_9416/VBIAS pixel_9416/NB2 pixel_9416/AMP_IN pixel_9416/SF_IB
+ pixel_9416/PIX_OUT pixel_9416/CSA_VREF pixel
Xpixel_8726 pixel_8726/gring pixel_8726/VDD pixel_8726/GND pixel_8726/VREF pixel_8726/ROW_SEL
+ pixel_8726/NB1 pixel_8726/VBIAS pixel_8726/NB2 pixel_8726/AMP_IN pixel_8726/SF_IB
+ pixel_8726/PIX_OUT pixel_8726/CSA_VREF pixel
Xpixel_8715 pixel_8715/gring pixel_8715/VDD pixel_8715/GND pixel_8715/VREF pixel_8715/ROW_SEL
+ pixel_8715/NB1 pixel_8715/VBIAS pixel_8715/NB2 pixel_8715/AMP_IN pixel_8715/SF_IB
+ pixel_8715/PIX_OUT pixel_8715/CSA_VREF pixel
Xpixel_8704 pixel_8704/gring pixel_8704/VDD pixel_8704/GND pixel_8704/VREF pixel_8704/ROW_SEL
+ pixel_8704/NB1 pixel_8704/VBIAS pixel_8704/NB2 pixel_8704/AMP_IN pixel_8704/SF_IB
+ pixel_8704/PIX_OUT pixel_8704/CSA_VREF pixel
Xpixel_9449 pixel_9449/gring pixel_9449/VDD pixel_9449/GND pixel_9449/VREF pixel_9449/ROW_SEL
+ pixel_9449/NB1 pixel_9449/VBIAS pixel_9449/NB2 pixel_9449/AMP_IN pixel_9449/SF_IB
+ pixel_9449/PIX_OUT pixel_9449/CSA_VREF pixel
Xpixel_8759 pixel_8759/gring pixel_8759/VDD pixel_8759/GND pixel_8759/VREF pixel_8759/ROW_SEL
+ pixel_8759/NB1 pixel_8759/VBIAS pixel_8759/NB2 pixel_8759/AMP_IN pixel_8759/SF_IB
+ pixel_8759/PIX_OUT pixel_8759/CSA_VREF pixel
Xpixel_8748 pixel_8748/gring pixel_8748/VDD pixel_8748/GND pixel_8748/VREF pixel_8748/ROW_SEL
+ pixel_8748/NB1 pixel_8748/VBIAS pixel_8748/NB2 pixel_8748/AMP_IN pixel_8748/SF_IB
+ pixel_8748/PIX_OUT pixel_8748/CSA_VREF pixel
Xpixel_8737 pixel_8737/gring pixel_8737/VDD pixel_8737/GND pixel_8737/VREF pixel_8737/ROW_SEL
+ pixel_8737/NB1 pixel_8737/VBIAS pixel_8737/NB2 pixel_8737/AMP_IN pixel_8737/SF_IB
+ pixel_8737/PIX_OUT pixel_8737/CSA_VREF pixel
Xpixel_3022 pixel_3022/gring pixel_3022/VDD pixel_3022/GND pixel_3022/VREF pixel_3022/ROW_SEL
+ pixel_3022/NB1 pixel_3022/VBIAS pixel_3022/NB2 pixel_3022/AMP_IN pixel_3022/SF_IB
+ pixel_3022/PIX_OUT pixel_3022/CSA_VREF pixel
Xpixel_3011 pixel_3011/gring pixel_3011/VDD pixel_3011/GND pixel_3011/VREF pixel_3011/ROW_SEL
+ pixel_3011/NB1 pixel_3011/VBIAS pixel_3011/NB2 pixel_3011/AMP_IN pixel_3011/SF_IB
+ pixel_3011/PIX_OUT pixel_3011/CSA_VREF pixel
Xpixel_3000 pixel_3000/gring pixel_3000/VDD pixel_3000/GND pixel_3000/VREF pixel_3000/ROW_SEL
+ pixel_3000/NB1 pixel_3000/VBIAS pixel_3000/NB2 pixel_3000/AMP_IN pixel_3000/SF_IB
+ pixel_3000/PIX_OUT pixel_3000/CSA_VREF pixel
Xpixel_2321 pixel_2321/gring pixel_2321/VDD pixel_2321/GND pixel_2321/VREF pixel_2321/ROW_SEL
+ pixel_2321/NB1 pixel_2321/VBIAS pixel_2321/NB2 pixel_2321/AMP_IN pixel_2321/SF_IB
+ pixel_2321/PIX_OUT pixel_2321/CSA_VREF pixel
Xpixel_2310 pixel_2310/gring pixel_2310/VDD pixel_2310/GND pixel_2310/VREF pixel_2310/ROW_SEL
+ pixel_2310/NB1 pixel_2310/VBIAS pixel_2310/NB2 pixel_2310/AMP_IN pixel_2310/SF_IB
+ pixel_2310/PIX_OUT pixel_2310/CSA_VREF pixel
Xpixel_3066 pixel_3066/gring pixel_3066/VDD pixel_3066/GND pixel_3066/VREF pixel_3066/ROW_SEL
+ pixel_3066/NB1 pixel_3066/VBIAS pixel_3066/NB2 pixel_3066/AMP_IN pixel_3066/SF_IB
+ pixel_3066/PIX_OUT pixel_3066/CSA_VREF pixel
Xpixel_3055 pixel_3055/gring pixel_3055/VDD pixel_3055/GND pixel_3055/VREF pixel_3055/ROW_SEL
+ pixel_3055/NB1 pixel_3055/VBIAS pixel_3055/NB2 pixel_3055/AMP_IN pixel_3055/SF_IB
+ pixel_3055/PIX_OUT pixel_3055/CSA_VREF pixel
Xpixel_3044 pixel_3044/gring pixel_3044/VDD pixel_3044/GND pixel_3044/VREF pixel_3044/ROW_SEL
+ pixel_3044/NB1 pixel_3044/VBIAS pixel_3044/NB2 pixel_3044/AMP_IN pixel_3044/SF_IB
+ pixel_3044/PIX_OUT pixel_3044/CSA_VREF pixel
Xpixel_3033 pixel_3033/gring pixel_3033/VDD pixel_3033/GND pixel_3033/VREF pixel_3033/ROW_SEL
+ pixel_3033/NB1 pixel_3033/VBIAS pixel_3033/NB2 pixel_3033/AMP_IN pixel_3033/SF_IB
+ pixel_3033/PIX_OUT pixel_3033/CSA_VREF pixel
Xpixel_2354 pixel_2354/gring pixel_2354/VDD pixel_2354/GND pixel_2354/VREF pixel_2354/ROW_SEL
+ pixel_2354/NB1 pixel_2354/VBIAS pixel_2354/NB2 pixel_2354/AMP_IN pixel_2354/SF_IB
+ pixel_2354/PIX_OUT pixel_2354/CSA_VREF pixel
Xpixel_2343 pixel_2343/gring pixel_2343/VDD pixel_2343/GND pixel_2343/VREF pixel_2343/ROW_SEL
+ pixel_2343/NB1 pixel_2343/VBIAS pixel_2343/NB2 pixel_2343/AMP_IN pixel_2343/SF_IB
+ pixel_2343/PIX_OUT pixel_2343/CSA_VREF pixel
Xpixel_2332 pixel_2332/gring pixel_2332/VDD pixel_2332/GND pixel_2332/VREF pixel_2332/ROW_SEL
+ pixel_2332/NB1 pixel_2332/VBIAS pixel_2332/NB2 pixel_2332/AMP_IN pixel_2332/SF_IB
+ pixel_2332/PIX_OUT pixel_2332/CSA_VREF pixel
Xpixel_3099 pixel_3099/gring pixel_3099/VDD pixel_3099/GND pixel_3099/VREF pixel_3099/ROW_SEL
+ pixel_3099/NB1 pixel_3099/VBIAS pixel_3099/NB2 pixel_3099/AMP_IN pixel_3099/SF_IB
+ pixel_3099/PIX_OUT pixel_3099/CSA_VREF pixel
Xpixel_3088 pixel_3088/gring pixel_3088/VDD pixel_3088/GND pixel_3088/VREF pixel_3088/ROW_SEL
+ pixel_3088/NB1 pixel_3088/VBIAS pixel_3088/NB2 pixel_3088/AMP_IN pixel_3088/SF_IB
+ pixel_3088/PIX_OUT pixel_3088/CSA_VREF pixel
Xpixel_3077 pixel_3077/gring pixel_3077/VDD pixel_3077/GND pixel_3077/VREF pixel_3077/ROW_SEL
+ pixel_3077/NB1 pixel_3077/VBIAS pixel_3077/NB2 pixel_3077/AMP_IN pixel_3077/SF_IB
+ pixel_3077/PIX_OUT pixel_3077/CSA_VREF pixel
Xpixel_1642 pixel_1642/gring pixel_1642/VDD pixel_1642/GND pixel_1642/VREF pixel_1642/ROW_SEL
+ pixel_1642/NB1 pixel_1642/VBIAS pixel_1642/NB2 pixel_1642/AMP_IN pixel_1642/SF_IB
+ pixel_1642/PIX_OUT pixel_1642/CSA_VREF pixel
Xpixel_1631 pixel_1631/gring pixel_1631/VDD pixel_1631/GND pixel_1631/VREF pixel_1631/ROW_SEL
+ pixel_1631/NB1 pixel_1631/VBIAS pixel_1631/NB2 pixel_1631/AMP_IN pixel_1631/SF_IB
+ pixel_1631/PIX_OUT pixel_1631/CSA_VREF pixel
Xpixel_1620 pixel_1620/gring pixel_1620/VDD pixel_1620/GND pixel_1620/VREF pixel_1620/ROW_SEL
+ pixel_1620/NB1 pixel_1620/VBIAS pixel_1620/NB2 pixel_1620/AMP_IN pixel_1620/SF_IB
+ pixel_1620/PIX_OUT pixel_1620/CSA_VREF pixel
Xpixel_2387 pixel_2387/gring pixel_2387/VDD pixel_2387/GND pixel_2387/VREF pixel_2387/ROW_SEL
+ pixel_2387/NB1 pixel_2387/VBIAS pixel_2387/NB2 pixel_2387/AMP_IN pixel_2387/SF_IB
+ pixel_2387/PIX_OUT pixel_2387/CSA_VREF pixel
Xpixel_2376 pixel_2376/gring pixel_2376/VDD pixel_2376/GND pixel_2376/VREF pixel_2376/ROW_SEL
+ pixel_2376/NB1 pixel_2376/VBIAS pixel_2376/NB2 pixel_2376/AMP_IN pixel_2376/SF_IB
+ pixel_2376/PIX_OUT pixel_2376/CSA_VREF pixel
Xpixel_2365 pixel_2365/gring pixel_2365/VDD pixel_2365/GND pixel_2365/VREF pixel_2365/ROW_SEL
+ pixel_2365/NB1 pixel_2365/VBIAS pixel_2365/NB2 pixel_2365/AMP_IN pixel_2365/SF_IB
+ pixel_2365/PIX_OUT pixel_2365/CSA_VREF pixel
Xpixel_1686 pixel_1686/gring pixel_1686/VDD pixel_1686/GND pixel_1686/VREF pixel_1686/ROW_SEL
+ pixel_1686/NB1 pixel_1686/VBIAS pixel_1686/NB2 pixel_1686/AMP_IN pixel_1686/SF_IB
+ pixel_1686/PIX_OUT pixel_1686/CSA_VREF pixel
Xpixel_1675 pixel_1675/gring pixel_1675/VDD pixel_1675/GND pixel_1675/VREF pixel_1675/ROW_SEL
+ pixel_1675/NB1 pixel_1675/VBIAS pixel_1675/NB2 pixel_1675/AMP_IN pixel_1675/SF_IB
+ pixel_1675/PIX_OUT pixel_1675/CSA_VREF pixel
Xpixel_1664 pixel_1664/gring pixel_1664/VDD pixel_1664/GND pixel_1664/VREF pixel_1664/ROW_SEL
+ pixel_1664/NB1 pixel_1664/VBIAS pixel_1664/NB2 pixel_1664/AMP_IN pixel_1664/SF_IB
+ pixel_1664/PIX_OUT pixel_1664/CSA_VREF pixel
Xpixel_1653 pixel_1653/gring pixel_1653/VDD pixel_1653/GND pixel_1653/VREF pixel_1653/ROW_SEL
+ pixel_1653/NB1 pixel_1653/VBIAS pixel_1653/NB2 pixel_1653/AMP_IN pixel_1653/SF_IB
+ pixel_1653/PIX_OUT pixel_1653/CSA_VREF pixel
Xpixel_2398 pixel_2398/gring pixel_2398/VDD pixel_2398/GND pixel_2398/VREF pixel_2398/ROW_SEL
+ pixel_2398/NB1 pixel_2398/VBIAS pixel_2398/NB2 pixel_2398/AMP_IN pixel_2398/SF_IB
+ pixel_2398/PIX_OUT pixel_2398/CSA_VREF pixel
Xpixel_1697 pixel_1697/gring pixel_1697/VDD pixel_1697/GND pixel_1697/VREF pixel_1697/ROW_SEL
+ pixel_1697/NB1 pixel_1697/VBIAS pixel_1697/NB2 pixel_1697/AMP_IN pixel_1697/SF_IB
+ pixel_1697/PIX_OUT pixel_1697/CSA_VREF pixel
Xpixel_9950 pixel_9950/gring pixel_9950/VDD pixel_9950/GND pixel_9950/VREF pixel_9950/ROW_SEL
+ pixel_9950/NB1 pixel_9950/VBIAS pixel_9950/NB2 pixel_9950/AMP_IN pixel_9950/SF_IB
+ pixel_9950/PIX_OUT pixel_9950/CSA_VREF pixel
Xpixel_9961 pixel_9961/gring pixel_9961/VDD pixel_9961/GND pixel_9961/VREF pixel_9961/ROW_SEL
+ pixel_9961/NB1 pixel_9961/VBIAS pixel_9961/NB2 pixel_9961/AMP_IN pixel_9961/SF_IB
+ pixel_9961/PIX_OUT pixel_9961/CSA_VREF pixel
Xpixel_9972 pixel_9972/gring pixel_9972/VDD pixel_9972/GND pixel_9972/VREF pixel_9972/ROW_SEL
+ pixel_9972/NB1 pixel_9972/VBIAS pixel_9972/NB2 pixel_9972/AMP_IN pixel_9972/SF_IB
+ pixel_9972/PIX_OUT pixel_9972/CSA_VREF pixel
Xpixel_9983 pixel_9983/gring pixel_9983/VDD pixel_9983/GND pixel_9983/VREF pixel_9983/ROW_SEL
+ pixel_9983/NB1 pixel_9983/VBIAS pixel_9983/NB2 pixel_9983/AMP_IN pixel_9983/SF_IB
+ pixel_9983/PIX_OUT pixel_9983/CSA_VREF pixel
Xpixel_9994 pixel_9994/gring pixel_9994/VDD pixel_9994/GND pixel_9994/VREF pixel_9994/ROW_SEL
+ pixel_9994/NB1 pixel_9994/VBIAS pixel_9994/NB2 pixel_9994/AMP_IN pixel_9994/SF_IB
+ pixel_9994/PIX_OUT pixel_9994/CSA_VREF pixel
Xpixel_4290 pixel_4290/gring pixel_4290/VDD pixel_4290/GND pixel_4290/VREF pixel_4290/ROW_SEL
+ pixel_4290/NB1 pixel_4290/VBIAS pixel_4290/NB2 pixel_4290/AMP_IN pixel_4290/SF_IB
+ pixel_4290/PIX_OUT pixel_4290/CSA_VREF pixel
Xpixel_6609 pixel_6609/gring pixel_6609/VDD pixel_6609/GND pixel_6609/VREF pixel_6609/ROW_SEL
+ pixel_6609/NB1 pixel_6609/VBIAS pixel_6609/NB2 pixel_6609/AMP_IN pixel_6609/SF_IB
+ pixel_6609/PIX_OUT pixel_6609/CSA_VREF pixel
Xpixel_5908 pixel_5908/gring pixel_5908/VDD pixel_5908/GND pixel_5908/VREF pixel_5908/ROW_SEL
+ pixel_5908/NB1 pixel_5908/VBIAS pixel_5908/NB2 pixel_5908/AMP_IN pixel_5908/SF_IB
+ pixel_5908/PIX_OUT pixel_5908/CSA_VREF pixel
Xpixel_5919 pixel_5919/gring pixel_5919/VDD pixel_5919/GND pixel_5919/VREF pixel_5919/ROW_SEL
+ pixel_5919/NB1 pixel_5919/VBIAS pixel_5919/NB2 pixel_5919/AMP_IN pixel_5919/SF_IB
+ pixel_5919/PIX_OUT pixel_5919/CSA_VREF pixel
Xpixel_9213 pixel_9213/gring pixel_9213/VDD pixel_9213/GND pixel_9213/VREF pixel_9213/ROW_SEL
+ pixel_9213/NB1 pixel_9213/VBIAS pixel_9213/NB2 pixel_9213/AMP_IN pixel_9213/SF_IB
+ pixel_9213/PIX_OUT pixel_9213/CSA_VREF pixel
Xpixel_9202 pixel_9202/gring pixel_9202/VDD pixel_9202/GND pixel_9202/VREF pixel_9202/ROW_SEL
+ pixel_9202/NB1 pixel_9202/VBIAS pixel_9202/NB2 pixel_9202/AMP_IN pixel_9202/SF_IB
+ pixel_9202/PIX_OUT pixel_9202/CSA_VREF pixel
Xpixel_8501 pixel_8501/gring pixel_8501/VDD pixel_8501/GND pixel_8501/VREF pixel_8501/ROW_SEL
+ pixel_8501/NB1 pixel_8501/VBIAS pixel_8501/NB2 pixel_8501/AMP_IN pixel_8501/SF_IB
+ pixel_8501/PIX_OUT pixel_8501/CSA_VREF pixel
Xpixel_9246 pixel_9246/gring pixel_9246/VDD pixel_9246/GND pixel_9246/VREF pixel_9246/ROW_SEL
+ pixel_9246/NB1 pixel_9246/VBIAS pixel_9246/NB2 pixel_9246/AMP_IN pixel_9246/SF_IB
+ pixel_9246/PIX_OUT pixel_9246/CSA_VREF pixel
Xpixel_9235 pixel_9235/gring pixel_9235/VDD pixel_9235/GND pixel_9235/VREF pixel_9235/ROW_SEL
+ pixel_9235/NB1 pixel_9235/VBIAS pixel_9235/NB2 pixel_9235/AMP_IN pixel_9235/SF_IB
+ pixel_9235/PIX_OUT pixel_9235/CSA_VREF pixel
Xpixel_9224 pixel_9224/gring pixel_9224/VDD pixel_9224/GND pixel_9224/VREF pixel_9224/ROW_SEL
+ pixel_9224/NB1 pixel_9224/VBIAS pixel_9224/NB2 pixel_9224/AMP_IN pixel_9224/SF_IB
+ pixel_9224/PIX_OUT pixel_9224/CSA_VREF pixel
Xpixel_8545 pixel_8545/gring pixel_8545/VDD pixel_8545/GND pixel_8545/VREF pixel_8545/ROW_SEL
+ pixel_8545/NB1 pixel_8545/VBIAS pixel_8545/NB2 pixel_8545/AMP_IN pixel_8545/SF_IB
+ pixel_8545/PIX_OUT pixel_8545/CSA_VREF pixel
Xpixel_8534 pixel_8534/gring pixel_8534/VDD pixel_8534/GND pixel_8534/VREF pixel_8534/ROW_SEL
+ pixel_8534/NB1 pixel_8534/VBIAS pixel_8534/NB2 pixel_8534/AMP_IN pixel_8534/SF_IB
+ pixel_8534/PIX_OUT pixel_8534/CSA_VREF pixel
Xpixel_8523 pixel_8523/gring pixel_8523/VDD pixel_8523/GND pixel_8523/VREF pixel_8523/ROW_SEL
+ pixel_8523/NB1 pixel_8523/VBIAS pixel_8523/NB2 pixel_8523/AMP_IN pixel_8523/SF_IB
+ pixel_8523/PIX_OUT pixel_8523/CSA_VREF pixel
Xpixel_8512 pixel_8512/gring pixel_8512/VDD pixel_8512/GND pixel_8512/VREF pixel_8512/ROW_SEL
+ pixel_8512/NB1 pixel_8512/VBIAS pixel_8512/NB2 pixel_8512/AMP_IN pixel_8512/SF_IB
+ pixel_8512/PIX_OUT pixel_8512/CSA_VREF pixel
Xpixel_9279 pixel_9279/gring pixel_9279/VDD pixel_9279/GND pixel_9279/VREF pixel_9279/ROW_SEL
+ pixel_9279/NB1 pixel_9279/VBIAS pixel_9279/NB2 pixel_9279/AMP_IN pixel_9279/SF_IB
+ pixel_9279/PIX_OUT pixel_9279/CSA_VREF pixel
Xpixel_9268 pixel_9268/gring pixel_9268/VDD pixel_9268/GND pixel_9268/VREF pixel_9268/ROW_SEL
+ pixel_9268/NB1 pixel_9268/VBIAS pixel_9268/NB2 pixel_9268/AMP_IN pixel_9268/SF_IB
+ pixel_9268/PIX_OUT pixel_9268/CSA_VREF pixel
Xpixel_9257 pixel_9257/gring pixel_9257/VDD pixel_9257/GND pixel_9257/VREF pixel_9257/ROW_SEL
+ pixel_9257/NB1 pixel_9257/VBIAS pixel_9257/NB2 pixel_9257/AMP_IN pixel_9257/SF_IB
+ pixel_9257/PIX_OUT pixel_9257/CSA_VREF pixel
Xpixel_7800 pixel_7800/gring pixel_7800/VDD pixel_7800/GND pixel_7800/VREF pixel_7800/ROW_SEL
+ pixel_7800/NB1 pixel_7800/VBIAS pixel_7800/NB2 pixel_7800/AMP_IN pixel_7800/SF_IB
+ pixel_7800/PIX_OUT pixel_7800/CSA_VREF pixel
Xpixel_8578 pixel_8578/gring pixel_8578/VDD pixel_8578/GND pixel_8578/VREF pixel_8578/ROW_SEL
+ pixel_8578/NB1 pixel_8578/VBIAS pixel_8578/NB2 pixel_8578/AMP_IN pixel_8578/SF_IB
+ pixel_8578/PIX_OUT pixel_8578/CSA_VREF pixel
Xpixel_8567 pixel_8567/gring pixel_8567/VDD pixel_8567/GND pixel_8567/VREF pixel_8567/ROW_SEL
+ pixel_8567/NB1 pixel_8567/VBIAS pixel_8567/NB2 pixel_8567/AMP_IN pixel_8567/SF_IB
+ pixel_8567/PIX_OUT pixel_8567/CSA_VREF pixel
Xpixel_8556 pixel_8556/gring pixel_8556/VDD pixel_8556/GND pixel_8556/VREF pixel_8556/ROW_SEL
+ pixel_8556/NB1 pixel_8556/VBIAS pixel_8556/NB2 pixel_8556/AMP_IN pixel_8556/SF_IB
+ pixel_8556/PIX_OUT pixel_8556/CSA_VREF pixel
Xpixel_7811 pixel_7811/gring pixel_7811/VDD pixel_7811/GND pixel_7811/VREF pixel_7811/ROW_SEL
+ pixel_7811/NB1 pixel_7811/VBIAS pixel_7811/NB2 pixel_7811/AMP_IN pixel_7811/SF_IB
+ pixel_7811/PIX_OUT pixel_7811/CSA_VREF pixel
Xpixel_7822 pixel_7822/gring pixel_7822/VDD pixel_7822/GND pixel_7822/VREF pixel_7822/ROW_SEL
+ pixel_7822/NB1 pixel_7822/VBIAS pixel_7822/NB2 pixel_7822/AMP_IN pixel_7822/SF_IB
+ pixel_7822/PIX_OUT pixel_7822/CSA_VREF pixel
Xpixel_7833 pixel_7833/gring pixel_7833/VDD pixel_7833/GND pixel_7833/VREF pixel_7833/ROW_SEL
+ pixel_7833/NB1 pixel_7833/VBIAS pixel_7833/NB2 pixel_7833/AMP_IN pixel_7833/SF_IB
+ pixel_7833/PIX_OUT pixel_7833/CSA_VREF pixel
Xpixel_8589 pixel_8589/gring pixel_8589/VDD pixel_8589/GND pixel_8589/VREF pixel_8589/ROW_SEL
+ pixel_8589/NB1 pixel_8589/VBIAS pixel_8589/NB2 pixel_8589/AMP_IN pixel_8589/SF_IB
+ pixel_8589/PIX_OUT pixel_8589/CSA_VREF pixel
Xpixel_7844 pixel_7844/gring pixel_7844/VDD pixel_7844/GND pixel_7844/VREF pixel_7844/ROW_SEL
+ pixel_7844/NB1 pixel_7844/VBIAS pixel_7844/NB2 pixel_7844/AMP_IN pixel_7844/SF_IB
+ pixel_7844/PIX_OUT pixel_7844/CSA_VREF pixel
Xpixel_7855 pixel_7855/gring pixel_7855/VDD pixel_7855/GND pixel_7855/VREF pixel_7855/ROW_SEL
+ pixel_7855/NB1 pixel_7855/VBIAS pixel_7855/NB2 pixel_7855/AMP_IN pixel_7855/SF_IB
+ pixel_7855/PIX_OUT pixel_7855/CSA_VREF pixel
Xpixel_7866 pixel_7866/gring pixel_7866/VDD pixel_7866/GND pixel_7866/VREF pixel_7866/ROW_SEL
+ pixel_7866/NB1 pixel_7866/VBIAS pixel_7866/NB2 pixel_7866/AMP_IN pixel_7866/SF_IB
+ pixel_7866/PIX_OUT pixel_7866/CSA_VREF pixel
Xpixel_7877 pixel_7877/gring pixel_7877/VDD pixel_7877/GND pixel_7877/VREF pixel_7877/ROW_SEL
+ pixel_7877/NB1 pixel_7877/VBIAS pixel_7877/NB2 pixel_7877/AMP_IN pixel_7877/SF_IB
+ pixel_7877/PIX_OUT pixel_7877/CSA_VREF pixel
Xpixel_7888 pixel_7888/gring pixel_7888/VDD pixel_7888/GND pixel_7888/VREF pixel_7888/ROW_SEL
+ pixel_7888/NB1 pixel_7888/VBIAS pixel_7888/NB2 pixel_7888/AMP_IN pixel_7888/SF_IB
+ pixel_7888/PIX_OUT pixel_7888/CSA_VREF pixel
Xpixel_7899 pixel_7899/gring pixel_7899/VDD pixel_7899/GND pixel_7899/VREF pixel_7899/ROW_SEL
+ pixel_7899/NB1 pixel_7899/VBIAS pixel_7899/NB2 pixel_7899/AMP_IN pixel_7899/SF_IB
+ pixel_7899/PIX_OUT pixel_7899/CSA_VREF pixel
Xpixel_2162 pixel_2162/gring pixel_2162/VDD pixel_2162/GND pixel_2162/VREF pixel_2162/ROW_SEL
+ pixel_2162/NB1 pixel_2162/VBIAS pixel_2162/NB2 pixel_2162/AMP_IN pixel_2162/SF_IB
+ pixel_2162/PIX_OUT pixel_2162/CSA_VREF pixel
Xpixel_2151 pixel_2151/gring pixel_2151/VDD pixel_2151/GND pixel_2151/VREF pixel_2151/ROW_SEL
+ pixel_2151/NB1 pixel_2151/VBIAS pixel_2151/NB2 pixel_2151/AMP_IN pixel_2151/SF_IB
+ pixel_2151/PIX_OUT pixel_2151/CSA_VREF pixel
Xpixel_2140 pixel_2140/gring pixel_2140/VDD pixel_2140/GND pixel_2140/VREF pixel_2140/ROW_SEL
+ pixel_2140/NB1 pixel_2140/VBIAS pixel_2140/NB2 pixel_2140/AMP_IN pixel_2140/SF_IB
+ pixel_2140/PIX_OUT pixel_2140/CSA_VREF pixel
Xpixel_1461 pixel_1461/gring pixel_1461/VDD pixel_1461/GND pixel_1461/VREF pixel_1461/ROW_SEL
+ pixel_1461/NB1 pixel_1461/VBIAS pixel_1461/NB2 pixel_1461/AMP_IN pixel_1461/SF_IB
+ pixel_1461/PIX_OUT pixel_1461/CSA_VREF pixel
Xpixel_1450 pixel_1450/gring pixel_1450/VDD pixel_1450/GND pixel_1450/VREF pixel_1450/ROW_SEL
+ pixel_1450/NB1 pixel_1450/VBIAS pixel_1450/NB2 pixel_1450/AMP_IN pixel_1450/SF_IB
+ pixel_1450/PIX_OUT pixel_1450/CSA_VREF pixel
Xpixel_2195 pixel_2195/gring pixel_2195/VDD pixel_2195/GND pixel_2195/VREF pixel_2195/ROW_SEL
+ pixel_2195/NB1 pixel_2195/VBIAS pixel_2195/NB2 pixel_2195/AMP_IN pixel_2195/SF_IB
+ pixel_2195/PIX_OUT pixel_2195/CSA_VREF pixel
Xpixel_2184 pixel_2184/gring pixel_2184/VDD pixel_2184/GND pixel_2184/VREF pixel_2184/ROW_SEL
+ pixel_2184/NB1 pixel_2184/VBIAS pixel_2184/NB2 pixel_2184/AMP_IN pixel_2184/SF_IB
+ pixel_2184/PIX_OUT pixel_2184/CSA_VREF pixel
Xpixel_2173 pixel_2173/gring pixel_2173/VDD pixel_2173/GND pixel_2173/VREF pixel_2173/ROW_SEL
+ pixel_2173/NB1 pixel_2173/VBIAS pixel_2173/NB2 pixel_2173/AMP_IN pixel_2173/SF_IB
+ pixel_2173/PIX_OUT pixel_2173/CSA_VREF pixel
Xpixel_1494 pixel_1494/gring pixel_1494/VDD pixel_1494/GND pixel_1494/VREF pixel_1494/ROW_SEL
+ pixel_1494/NB1 pixel_1494/VBIAS pixel_1494/NB2 pixel_1494/AMP_IN pixel_1494/SF_IB
+ pixel_1494/PIX_OUT pixel_1494/CSA_VREF pixel
Xpixel_1483 pixel_1483/gring pixel_1483/VDD pixel_1483/GND pixel_1483/VREF pixel_1483/ROW_SEL
+ pixel_1483/NB1 pixel_1483/VBIAS pixel_1483/NB2 pixel_1483/AMP_IN pixel_1483/SF_IB
+ pixel_1483/PIX_OUT pixel_1483/CSA_VREF pixel
Xpixel_1472 pixel_1472/gring pixel_1472/VDD pixel_1472/GND pixel_1472/VREF pixel_1472/ROW_SEL
+ pixel_1472/NB1 pixel_1472/VBIAS pixel_1472/NB2 pixel_1472/AMP_IN pixel_1472/SF_IB
+ pixel_1472/PIX_OUT pixel_1472/CSA_VREF pixel
Xpixel_9780 pixel_9780/gring pixel_9780/VDD pixel_9780/GND pixel_9780/VREF pixel_9780/ROW_SEL
+ pixel_9780/NB1 pixel_9780/VBIAS pixel_9780/NB2 pixel_9780/AMP_IN pixel_9780/SF_IB
+ pixel_9780/PIX_OUT pixel_9780/CSA_VREF pixel
Xpixel_9791 pixel_9791/gring pixel_9791/VDD pixel_9791/GND pixel_9791/VREF pixel_9791/ROW_SEL
+ pixel_9791/NB1 pixel_9791/VBIAS pixel_9791/NB2 pixel_9791/AMP_IN pixel_9791/SF_IB
+ pixel_9791/PIX_OUT pixel_9791/CSA_VREF pixel
Xpixel_509 pixel_509/gring pixel_509/VDD pixel_509/GND pixel_509/VREF pixel_509/ROW_SEL
+ pixel_509/NB1 pixel_509/VBIAS pixel_509/NB2 pixel_509/AMP_IN pixel_509/SF_IB pixel_509/PIX_OUT
+ pixel_509/CSA_VREF pixel
Xpixel_7107 pixel_7107/gring pixel_7107/VDD pixel_7107/GND pixel_7107/VREF pixel_7107/ROW_SEL
+ pixel_7107/NB1 pixel_7107/VBIAS pixel_7107/NB2 pixel_7107/AMP_IN pixel_7107/SF_IB
+ pixel_7107/PIX_OUT pixel_7107/CSA_VREF pixel
Xpixel_7118 pixel_7118/gring pixel_7118/VDD pixel_7118/GND pixel_7118/VREF pixel_7118/ROW_SEL
+ pixel_7118/NB1 pixel_7118/VBIAS pixel_7118/NB2 pixel_7118/AMP_IN pixel_7118/SF_IB
+ pixel_7118/PIX_OUT pixel_7118/CSA_VREF pixel
Xpixel_7129 pixel_7129/gring pixel_7129/VDD pixel_7129/GND pixel_7129/VREF pixel_7129/ROW_SEL
+ pixel_7129/NB1 pixel_7129/VBIAS pixel_7129/NB2 pixel_7129/AMP_IN pixel_7129/SF_IB
+ pixel_7129/PIX_OUT pixel_7129/CSA_VREF pixel
Xpixel_6406 pixel_6406/gring pixel_6406/VDD pixel_6406/GND pixel_6406/VREF pixel_6406/ROW_SEL
+ pixel_6406/NB1 pixel_6406/VBIAS pixel_6406/NB2 pixel_6406/AMP_IN pixel_6406/SF_IB
+ pixel_6406/PIX_OUT pixel_6406/CSA_VREF pixel
Xpixel_6417 pixel_6417/gring pixel_6417/VDD pixel_6417/GND pixel_6417/VREF pixel_6417/ROW_SEL
+ pixel_6417/NB1 pixel_6417/VBIAS pixel_6417/NB2 pixel_6417/AMP_IN pixel_6417/SF_IB
+ pixel_6417/PIX_OUT pixel_6417/CSA_VREF pixel
Xpixel_6428 pixel_6428/gring pixel_6428/VDD pixel_6428/GND pixel_6428/VREF pixel_6428/ROW_SEL
+ pixel_6428/NB1 pixel_6428/VBIAS pixel_6428/NB2 pixel_6428/AMP_IN pixel_6428/SF_IB
+ pixel_6428/PIX_OUT pixel_6428/CSA_VREF pixel
Xpixel_6439 pixel_6439/gring pixel_6439/VDD pixel_6439/GND pixel_6439/VREF pixel_6439/ROW_SEL
+ pixel_6439/NB1 pixel_6439/VBIAS pixel_6439/NB2 pixel_6439/AMP_IN pixel_6439/SF_IB
+ pixel_6439/PIX_OUT pixel_6439/CSA_VREF pixel
Xpixel_5705 pixel_5705/gring pixel_5705/VDD pixel_5705/GND pixel_5705/VREF pixel_5705/ROW_SEL
+ pixel_5705/NB1 pixel_5705/VBIAS pixel_5705/NB2 pixel_5705/AMP_IN pixel_5705/SF_IB
+ pixel_5705/PIX_OUT pixel_5705/CSA_VREF pixel
Xpixel_5716 pixel_5716/gring pixel_5716/VDD pixel_5716/GND pixel_5716/VREF pixel_5716/ROW_SEL
+ pixel_5716/NB1 pixel_5716/VBIAS pixel_5716/NB2 pixel_5716/AMP_IN pixel_5716/SF_IB
+ pixel_5716/PIX_OUT pixel_5716/CSA_VREF pixel
Xpixel_5727 pixel_5727/gring pixel_5727/VDD pixel_5727/GND pixel_5727/VREF pixel_5727/ROW_SEL
+ pixel_5727/NB1 pixel_5727/VBIAS pixel_5727/NB2 pixel_5727/AMP_IN pixel_5727/SF_IB
+ pixel_5727/PIX_OUT pixel_5727/CSA_VREF pixel
Xpixel_5738 pixel_5738/gring pixel_5738/VDD pixel_5738/GND pixel_5738/VREF pixel_5738/ROW_SEL
+ pixel_5738/NB1 pixel_5738/VBIAS pixel_5738/NB2 pixel_5738/AMP_IN pixel_5738/SF_IB
+ pixel_5738/PIX_OUT pixel_5738/CSA_VREF pixel
Xpixel_5749 pixel_5749/gring pixel_5749/VDD pixel_5749/GND pixel_5749/VREF pixel_5749/ROW_SEL
+ pixel_5749/NB1 pixel_5749/VBIAS pixel_5749/NB2 pixel_5749/AMP_IN pixel_5749/SF_IB
+ pixel_5749/PIX_OUT pixel_5749/CSA_VREF pixel
Xpixel_9021 pixel_9021/gring pixel_9021/VDD pixel_9021/GND pixel_9021/VREF pixel_9021/ROW_SEL
+ pixel_9021/NB1 pixel_9021/VBIAS pixel_9021/NB2 pixel_9021/AMP_IN pixel_9021/SF_IB
+ pixel_9021/PIX_OUT pixel_9021/CSA_VREF pixel
Xpixel_9010 pixel_9010/gring pixel_9010/VDD pixel_9010/GND pixel_9010/VREF pixel_9010/ROW_SEL
+ pixel_9010/NB1 pixel_9010/VBIAS pixel_9010/NB2 pixel_9010/AMP_IN pixel_9010/SF_IB
+ pixel_9010/PIX_OUT pixel_9010/CSA_VREF pixel
Xpixel_9054 pixel_9054/gring pixel_9054/VDD pixel_9054/GND pixel_9054/VREF pixel_9054/ROW_SEL
+ pixel_9054/NB1 pixel_9054/VBIAS pixel_9054/NB2 pixel_9054/AMP_IN pixel_9054/SF_IB
+ pixel_9054/PIX_OUT pixel_9054/CSA_VREF pixel
Xpixel_9043 pixel_9043/gring pixel_9043/VDD pixel_9043/GND pixel_9043/VREF pixel_9043/ROW_SEL
+ pixel_9043/NB1 pixel_9043/VBIAS pixel_9043/NB2 pixel_9043/AMP_IN pixel_9043/SF_IB
+ pixel_9043/PIX_OUT pixel_9043/CSA_VREF pixel
Xpixel_9032 pixel_9032/gring pixel_9032/VDD pixel_9032/GND pixel_9032/VREF pixel_9032/ROW_SEL
+ pixel_9032/NB1 pixel_9032/VBIAS pixel_9032/NB2 pixel_9032/AMP_IN pixel_9032/SF_IB
+ pixel_9032/PIX_OUT pixel_9032/CSA_VREF pixel
Xpixel_9098 pixel_9098/gring pixel_9098/VDD pixel_9098/GND pixel_9098/VREF pixel_9098/ROW_SEL
+ pixel_9098/NB1 pixel_9098/VBIAS pixel_9098/NB2 pixel_9098/AMP_IN pixel_9098/SF_IB
+ pixel_9098/PIX_OUT pixel_9098/CSA_VREF pixel
Xpixel_9087 pixel_9087/gring pixel_9087/VDD pixel_9087/GND pixel_9087/VREF pixel_9087/ROW_SEL
+ pixel_9087/NB1 pixel_9087/VBIAS pixel_9087/NB2 pixel_9087/AMP_IN pixel_9087/SF_IB
+ pixel_9087/PIX_OUT pixel_9087/CSA_VREF pixel
Xpixel_9076 pixel_9076/gring pixel_9076/VDD pixel_9076/GND pixel_9076/VREF pixel_9076/ROW_SEL
+ pixel_9076/NB1 pixel_9076/VBIAS pixel_9076/NB2 pixel_9076/AMP_IN pixel_9076/SF_IB
+ pixel_9076/PIX_OUT pixel_9076/CSA_VREF pixel
Xpixel_9065 pixel_9065/gring pixel_9065/VDD pixel_9065/GND pixel_9065/VREF pixel_9065/ROW_SEL
+ pixel_9065/NB1 pixel_9065/VBIAS pixel_9065/NB2 pixel_9065/AMP_IN pixel_9065/SF_IB
+ pixel_9065/PIX_OUT pixel_9065/CSA_VREF pixel
Xpixel_8320 pixel_8320/gring pixel_8320/VDD pixel_8320/GND pixel_8320/VREF pixel_8320/ROW_SEL
+ pixel_8320/NB1 pixel_8320/VBIAS pixel_8320/NB2 pixel_8320/AMP_IN pixel_8320/SF_IB
+ pixel_8320/PIX_OUT pixel_8320/CSA_VREF pixel
Xpixel_8331 pixel_8331/gring pixel_8331/VDD pixel_8331/GND pixel_8331/VREF pixel_8331/ROW_SEL
+ pixel_8331/NB1 pixel_8331/VBIAS pixel_8331/NB2 pixel_8331/AMP_IN pixel_8331/SF_IB
+ pixel_8331/PIX_OUT pixel_8331/CSA_VREF pixel
Xpixel_8342 pixel_8342/gring pixel_8342/VDD pixel_8342/GND pixel_8342/VREF pixel_8342/ROW_SEL
+ pixel_8342/NB1 pixel_8342/VBIAS pixel_8342/NB2 pixel_8342/AMP_IN pixel_8342/SF_IB
+ pixel_8342/PIX_OUT pixel_8342/CSA_VREF pixel
Xpixel_8353 pixel_8353/gring pixel_8353/VDD pixel_8353/GND pixel_8353/VREF pixel_8353/ROW_SEL
+ pixel_8353/NB1 pixel_8353/VBIAS pixel_8353/NB2 pixel_8353/AMP_IN pixel_8353/SF_IB
+ pixel_8353/PIX_OUT pixel_8353/CSA_VREF pixel
Xpixel_8364 pixel_8364/gring pixel_8364/VDD pixel_8364/GND pixel_8364/VREF pixel_8364/ROW_SEL
+ pixel_8364/NB1 pixel_8364/VBIAS pixel_8364/NB2 pixel_8364/AMP_IN pixel_8364/SF_IB
+ pixel_8364/PIX_OUT pixel_8364/CSA_VREF pixel
Xpixel_8375 pixel_8375/gring pixel_8375/VDD pixel_8375/GND pixel_8375/VREF pixel_8375/ROW_SEL
+ pixel_8375/NB1 pixel_8375/VBIAS pixel_8375/NB2 pixel_8375/AMP_IN pixel_8375/SF_IB
+ pixel_8375/PIX_OUT pixel_8375/CSA_VREF pixel
Xpixel_8386 pixel_8386/gring pixel_8386/VDD pixel_8386/GND pixel_8386/VREF pixel_8386/ROW_SEL
+ pixel_8386/NB1 pixel_8386/VBIAS pixel_8386/NB2 pixel_8386/AMP_IN pixel_8386/SF_IB
+ pixel_8386/PIX_OUT pixel_8386/CSA_VREF pixel
Xpixel_7630 pixel_7630/gring pixel_7630/VDD pixel_7630/GND pixel_7630/VREF pixel_7630/ROW_SEL
+ pixel_7630/NB1 pixel_7630/VBIAS pixel_7630/NB2 pixel_7630/AMP_IN pixel_7630/SF_IB
+ pixel_7630/PIX_OUT pixel_7630/CSA_VREF pixel
Xpixel_7641 pixel_7641/gring pixel_7641/VDD pixel_7641/GND pixel_7641/VREF pixel_7641/ROW_SEL
+ pixel_7641/NB1 pixel_7641/VBIAS pixel_7641/NB2 pixel_7641/AMP_IN pixel_7641/SF_IB
+ pixel_7641/PIX_OUT pixel_7641/CSA_VREF pixel
Xpixel_8397 pixel_8397/gring pixel_8397/VDD pixel_8397/GND pixel_8397/VREF pixel_8397/ROW_SEL
+ pixel_8397/NB1 pixel_8397/VBIAS pixel_8397/NB2 pixel_8397/AMP_IN pixel_8397/SF_IB
+ pixel_8397/PIX_OUT pixel_8397/CSA_VREF pixel
Xpixel_7652 pixel_7652/gring pixel_7652/VDD pixel_7652/GND pixel_7652/VREF pixel_7652/ROW_SEL
+ pixel_7652/NB1 pixel_7652/VBIAS pixel_7652/NB2 pixel_7652/AMP_IN pixel_7652/SF_IB
+ pixel_7652/PIX_OUT pixel_7652/CSA_VREF pixel
Xpixel_7663 pixel_7663/gring pixel_7663/VDD pixel_7663/GND pixel_7663/VREF pixel_7663/ROW_SEL
+ pixel_7663/NB1 pixel_7663/VBIAS pixel_7663/NB2 pixel_7663/AMP_IN pixel_7663/SF_IB
+ pixel_7663/PIX_OUT pixel_7663/CSA_VREF pixel
Xpixel_7674 pixel_7674/gring pixel_7674/VDD pixel_7674/GND pixel_7674/VREF pixel_7674/ROW_SEL
+ pixel_7674/NB1 pixel_7674/VBIAS pixel_7674/NB2 pixel_7674/AMP_IN pixel_7674/SF_IB
+ pixel_7674/PIX_OUT pixel_7674/CSA_VREF pixel
Xpixel_7685 pixel_7685/gring pixel_7685/VDD pixel_7685/GND pixel_7685/VREF pixel_7685/ROW_SEL
+ pixel_7685/NB1 pixel_7685/VBIAS pixel_7685/NB2 pixel_7685/AMP_IN pixel_7685/SF_IB
+ pixel_7685/PIX_OUT pixel_7685/CSA_VREF pixel
Xpixel_6940 pixel_6940/gring pixel_6940/VDD pixel_6940/GND pixel_6940/VREF pixel_6940/ROW_SEL
+ pixel_6940/NB1 pixel_6940/VBIAS pixel_6940/NB2 pixel_6940/AMP_IN pixel_6940/SF_IB
+ pixel_6940/PIX_OUT pixel_6940/CSA_VREF pixel
Xpixel_21 pixel_21/gring pixel_21/VDD pixel_21/GND pixel_21/VREF pixel_21/ROW_SEL
+ pixel_21/NB1 pixel_21/VBIAS pixel_21/NB2 pixel_21/AMP_IN pixel_21/SF_IB pixel_21/PIX_OUT
+ pixel_21/CSA_VREF pixel
Xpixel_10 pixel_10/gring pixel_10/VDD pixel_10/GND pixel_10/VREF pixel_10/ROW_SEL
+ pixel_10/NB1 pixel_10/VBIAS pixel_10/NB2 pixel_10/AMP_IN pixel_10/SF_IB pixel_10/PIX_OUT
+ pixel_10/CSA_VREF pixel
Xpixel_7696 pixel_7696/gring pixel_7696/VDD pixel_7696/GND pixel_7696/VREF pixel_7696/ROW_SEL
+ pixel_7696/NB1 pixel_7696/VBIAS pixel_7696/NB2 pixel_7696/AMP_IN pixel_7696/SF_IB
+ pixel_7696/PIX_OUT pixel_7696/CSA_VREF pixel
Xpixel_6951 pixel_6951/gring pixel_6951/VDD pixel_6951/GND pixel_6951/VREF pixel_6951/ROW_SEL
+ pixel_6951/NB1 pixel_6951/VBIAS pixel_6951/NB2 pixel_6951/AMP_IN pixel_6951/SF_IB
+ pixel_6951/PIX_OUT pixel_6951/CSA_VREF pixel
Xpixel_6962 pixel_6962/gring pixel_6962/VDD pixel_6962/GND pixel_6962/VREF pixel_6962/ROW_SEL
+ pixel_6962/NB1 pixel_6962/VBIAS pixel_6962/NB2 pixel_6962/AMP_IN pixel_6962/SF_IB
+ pixel_6962/PIX_OUT pixel_6962/CSA_VREF pixel
Xpixel_6973 pixel_6973/gring pixel_6973/VDD pixel_6973/GND pixel_6973/VREF pixel_6973/ROW_SEL
+ pixel_6973/NB1 pixel_6973/VBIAS pixel_6973/NB2 pixel_6973/AMP_IN pixel_6973/SF_IB
+ pixel_6973/PIX_OUT pixel_6973/CSA_VREF pixel
Xpixel_54 pixel_54/gring pixel_54/VDD pixel_54/GND pixel_54/VREF pixel_54/ROW_SEL
+ pixel_54/NB1 pixel_54/VBIAS pixel_54/NB2 pixel_54/AMP_IN pixel_54/SF_IB pixel_54/PIX_OUT
+ pixel_54/CSA_VREF pixel
Xpixel_43 pixel_43/gring pixel_43/VDD pixel_43/GND pixel_43/VREF pixel_43/ROW_SEL
+ pixel_43/NB1 pixel_43/VBIAS pixel_43/NB2 pixel_43/AMP_IN pixel_43/SF_IB pixel_43/PIX_OUT
+ pixel_43/CSA_VREF pixel
Xpixel_32 pixel_32/gring pixel_32/VDD pixel_32/GND pixel_32/VREF pixel_32/ROW_SEL
+ pixel_32/NB1 pixel_32/VBIAS pixel_32/NB2 pixel_32/AMP_IN pixel_32/SF_IB pixel_32/PIX_OUT
+ pixel_32/CSA_VREF pixel
Xpixel_6984 pixel_6984/gring pixel_6984/VDD pixel_6984/GND pixel_6984/VREF pixel_6984/ROW_SEL
+ pixel_6984/NB1 pixel_6984/VBIAS pixel_6984/NB2 pixel_6984/AMP_IN pixel_6984/SF_IB
+ pixel_6984/PIX_OUT pixel_6984/CSA_VREF pixel
Xpixel_6995 pixel_6995/gring pixel_6995/VDD pixel_6995/GND pixel_6995/VREF pixel_6995/ROW_SEL
+ pixel_6995/NB1 pixel_6995/VBIAS pixel_6995/NB2 pixel_6995/AMP_IN pixel_6995/SF_IB
+ pixel_6995/PIX_OUT pixel_6995/CSA_VREF pixel
Xpixel_87 pixel_87/gring pixel_87/VDD pixel_87/GND pixel_87/VREF pixel_87/ROW_SEL
+ pixel_87/NB1 pixel_87/VBIAS pixel_87/NB2 pixel_87/AMP_IN pixel_87/SF_IB pixel_87/PIX_OUT
+ pixel_87/CSA_VREF pixel
Xpixel_76 pixel_76/gring pixel_76/VDD pixel_76/GND pixel_76/VREF pixel_76/ROW_SEL
+ pixel_76/NB1 pixel_76/VBIAS pixel_76/NB2 pixel_76/AMP_IN pixel_76/SF_IB pixel_76/PIX_OUT
+ pixel_76/CSA_VREF pixel
Xpixel_65 pixel_65/gring pixel_65/VDD pixel_65/GND pixel_65/VREF pixel_65/ROW_SEL
+ pixel_65/NB1 pixel_65/VBIAS pixel_65/NB2 pixel_65/AMP_IN pixel_65/SF_IB pixel_65/PIX_OUT
+ pixel_65/CSA_VREF pixel
Xpixel_98 pixel_98/gring pixel_98/VDD pixel_98/GND pixel_98/VREF pixel_98/ROW_SEL
+ pixel_98/NB1 pixel_98/VBIAS pixel_98/NB2 pixel_98/AMP_IN pixel_98/SF_IB pixel_98/PIX_OUT
+ pixel_98/CSA_VREF pixel
Xpixel_1291 pixel_1291/gring pixel_1291/VDD pixel_1291/GND pixel_1291/VREF pixel_1291/ROW_SEL
+ pixel_1291/NB1 pixel_1291/VBIAS pixel_1291/NB2 pixel_1291/AMP_IN pixel_1291/SF_IB
+ pixel_1291/PIX_OUT pixel_1291/CSA_VREF pixel
Xpixel_1280 pixel_1280/gring pixel_1280/VDD pixel_1280/GND pixel_1280/VREF pixel_1280/ROW_SEL
+ pixel_1280/NB1 pixel_1280/VBIAS pixel_1280/NB2 pixel_1280/AMP_IN pixel_1280/SF_IB
+ pixel_1280/PIX_OUT pixel_1280/CSA_VREF pixel
Xpixel_328 pixel_328/gring pixel_328/VDD pixel_328/GND pixel_328/VREF pixel_328/ROW_SEL
+ pixel_328/NB1 pixel_328/VBIAS pixel_328/NB2 pixel_328/AMP_IN pixel_328/SF_IB pixel_328/PIX_OUT
+ pixel_328/CSA_VREF pixel
Xpixel_317 pixel_317/gring pixel_317/VDD pixel_317/GND pixel_317/VREF pixel_317/ROW_SEL
+ pixel_317/NB1 pixel_317/VBIAS pixel_317/NB2 pixel_317/AMP_IN pixel_317/SF_IB pixel_317/PIX_OUT
+ pixel_317/CSA_VREF pixel
Xpixel_306 pixel_306/gring pixel_306/VDD pixel_306/GND pixel_306/VREF pixel_306/ROW_SEL
+ pixel_306/NB1 pixel_306/VBIAS pixel_306/NB2 pixel_306/AMP_IN pixel_306/SF_IB pixel_306/PIX_OUT
+ pixel_306/CSA_VREF pixel
Xpixel_339 pixel_339/gring pixel_339/VDD pixel_339/GND pixel_339/VREF pixel_339/ROW_SEL
+ pixel_339/NB1 pixel_339/VBIAS pixel_339/NB2 pixel_339/AMP_IN pixel_339/SF_IB pixel_339/PIX_OUT
+ pixel_339/CSA_VREF pixel
Xpixel_2909 pixel_2909/gring pixel_2909/VDD pixel_2909/GND pixel_2909/VREF pixel_2909/ROW_SEL
+ pixel_2909/NB1 pixel_2909/VBIAS pixel_2909/NB2 pixel_2909/AMP_IN pixel_2909/SF_IB
+ pixel_2909/PIX_OUT pixel_2909/CSA_VREF pixel
Xpixel_6203 pixel_6203/gring pixel_6203/VDD pixel_6203/GND pixel_6203/VREF pixel_6203/ROW_SEL
+ pixel_6203/NB1 pixel_6203/VBIAS pixel_6203/NB2 pixel_6203/AMP_IN pixel_6203/SF_IB
+ pixel_6203/PIX_OUT pixel_6203/CSA_VREF pixel
Xpixel_6214 pixel_6214/gring pixel_6214/VDD pixel_6214/GND pixel_6214/VREF pixel_6214/ROW_SEL
+ pixel_6214/NB1 pixel_6214/VBIAS pixel_6214/NB2 pixel_6214/AMP_IN pixel_6214/SF_IB
+ pixel_6214/PIX_OUT pixel_6214/CSA_VREF pixel
Xpixel_6225 pixel_6225/gring pixel_6225/VDD pixel_6225/GND pixel_6225/VREF pixel_6225/ROW_SEL
+ pixel_6225/NB1 pixel_6225/VBIAS pixel_6225/NB2 pixel_6225/AMP_IN pixel_6225/SF_IB
+ pixel_6225/PIX_OUT pixel_6225/CSA_VREF pixel
Xpixel_6236 pixel_6236/gring pixel_6236/VDD pixel_6236/GND pixel_6236/VREF pixel_6236/ROW_SEL
+ pixel_6236/NB1 pixel_6236/VBIAS pixel_6236/NB2 pixel_6236/AMP_IN pixel_6236/SF_IB
+ pixel_6236/PIX_OUT pixel_6236/CSA_VREF pixel
Xpixel_6247 pixel_6247/gring pixel_6247/VDD pixel_6247/GND pixel_6247/VREF pixel_6247/ROW_SEL
+ pixel_6247/NB1 pixel_6247/VBIAS pixel_6247/NB2 pixel_6247/AMP_IN pixel_6247/SF_IB
+ pixel_6247/PIX_OUT pixel_6247/CSA_VREF pixel
Xpixel_6258 pixel_6258/gring pixel_6258/VDD pixel_6258/GND pixel_6258/VREF pixel_6258/ROW_SEL
+ pixel_6258/NB1 pixel_6258/VBIAS pixel_6258/NB2 pixel_6258/AMP_IN pixel_6258/SF_IB
+ pixel_6258/PIX_OUT pixel_6258/CSA_VREF pixel
Xpixel_6269 pixel_6269/gring pixel_6269/VDD pixel_6269/GND pixel_6269/VREF pixel_6269/ROW_SEL
+ pixel_6269/NB1 pixel_6269/VBIAS pixel_6269/NB2 pixel_6269/AMP_IN pixel_6269/SF_IB
+ pixel_6269/PIX_OUT pixel_6269/CSA_VREF pixel
Xpixel_5502 pixel_5502/gring pixel_5502/VDD pixel_5502/GND pixel_5502/VREF pixel_5502/ROW_SEL
+ pixel_5502/NB1 pixel_5502/VBIAS pixel_5502/NB2 pixel_5502/AMP_IN pixel_5502/SF_IB
+ pixel_5502/PIX_OUT pixel_5502/CSA_VREF pixel
Xpixel_5513 pixel_5513/gring pixel_5513/VDD pixel_5513/GND pixel_5513/VREF pixel_5513/ROW_SEL
+ pixel_5513/NB1 pixel_5513/VBIAS pixel_5513/NB2 pixel_5513/AMP_IN pixel_5513/SF_IB
+ pixel_5513/PIX_OUT pixel_5513/CSA_VREF pixel
Xpixel_5524 pixel_5524/gring pixel_5524/VDD pixel_5524/GND pixel_5524/VREF pixel_5524/ROW_SEL
+ pixel_5524/NB1 pixel_5524/VBIAS pixel_5524/NB2 pixel_5524/AMP_IN pixel_5524/SF_IB
+ pixel_5524/PIX_OUT pixel_5524/CSA_VREF pixel
Xpixel_5535 pixel_5535/gring pixel_5535/VDD pixel_5535/GND pixel_5535/VREF pixel_5535/ROW_SEL
+ pixel_5535/NB1 pixel_5535/VBIAS pixel_5535/NB2 pixel_5535/AMP_IN pixel_5535/SF_IB
+ pixel_5535/PIX_OUT pixel_5535/CSA_VREF pixel
Xpixel_5546 pixel_5546/gring pixel_5546/VDD pixel_5546/GND pixel_5546/VREF pixel_5546/ROW_SEL
+ pixel_5546/NB1 pixel_5546/VBIAS pixel_5546/NB2 pixel_5546/AMP_IN pixel_5546/SF_IB
+ pixel_5546/PIX_OUT pixel_5546/CSA_VREF pixel
Xpixel_5557 pixel_5557/gring pixel_5557/VDD pixel_5557/GND pixel_5557/VREF pixel_5557/ROW_SEL
+ pixel_5557/NB1 pixel_5557/VBIAS pixel_5557/NB2 pixel_5557/AMP_IN pixel_5557/SF_IB
+ pixel_5557/PIX_OUT pixel_5557/CSA_VREF pixel
Xpixel_4801 pixel_4801/gring pixel_4801/VDD pixel_4801/GND pixel_4801/VREF pixel_4801/ROW_SEL
+ pixel_4801/NB1 pixel_4801/VBIAS pixel_4801/NB2 pixel_4801/AMP_IN pixel_4801/SF_IB
+ pixel_4801/PIX_OUT pixel_4801/CSA_VREF pixel
Xpixel_4812 pixel_4812/gring pixel_4812/VDD pixel_4812/GND pixel_4812/VREF pixel_4812/ROW_SEL
+ pixel_4812/NB1 pixel_4812/VBIAS pixel_4812/NB2 pixel_4812/AMP_IN pixel_4812/SF_IB
+ pixel_4812/PIX_OUT pixel_4812/CSA_VREF pixel
Xpixel_851 pixel_851/gring pixel_851/VDD pixel_851/GND pixel_851/VREF pixel_851/ROW_SEL
+ pixel_851/NB1 pixel_851/VBIAS pixel_851/NB2 pixel_851/AMP_IN pixel_851/SF_IB pixel_851/PIX_OUT
+ pixel_851/CSA_VREF pixel
Xpixel_840 pixel_840/gring pixel_840/VDD pixel_840/GND pixel_840/VREF pixel_840/ROW_SEL
+ pixel_840/NB1 pixel_840/VBIAS pixel_840/NB2 pixel_840/AMP_IN pixel_840/SF_IB pixel_840/PIX_OUT
+ pixel_840/CSA_VREF pixel
Xpixel_5568 pixel_5568/gring pixel_5568/VDD pixel_5568/GND pixel_5568/VREF pixel_5568/ROW_SEL
+ pixel_5568/NB1 pixel_5568/VBIAS pixel_5568/NB2 pixel_5568/AMP_IN pixel_5568/SF_IB
+ pixel_5568/PIX_OUT pixel_5568/CSA_VREF pixel
Xpixel_5579 pixel_5579/gring pixel_5579/VDD pixel_5579/GND pixel_5579/VREF pixel_5579/ROW_SEL
+ pixel_5579/NB1 pixel_5579/VBIAS pixel_5579/NB2 pixel_5579/AMP_IN pixel_5579/SF_IB
+ pixel_5579/PIX_OUT pixel_5579/CSA_VREF pixel
Xpixel_4823 pixel_4823/gring pixel_4823/VDD pixel_4823/GND pixel_4823/VREF pixel_4823/ROW_SEL
+ pixel_4823/NB1 pixel_4823/VBIAS pixel_4823/NB2 pixel_4823/AMP_IN pixel_4823/SF_IB
+ pixel_4823/PIX_OUT pixel_4823/CSA_VREF pixel
Xpixel_4834 pixel_4834/gring pixel_4834/VDD pixel_4834/GND pixel_4834/VREF pixel_4834/ROW_SEL
+ pixel_4834/NB1 pixel_4834/VBIAS pixel_4834/NB2 pixel_4834/AMP_IN pixel_4834/SF_IB
+ pixel_4834/PIX_OUT pixel_4834/CSA_VREF pixel
Xpixel_4845 pixel_4845/gring pixel_4845/VDD pixel_4845/GND pixel_4845/VREF pixel_4845/ROW_SEL
+ pixel_4845/NB1 pixel_4845/VBIAS pixel_4845/NB2 pixel_4845/AMP_IN pixel_4845/SF_IB
+ pixel_4845/PIX_OUT pixel_4845/CSA_VREF pixel
Xpixel_4856 pixel_4856/gring pixel_4856/VDD pixel_4856/GND pixel_4856/VREF pixel_4856/ROW_SEL
+ pixel_4856/NB1 pixel_4856/VBIAS pixel_4856/NB2 pixel_4856/AMP_IN pixel_4856/SF_IB
+ pixel_4856/PIX_OUT pixel_4856/CSA_VREF pixel
Xpixel_884 pixel_884/gring pixel_884/VDD pixel_884/GND pixel_884/VREF pixel_884/ROW_SEL
+ pixel_884/NB1 pixel_884/VBIAS pixel_884/NB2 pixel_884/AMP_IN pixel_884/SF_IB pixel_884/PIX_OUT
+ pixel_884/CSA_VREF pixel
Xpixel_873 pixel_873/gring pixel_873/VDD pixel_873/GND pixel_873/VREF pixel_873/ROW_SEL
+ pixel_873/NB1 pixel_873/VBIAS pixel_873/NB2 pixel_873/AMP_IN pixel_873/SF_IB pixel_873/PIX_OUT
+ pixel_873/CSA_VREF pixel
Xpixel_862 pixel_862/gring pixel_862/VDD pixel_862/GND pixel_862/VREF pixel_862/ROW_SEL
+ pixel_862/NB1 pixel_862/VBIAS pixel_862/NB2 pixel_862/AMP_IN pixel_862/SF_IB pixel_862/PIX_OUT
+ pixel_862/CSA_VREF pixel
Xpixel_4867 pixel_4867/gring pixel_4867/VDD pixel_4867/GND pixel_4867/VREF pixel_4867/ROW_SEL
+ pixel_4867/NB1 pixel_4867/VBIAS pixel_4867/NB2 pixel_4867/AMP_IN pixel_4867/SF_IB
+ pixel_4867/PIX_OUT pixel_4867/CSA_VREF pixel
Xpixel_4878 pixel_4878/gring pixel_4878/VDD pixel_4878/GND pixel_4878/VREF pixel_4878/ROW_SEL
+ pixel_4878/NB1 pixel_4878/VBIAS pixel_4878/NB2 pixel_4878/AMP_IN pixel_4878/SF_IB
+ pixel_4878/PIX_OUT pixel_4878/CSA_VREF pixel
Xpixel_4889 pixel_4889/gring pixel_4889/VDD pixel_4889/GND pixel_4889/VREF pixel_4889/ROW_SEL
+ pixel_4889/NB1 pixel_4889/VBIAS pixel_4889/NB2 pixel_4889/AMP_IN pixel_4889/SF_IB
+ pixel_4889/PIX_OUT pixel_4889/CSA_VREF pixel
Xpixel_895 pixel_895/gring pixel_895/VDD pixel_895/GND pixel_895/VREF pixel_895/ROW_SEL
+ pixel_895/NB1 pixel_895/VBIAS pixel_895/NB2 pixel_895/AMP_IN pixel_895/SF_IB pixel_895/PIX_OUT
+ pixel_895/CSA_VREF pixel
Xpixel_8150 pixel_8150/gring pixel_8150/VDD pixel_8150/GND pixel_8150/VREF pixel_8150/ROW_SEL
+ pixel_8150/NB1 pixel_8150/VBIAS pixel_8150/NB2 pixel_8150/AMP_IN pixel_8150/SF_IB
+ pixel_8150/PIX_OUT pixel_8150/CSA_VREF pixel
Xpixel_8161 pixel_8161/gring pixel_8161/VDD pixel_8161/GND pixel_8161/VREF pixel_8161/ROW_SEL
+ pixel_8161/NB1 pixel_8161/VBIAS pixel_8161/NB2 pixel_8161/AMP_IN pixel_8161/SF_IB
+ pixel_8161/PIX_OUT pixel_8161/CSA_VREF pixel
Xpixel_8172 pixel_8172/gring pixel_8172/VDD pixel_8172/GND pixel_8172/VREF pixel_8172/ROW_SEL
+ pixel_8172/NB1 pixel_8172/VBIAS pixel_8172/NB2 pixel_8172/AMP_IN pixel_8172/SF_IB
+ pixel_8172/PIX_OUT pixel_8172/CSA_VREF pixel
Xpixel_8183 pixel_8183/gring pixel_8183/VDD pixel_8183/GND pixel_8183/VREF pixel_8183/ROW_SEL
+ pixel_8183/NB1 pixel_8183/VBIAS pixel_8183/NB2 pixel_8183/AMP_IN pixel_8183/SF_IB
+ pixel_8183/PIX_OUT pixel_8183/CSA_VREF pixel
Xpixel_8194 pixel_8194/gring pixel_8194/VDD pixel_8194/GND pixel_8194/VREF pixel_8194/ROW_SEL
+ pixel_8194/NB1 pixel_8194/VBIAS pixel_8194/NB2 pixel_8194/AMP_IN pixel_8194/SF_IB
+ pixel_8194/PIX_OUT pixel_8194/CSA_VREF pixel
Xpixel_7460 pixel_7460/gring pixel_7460/VDD pixel_7460/GND pixel_7460/VREF pixel_7460/ROW_SEL
+ pixel_7460/NB1 pixel_7460/VBIAS pixel_7460/NB2 pixel_7460/AMP_IN pixel_7460/SF_IB
+ pixel_7460/PIX_OUT pixel_7460/CSA_VREF pixel
Xpixel_7471 pixel_7471/gring pixel_7471/VDD pixel_7471/GND pixel_7471/VREF pixel_7471/ROW_SEL
+ pixel_7471/NB1 pixel_7471/VBIAS pixel_7471/NB2 pixel_7471/AMP_IN pixel_7471/SF_IB
+ pixel_7471/PIX_OUT pixel_7471/CSA_VREF pixel
Xpixel_7482 pixel_7482/gring pixel_7482/VDD pixel_7482/GND pixel_7482/VREF pixel_7482/ROW_SEL
+ pixel_7482/NB1 pixel_7482/VBIAS pixel_7482/NB2 pixel_7482/AMP_IN pixel_7482/SF_IB
+ pixel_7482/PIX_OUT pixel_7482/CSA_VREF pixel
Xpixel_7493 pixel_7493/gring pixel_7493/VDD pixel_7493/GND pixel_7493/VREF pixel_7493/ROW_SEL
+ pixel_7493/NB1 pixel_7493/VBIAS pixel_7493/NB2 pixel_7493/AMP_IN pixel_7493/SF_IB
+ pixel_7493/PIX_OUT pixel_7493/CSA_VREF pixel
Xpixel_6770 pixel_6770/gring pixel_6770/VDD pixel_6770/GND pixel_6770/VREF pixel_6770/ROW_SEL
+ pixel_6770/NB1 pixel_6770/VBIAS pixel_6770/NB2 pixel_6770/AMP_IN pixel_6770/SF_IB
+ pixel_6770/PIX_OUT pixel_6770/CSA_VREF pixel
Xpixel_6781 pixel_6781/gring pixel_6781/VDD pixel_6781/GND pixel_6781/VREF pixel_6781/ROW_SEL
+ pixel_6781/NB1 pixel_6781/VBIAS pixel_6781/NB2 pixel_6781/AMP_IN pixel_6781/SF_IB
+ pixel_6781/PIX_OUT pixel_6781/CSA_VREF pixel
Xpixel_6792 pixel_6792/gring pixel_6792/VDD pixel_6792/GND pixel_6792/VREF pixel_6792/ROW_SEL
+ pixel_6792/NB1 pixel_6792/VBIAS pixel_6792/NB2 pixel_6792/AMP_IN pixel_6792/SF_IB
+ pixel_6792/PIX_OUT pixel_6792/CSA_VREF pixel
Xpixel_103 pixel_103/gring pixel_103/VDD pixel_103/GND pixel_103/VREF pixel_103/ROW_SEL
+ pixel_103/NB1 pixel_103/VBIAS pixel_103/NB2 pixel_103/AMP_IN pixel_103/SF_IB pixel_103/PIX_OUT
+ pixel_103/CSA_VREF pixel
Xpixel_4108 pixel_4108/gring pixel_4108/VDD pixel_4108/GND pixel_4108/VREF pixel_4108/ROW_SEL
+ pixel_4108/NB1 pixel_4108/VBIAS pixel_4108/NB2 pixel_4108/AMP_IN pixel_4108/SF_IB
+ pixel_4108/PIX_OUT pixel_4108/CSA_VREF pixel
Xpixel_136 pixel_136/gring pixel_136/VDD pixel_136/GND pixel_136/VREF pixel_136/ROW_SEL
+ pixel_136/NB1 pixel_136/VBIAS pixel_136/NB2 pixel_136/AMP_IN pixel_136/SF_IB pixel_136/PIX_OUT
+ pixel_136/CSA_VREF pixel
Xpixel_125 pixel_125/gring pixel_125/VDD pixel_125/GND pixel_125/VREF pixel_125/ROW_SEL
+ pixel_125/NB1 pixel_125/VBIAS pixel_125/NB2 pixel_125/AMP_IN pixel_125/SF_IB pixel_125/PIX_OUT
+ pixel_125/CSA_VREF pixel
Xpixel_114 pixel_114/gring pixel_114/VDD pixel_114/GND pixel_114/VREF pixel_114/ROW_SEL
+ pixel_114/NB1 pixel_114/VBIAS pixel_114/NB2 pixel_114/AMP_IN pixel_114/SF_IB pixel_114/PIX_OUT
+ pixel_114/CSA_VREF pixel
Xpixel_4119 pixel_4119/gring pixel_4119/VDD pixel_4119/GND pixel_4119/VREF pixel_4119/ROW_SEL
+ pixel_4119/NB1 pixel_4119/VBIAS pixel_4119/NB2 pixel_4119/AMP_IN pixel_4119/SF_IB
+ pixel_4119/PIX_OUT pixel_4119/CSA_VREF pixel
Xpixel_169 pixel_169/gring pixel_169/VDD pixel_169/GND pixel_169/VREF pixel_169/ROW_SEL
+ pixel_169/NB1 pixel_169/VBIAS pixel_169/NB2 pixel_169/AMP_IN pixel_169/SF_IB pixel_169/PIX_OUT
+ pixel_169/CSA_VREF pixel
Xpixel_158 pixel_158/gring pixel_158/VDD pixel_158/GND pixel_158/VREF pixel_158/ROW_SEL
+ pixel_158/NB1 pixel_158/VBIAS pixel_158/NB2 pixel_158/AMP_IN pixel_158/SF_IB pixel_158/PIX_OUT
+ pixel_158/CSA_VREF pixel
Xpixel_147 pixel_147/gring pixel_147/VDD pixel_147/GND pixel_147/VREF pixel_147/ROW_SEL
+ pixel_147/NB1 pixel_147/VBIAS pixel_147/NB2 pixel_147/AMP_IN pixel_147/SF_IB pixel_147/PIX_OUT
+ pixel_147/CSA_VREF pixel
Xpixel_3429 pixel_3429/gring pixel_3429/VDD pixel_3429/GND pixel_3429/VREF pixel_3429/ROW_SEL
+ pixel_3429/NB1 pixel_3429/VBIAS pixel_3429/NB2 pixel_3429/AMP_IN pixel_3429/SF_IB
+ pixel_3429/PIX_OUT pixel_3429/CSA_VREF pixel
Xpixel_3418 pixel_3418/gring pixel_3418/VDD pixel_3418/GND pixel_3418/VREF pixel_3418/ROW_SEL
+ pixel_3418/NB1 pixel_3418/VBIAS pixel_3418/NB2 pixel_3418/AMP_IN pixel_3418/SF_IB
+ pixel_3418/PIX_OUT pixel_3418/CSA_VREF pixel
Xpixel_3407 pixel_3407/gring pixel_3407/VDD pixel_3407/GND pixel_3407/VREF pixel_3407/ROW_SEL
+ pixel_3407/NB1 pixel_3407/VBIAS pixel_3407/NB2 pixel_3407/AMP_IN pixel_3407/SF_IB
+ pixel_3407/PIX_OUT pixel_3407/CSA_VREF pixel
Xpixel_2728 pixel_2728/gring pixel_2728/VDD pixel_2728/GND pixel_2728/VREF pixel_2728/ROW_SEL
+ pixel_2728/NB1 pixel_2728/VBIAS pixel_2728/NB2 pixel_2728/AMP_IN pixel_2728/SF_IB
+ pixel_2728/PIX_OUT pixel_2728/CSA_VREF pixel
Xpixel_2717 pixel_2717/gring pixel_2717/VDD pixel_2717/GND pixel_2717/VREF pixel_2717/ROW_SEL
+ pixel_2717/NB1 pixel_2717/VBIAS pixel_2717/NB2 pixel_2717/AMP_IN pixel_2717/SF_IB
+ pixel_2717/PIX_OUT pixel_2717/CSA_VREF pixel
Xpixel_2706 pixel_2706/gring pixel_2706/VDD pixel_2706/GND pixel_2706/VREF pixel_2706/ROW_SEL
+ pixel_2706/NB1 pixel_2706/VBIAS pixel_2706/NB2 pixel_2706/AMP_IN pixel_2706/SF_IB
+ pixel_2706/PIX_OUT pixel_2706/CSA_VREF pixel
Xpixel_2739 pixel_2739/gring pixel_2739/VDD pixel_2739/GND pixel_2739/VREF pixel_2739/ROW_SEL
+ pixel_2739/NB1 pixel_2739/VBIAS pixel_2739/NB2 pixel_2739/AMP_IN pixel_2739/SF_IB
+ pixel_2739/PIX_OUT pixel_2739/CSA_VREF pixel
Xpixel_6000 pixel_6000/gring pixel_6000/VDD pixel_6000/GND pixel_6000/VREF pixel_6000/ROW_SEL
+ pixel_6000/NB1 pixel_6000/VBIAS pixel_6000/NB2 pixel_6000/AMP_IN pixel_6000/SF_IB
+ pixel_6000/PIX_OUT pixel_6000/CSA_VREF pixel
Xpixel_6011 pixel_6011/gring pixel_6011/VDD pixel_6011/GND pixel_6011/VREF pixel_6011/ROW_SEL
+ pixel_6011/NB1 pixel_6011/VBIAS pixel_6011/NB2 pixel_6011/AMP_IN pixel_6011/SF_IB
+ pixel_6011/PIX_OUT pixel_6011/CSA_VREF pixel
Xpixel_6022 pixel_6022/gring pixel_6022/VDD pixel_6022/GND pixel_6022/VREF pixel_6022/ROW_SEL
+ pixel_6022/NB1 pixel_6022/VBIAS pixel_6022/NB2 pixel_6022/AMP_IN pixel_6022/SF_IB
+ pixel_6022/PIX_OUT pixel_6022/CSA_VREF pixel
Xpixel_6033 pixel_6033/gring pixel_6033/VDD pixel_6033/GND pixel_6033/VREF pixel_6033/ROW_SEL
+ pixel_6033/NB1 pixel_6033/VBIAS pixel_6033/NB2 pixel_6033/AMP_IN pixel_6033/SF_IB
+ pixel_6033/PIX_OUT pixel_6033/CSA_VREF pixel
Xpixel_6044 pixel_6044/gring pixel_6044/VDD pixel_6044/GND pixel_6044/VREF pixel_6044/ROW_SEL
+ pixel_6044/NB1 pixel_6044/VBIAS pixel_6044/NB2 pixel_6044/AMP_IN pixel_6044/SF_IB
+ pixel_6044/PIX_OUT pixel_6044/CSA_VREF pixel
Xpixel_6055 pixel_6055/gring pixel_6055/VDD pixel_6055/GND pixel_6055/VREF pixel_6055/ROW_SEL
+ pixel_6055/NB1 pixel_6055/VBIAS pixel_6055/NB2 pixel_6055/AMP_IN pixel_6055/SF_IB
+ pixel_6055/PIX_OUT pixel_6055/CSA_VREF pixel
Xpixel_6066 pixel_6066/gring pixel_6066/VDD pixel_6066/GND pixel_6066/VREF pixel_6066/ROW_SEL
+ pixel_6066/NB1 pixel_6066/VBIAS pixel_6066/NB2 pixel_6066/AMP_IN pixel_6066/SF_IB
+ pixel_6066/PIX_OUT pixel_6066/CSA_VREF pixel
Xpixel_6077 pixel_6077/gring pixel_6077/VDD pixel_6077/GND pixel_6077/VREF pixel_6077/ROW_SEL
+ pixel_6077/NB1 pixel_6077/VBIAS pixel_6077/NB2 pixel_6077/AMP_IN pixel_6077/SF_IB
+ pixel_6077/PIX_OUT pixel_6077/CSA_VREF pixel
Xpixel_5310 pixel_5310/gring pixel_5310/VDD pixel_5310/GND pixel_5310/VREF pixel_5310/ROW_SEL
+ pixel_5310/NB1 pixel_5310/VBIAS pixel_5310/NB2 pixel_5310/AMP_IN pixel_5310/SF_IB
+ pixel_5310/PIX_OUT pixel_5310/CSA_VREF pixel
Xpixel_5321 pixel_5321/gring pixel_5321/VDD pixel_5321/GND pixel_5321/VREF pixel_5321/ROW_SEL
+ pixel_5321/NB1 pixel_5321/VBIAS pixel_5321/NB2 pixel_5321/AMP_IN pixel_5321/SF_IB
+ pixel_5321/PIX_OUT pixel_5321/CSA_VREF pixel
Xpixel_5332 pixel_5332/gring pixel_5332/VDD pixel_5332/GND pixel_5332/VREF pixel_5332/ROW_SEL
+ pixel_5332/NB1 pixel_5332/VBIAS pixel_5332/NB2 pixel_5332/AMP_IN pixel_5332/SF_IB
+ pixel_5332/PIX_OUT pixel_5332/CSA_VREF pixel
Xpixel_6088 pixel_6088/gring pixel_6088/VDD pixel_6088/GND pixel_6088/VREF pixel_6088/ROW_SEL
+ pixel_6088/NB1 pixel_6088/VBIAS pixel_6088/NB2 pixel_6088/AMP_IN pixel_6088/SF_IB
+ pixel_6088/PIX_OUT pixel_6088/CSA_VREF pixel
Xpixel_6099 pixel_6099/gring pixel_6099/VDD pixel_6099/GND pixel_6099/VREF pixel_6099/ROW_SEL
+ pixel_6099/NB1 pixel_6099/VBIAS pixel_6099/NB2 pixel_6099/AMP_IN pixel_6099/SF_IB
+ pixel_6099/PIX_OUT pixel_6099/CSA_VREF pixel
Xpixel_5343 pixel_5343/gring pixel_5343/VDD pixel_5343/GND pixel_5343/VREF pixel_5343/ROW_SEL
+ pixel_5343/NB1 pixel_5343/VBIAS pixel_5343/NB2 pixel_5343/AMP_IN pixel_5343/SF_IB
+ pixel_5343/PIX_OUT pixel_5343/CSA_VREF pixel
Xpixel_5354 pixel_5354/gring pixel_5354/VDD pixel_5354/GND pixel_5354/VREF pixel_5354/ROW_SEL
+ pixel_5354/NB1 pixel_5354/VBIAS pixel_5354/NB2 pixel_5354/AMP_IN pixel_5354/SF_IB
+ pixel_5354/PIX_OUT pixel_5354/CSA_VREF pixel
Xpixel_5365 pixel_5365/gring pixel_5365/VDD pixel_5365/GND pixel_5365/VREF pixel_5365/ROW_SEL
+ pixel_5365/NB1 pixel_5365/VBIAS pixel_5365/NB2 pixel_5365/AMP_IN pixel_5365/SF_IB
+ pixel_5365/PIX_OUT pixel_5365/CSA_VREF pixel
Xpixel_4620 pixel_4620/gring pixel_4620/VDD pixel_4620/GND pixel_4620/VREF pixel_4620/ROW_SEL
+ pixel_4620/NB1 pixel_4620/VBIAS pixel_4620/NB2 pixel_4620/AMP_IN pixel_4620/SF_IB
+ pixel_4620/PIX_OUT pixel_4620/CSA_VREF pixel
Xpixel_5376 pixel_5376/gring pixel_5376/VDD pixel_5376/GND pixel_5376/VREF pixel_5376/ROW_SEL
+ pixel_5376/NB1 pixel_5376/VBIAS pixel_5376/NB2 pixel_5376/AMP_IN pixel_5376/SF_IB
+ pixel_5376/PIX_OUT pixel_5376/CSA_VREF pixel
Xpixel_5387 pixel_5387/gring pixel_5387/VDD pixel_5387/GND pixel_5387/VREF pixel_5387/ROW_SEL
+ pixel_5387/NB1 pixel_5387/VBIAS pixel_5387/NB2 pixel_5387/AMP_IN pixel_5387/SF_IB
+ pixel_5387/PIX_OUT pixel_5387/CSA_VREF pixel
Xpixel_5398 pixel_5398/gring pixel_5398/VDD pixel_5398/GND pixel_5398/VREF pixel_5398/ROW_SEL
+ pixel_5398/NB1 pixel_5398/VBIAS pixel_5398/NB2 pixel_5398/AMP_IN pixel_5398/SF_IB
+ pixel_5398/PIX_OUT pixel_5398/CSA_VREF pixel
Xpixel_4631 pixel_4631/gring pixel_4631/VDD pixel_4631/GND pixel_4631/VREF pixel_4631/ROW_SEL
+ pixel_4631/NB1 pixel_4631/VBIAS pixel_4631/NB2 pixel_4631/AMP_IN pixel_4631/SF_IB
+ pixel_4631/PIX_OUT pixel_4631/CSA_VREF pixel
Xpixel_4642 pixel_4642/gring pixel_4642/VDD pixel_4642/GND pixel_4642/VREF pixel_4642/ROW_SEL
+ pixel_4642/NB1 pixel_4642/VBIAS pixel_4642/NB2 pixel_4642/AMP_IN pixel_4642/SF_IB
+ pixel_4642/PIX_OUT pixel_4642/CSA_VREF pixel
Xpixel_4653 pixel_4653/gring pixel_4653/VDD pixel_4653/GND pixel_4653/VREF pixel_4653/ROW_SEL
+ pixel_4653/NB1 pixel_4653/VBIAS pixel_4653/NB2 pixel_4653/AMP_IN pixel_4653/SF_IB
+ pixel_4653/PIX_OUT pixel_4653/CSA_VREF pixel
Xpixel_4664 pixel_4664/gring pixel_4664/VDD pixel_4664/GND pixel_4664/VREF pixel_4664/ROW_SEL
+ pixel_4664/NB1 pixel_4664/VBIAS pixel_4664/NB2 pixel_4664/AMP_IN pixel_4664/SF_IB
+ pixel_4664/PIX_OUT pixel_4664/CSA_VREF pixel
Xpixel_692 pixel_692/gring pixel_692/VDD pixel_692/GND pixel_692/VREF pixel_692/ROW_SEL
+ pixel_692/NB1 pixel_692/VBIAS pixel_692/NB2 pixel_692/AMP_IN pixel_692/SF_IB pixel_692/PIX_OUT
+ pixel_692/CSA_VREF pixel
Xpixel_681 pixel_681/gring pixel_681/VDD pixel_681/GND pixel_681/VREF pixel_681/ROW_SEL
+ pixel_681/NB1 pixel_681/VBIAS pixel_681/NB2 pixel_681/AMP_IN pixel_681/SF_IB pixel_681/PIX_OUT
+ pixel_681/CSA_VREF pixel
Xpixel_670 pixel_670/gring pixel_670/VDD pixel_670/GND pixel_670/VREF pixel_670/ROW_SEL
+ pixel_670/NB1 pixel_670/VBIAS pixel_670/NB2 pixel_670/AMP_IN pixel_670/SF_IB pixel_670/PIX_OUT
+ pixel_670/CSA_VREF pixel
Xpixel_4675 pixel_4675/gring pixel_4675/VDD pixel_4675/GND pixel_4675/VREF pixel_4675/ROW_SEL
+ pixel_4675/NB1 pixel_4675/VBIAS pixel_4675/NB2 pixel_4675/AMP_IN pixel_4675/SF_IB
+ pixel_4675/PIX_OUT pixel_4675/CSA_VREF pixel
Xpixel_4686 pixel_4686/gring pixel_4686/VDD pixel_4686/GND pixel_4686/VREF pixel_4686/ROW_SEL
+ pixel_4686/NB1 pixel_4686/VBIAS pixel_4686/NB2 pixel_4686/AMP_IN pixel_4686/SF_IB
+ pixel_4686/PIX_OUT pixel_4686/CSA_VREF pixel
Xpixel_4697 pixel_4697/gring pixel_4697/VDD pixel_4697/GND pixel_4697/VREF pixel_4697/ROW_SEL
+ pixel_4697/NB1 pixel_4697/VBIAS pixel_4697/NB2 pixel_4697/AMP_IN pixel_4697/SF_IB
+ pixel_4697/PIX_OUT pixel_4697/CSA_VREF pixel
Xpixel_3930 pixel_3930/gring pixel_3930/VDD pixel_3930/GND pixel_3930/VREF pixel_3930/ROW_SEL
+ pixel_3930/NB1 pixel_3930/VBIAS pixel_3930/NB2 pixel_3930/AMP_IN pixel_3930/SF_IB
+ pixel_3930/PIX_OUT pixel_3930/CSA_VREF pixel
Xpixel_3941 pixel_3941/gring pixel_3941/VDD pixel_3941/GND pixel_3941/VREF pixel_3941/ROW_SEL
+ pixel_3941/NB1 pixel_3941/VBIAS pixel_3941/NB2 pixel_3941/AMP_IN pixel_3941/SF_IB
+ pixel_3941/PIX_OUT pixel_3941/CSA_VREF pixel
Xpixel_3952 pixel_3952/gring pixel_3952/VDD pixel_3952/GND pixel_3952/VREF pixel_3952/ROW_SEL
+ pixel_3952/NB1 pixel_3952/VBIAS pixel_3952/NB2 pixel_3952/AMP_IN pixel_3952/SF_IB
+ pixel_3952/PIX_OUT pixel_3952/CSA_VREF pixel
Xpixel_3963 pixel_3963/gring pixel_3963/VDD pixel_3963/GND pixel_3963/VREF pixel_3963/ROW_SEL
+ pixel_3963/NB1 pixel_3963/VBIAS pixel_3963/NB2 pixel_3963/AMP_IN pixel_3963/SF_IB
+ pixel_3963/PIX_OUT pixel_3963/CSA_VREF pixel
Xpixel_3974 pixel_3974/gring pixel_3974/VDD pixel_3974/GND pixel_3974/VREF pixel_3974/ROW_SEL
+ pixel_3974/NB1 pixel_3974/VBIAS pixel_3974/NB2 pixel_3974/AMP_IN pixel_3974/SF_IB
+ pixel_3974/PIX_OUT pixel_3974/CSA_VREF pixel
Xpixel_3985 pixel_3985/gring pixel_3985/VDD pixel_3985/GND pixel_3985/VREF pixel_3985/ROW_SEL
+ pixel_3985/NB1 pixel_3985/VBIAS pixel_3985/NB2 pixel_3985/AMP_IN pixel_3985/SF_IB
+ pixel_3985/PIX_OUT pixel_3985/CSA_VREF pixel
Xpixel_3996 pixel_3996/gring pixel_3996/VDD pixel_3996/GND pixel_3996/VREF pixel_3996/ROW_SEL
+ pixel_3996/NB1 pixel_3996/VBIAS pixel_3996/NB2 pixel_3996/AMP_IN pixel_3996/SF_IB
+ pixel_3996/PIX_OUT pixel_3996/CSA_VREF pixel
Xpixel_6 pixel_6/gring pixel_6/VDD pixel_6/GND pixel_6/VREF pixel_6/ROW_SEL pixel_6/NB1
+ pixel_6/VBIAS pixel_6/NB2 pixel_6/AMP_IN pixel_6/SF_IB pixel_6/PIX_OUT pixel_6/CSA_VREF
+ pixel
Xpixel_7290 pixel_7290/gring pixel_7290/VDD pixel_7290/GND pixel_7290/VREF pixel_7290/ROW_SEL
+ pixel_7290/NB1 pixel_7290/VBIAS pixel_7290/NB2 pixel_7290/AMP_IN pixel_7290/SF_IB
+ pixel_7290/PIX_OUT pixel_7290/CSA_VREF pixel
Xpixel_9609 pixel_9609/gring pixel_9609/VDD pixel_9609/GND pixel_9609/VREF pixel_9609/ROW_SEL
+ pixel_9609/NB1 pixel_9609/VBIAS pixel_9609/NB2 pixel_9609/AMP_IN pixel_9609/SF_IB
+ pixel_9609/PIX_OUT pixel_9609/CSA_VREF pixel
Xpixel_8919 pixel_8919/gring pixel_8919/VDD pixel_8919/GND pixel_8919/VREF pixel_8919/ROW_SEL
+ pixel_8919/NB1 pixel_8919/VBIAS pixel_8919/NB2 pixel_8919/AMP_IN pixel_8919/SF_IB
+ pixel_8919/PIX_OUT pixel_8919/CSA_VREF pixel
Xpixel_8908 pixel_8908/gring pixel_8908/VDD pixel_8908/GND pixel_8908/VREF pixel_8908/ROW_SEL
+ pixel_8908/NB1 pixel_8908/VBIAS pixel_8908/NB2 pixel_8908/AMP_IN pixel_8908/SF_IB
+ pixel_8908/PIX_OUT pixel_8908/CSA_VREF pixel
Xpixel_3215 pixel_3215/gring pixel_3215/VDD pixel_3215/GND pixel_3215/VREF pixel_3215/ROW_SEL
+ pixel_3215/NB1 pixel_3215/VBIAS pixel_3215/NB2 pixel_3215/AMP_IN pixel_3215/SF_IB
+ pixel_3215/PIX_OUT pixel_3215/CSA_VREF pixel
Xpixel_3204 pixel_3204/gring pixel_3204/VDD pixel_3204/GND pixel_3204/VREF pixel_3204/ROW_SEL
+ pixel_3204/NB1 pixel_3204/VBIAS pixel_3204/NB2 pixel_3204/AMP_IN pixel_3204/SF_IB
+ pixel_3204/PIX_OUT pixel_3204/CSA_VREF pixel
Xpixel_2503 pixel_2503/gring pixel_2503/VDD pixel_2503/GND pixel_2503/VREF pixel_2503/ROW_SEL
+ pixel_2503/NB1 pixel_2503/VBIAS pixel_2503/NB2 pixel_2503/AMP_IN pixel_2503/SF_IB
+ pixel_2503/PIX_OUT pixel_2503/CSA_VREF pixel
Xpixel_3248 pixel_3248/gring pixel_3248/VDD pixel_3248/GND pixel_3248/VREF pixel_3248/ROW_SEL
+ pixel_3248/NB1 pixel_3248/VBIAS pixel_3248/NB2 pixel_3248/AMP_IN pixel_3248/SF_IB
+ pixel_3248/PIX_OUT pixel_3248/CSA_VREF pixel
Xpixel_3237 pixel_3237/gring pixel_3237/VDD pixel_3237/GND pixel_3237/VREF pixel_3237/ROW_SEL
+ pixel_3237/NB1 pixel_3237/VBIAS pixel_3237/NB2 pixel_3237/AMP_IN pixel_3237/SF_IB
+ pixel_3237/PIX_OUT pixel_3237/CSA_VREF pixel
Xpixel_3226 pixel_3226/gring pixel_3226/VDD pixel_3226/GND pixel_3226/VREF pixel_3226/ROW_SEL
+ pixel_3226/NB1 pixel_3226/VBIAS pixel_3226/NB2 pixel_3226/AMP_IN pixel_3226/SF_IB
+ pixel_3226/PIX_OUT pixel_3226/CSA_VREF pixel
Xpixel_2536 pixel_2536/gring pixel_2536/VDD pixel_2536/GND pixel_2536/VREF pixel_2536/ROW_SEL
+ pixel_2536/NB1 pixel_2536/VBIAS pixel_2536/NB2 pixel_2536/AMP_IN pixel_2536/SF_IB
+ pixel_2536/PIX_OUT pixel_2536/CSA_VREF pixel
Xpixel_2525 pixel_2525/gring pixel_2525/VDD pixel_2525/GND pixel_2525/VREF pixel_2525/ROW_SEL
+ pixel_2525/NB1 pixel_2525/VBIAS pixel_2525/NB2 pixel_2525/AMP_IN pixel_2525/SF_IB
+ pixel_2525/PIX_OUT pixel_2525/CSA_VREF pixel
Xpixel_2514 pixel_2514/gring pixel_2514/VDD pixel_2514/GND pixel_2514/VREF pixel_2514/ROW_SEL
+ pixel_2514/NB1 pixel_2514/VBIAS pixel_2514/NB2 pixel_2514/AMP_IN pixel_2514/SF_IB
+ pixel_2514/PIX_OUT pixel_2514/CSA_VREF pixel
Xpixel_3259 pixel_3259/gring pixel_3259/VDD pixel_3259/GND pixel_3259/VREF pixel_3259/ROW_SEL
+ pixel_3259/NB1 pixel_3259/VBIAS pixel_3259/NB2 pixel_3259/AMP_IN pixel_3259/SF_IB
+ pixel_3259/PIX_OUT pixel_3259/CSA_VREF pixel
Xpixel_1835 pixel_1835/gring pixel_1835/VDD pixel_1835/GND pixel_1835/VREF pixel_1835/ROW_SEL
+ pixel_1835/NB1 pixel_1835/VBIAS pixel_1835/NB2 pixel_1835/AMP_IN pixel_1835/SF_IB
+ pixel_1835/PIX_OUT pixel_1835/CSA_VREF pixel
Xpixel_1824 pixel_1824/gring pixel_1824/VDD pixel_1824/GND pixel_1824/VREF pixel_1824/ROW_SEL
+ pixel_1824/NB1 pixel_1824/VBIAS pixel_1824/NB2 pixel_1824/AMP_IN pixel_1824/SF_IB
+ pixel_1824/PIX_OUT pixel_1824/CSA_VREF pixel
Xpixel_1813 pixel_1813/gring pixel_1813/VDD pixel_1813/GND pixel_1813/VREF pixel_1813/ROW_SEL
+ pixel_1813/NB1 pixel_1813/VBIAS pixel_1813/NB2 pixel_1813/AMP_IN pixel_1813/SF_IB
+ pixel_1813/PIX_OUT pixel_1813/CSA_VREF pixel
Xpixel_1802 pixel_1802/gring pixel_1802/VDD pixel_1802/GND pixel_1802/VREF pixel_1802/ROW_SEL
+ pixel_1802/NB1 pixel_1802/VBIAS pixel_1802/NB2 pixel_1802/AMP_IN pixel_1802/SF_IB
+ pixel_1802/PIX_OUT pixel_1802/CSA_VREF pixel
Xpixel_2569 pixel_2569/gring pixel_2569/VDD pixel_2569/GND pixel_2569/VREF pixel_2569/ROW_SEL
+ pixel_2569/NB1 pixel_2569/VBIAS pixel_2569/NB2 pixel_2569/AMP_IN pixel_2569/SF_IB
+ pixel_2569/PIX_OUT pixel_2569/CSA_VREF pixel
Xpixel_2558 pixel_2558/gring pixel_2558/VDD pixel_2558/GND pixel_2558/VREF pixel_2558/ROW_SEL
+ pixel_2558/NB1 pixel_2558/VBIAS pixel_2558/NB2 pixel_2558/AMP_IN pixel_2558/SF_IB
+ pixel_2558/PIX_OUT pixel_2558/CSA_VREF pixel
Xpixel_2547 pixel_2547/gring pixel_2547/VDD pixel_2547/GND pixel_2547/VREF pixel_2547/ROW_SEL
+ pixel_2547/NB1 pixel_2547/VBIAS pixel_2547/NB2 pixel_2547/AMP_IN pixel_2547/SF_IB
+ pixel_2547/PIX_OUT pixel_2547/CSA_VREF pixel
Xpixel_1868 pixel_1868/gring pixel_1868/VDD pixel_1868/GND pixel_1868/VREF pixel_1868/ROW_SEL
+ pixel_1868/NB1 pixel_1868/VBIAS pixel_1868/NB2 pixel_1868/AMP_IN pixel_1868/SF_IB
+ pixel_1868/PIX_OUT pixel_1868/CSA_VREF pixel
Xpixel_1857 pixel_1857/gring pixel_1857/VDD pixel_1857/GND pixel_1857/VREF pixel_1857/ROW_SEL
+ pixel_1857/NB1 pixel_1857/VBIAS pixel_1857/NB2 pixel_1857/AMP_IN pixel_1857/SF_IB
+ pixel_1857/PIX_OUT pixel_1857/CSA_VREF pixel
Xpixel_1846 pixel_1846/gring pixel_1846/VDD pixel_1846/GND pixel_1846/VREF pixel_1846/ROW_SEL
+ pixel_1846/NB1 pixel_1846/VBIAS pixel_1846/NB2 pixel_1846/AMP_IN pixel_1846/SF_IB
+ pixel_1846/PIX_OUT pixel_1846/CSA_VREF pixel
Xpixel_1879 pixel_1879/gring pixel_1879/VDD pixel_1879/GND pixel_1879/VREF pixel_1879/ROW_SEL
+ pixel_1879/NB1 pixel_1879/VBIAS pixel_1879/NB2 pixel_1879/AMP_IN pixel_1879/SF_IB
+ pixel_1879/PIX_OUT pixel_1879/CSA_VREF pixel
Xpixel_5140 pixel_5140/gring pixel_5140/VDD pixel_5140/GND pixel_5140/VREF pixel_5140/ROW_SEL
+ pixel_5140/NB1 pixel_5140/VBIAS pixel_5140/NB2 pixel_5140/AMP_IN pixel_5140/SF_IB
+ pixel_5140/PIX_OUT pixel_5140/CSA_VREF pixel
Xpixel_5151 pixel_5151/gring pixel_5151/VDD pixel_5151/GND pixel_5151/VREF pixel_5151/ROW_SEL
+ pixel_5151/NB1 pixel_5151/VBIAS pixel_5151/NB2 pixel_5151/AMP_IN pixel_5151/SF_IB
+ pixel_5151/PIX_OUT pixel_5151/CSA_VREF pixel
Xpixel_5162 pixel_5162/gring pixel_5162/VDD pixel_5162/GND pixel_5162/VREF pixel_5162/ROW_SEL
+ pixel_5162/NB1 pixel_5162/VBIAS pixel_5162/NB2 pixel_5162/AMP_IN pixel_5162/SF_IB
+ pixel_5162/PIX_OUT pixel_5162/CSA_VREF pixel
Xpixel_5173 pixel_5173/gring pixel_5173/VDD pixel_5173/GND pixel_5173/VREF pixel_5173/ROW_SEL
+ pixel_5173/NB1 pixel_5173/VBIAS pixel_5173/NB2 pixel_5173/AMP_IN pixel_5173/SF_IB
+ pixel_5173/PIX_OUT pixel_5173/CSA_VREF pixel
Xpixel_5184 pixel_5184/gring pixel_5184/VDD pixel_5184/GND pixel_5184/VREF pixel_5184/ROW_SEL
+ pixel_5184/NB1 pixel_5184/VBIAS pixel_5184/NB2 pixel_5184/AMP_IN pixel_5184/SF_IB
+ pixel_5184/PIX_OUT pixel_5184/CSA_VREF pixel
Xpixel_5195 pixel_5195/gring pixel_5195/VDD pixel_5195/GND pixel_5195/VREF pixel_5195/ROW_SEL
+ pixel_5195/NB1 pixel_5195/VBIAS pixel_5195/NB2 pixel_5195/AMP_IN pixel_5195/SF_IB
+ pixel_5195/PIX_OUT pixel_5195/CSA_VREF pixel
Xpixel_4450 pixel_4450/gring pixel_4450/VDD pixel_4450/GND pixel_4450/VREF pixel_4450/ROW_SEL
+ pixel_4450/NB1 pixel_4450/VBIAS pixel_4450/NB2 pixel_4450/AMP_IN pixel_4450/SF_IB
+ pixel_4450/PIX_OUT pixel_4450/CSA_VREF pixel
Xpixel_4461 pixel_4461/gring pixel_4461/VDD pixel_4461/GND pixel_4461/VREF pixel_4461/ROW_SEL
+ pixel_4461/NB1 pixel_4461/VBIAS pixel_4461/NB2 pixel_4461/AMP_IN pixel_4461/SF_IB
+ pixel_4461/PIX_OUT pixel_4461/CSA_VREF pixel
Xpixel_4472 pixel_4472/gring pixel_4472/VDD pixel_4472/GND pixel_4472/VREF pixel_4472/ROW_SEL
+ pixel_4472/NB1 pixel_4472/VBIAS pixel_4472/NB2 pixel_4472/AMP_IN pixel_4472/SF_IB
+ pixel_4472/PIX_OUT pixel_4472/CSA_VREF pixel
Xpixel_3760 pixel_3760/gring pixel_3760/VDD pixel_3760/GND pixel_3760/VREF pixel_3760/ROW_SEL
+ pixel_3760/NB1 pixel_3760/VBIAS pixel_3760/NB2 pixel_3760/AMP_IN pixel_3760/SF_IB
+ pixel_3760/PIX_OUT pixel_3760/CSA_VREF pixel
Xpixel_4483 pixel_4483/gring pixel_4483/VDD pixel_4483/GND pixel_4483/VREF pixel_4483/ROW_SEL
+ pixel_4483/NB1 pixel_4483/VBIAS pixel_4483/NB2 pixel_4483/AMP_IN pixel_4483/SF_IB
+ pixel_4483/PIX_OUT pixel_4483/CSA_VREF pixel
Xpixel_4494 pixel_4494/gring pixel_4494/VDD pixel_4494/GND pixel_4494/VREF pixel_4494/ROW_SEL
+ pixel_4494/NB1 pixel_4494/VBIAS pixel_4494/NB2 pixel_4494/AMP_IN pixel_4494/SF_IB
+ pixel_4494/PIX_OUT pixel_4494/CSA_VREF pixel
Xpixel_3793 pixel_3793/gring pixel_3793/VDD pixel_3793/GND pixel_3793/VREF pixel_3793/ROW_SEL
+ pixel_3793/NB1 pixel_3793/VBIAS pixel_3793/NB2 pixel_3793/AMP_IN pixel_3793/SF_IB
+ pixel_3793/PIX_OUT pixel_3793/CSA_VREF pixel
Xpixel_3782 pixel_3782/gring pixel_3782/VDD pixel_3782/GND pixel_3782/VREF pixel_3782/ROW_SEL
+ pixel_3782/NB1 pixel_3782/VBIAS pixel_3782/NB2 pixel_3782/AMP_IN pixel_3782/SF_IB
+ pixel_3782/PIX_OUT pixel_3782/CSA_VREF pixel
Xpixel_3771 pixel_3771/gring pixel_3771/VDD pixel_3771/GND pixel_3771/VREF pixel_3771/ROW_SEL
+ pixel_3771/NB1 pixel_3771/VBIAS pixel_3771/NB2 pixel_3771/AMP_IN pixel_3771/SF_IB
+ pixel_3771/PIX_OUT pixel_3771/CSA_VREF pixel
Xpixel_1109 pixel_1109/gring pixel_1109/VDD pixel_1109/GND pixel_1109/VREF pixel_1109/ROW_SEL
+ pixel_1109/NB1 pixel_1109/VBIAS pixel_1109/NB2 pixel_1109/AMP_IN pixel_1109/SF_IB
+ pixel_1109/PIX_OUT pixel_1109/CSA_VREF pixel
Xpixel_9428 pixel_9428/gring pixel_9428/VDD pixel_9428/GND pixel_9428/VREF pixel_9428/ROW_SEL
+ pixel_9428/NB1 pixel_9428/VBIAS pixel_9428/NB2 pixel_9428/AMP_IN pixel_9428/SF_IB
+ pixel_9428/PIX_OUT pixel_9428/CSA_VREF pixel
Xpixel_9417 pixel_9417/gring pixel_9417/VDD pixel_9417/GND pixel_9417/VREF pixel_9417/ROW_SEL
+ pixel_9417/NB1 pixel_9417/VBIAS pixel_9417/NB2 pixel_9417/AMP_IN pixel_9417/SF_IB
+ pixel_9417/PIX_OUT pixel_9417/CSA_VREF pixel
Xpixel_9406 pixel_9406/gring pixel_9406/VDD pixel_9406/GND pixel_9406/VREF pixel_9406/ROW_SEL
+ pixel_9406/NB1 pixel_9406/VBIAS pixel_9406/NB2 pixel_9406/AMP_IN pixel_9406/SF_IB
+ pixel_9406/PIX_OUT pixel_9406/CSA_VREF pixel
Xpixel_8727 pixel_8727/gring pixel_8727/VDD pixel_8727/GND pixel_8727/VREF pixel_8727/ROW_SEL
+ pixel_8727/NB1 pixel_8727/VBIAS pixel_8727/NB2 pixel_8727/AMP_IN pixel_8727/SF_IB
+ pixel_8727/PIX_OUT pixel_8727/CSA_VREF pixel
Xpixel_8716 pixel_8716/gring pixel_8716/VDD pixel_8716/GND pixel_8716/VREF pixel_8716/ROW_SEL
+ pixel_8716/NB1 pixel_8716/VBIAS pixel_8716/NB2 pixel_8716/AMP_IN pixel_8716/SF_IB
+ pixel_8716/PIX_OUT pixel_8716/CSA_VREF pixel
Xpixel_8705 pixel_8705/gring pixel_8705/VDD pixel_8705/GND pixel_8705/VREF pixel_8705/ROW_SEL
+ pixel_8705/NB1 pixel_8705/VBIAS pixel_8705/NB2 pixel_8705/AMP_IN pixel_8705/SF_IB
+ pixel_8705/PIX_OUT pixel_8705/CSA_VREF pixel
Xpixel_9439 pixel_9439/gring pixel_9439/VDD pixel_9439/GND pixel_9439/VREF pixel_9439/ROW_SEL
+ pixel_9439/NB1 pixel_9439/VBIAS pixel_9439/NB2 pixel_9439/AMP_IN pixel_9439/SF_IB
+ pixel_9439/PIX_OUT pixel_9439/CSA_VREF pixel
Xpixel_8749 pixel_8749/gring pixel_8749/VDD pixel_8749/GND pixel_8749/VREF pixel_8749/ROW_SEL
+ pixel_8749/NB1 pixel_8749/VBIAS pixel_8749/NB2 pixel_8749/AMP_IN pixel_8749/SF_IB
+ pixel_8749/PIX_OUT pixel_8749/CSA_VREF pixel
Xpixel_8738 pixel_8738/gring pixel_8738/VDD pixel_8738/GND pixel_8738/VREF pixel_8738/ROW_SEL
+ pixel_8738/NB1 pixel_8738/VBIAS pixel_8738/NB2 pixel_8738/AMP_IN pixel_8738/SF_IB
+ pixel_8738/PIX_OUT pixel_8738/CSA_VREF pixel
Xpixel_3023 pixel_3023/gring pixel_3023/VDD pixel_3023/GND pixel_3023/VREF pixel_3023/ROW_SEL
+ pixel_3023/NB1 pixel_3023/VBIAS pixel_3023/NB2 pixel_3023/AMP_IN pixel_3023/SF_IB
+ pixel_3023/PIX_OUT pixel_3023/CSA_VREF pixel
Xpixel_3012 pixel_3012/gring pixel_3012/VDD pixel_3012/GND pixel_3012/VREF pixel_3012/ROW_SEL
+ pixel_3012/NB1 pixel_3012/VBIAS pixel_3012/NB2 pixel_3012/AMP_IN pixel_3012/SF_IB
+ pixel_3012/PIX_OUT pixel_3012/CSA_VREF pixel
Xpixel_3001 pixel_3001/gring pixel_3001/VDD pixel_3001/GND pixel_3001/VREF pixel_3001/ROW_SEL
+ pixel_3001/NB1 pixel_3001/VBIAS pixel_3001/NB2 pixel_3001/AMP_IN pixel_3001/SF_IB
+ pixel_3001/PIX_OUT pixel_3001/CSA_VREF pixel
Xpixel_2311 pixel_2311/gring pixel_2311/VDD pixel_2311/GND pixel_2311/VREF pixel_2311/ROW_SEL
+ pixel_2311/NB1 pixel_2311/VBIAS pixel_2311/NB2 pixel_2311/AMP_IN pixel_2311/SF_IB
+ pixel_2311/PIX_OUT pixel_2311/CSA_VREF pixel
Xpixel_2300 pixel_2300/gring pixel_2300/VDD pixel_2300/GND pixel_2300/VREF pixel_2300/ROW_SEL
+ pixel_2300/NB1 pixel_2300/VBIAS pixel_2300/NB2 pixel_2300/AMP_IN pixel_2300/SF_IB
+ pixel_2300/PIX_OUT pixel_2300/CSA_VREF pixel
Xpixel_3056 pixel_3056/gring pixel_3056/VDD pixel_3056/GND pixel_3056/VREF pixel_3056/ROW_SEL
+ pixel_3056/NB1 pixel_3056/VBIAS pixel_3056/NB2 pixel_3056/AMP_IN pixel_3056/SF_IB
+ pixel_3056/PIX_OUT pixel_3056/CSA_VREF pixel
Xpixel_3045 pixel_3045/gring pixel_3045/VDD pixel_3045/GND pixel_3045/VREF pixel_3045/ROW_SEL
+ pixel_3045/NB1 pixel_3045/VBIAS pixel_3045/NB2 pixel_3045/AMP_IN pixel_3045/SF_IB
+ pixel_3045/PIX_OUT pixel_3045/CSA_VREF pixel
Xpixel_3034 pixel_3034/gring pixel_3034/VDD pixel_3034/GND pixel_3034/VREF pixel_3034/ROW_SEL
+ pixel_3034/NB1 pixel_3034/VBIAS pixel_3034/NB2 pixel_3034/AMP_IN pixel_3034/SF_IB
+ pixel_3034/PIX_OUT pixel_3034/CSA_VREF pixel
Xpixel_1610 pixel_1610/gring pixel_1610/VDD pixel_1610/GND pixel_1610/VREF pixel_1610/ROW_SEL
+ pixel_1610/NB1 pixel_1610/VBIAS pixel_1610/NB2 pixel_1610/AMP_IN pixel_1610/SF_IB
+ pixel_1610/PIX_OUT pixel_1610/CSA_VREF pixel
Xpixel_2355 pixel_2355/gring pixel_2355/VDD pixel_2355/GND pixel_2355/VREF pixel_2355/ROW_SEL
+ pixel_2355/NB1 pixel_2355/VBIAS pixel_2355/NB2 pixel_2355/AMP_IN pixel_2355/SF_IB
+ pixel_2355/PIX_OUT pixel_2355/CSA_VREF pixel
Xpixel_2344 pixel_2344/gring pixel_2344/VDD pixel_2344/GND pixel_2344/VREF pixel_2344/ROW_SEL
+ pixel_2344/NB1 pixel_2344/VBIAS pixel_2344/NB2 pixel_2344/AMP_IN pixel_2344/SF_IB
+ pixel_2344/PIX_OUT pixel_2344/CSA_VREF pixel
Xpixel_2333 pixel_2333/gring pixel_2333/VDD pixel_2333/GND pixel_2333/VREF pixel_2333/ROW_SEL
+ pixel_2333/NB1 pixel_2333/VBIAS pixel_2333/NB2 pixel_2333/AMP_IN pixel_2333/SF_IB
+ pixel_2333/PIX_OUT pixel_2333/CSA_VREF pixel
Xpixel_2322 pixel_2322/gring pixel_2322/VDD pixel_2322/GND pixel_2322/VREF pixel_2322/ROW_SEL
+ pixel_2322/NB1 pixel_2322/VBIAS pixel_2322/NB2 pixel_2322/AMP_IN pixel_2322/SF_IB
+ pixel_2322/PIX_OUT pixel_2322/CSA_VREF pixel
Xpixel_3089 pixel_3089/gring pixel_3089/VDD pixel_3089/GND pixel_3089/VREF pixel_3089/ROW_SEL
+ pixel_3089/NB1 pixel_3089/VBIAS pixel_3089/NB2 pixel_3089/AMP_IN pixel_3089/SF_IB
+ pixel_3089/PIX_OUT pixel_3089/CSA_VREF pixel
Xpixel_3078 pixel_3078/gring pixel_3078/VDD pixel_3078/GND pixel_3078/VREF pixel_3078/ROW_SEL
+ pixel_3078/NB1 pixel_3078/VBIAS pixel_3078/NB2 pixel_3078/AMP_IN pixel_3078/SF_IB
+ pixel_3078/PIX_OUT pixel_3078/CSA_VREF pixel
Xpixel_3067 pixel_3067/gring pixel_3067/VDD pixel_3067/GND pixel_3067/VREF pixel_3067/ROW_SEL
+ pixel_3067/NB1 pixel_3067/VBIAS pixel_3067/NB2 pixel_3067/AMP_IN pixel_3067/SF_IB
+ pixel_3067/PIX_OUT pixel_3067/CSA_VREF pixel
Xpixel_1643 pixel_1643/gring pixel_1643/VDD pixel_1643/GND pixel_1643/VREF pixel_1643/ROW_SEL
+ pixel_1643/NB1 pixel_1643/VBIAS pixel_1643/NB2 pixel_1643/AMP_IN pixel_1643/SF_IB
+ pixel_1643/PIX_OUT pixel_1643/CSA_VREF pixel
Xpixel_1632 pixel_1632/gring pixel_1632/VDD pixel_1632/GND pixel_1632/VREF pixel_1632/ROW_SEL
+ pixel_1632/NB1 pixel_1632/VBIAS pixel_1632/NB2 pixel_1632/AMP_IN pixel_1632/SF_IB
+ pixel_1632/PIX_OUT pixel_1632/CSA_VREF pixel
Xpixel_1621 pixel_1621/gring pixel_1621/VDD pixel_1621/GND pixel_1621/VREF pixel_1621/ROW_SEL
+ pixel_1621/NB1 pixel_1621/VBIAS pixel_1621/NB2 pixel_1621/AMP_IN pixel_1621/SF_IB
+ pixel_1621/PIX_OUT pixel_1621/CSA_VREF pixel
Xpixel_2388 pixel_2388/gring pixel_2388/VDD pixel_2388/GND pixel_2388/VREF pixel_2388/ROW_SEL
+ pixel_2388/NB1 pixel_2388/VBIAS pixel_2388/NB2 pixel_2388/AMP_IN pixel_2388/SF_IB
+ pixel_2388/PIX_OUT pixel_2388/CSA_VREF pixel
Xpixel_2377 pixel_2377/gring pixel_2377/VDD pixel_2377/GND pixel_2377/VREF pixel_2377/ROW_SEL
+ pixel_2377/NB1 pixel_2377/VBIAS pixel_2377/NB2 pixel_2377/AMP_IN pixel_2377/SF_IB
+ pixel_2377/PIX_OUT pixel_2377/CSA_VREF pixel
Xpixel_2366 pixel_2366/gring pixel_2366/VDD pixel_2366/GND pixel_2366/VREF pixel_2366/ROW_SEL
+ pixel_2366/NB1 pixel_2366/VBIAS pixel_2366/NB2 pixel_2366/AMP_IN pixel_2366/SF_IB
+ pixel_2366/PIX_OUT pixel_2366/CSA_VREF pixel
Xpixel_1676 pixel_1676/gring pixel_1676/VDD pixel_1676/GND pixel_1676/VREF pixel_1676/ROW_SEL
+ pixel_1676/NB1 pixel_1676/VBIAS pixel_1676/NB2 pixel_1676/AMP_IN pixel_1676/SF_IB
+ pixel_1676/PIX_OUT pixel_1676/CSA_VREF pixel
Xpixel_1665 pixel_1665/gring pixel_1665/VDD pixel_1665/GND pixel_1665/VREF pixel_1665/ROW_SEL
+ pixel_1665/NB1 pixel_1665/VBIAS pixel_1665/NB2 pixel_1665/AMP_IN pixel_1665/SF_IB
+ pixel_1665/PIX_OUT pixel_1665/CSA_VREF pixel
Xpixel_1654 pixel_1654/gring pixel_1654/VDD pixel_1654/GND pixel_1654/VREF pixel_1654/ROW_SEL
+ pixel_1654/NB1 pixel_1654/VBIAS pixel_1654/NB2 pixel_1654/AMP_IN pixel_1654/SF_IB
+ pixel_1654/PIX_OUT pixel_1654/CSA_VREF pixel
Xpixel_2399 pixel_2399/gring pixel_2399/VDD pixel_2399/GND pixel_2399/VREF pixel_2399/ROW_SEL
+ pixel_2399/NB1 pixel_2399/VBIAS pixel_2399/NB2 pixel_2399/AMP_IN pixel_2399/SF_IB
+ pixel_2399/PIX_OUT pixel_2399/CSA_VREF pixel
Xpixel_1698 pixel_1698/gring pixel_1698/VDD pixel_1698/GND pixel_1698/VREF pixel_1698/ROW_SEL
+ pixel_1698/NB1 pixel_1698/VBIAS pixel_1698/NB2 pixel_1698/AMP_IN pixel_1698/SF_IB
+ pixel_1698/PIX_OUT pixel_1698/CSA_VREF pixel
Xpixel_1687 pixel_1687/gring pixel_1687/VDD pixel_1687/GND pixel_1687/VREF pixel_1687/ROW_SEL
+ pixel_1687/NB1 pixel_1687/VBIAS pixel_1687/NB2 pixel_1687/AMP_IN pixel_1687/SF_IB
+ pixel_1687/PIX_OUT pixel_1687/CSA_VREF pixel
Xpixel_9940 pixel_9940/gring pixel_9940/VDD pixel_9940/GND pixel_9940/VREF pixel_9940/ROW_SEL
+ pixel_9940/NB1 pixel_9940/VBIAS pixel_9940/NB2 pixel_9940/AMP_IN pixel_9940/SF_IB
+ pixel_9940/PIX_OUT pixel_9940/CSA_VREF pixel
Xpixel_9951 pixel_9951/gring pixel_9951/VDD pixel_9951/GND pixel_9951/VREF pixel_9951/ROW_SEL
+ pixel_9951/NB1 pixel_9951/VBIAS pixel_9951/NB2 pixel_9951/AMP_IN pixel_9951/SF_IB
+ pixel_9951/PIX_OUT pixel_9951/CSA_VREF pixel
Xpixel_9962 pixel_9962/gring pixel_9962/VDD pixel_9962/GND pixel_9962/VREF pixel_9962/ROW_SEL
+ pixel_9962/NB1 pixel_9962/VBIAS pixel_9962/NB2 pixel_9962/AMP_IN pixel_9962/SF_IB
+ pixel_9962/PIX_OUT pixel_9962/CSA_VREF pixel
Xpixel_9973 pixel_9973/gring pixel_9973/VDD pixel_9973/GND pixel_9973/VREF pixel_9973/ROW_SEL
+ pixel_9973/NB1 pixel_9973/VBIAS pixel_9973/NB2 pixel_9973/AMP_IN pixel_9973/SF_IB
+ pixel_9973/PIX_OUT pixel_9973/CSA_VREF pixel
Xpixel_9984 pixel_9984/gring pixel_9984/VDD pixel_9984/GND pixel_9984/VREF pixel_9984/ROW_SEL
+ pixel_9984/NB1 pixel_9984/VBIAS pixel_9984/NB2 pixel_9984/AMP_IN pixel_9984/SF_IB
+ pixel_9984/PIX_OUT pixel_9984/CSA_VREF pixel
Xpixel_9995 pixel_9995/gring pixel_9995/VDD pixel_9995/GND pixel_9995/VREF pixel_9995/ROW_SEL
+ pixel_9995/NB1 pixel_9995/VBIAS pixel_9995/NB2 pixel_9995/AMP_IN pixel_9995/SF_IB
+ pixel_9995/PIX_OUT pixel_9995/CSA_VREF pixel
Xpixel_4280 pixel_4280/gring pixel_4280/VDD pixel_4280/GND pixel_4280/VREF pixel_4280/ROW_SEL
+ pixel_4280/NB1 pixel_4280/VBIAS pixel_4280/NB2 pixel_4280/AMP_IN pixel_4280/SF_IB
+ pixel_4280/PIX_OUT pixel_4280/CSA_VREF pixel
Xpixel_4291 pixel_4291/gring pixel_4291/VDD pixel_4291/GND pixel_4291/VREF pixel_4291/ROW_SEL
+ pixel_4291/NB1 pixel_4291/VBIAS pixel_4291/NB2 pixel_4291/AMP_IN pixel_4291/SF_IB
+ pixel_4291/PIX_OUT pixel_4291/CSA_VREF pixel
Xpixel_3590 pixel_3590/gring pixel_3590/VDD pixel_3590/GND pixel_3590/VREF pixel_3590/ROW_SEL
+ pixel_3590/NB1 pixel_3590/VBIAS pixel_3590/NB2 pixel_3590/AMP_IN pixel_3590/SF_IB
+ pixel_3590/PIX_OUT pixel_3590/CSA_VREF pixel
Xpixel_5909 pixel_5909/gring pixel_5909/VDD pixel_5909/GND pixel_5909/VREF pixel_5909/ROW_SEL
+ pixel_5909/NB1 pixel_5909/VBIAS pixel_5909/NB2 pixel_5909/AMP_IN pixel_5909/SF_IB
+ pixel_5909/PIX_OUT pixel_5909/CSA_VREF pixel
Xpixel_9203 pixel_9203/gring pixel_9203/VDD pixel_9203/GND pixel_9203/VREF pixel_9203/ROW_SEL
+ pixel_9203/NB1 pixel_9203/VBIAS pixel_9203/NB2 pixel_9203/AMP_IN pixel_9203/SF_IB
+ pixel_9203/PIX_OUT pixel_9203/CSA_VREF pixel
Xpixel_8502 pixel_8502/gring pixel_8502/VDD pixel_8502/GND pixel_8502/VREF pixel_8502/ROW_SEL
+ pixel_8502/NB1 pixel_8502/VBIAS pixel_8502/NB2 pixel_8502/AMP_IN pixel_8502/SF_IB
+ pixel_8502/PIX_OUT pixel_8502/CSA_VREF pixel
Xpixel_9247 pixel_9247/gring pixel_9247/VDD pixel_9247/GND pixel_9247/VREF pixel_9247/ROW_SEL
+ pixel_9247/NB1 pixel_9247/VBIAS pixel_9247/NB2 pixel_9247/AMP_IN pixel_9247/SF_IB
+ pixel_9247/PIX_OUT pixel_9247/CSA_VREF pixel
Xpixel_9236 pixel_9236/gring pixel_9236/VDD pixel_9236/GND pixel_9236/VREF pixel_9236/ROW_SEL
+ pixel_9236/NB1 pixel_9236/VBIAS pixel_9236/NB2 pixel_9236/AMP_IN pixel_9236/SF_IB
+ pixel_9236/PIX_OUT pixel_9236/CSA_VREF pixel
Xpixel_9225 pixel_9225/gring pixel_9225/VDD pixel_9225/GND pixel_9225/VREF pixel_9225/ROW_SEL
+ pixel_9225/NB1 pixel_9225/VBIAS pixel_9225/NB2 pixel_9225/AMP_IN pixel_9225/SF_IB
+ pixel_9225/PIX_OUT pixel_9225/CSA_VREF pixel
Xpixel_9214 pixel_9214/gring pixel_9214/VDD pixel_9214/GND pixel_9214/VREF pixel_9214/ROW_SEL
+ pixel_9214/NB1 pixel_9214/VBIAS pixel_9214/NB2 pixel_9214/AMP_IN pixel_9214/SF_IB
+ pixel_9214/PIX_OUT pixel_9214/CSA_VREF pixel
Xpixel_8535 pixel_8535/gring pixel_8535/VDD pixel_8535/GND pixel_8535/VREF pixel_8535/ROW_SEL
+ pixel_8535/NB1 pixel_8535/VBIAS pixel_8535/NB2 pixel_8535/AMP_IN pixel_8535/SF_IB
+ pixel_8535/PIX_OUT pixel_8535/CSA_VREF pixel
Xpixel_8524 pixel_8524/gring pixel_8524/VDD pixel_8524/GND pixel_8524/VREF pixel_8524/ROW_SEL
+ pixel_8524/NB1 pixel_8524/VBIAS pixel_8524/NB2 pixel_8524/AMP_IN pixel_8524/SF_IB
+ pixel_8524/PIX_OUT pixel_8524/CSA_VREF pixel
Xpixel_8513 pixel_8513/gring pixel_8513/VDD pixel_8513/GND pixel_8513/VREF pixel_8513/ROW_SEL
+ pixel_8513/NB1 pixel_8513/VBIAS pixel_8513/NB2 pixel_8513/AMP_IN pixel_8513/SF_IB
+ pixel_8513/PIX_OUT pixel_8513/CSA_VREF pixel
Xpixel_9269 pixel_9269/gring pixel_9269/VDD pixel_9269/GND pixel_9269/VREF pixel_9269/ROW_SEL
+ pixel_9269/NB1 pixel_9269/VBIAS pixel_9269/NB2 pixel_9269/AMP_IN pixel_9269/SF_IB
+ pixel_9269/PIX_OUT pixel_9269/CSA_VREF pixel
Xpixel_9258 pixel_9258/gring pixel_9258/VDD pixel_9258/GND pixel_9258/VREF pixel_9258/ROW_SEL
+ pixel_9258/NB1 pixel_9258/VBIAS pixel_9258/NB2 pixel_9258/AMP_IN pixel_9258/SF_IB
+ pixel_9258/PIX_OUT pixel_9258/CSA_VREF pixel
Xpixel_8568 pixel_8568/gring pixel_8568/VDD pixel_8568/GND pixel_8568/VREF pixel_8568/ROW_SEL
+ pixel_8568/NB1 pixel_8568/VBIAS pixel_8568/NB2 pixel_8568/AMP_IN pixel_8568/SF_IB
+ pixel_8568/PIX_OUT pixel_8568/CSA_VREF pixel
Xpixel_8557 pixel_8557/gring pixel_8557/VDD pixel_8557/GND pixel_8557/VREF pixel_8557/ROW_SEL
+ pixel_8557/NB1 pixel_8557/VBIAS pixel_8557/NB2 pixel_8557/AMP_IN pixel_8557/SF_IB
+ pixel_8557/PIX_OUT pixel_8557/CSA_VREF pixel
Xpixel_8546 pixel_8546/gring pixel_8546/VDD pixel_8546/GND pixel_8546/VREF pixel_8546/ROW_SEL
+ pixel_8546/NB1 pixel_8546/VBIAS pixel_8546/NB2 pixel_8546/AMP_IN pixel_8546/SF_IB
+ pixel_8546/PIX_OUT pixel_8546/CSA_VREF pixel
Xpixel_7801 pixel_7801/gring pixel_7801/VDD pixel_7801/GND pixel_7801/VREF pixel_7801/ROW_SEL
+ pixel_7801/NB1 pixel_7801/VBIAS pixel_7801/NB2 pixel_7801/AMP_IN pixel_7801/SF_IB
+ pixel_7801/PIX_OUT pixel_7801/CSA_VREF pixel
Xpixel_7812 pixel_7812/gring pixel_7812/VDD pixel_7812/GND pixel_7812/VREF pixel_7812/ROW_SEL
+ pixel_7812/NB1 pixel_7812/VBIAS pixel_7812/NB2 pixel_7812/AMP_IN pixel_7812/SF_IB
+ pixel_7812/PIX_OUT pixel_7812/CSA_VREF pixel
Xpixel_7823 pixel_7823/gring pixel_7823/VDD pixel_7823/GND pixel_7823/VREF pixel_7823/ROW_SEL
+ pixel_7823/NB1 pixel_7823/VBIAS pixel_7823/NB2 pixel_7823/AMP_IN pixel_7823/SF_IB
+ pixel_7823/PIX_OUT pixel_7823/CSA_VREF pixel
Xpixel_7834 pixel_7834/gring pixel_7834/VDD pixel_7834/GND pixel_7834/VREF pixel_7834/ROW_SEL
+ pixel_7834/NB1 pixel_7834/VBIAS pixel_7834/NB2 pixel_7834/AMP_IN pixel_7834/SF_IB
+ pixel_7834/PIX_OUT pixel_7834/CSA_VREF pixel
Xpixel_8579 pixel_8579/gring pixel_8579/VDD pixel_8579/GND pixel_8579/VREF pixel_8579/ROW_SEL
+ pixel_8579/NB1 pixel_8579/VBIAS pixel_8579/NB2 pixel_8579/AMP_IN pixel_8579/SF_IB
+ pixel_8579/PIX_OUT pixel_8579/CSA_VREF pixel
Xpixel_7845 pixel_7845/gring pixel_7845/VDD pixel_7845/GND pixel_7845/VREF pixel_7845/ROW_SEL
+ pixel_7845/NB1 pixel_7845/VBIAS pixel_7845/NB2 pixel_7845/AMP_IN pixel_7845/SF_IB
+ pixel_7845/PIX_OUT pixel_7845/CSA_VREF pixel
Xpixel_7856 pixel_7856/gring pixel_7856/VDD pixel_7856/GND pixel_7856/VREF pixel_7856/ROW_SEL
+ pixel_7856/NB1 pixel_7856/VBIAS pixel_7856/NB2 pixel_7856/AMP_IN pixel_7856/SF_IB
+ pixel_7856/PIX_OUT pixel_7856/CSA_VREF pixel
Xpixel_7867 pixel_7867/gring pixel_7867/VDD pixel_7867/GND pixel_7867/VREF pixel_7867/ROW_SEL
+ pixel_7867/NB1 pixel_7867/VBIAS pixel_7867/NB2 pixel_7867/AMP_IN pixel_7867/SF_IB
+ pixel_7867/PIX_OUT pixel_7867/CSA_VREF pixel
Xpixel_7878 pixel_7878/gring pixel_7878/VDD pixel_7878/GND pixel_7878/VREF pixel_7878/ROW_SEL
+ pixel_7878/NB1 pixel_7878/VBIAS pixel_7878/NB2 pixel_7878/AMP_IN pixel_7878/SF_IB
+ pixel_7878/PIX_OUT pixel_7878/CSA_VREF pixel
Xpixel_7889 pixel_7889/gring pixel_7889/VDD pixel_7889/GND pixel_7889/VREF pixel_7889/ROW_SEL
+ pixel_7889/NB1 pixel_7889/VBIAS pixel_7889/NB2 pixel_7889/AMP_IN pixel_7889/SF_IB
+ pixel_7889/PIX_OUT pixel_7889/CSA_VREF pixel
Xpixel_2163 pixel_2163/gring pixel_2163/VDD pixel_2163/GND pixel_2163/VREF pixel_2163/ROW_SEL
+ pixel_2163/NB1 pixel_2163/VBIAS pixel_2163/NB2 pixel_2163/AMP_IN pixel_2163/SF_IB
+ pixel_2163/PIX_OUT pixel_2163/CSA_VREF pixel
Xpixel_2152 pixel_2152/gring pixel_2152/VDD pixel_2152/GND pixel_2152/VREF pixel_2152/ROW_SEL
+ pixel_2152/NB1 pixel_2152/VBIAS pixel_2152/NB2 pixel_2152/AMP_IN pixel_2152/SF_IB
+ pixel_2152/PIX_OUT pixel_2152/CSA_VREF pixel
Xpixel_2141 pixel_2141/gring pixel_2141/VDD pixel_2141/GND pixel_2141/VREF pixel_2141/ROW_SEL
+ pixel_2141/NB1 pixel_2141/VBIAS pixel_2141/NB2 pixel_2141/AMP_IN pixel_2141/SF_IB
+ pixel_2141/PIX_OUT pixel_2141/CSA_VREF pixel
Xpixel_2130 pixel_2130/gring pixel_2130/VDD pixel_2130/GND pixel_2130/VREF pixel_2130/ROW_SEL
+ pixel_2130/NB1 pixel_2130/VBIAS pixel_2130/NB2 pixel_2130/AMP_IN pixel_2130/SF_IB
+ pixel_2130/PIX_OUT pixel_2130/CSA_VREF pixel
Xpixel_1451 pixel_1451/gring pixel_1451/VDD pixel_1451/GND pixel_1451/VREF pixel_1451/ROW_SEL
+ pixel_1451/NB1 pixel_1451/VBIAS pixel_1451/NB2 pixel_1451/AMP_IN pixel_1451/SF_IB
+ pixel_1451/PIX_OUT pixel_1451/CSA_VREF pixel
Xpixel_1440 pixel_1440/gring pixel_1440/VDD pixel_1440/GND pixel_1440/VREF pixel_1440/ROW_SEL
+ pixel_1440/NB1 pixel_1440/VBIAS pixel_1440/NB2 pixel_1440/AMP_IN pixel_1440/SF_IB
+ pixel_1440/PIX_OUT pixel_1440/CSA_VREF pixel
Xpixel_2196 pixel_2196/gring pixel_2196/VDD pixel_2196/GND pixel_2196/VREF pixel_2196/ROW_SEL
+ pixel_2196/NB1 pixel_2196/VBIAS pixel_2196/NB2 pixel_2196/AMP_IN pixel_2196/SF_IB
+ pixel_2196/PIX_OUT pixel_2196/CSA_VREF pixel
Xpixel_2185 pixel_2185/gring pixel_2185/VDD pixel_2185/GND pixel_2185/VREF pixel_2185/ROW_SEL
+ pixel_2185/NB1 pixel_2185/VBIAS pixel_2185/NB2 pixel_2185/AMP_IN pixel_2185/SF_IB
+ pixel_2185/PIX_OUT pixel_2185/CSA_VREF pixel
Xpixel_2174 pixel_2174/gring pixel_2174/VDD pixel_2174/GND pixel_2174/VREF pixel_2174/ROW_SEL
+ pixel_2174/NB1 pixel_2174/VBIAS pixel_2174/NB2 pixel_2174/AMP_IN pixel_2174/SF_IB
+ pixel_2174/PIX_OUT pixel_2174/CSA_VREF pixel
Xpixel_1484 pixel_1484/gring pixel_1484/VDD pixel_1484/GND pixel_1484/VREF pixel_1484/ROW_SEL
+ pixel_1484/NB1 pixel_1484/VBIAS pixel_1484/NB2 pixel_1484/AMP_IN pixel_1484/SF_IB
+ pixel_1484/PIX_OUT pixel_1484/CSA_VREF pixel
Xpixel_1473 pixel_1473/gring pixel_1473/VDD pixel_1473/GND pixel_1473/VREF pixel_1473/ROW_SEL
+ pixel_1473/NB1 pixel_1473/VBIAS pixel_1473/NB2 pixel_1473/AMP_IN pixel_1473/SF_IB
+ pixel_1473/PIX_OUT pixel_1473/CSA_VREF pixel
Xpixel_1462 pixel_1462/gring pixel_1462/VDD pixel_1462/GND pixel_1462/VREF pixel_1462/ROW_SEL
+ pixel_1462/NB1 pixel_1462/VBIAS pixel_1462/NB2 pixel_1462/AMP_IN pixel_1462/SF_IB
+ pixel_1462/PIX_OUT pixel_1462/CSA_VREF pixel
Xpixel_1495 pixel_1495/gring pixel_1495/VDD pixel_1495/GND pixel_1495/VREF pixel_1495/ROW_SEL
+ pixel_1495/NB1 pixel_1495/VBIAS pixel_1495/NB2 pixel_1495/AMP_IN pixel_1495/SF_IB
+ pixel_1495/PIX_OUT pixel_1495/CSA_VREF pixel
Xpixel_9770 pixel_9770/gring pixel_9770/VDD pixel_9770/GND pixel_9770/VREF pixel_9770/ROW_SEL
+ pixel_9770/NB1 pixel_9770/VBIAS pixel_9770/NB2 pixel_9770/AMP_IN pixel_9770/SF_IB
+ pixel_9770/PIX_OUT pixel_9770/CSA_VREF pixel
Xpixel_9781 pixel_9781/gring pixel_9781/VDD pixel_9781/GND pixel_9781/VREF pixel_9781/ROW_SEL
+ pixel_9781/NB1 pixel_9781/VBIAS pixel_9781/NB2 pixel_9781/AMP_IN pixel_9781/SF_IB
+ pixel_9781/PIX_OUT pixel_9781/CSA_VREF pixel
Xpixel_9792 pixel_9792/gring pixel_9792/VDD pixel_9792/GND pixel_9792/VREF pixel_9792/ROW_SEL
+ pixel_9792/NB1 pixel_9792/VBIAS pixel_9792/NB2 pixel_9792/AMP_IN pixel_9792/SF_IB
+ pixel_9792/PIX_OUT pixel_9792/CSA_VREF pixel
Xpixel_7108 pixel_7108/gring pixel_7108/VDD pixel_7108/GND pixel_7108/VREF pixel_7108/ROW_SEL
+ pixel_7108/NB1 pixel_7108/VBIAS pixel_7108/NB2 pixel_7108/AMP_IN pixel_7108/SF_IB
+ pixel_7108/PIX_OUT pixel_7108/CSA_VREF pixel
Xpixel_7119 pixel_7119/gring pixel_7119/VDD pixel_7119/GND pixel_7119/VREF pixel_7119/ROW_SEL
+ pixel_7119/NB1 pixel_7119/VBIAS pixel_7119/NB2 pixel_7119/AMP_IN pixel_7119/SF_IB
+ pixel_7119/PIX_OUT pixel_7119/CSA_VREF pixel
Xpixel_6407 pixel_6407/gring pixel_6407/VDD pixel_6407/GND pixel_6407/VREF pixel_6407/ROW_SEL
+ pixel_6407/NB1 pixel_6407/VBIAS pixel_6407/NB2 pixel_6407/AMP_IN pixel_6407/SF_IB
+ pixel_6407/PIX_OUT pixel_6407/CSA_VREF pixel
Xpixel_6418 pixel_6418/gring pixel_6418/VDD pixel_6418/GND pixel_6418/VREF pixel_6418/ROW_SEL
+ pixel_6418/NB1 pixel_6418/VBIAS pixel_6418/NB2 pixel_6418/AMP_IN pixel_6418/SF_IB
+ pixel_6418/PIX_OUT pixel_6418/CSA_VREF pixel
Xpixel_6429 pixel_6429/gring pixel_6429/VDD pixel_6429/GND pixel_6429/VREF pixel_6429/ROW_SEL
+ pixel_6429/NB1 pixel_6429/VBIAS pixel_6429/NB2 pixel_6429/AMP_IN pixel_6429/SF_IB
+ pixel_6429/PIX_OUT pixel_6429/CSA_VREF pixel
Xpixel_5706 pixel_5706/gring pixel_5706/VDD pixel_5706/GND pixel_5706/VREF pixel_5706/ROW_SEL
+ pixel_5706/NB1 pixel_5706/VBIAS pixel_5706/NB2 pixel_5706/AMP_IN pixel_5706/SF_IB
+ pixel_5706/PIX_OUT pixel_5706/CSA_VREF pixel
Xpixel_5717 pixel_5717/gring pixel_5717/VDD pixel_5717/GND pixel_5717/VREF pixel_5717/ROW_SEL
+ pixel_5717/NB1 pixel_5717/VBIAS pixel_5717/NB2 pixel_5717/AMP_IN pixel_5717/SF_IB
+ pixel_5717/PIX_OUT pixel_5717/CSA_VREF pixel
Xpixel_5728 pixel_5728/gring pixel_5728/VDD pixel_5728/GND pixel_5728/VREF pixel_5728/ROW_SEL
+ pixel_5728/NB1 pixel_5728/VBIAS pixel_5728/NB2 pixel_5728/AMP_IN pixel_5728/SF_IB
+ pixel_5728/PIX_OUT pixel_5728/CSA_VREF pixel
Xpixel_5739 pixel_5739/gring pixel_5739/VDD pixel_5739/GND pixel_5739/VREF pixel_5739/ROW_SEL
+ pixel_5739/NB1 pixel_5739/VBIAS pixel_5739/NB2 pixel_5739/AMP_IN pixel_5739/SF_IB
+ pixel_5739/PIX_OUT pixel_5739/CSA_VREF pixel
Xpixel_9022 pixel_9022/gring pixel_9022/VDD pixel_9022/GND pixel_9022/VREF pixel_9022/ROW_SEL
+ pixel_9022/NB1 pixel_9022/VBIAS pixel_9022/NB2 pixel_9022/AMP_IN pixel_9022/SF_IB
+ pixel_9022/PIX_OUT pixel_9022/CSA_VREF pixel
Xpixel_9011 pixel_9011/gring pixel_9011/VDD pixel_9011/GND pixel_9011/VREF pixel_9011/ROW_SEL
+ pixel_9011/NB1 pixel_9011/VBIAS pixel_9011/NB2 pixel_9011/AMP_IN pixel_9011/SF_IB
+ pixel_9011/PIX_OUT pixel_9011/CSA_VREF pixel
Xpixel_9000 pixel_9000/gring pixel_9000/VDD pixel_9000/GND pixel_9000/VREF pixel_9000/ROW_SEL
+ pixel_9000/NB1 pixel_9000/VBIAS pixel_9000/NB2 pixel_9000/AMP_IN pixel_9000/SF_IB
+ pixel_9000/PIX_OUT pixel_9000/CSA_VREF pixel
Xpixel_9055 pixel_9055/gring pixel_9055/VDD pixel_9055/GND pixel_9055/VREF pixel_9055/ROW_SEL
+ pixel_9055/NB1 pixel_9055/VBIAS pixel_9055/NB2 pixel_9055/AMP_IN pixel_9055/SF_IB
+ pixel_9055/PIX_OUT pixel_9055/CSA_VREF pixel
Xpixel_9044 pixel_9044/gring pixel_9044/VDD pixel_9044/GND pixel_9044/VREF pixel_9044/ROW_SEL
+ pixel_9044/NB1 pixel_9044/VBIAS pixel_9044/NB2 pixel_9044/AMP_IN pixel_9044/SF_IB
+ pixel_9044/PIX_OUT pixel_9044/CSA_VREF pixel
Xpixel_9033 pixel_9033/gring pixel_9033/VDD pixel_9033/GND pixel_9033/VREF pixel_9033/ROW_SEL
+ pixel_9033/NB1 pixel_9033/VBIAS pixel_9033/NB2 pixel_9033/AMP_IN pixel_9033/SF_IB
+ pixel_9033/PIX_OUT pixel_9033/CSA_VREF pixel
Xpixel_8310 pixel_8310/gring pixel_8310/VDD pixel_8310/GND pixel_8310/VREF pixel_8310/ROW_SEL
+ pixel_8310/NB1 pixel_8310/VBIAS pixel_8310/NB2 pixel_8310/AMP_IN pixel_8310/SF_IB
+ pixel_8310/PIX_OUT pixel_8310/CSA_VREF pixel
Xpixel_9088 pixel_9088/gring pixel_9088/VDD pixel_9088/GND pixel_9088/VREF pixel_9088/ROW_SEL
+ pixel_9088/NB1 pixel_9088/VBIAS pixel_9088/NB2 pixel_9088/AMP_IN pixel_9088/SF_IB
+ pixel_9088/PIX_OUT pixel_9088/CSA_VREF pixel
Xpixel_9077 pixel_9077/gring pixel_9077/VDD pixel_9077/GND pixel_9077/VREF pixel_9077/ROW_SEL
+ pixel_9077/NB1 pixel_9077/VBIAS pixel_9077/NB2 pixel_9077/AMP_IN pixel_9077/SF_IB
+ pixel_9077/PIX_OUT pixel_9077/CSA_VREF pixel
Xpixel_9066 pixel_9066/gring pixel_9066/VDD pixel_9066/GND pixel_9066/VREF pixel_9066/ROW_SEL
+ pixel_9066/NB1 pixel_9066/VBIAS pixel_9066/NB2 pixel_9066/AMP_IN pixel_9066/SF_IB
+ pixel_9066/PIX_OUT pixel_9066/CSA_VREF pixel
Xpixel_8321 pixel_8321/gring pixel_8321/VDD pixel_8321/GND pixel_8321/VREF pixel_8321/ROW_SEL
+ pixel_8321/NB1 pixel_8321/VBIAS pixel_8321/NB2 pixel_8321/AMP_IN pixel_8321/SF_IB
+ pixel_8321/PIX_OUT pixel_8321/CSA_VREF pixel
Xpixel_8332 pixel_8332/gring pixel_8332/VDD pixel_8332/GND pixel_8332/VREF pixel_8332/ROW_SEL
+ pixel_8332/NB1 pixel_8332/VBIAS pixel_8332/NB2 pixel_8332/AMP_IN pixel_8332/SF_IB
+ pixel_8332/PIX_OUT pixel_8332/CSA_VREF pixel
Xpixel_8343 pixel_8343/gring pixel_8343/VDD pixel_8343/GND pixel_8343/VREF pixel_8343/ROW_SEL
+ pixel_8343/NB1 pixel_8343/VBIAS pixel_8343/NB2 pixel_8343/AMP_IN pixel_8343/SF_IB
+ pixel_8343/PIX_OUT pixel_8343/CSA_VREF pixel
Xpixel_9099 pixel_9099/gring pixel_9099/VDD pixel_9099/GND pixel_9099/VREF pixel_9099/ROW_SEL
+ pixel_9099/NB1 pixel_9099/VBIAS pixel_9099/NB2 pixel_9099/AMP_IN pixel_9099/SF_IB
+ pixel_9099/PIX_OUT pixel_9099/CSA_VREF pixel
Xpixel_8354 pixel_8354/gring pixel_8354/VDD pixel_8354/GND pixel_8354/VREF pixel_8354/ROW_SEL
+ pixel_8354/NB1 pixel_8354/VBIAS pixel_8354/NB2 pixel_8354/AMP_IN pixel_8354/SF_IB
+ pixel_8354/PIX_OUT pixel_8354/CSA_VREF pixel
Xpixel_8365 pixel_8365/gring pixel_8365/VDD pixel_8365/GND pixel_8365/VREF pixel_8365/ROW_SEL
+ pixel_8365/NB1 pixel_8365/VBIAS pixel_8365/NB2 pixel_8365/AMP_IN pixel_8365/SF_IB
+ pixel_8365/PIX_OUT pixel_8365/CSA_VREF pixel
Xpixel_8376 pixel_8376/gring pixel_8376/VDD pixel_8376/GND pixel_8376/VREF pixel_8376/ROW_SEL
+ pixel_8376/NB1 pixel_8376/VBIAS pixel_8376/NB2 pixel_8376/AMP_IN pixel_8376/SF_IB
+ pixel_8376/PIX_OUT pixel_8376/CSA_VREF pixel
Xpixel_8387 pixel_8387/gring pixel_8387/VDD pixel_8387/GND pixel_8387/VREF pixel_8387/ROW_SEL
+ pixel_8387/NB1 pixel_8387/VBIAS pixel_8387/NB2 pixel_8387/AMP_IN pixel_8387/SF_IB
+ pixel_8387/PIX_OUT pixel_8387/CSA_VREF pixel
Xpixel_7620 pixel_7620/gring pixel_7620/VDD pixel_7620/GND pixel_7620/VREF pixel_7620/ROW_SEL
+ pixel_7620/NB1 pixel_7620/VBIAS pixel_7620/NB2 pixel_7620/AMP_IN pixel_7620/SF_IB
+ pixel_7620/PIX_OUT pixel_7620/CSA_VREF pixel
Xpixel_7631 pixel_7631/gring pixel_7631/VDD pixel_7631/GND pixel_7631/VREF pixel_7631/ROW_SEL
+ pixel_7631/NB1 pixel_7631/VBIAS pixel_7631/NB2 pixel_7631/AMP_IN pixel_7631/SF_IB
+ pixel_7631/PIX_OUT pixel_7631/CSA_VREF pixel
Xpixel_7642 pixel_7642/gring pixel_7642/VDD pixel_7642/GND pixel_7642/VREF pixel_7642/ROW_SEL
+ pixel_7642/NB1 pixel_7642/VBIAS pixel_7642/NB2 pixel_7642/AMP_IN pixel_7642/SF_IB
+ pixel_7642/PIX_OUT pixel_7642/CSA_VREF pixel
Xpixel_8398 pixel_8398/gring pixel_8398/VDD pixel_8398/GND pixel_8398/VREF pixel_8398/ROW_SEL
+ pixel_8398/NB1 pixel_8398/VBIAS pixel_8398/NB2 pixel_8398/AMP_IN pixel_8398/SF_IB
+ pixel_8398/PIX_OUT pixel_8398/CSA_VREF pixel
Xpixel_7653 pixel_7653/gring pixel_7653/VDD pixel_7653/GND pixel_7653/VREF pixel_7653/ROW_SEL
+ pixel_7653/NB1 pixel_7653/VBIAS pixel_7653/NB2 pixel_7653/AMP_IN pixel_7653/SF_IB
+ pixel_7653/PIX_OUT pixel_7653/CSA_VREF pixel
Xpixel_7664 pixel_7664/gring pixel_7664/VDD pixel_7664/GND pixel_7664/VREF pixel_7664/ROW_SEL
+ pixel_7664/NB1 pixel_7664/VBIAS pixel_7664/NB2 pixel_7664/AMP_IN pixel_7664/SF_IB
+ pixel_7664/PIX_OUT pixel_7664/CSA_VREF pixel
Xpixel_7675 pixel_7675/gring pixel_7675/VDD pixel_7675/GND pixel_7675/VREF pixel_7675/ROW_SEL
+ pixel_7675/NB1 pixel_7675/VBIAS pixel_7675/NB2 pixel_7675/AMP_IN pixel_7675/SF_IB
+ pixel_7675/PIX_OUT pixel_7675/CSA_VREF pixel
Xpixel_6930 pixel_6930/gring pixel_6930/VDD pixel_6930/GND pixel_6930/VREF pixel_6930/ROW_SEL
+ pixel_6930/NB1 pixel_6930/VBIAS pixel_6930/NB2 pixel_6930/AMP_IN pixel_6930/SF_IB
+ pixel_6930/PIX_OUT pixel_6930/CSA_VREF pixel
Xpixel_11 pixel_11/gring pixel_11/VDD pixel_11/GND pixel_11/VREF pixel_11/ROW_SEL
+ pixel_11/NB1 pixel_11/VBIAS pixel_11/NB2 pixel_11/AMP_IN pixel_11/SF_IB pixel_11/PIX_OUT
+ pixel_11/CSA_VREF pixel
Xpixel_7686 pixel_7686/gring pixel_7686/VDD pixel_7686/GND pixel_7686/VREF pixel_7686/ROW_SEL
+ pixel_7686/NB1 pixel_7686/VBIAS pixel_7686/NB2 pixel_7686/AMP_IN pixel_7686/SF_IB
+ pixel_7686/PIX_OUT pixel_7686/CSA_VREF pixel
Xpixel_7697 pixel_7697/gring pixel_7697/VDD pixel_7697/GND pixel_7697/VREF pixel_7697/ROW_SEL
+ pixel_7697/NB1 pixel_7697/VBIAS pixel_7697/NB2 pixel_7697/AMP_IN pixel_7697/SF_IB
+ pixel_7697/PIX_OUT pixel_7697/CSA_VREF pixel
Xpixel_6941 pixel_6941/gring pixel_6941/VDD pixel_6941/GND pixel_6941/VREF pixel_6941/ROW_SEL
+ pixel_6941/NB1 pixel_6941/VBIAS pixel_6941/NB2 pixel_6941/AMP_IN pixel_6941/SF_IB
+ pixel_6941/PIX_OUT pixel_6941/CSA_VREF pixel
Xpixel_6952 pixel_6952/gring pixel_6952/VDD pixel_6952/GND pixel_6952/VREF pixel_6952/ROW_SEL
+ pixel_6952/NB1 pixel_6952/VBIAS pixel_6952/NB2 pixel_6952/AMP_IN pixel_6952/SF_IB
+ pixel_6952/PIX_OUT pixel_6952/CSA_VREF pixel
Xpixel_6963 pixel_6963/gring pixel_6963/VDD pixel_6963/GND pixel_6963/VREF pixel_6963/ROW_SEL
+ pixel_6963/NB1 pixel_6963/VBIAS pixel_6963/NB2 pixel_6963/AMP_IN pixel_6963/SF_IB
+ pixel_6963/PIX_OUT pixel_6963/CSA_VREF pixel
Xpixel_55 pixel_55/gring pixel_55/VDD pixel_55/GND pixel_55/VREF pixel_55/ROW_SEL
+ pixel_55/NB1 pixel_55/VBIAS pixel_55/NB2 pixel_55/AMP_IN pixel_55/SF_IB pixel_55/PIX_OUT
+ pixel_55/CSA_VREF pixel
Xpixel_44 pixel_44/gring pixel_44/VDD pixel_44/GND pixel_44/VREF pixel_44/ROW_SEL
+ pixel_44/NB1 pixel_44/VBIAS pixel_44/NB2 pixel_44/AMP_IN pixel_44/SF_IB pixel_44/PIX_OUT
+ pixel_44/CSA_VREF pixel
Xpixel_33 pixel_33/gring pixel_33/VDD pixel_33/GND pixel_33/VREF pixel_33/ROW_SEL
+ pixel_33/NB1 pixel_33/VBIAS pixel_33/NB2 pixel_33/AMP_IN pixel_33/SF_IB pixel_33/PIX_OUT
+ pixel_33/CSA_VREF pixel
Xpixel_22 pixel_22/gring pixel_22/VDD pixel_22/GND pixel_22/VREF pixel_22/ROW_SEL
+ pixel_22/NB1 pixel_22/VBIAS pixel_22/NB2 pixel_22/AMP_IN pixel_22/SF_IB pixel_22/PIX_OUT
+ pixel_22/CSA_VREF pixel
Xpixel_6974 pixel_6974/gring pixel_6974/VDD pixel_6974/GND pixel_6974/VREF pixel_6974/ROW_SEL
+ pixel_6974/NB1 pixel_6974/VBIAS pixel_6974/NB2 pixel_6974/AMP_IN pixel_6974/SF_IB
+ pixel_6974/PIX_OUT pixel_6974/CSA_VREF pixel
Xpixel_6985 pixel_6985/gring pixel_6985/VDD pixel_6985/GND pixel_6985/VREF pixel_6985/ROW_SEL
+ pixel_6985/NB1 pixel_6985/VBIAS pixel_6985/NB2 pixel_6985/AMP_IN pixel_6985/SF_IB
+ pixel_6985/PIX_OUT pixel_6985/CSA_VREF pixel
Xpixel_6996 pixel_6996/gring pixel_6996/VDD pixel_6996/GND pixel_6996/VREF pixel_6996/ROW_SEL
+ pixel_6996/NB1 pixel_6996/VBIAS pixel_6996/NB2 pixel_6996/AMP_IN pixel_6996/SF_IB
+ pixel_6996/PIX_OUT pixel_6996/CSA_VREF pixel
Xpixel_88 pixel_88/gring pixel_88/VDD pixel_88/GND pixel_88/VREF pixel_88/ROW_SEL
+ pixel_88/NB1 pixel_88/VBIAS pixel_88/NB2 pixel_88/AMP_IN pixel_88/SF_IB pixel_88/PIX_OUT
+ pixel_88/CSA_VREF pixel
Xpixel_77 pixel_77/gring pixel_77/VDD pixel_77/GND pixel_77/VREF pixel_77/ROW_SEL
+ pixel_77/NB1 pixel_77/VBIAS pixel_77/NB2 pixel_77/AMP_IN pixel_77/SF_IB pixel_77/PIX_OUT
+ pixel_77/CSA_VREF pixel
Xpixel_66 pixel_66/gring pixel_66/VDD pixel_66/GND pixel_66/VREF pixel_66/ROW_SEL
+ pixel_66/NB1 pixel_66/VBIAS pixel_66/NB2 pixel_66/AMP_IN pixel_66/SF_IB pixel_66/PIX_OUT
+ pixel_66/CSA_VREF pixel
Xpixel_99 pixel_99/gring pixel_99/VDD pixel_99/GND pixel_99/VREF pixel_99/ROW_SEL
+ pixel_99/NB1 pixel_99/VBIAS pixel_99/NB2 pixel_99/AMP_IN pixel_99/SF_IB pixel_99/PIX_OUT
+ pixel_99/CSA_VREF pixel
Xpixel_1292 pixel_1292/gring pixel_1292/VDD pixel_1292/GND pixel_1292/VREF pixel_1292/ROW_SEL
+ pixel_1292/NB1 pixel_1292/VBIAS pixel_1292/NB2 pixel_1292/AMP_IN pixel_1292/SF_IB
+ pixel_1292/PIX_OUT pixel_1292/CSA_VREF pixel
Xpixel_1281 pixel_1281/gring pixel_1281/VDD pixel_1281/GND pixel_1281/VREF pixel_1281/ROW_SEL
+ pixel_1281/NB1 pixel_1281/VBIAS pixel_1281/NB2 pixel_1281/AMP_IN pixel_1281/SF_IB
+ pixel_1281/PIX_OUT pixel_1281/CSA_VREF pixel
Xpixel_1270 pixel_1270/gring pixel_1270/VDD pixel_1270/GND pixel_1270/VREF pixel_1270/ROW_SEL
+ pixel_1270/NB1 pixel_1270/VBIAS pixel_1270/NB2 pixel_1270/AMP_IN pixel_1270/SF_IB
+ pixel_1270/PIX_OUT pixel_1270/CSA_VREF pixel
Xpixel_329 pixel_329/gring pixel_329/VDD pixel_329/GND pixel_329/VREF pixel_329/ROW_SEL
+ pixel_329/NB1 pixel_329/VBIAS pixel_329/NB2 pixel_329/AMP_IN pixel_329/SF_IB pixel_329/PIX_OUT
+ pixel_329/CSA_VREF pixel
Xpixel_318 pixel_318/gring pixel_318/VDD pixel_318/GND pixel_318/VREF pixel_318/ROW_SEL
+ pixel_318/NB1 pixel_318/VBIAS pixel_318/NB2 pixel_318/AMP_IN pixel_318/SF_IB pixel_318/PIX_OUT
+ pixel_318/CSA_VREF pixel
Xpixel_307 pixel_307/gring pixel_307/VDD pixel_307/GND pixel_307/VREF pixel_307/ROW_SEL
+ pixel_307/NB1 pixel_307/VBIAS pixel_307/NB2 pixel_307/AMP_IN pixel_307/SF_IB pixel_307/PIX_OUT
+ pixel_307/CSA_VREF pixel
Xpixel_6204 pixel_6204/gring pixel_6204/VDD pixel_6204/GND pixel_6204/VREF pixel_6204/ROW_SEL
+ pixel_6204/NB1 pixel_6204/VBIAS pixel_6204/NB2 pixel_6204/AMP_IN pixel_6204/SF_IB
+ pixel_6204/PIX_OUT pixel_6204/CSA_VREF pixel
Xpixel_6215 pixel_6215/gring pixel_6215/VDD pixel_6215/GND pixel_6215/VREF pixel_6215/ROW_SEL
+ pixel_6215/NB1 pixel_6215/VBIAS pixel_6215/NB2 pixel_6215/AMP_IN pixel_6215/SF_IB
+ pixel_6215/PIX_OUT pixel_6215/CSA_VREF pixel
Xpixel_6226 pixel_6226/gring pixel_6226/VDD pixel_6226/GND pixel_6226/VREF pixel_6226/ROW_SEL
+ pixel_6226/NB1 pixel_6226/VBIAS pixel_6226/NB2 pixel_6226/AMP_IN pixel_6226/SF_IB
+ pixel_6226/PIX_OUT pixel_6226/CSA_VREF pixel
Xpixel_6237 pixel_6237/gring pixel_6237/VDD pixel_6237/GND pixel_6237/VREF pixel_6237/ROW_SEL
+ pixel_6237/NB1 pixel_6237/VBIAS pixel_6237/NB2 pixel_6237/AMP_IN pixel_6237/SF_IB
+ pixel_6237/PIX_OUT pixel_6237/CSA_VREF pixel
Xpixel_6248 pixel_6248/gring pixel_6248/VDD pixel_6248/GND pixel_6248/VREF pixel_6248/ROW_SEL
+ pixel_6248/NB1 pixel_6248/VBIAS pixel_6248/NB2 pixel_6248/AMP_IN pixel_6248/SF_IB
+ pixel_6248/PIX_OUT pixel_6248/CSA_VREF pixel
Xpixel_6259 pixel_6259/gring pixel_6259/VDD pixel_6259/GND pixel_6259/VREF pixel_6259/ROW_SEL
+ pixel_6259/NB1 pixel_6259/VBIAS pixel_6259/NB2 pixel_6259/AMP_IN pixel_6259/SF_IB
+ pixel_6259/PIX_OUT pixel_6259/CSA_VREF pixel
Xpixel_5503 pixel_5503/gring pixel_5503/VDD pixel_5503/GND pixel_5503/VREF pixel_5503/ROW_SEL
+ pixel_5503/NB1 pixel_5503/VBIAS pixel_5503/NB2 pixel_5503/AMP_IN pixel_5503/SF_IB
+ pixel_5503/PIX_OUT pixel_5503/CSA_VREF pixel
Xpixel_5514 pixel_5514/gring pixel_5514/VDD pixel_5514/GND pixel_5514/VREF pixel_5514/ROW_SEL
+ pixel_5514/NB1 pixel_5514/VBIAS pixel_5514/NB2 pixel_5514/AMP_IN pixel_5514/SF_IB
+ pixel_5514/PIX_OUT pixel_5514/CSA_VREF pixel
Xpixel_5525 pixel_5525/gring pixel_5525/VDD pixel_5525/GND pixel_5525/VREF pixel_5525/ROW_SEL
+ pixel_5525/NB1 pixel_5525/VBIAS pixel_5525/NB2 pixel_5525/AMP_IN pixel_5525/SF_IB
+ pixel_5525/PIX_OUT pixel_5525/CSA_VREF pixel
Xpixel_5536 pixel_5536/gring pixel_5536/VDD pixel_5536/GND pixel_5536/VREF pixel_5536/ROW_SEL
+ pixel_5536/NB1 pixel_5536/VBIAS pixel_5536/NB2 pixel_5536/AMP_IN pixel_5536/SF_IB
+ pixel_5536/PIX_OUT pixel_5536/CSA_VREF pixel
Xpixel_5547 pixel_5547/gring pixel_5547/VDD pixel_5547/GND pixel_5547/VREF pixel_5547/ROW_SEL
+ pixel_5547/NB1 pixel_5547/VBIAS pixel_5547/NB2 pixel_5547/AMP_IN pixel_5547/SF_IB
+ pixel_5547/PIX_OUT pixel_5547/CSA_VREF pixel
Xpixel_5558 pixel_5558/gring pixel_5558/VDD pixel_5558/GND pixel_5558/VREF pixel_5558/ROW_SEL
+ pixel_5558/NB1 pixel_5558/VBIAS pixel_5558/NB2 pixel_5558/AMP_IN pixel_5558/SF_IB
+ pixel_5558/PIX_OUT pixel_5558/CSA_VREF pixel
Xpixel_4802 pixel_4802/gring pixel_4802/VDD pixel_4802/GND pixel_4802/VREF pixel_4802/ROW_SEL
+ pixel_4802/NB1 pixel_4802/VBIAS pixel_4802/NB2 pixel_4802/AMP_IN pixel_4802/SF_IB
+ pixel_4802/PIX_OUT pixel_4802/CSA_VREF pixel
Xpixel_4813 pixel_4813/gring pixel_4813/VDD pixel_4813/GND pixel_4813/VREF pixel_4813/ROW_SEL
+ pixel_4813/NB1 pixel_4813/VBIAS pixel_4813/NB2 pixel_4813/AMP_IN pixel_4813/SF_IB
+ pixel_4813/PIX_OUT pixel_4813/CSA_VREF pixel
Xpixel_841 pixel_841/gring pixel_841/VDD pixel_841/GND pixel_841/VREF pixel_841/ROW_SEL
+ pixel_841/NB1 pixel_841/VBIAS pixel_841/NB2 pixel_841/AMP_IN pixel_841/SF_IB pixel_841/PIX_OUT
+ pixel_841/CSA_VREF pixel
Xpixel_830 pixel_830/gring pixel_830/VDD pixel_830/GND pixel_830/VREF pixel_830/ROW_SEL
+ pixel_830/NB1 pixel_830/VBIAS pixel_830/NB2 pixel_830/AMP_IN pixel_830/SF_IB pixel_830/PIX_OUT
+ pixel_830/CSA_VREF pixel
Xpixel_5569 pixel_5569/gring pixel_5569/VDD pixel_5569/GND pixel_5569/VREF pixel_5569/ROW_SEL
+ pixel_5569/NB1 pixel_5569/VBIAS pixel_5569/NB2 pixel_5569/AMP_IN pixel_5569/SF_IB
+ pixel_5569/PIX_OUT pixel_5569/CSA_VREF pixel
Xpixel_4824 pixel_4824/gring pixel_4824/VDD pixel_4824/GND pixel_4824/VREF pixel_4824/ROW_SEL
+ pixel_4824/NB1 pixel_4824/VBIAS pixel_4824/NB2 pixel_4824/AMP_IN pixel_4824/SF_IB
+ pixel_4824/PIX_OUT pixel_4824/CSA_VREF pixel
Xpixel_4835 pixel_4835/gring pixel_4835/VDD pixel_4835/GND pixel_4835/VREF pixel_4835/ROW_SEL
+ pixel_4835/NB1 pixel_4835/VBIAS pixel_4835/NB2 pixel_4835/AMP_IN pixel_4835/SF_IB
+ pixel_4835/PIX_OUT pixel_4835/CSA_VREF pixel
Xpixel_4846 pixel_4846/gring pixel_4846/VDD pixel_4846/GND pixel_4846/VREF pixel_4846/ROW_SEL
+ pixel_4846/NB1 pixel_4846/VBIAS pixel_4846/NB2 pixel_4846/AMP_IN pixel_4846/SF_IB
+ pixel_4846/PIX_OUT pixel_4846/CSA_VREF pixel
Xpixel_885 pixel_885/gring pixel_885/VDD pixel_885/GND pixel_885/VREF pixel_885/ROW_SEL
+ pixel_885/NB1 pixel_885/VBIAS pixel_885/NB2 pixel_885/AMP_IN pixel_885/SF_IB pixel_885/PIX_OUT
+ pixel_885/CSA_VREF pixel
Xpixel_874 pixel_874/gring pixel_874/VDD pixel_874/GND pixel_874/VREF pixel_874/ROW_SEL
+ pixel_874/NB1 pixel_874/VBIAS pixel_874/NB2 pixel_874/AMP_IN pixel_874/SF_IB pixel_874/PIX_OUT
+ pixel_874/CSA_VREF pixel
Xpixel_863 pixel_863/gring pixel_863/VDD pixel_863/GND pixel_863/VREF pixel_863/ROW_SEL
+ pixel_863/NB1 pixel_863/VBIAS pixel_863/NB2 pixel_863/AMP_IN pixel_863/SF_IB pixel_863/PIX_OUT
+ pixel_863/CSA_VREF pixel
Xpixel_852 pixel_852/gring pixel_852/VDD pixel_852/GND pixel_852/VREF pixel_852/ROW_SEL
+ pixel_852/NB1 pixel_852/VBIAS pixel_852/NB2 pixel_852/AMP_IN pixel_852/SF_IB pixel_852/PIX_OUT
+ pixel_852/CSA_VREF pixel
Xpixel_4857 pixel_4857/gring pixel_4857/VDD pixel_4857/GND pixel_4857/VREF pixel_4857/ROW_SEL
+ pixel_4857/NB1 pixel_4857/VBIAS pixel_4857/NB2 pixel_4857/AMP_IN pixel_4857/SF_IB
+ pixel_4857/PIX_OUT pixel_4857/CSA_VREF pixel
Xpixel_4868 pixel_4868/gring pixel_4868/VDD pixel_4868/GND pixel_4868/VREF pixel_4868/ROW_SEL
+ pixel_4868/NB1 pixel_4868/VBIAS pixel_4868/NB2 pixel_4868/AMP_IN pixel_4868/SF_IB
+ pixel_4868/PIX_OUT pixel_4868/CSA_VREF pixel
Xpixel_4879 pixel_4879/gring pixel_4879/VDD pixel_4879/GND pixel_4879/VREF pixel_4879/ROW_SEL
+ pixel_4879/NB1 pixel_4879/VBIAS pixel_4879/NB2 pixel_4879/AMP_IN pixel_4879/SF_IB
+ pixel_4879/PIX_OUT pixel_4879/CSA_VREF pixel
Xpixel_896 pixel_896/gring pixel_896/VDD pixel_896/GND pixel_896/VREF pixel_896/ROW_SEL
+ pixel_896/NB1 pixel_896/VBIAS pixel_896/NB2 pixel_896/AMP_IN pixel_896/SF_IB pixel_896/PIX_OUT
+ pixel_896/CSA_VREF pixel
Xpixel_8140 pixel_8140/gring pixel_8140/VDD pixel_8140/GND pixel_8140/VREF pixel_8140/ROW_SEL
+ pixel_8140/NB1 pixel_8140/VBIAS pixel_8140/NB2 pixel_8140/AMP_IN pixel_8140/SF_IB
+ pixel_8140/PIX_OUT pixel_8140/CSA_VREF pixel
Xpixel_8151 pixel_8151/gring pixel_8151/VDD pixel_8151/GND pixel_8151/VREF pixel_8151/ROW_SEL
+ pixel_8151/NB1 pixel_8151/VBIAS pixel_8151/NB2 pixel_8151/AMP_IN pixel_8151/SF_IB
+ pixel_8151/PIX_OUT pixel_8151/CSA_VREF pixel
Xpixel_8162 pixel_8162/gring pixel_8162/VDD pixel_8162/GND pixel_8162/VREF pixel_8162/ROW_SEL
+ pixel_8162/NB1 pixel_8162/VBIAS pixel_8162/NB2 pixel_8162/AMP_IN pixel_8162/SF_IB
+ pixel_8162/PIX_OUT pixel_8162/CSA_VREF pixel
Xpixel_8173 pixel_8173/gring pixel_8173/VDD pixel_8173/GND pixel_8173/VREF pixel_8173/ROW_SEL
+ pixel_8173/NB1 pixel_8173/VBIAS pixel_8173/NB2 pixel_8173/AMP_IN pixel_8173/SF_IB
+ pixel_8173/PIX_OUT pixel_8173/CSA_VREF pixel
Xpixel_8184 pixel_8184/gring pixel_8184/VDD pixel_8184/GND pixel_8184/VREF pixel_8184/ROW_SEL
+ pixel_8184/NB1 pixel_8184/VBIAS pixel_8184/NB2 pixel_8184/AMP_IN pixel_8184/SF_IB
+ pixel_8184/PIX_OUT pixel_8184/CSA_VREF pixel
Xpixel_8195 pixel_8195/gring pixel_8195/VDD pixel_8195/GND pixel_8195/VREF pixel_8195/ROW_SEL
+ pixel_8195/NB1 pixel_8195/VBIAS pixel_8195/NB2 pixel_8195/AMP_IN pixel_8195/SF_IB
+ pixel_8195/PIX_OUT pixel_8195/CSA_VREF pixel
Xpixel_7450 pixel_7450/gring pixel_7450/VDD pixel_7450/GND pixel_7450/VREF pixel_7450/ROW_SEL
+ pixel_7450/NB1 pixel_7450/VBIAS pixel_7450/NB2 pixel_7450/AMP_IN pixel_7450/SF_IB
+ pixel_7450/PIX_OUT pixel_7450/CSA_VREF pixel
Xpixel_7461 pixel_7461/gring pixel_7461/VDD pixel_7461/GND pixel_7461/VREF pixel_7461/ROW_SEL
+ pixel_7461/NB1 pixel_7461/VBIAS pixel_7461/NB2 pixel_7461/AMP_IN pixel_7461/SF_IB
+ pixel_7461/PIX_OUT pixel_7461/CSA_VREF pixel
Xpixel_7472 pixel_7472/gring pixel_7472/VDD pixel_7472/GND pixel_7472/VREF pixel_7472/ROW_SEL
+ pixel_7472/NB1 pixel_7472/VBIAS pixel_7472/NB2 pixel_7472/AMP_IN pixel_7472/SF_IB
+ pixel_7472/PIX_OUT pixel_7472/CSA_VREF pixel
Xpixel_7483 pixel_7483/gring pixel_7483/VDD pixel_7483/GND pixel_7483/VREF pixel_7483/ROW_SEL
+ pixel_7483/NB1 pixel_7483/VBIAS pixel_7483/NB2 pixel_7483/AMP_IN pixel_7483/SF_IB
+ pixel_7483/PIX_OUT pixel_7483/CSA_VREF pixel
Xpixel_7494 pixel_7494/gring pixel_7494/VDD pixel_7494/GND pixel_7494/VREF pixel_7494/ROW_SEL
+ pixel_7494/NB1 pixel_7494/VBIAS pixel_7494/NB2 pixel_7494/AMP_IN pixel_7494/SF_IB
+ pixel_7494/PIX_OUT pixel_7494/CSA_VREF pixel
Xpixel_6760 pixel_6760/gring pixel_6760/VDD pixel_6760/GND pixel_6760/VREF pixel_6760/ROW_SEL
+ pixel_6760/NB1 pixel_6760/VBIAS pixel_6760/NB2 pixel_6760/AMP_IN pixel_6760/SF_IB
+ pixel_6760/PIX_OUT pixel_6760/CSA_VREF pixel
Xpixel_6771 pixel_6771/gring pixel_6771/VDD pixel_6771/GND pixel_6771/VREF pixel_6771/ROW_SEL
+ pixel_6771/NB1 pixel_6771/VBIAS pixel_6771/NB2 pixel_6771/AMP_IN pixel_6771/SF_IB
+ pixel_6771/PIX_OUT pixel_6771/CSA_VREF pixel
Xpixel_6782 pixel_6782/gring pixel_6782/VDD pixel_6782/GND pixel_6782/VREF pixel_6782/ROW_SEL
+ pixel_6782/NB1 pixel_6782/VBIAS pixel_6782/NB2 pixel_6782/AMP_IN pixel_6782/SF_IB
+ pixel_6782/PIX_OUT pixel_6782/CSA_VREF pixel
Xpixel_6793 pixel_6793/gring pixel_6793/VDD pixel_6793/GND pixel_6793/VREF pixel_6793/ROW_SEL
+ pixel_6793/NB1 pixel_6793/VBIAS pixel_6793/NB2 pixel_6793/AMP_IN pixel_6793/SF_IB
+ pixel_6793/PIX_OUT pixel_6793/CSA_VREF pixel
Xpixel_104 pixel_104/gring pixel_104/VDD pixel_104/GND pixel_104/VREF pixel_104/ROW_SEL
+ pixel_104/NB1 pixel_104/VBIAS pixel_104/NB2 pixel_104/AMP_IN pixel_104/SF_IB pixel_104/PIX_OUT
+ pixel_104/CSA_VREF pixel
Xpixel_137 pixel_137/gring pixel_137/VDD pixel_137/GND pixel_137/VREF pixel_137/ROW_SEL
+ pixel_137/NB1 pixel_137/VBIAS pixel_137/NB2 pixel_137/AMP_IN pixel_137/SF_IB pixel_137/PIX_OUT
+ pixel_137/CSA_VREF pixel
Xpixel_126 pixel_126/gring pixel_126/VDD pixel_126/GND pixel_126/VREF pixel_126/ROW_SEL
+ pixel_126/NB1 pixel_126/VBIAS pixel_126/NB2 pixel_126/AMP_IN pixel_126/SF_IB pixel_126/PIX_OUT
+ pixel_126/CSA_VREF pixel
Xpixel_115 pixel_115/gring pixel_115/VDD pixel_115/GND pixel_115/VREF pixel_115/ROW_SEL
+ pixel_115/NB1 pixel_115/VBIAS pixel_115/NB2 pixel_115/AMP_IN pixel_115/SF_IB pixel_115/PIX_OUT
+ pixel_115/CSA_VREF pixel
Xpixel_4109 pixel_4109/gring pixel_4109/VDD pixel_4109/GND pixel_4109/VREF pixel_4109/ROW_SEL
+ pixel_4109/NB1 pixel_4109/VBIAS pixel_4109/NB2 pixel_4109/AMP_IN pixel_4109/SF_IB
+ pixel_4109/PIX_OUT pixel_4109/CSA_VREF pixel
Xpixel_159 pixel_159/gring pixel_159/VDD pixel_159/GND pixel_159/VREF pixel_159/ROW_SEL
+ pixel_159/NB1 pixel_159/VBIAS pixel_159/NB2 pixel_159/AMP_IN pixel_159/SF_IB pixel_159/PIX_OUT
+ pixel_159/CSA_VREF pixel
Xpixel_148 pixel_148/gring pixel_148/VDD pixel_148/GND pixel_148/VREF pixel_148/ROW_SEL
+ pixel_148/NB1 pixel_148/VBIAS pixel_148/NB2 pixel_148/AMP_IN pixel_148/SF_IB pixel_148/PIX_OUT
+ pixel_148/CSA_VREF pixel
Xpixel_3419 pixel_3419/gring pixel_3419/VDD pixel_3419/GND pixel_3419/VREF pixel_3419/ROW_SEL
+ pixel_3419/NB1 pixel_3419/VBIAS pixel_3419/NB2 pixel_3419/AMP_IN pixel_3419/SF_IB
+ pixel_3419/PIX_OUT pixel_3419/CSA_VREF pixel
Xpixel_3408 pixel_3408/gring pixel_3408/VDD pixel_3408/GND pixel_3408/VREF pixel_3408/ROW_SEL
+ pixel_3408/NB1 pixel_3408/VBIAS pixel_3408/NB2 pixel_3408/AMP_IN pixel_3408/SF_IB
+ pixel_3408/PIX_OUT pixel_3408/CSA_VREF pixel
Xpixel_2729 pixel_2729/gring pixel_2729/VDD pixel_2729/GND pixel_2729/VREF pixel_2729/ROW_SEL
+ pixel_2729/NB1 pixel_2729/VBIAS pixel_2729/NB2 pixel_2729/AMP_IN pixel_2729/SF_IB
+ pixel_2729/PIX_OUT pixel_2729/CSA_VREF pixel
Xpixel_2718 pixel_2718/gring pixel_2718/VDD pixel_2718/GND pixel_2718/VREF pixel_2718/ROW_SEL
+ pixel_2718/NB1 pixel_2718/VBIAS pixel_2718/NB2 pixel_2718/AMP_IN pixel_2718/SF_IB
+ pixel_2718/PIX_OUT pixel_2718/CSA_VREF pixel
Xpixel_2707 pixel_2707/gring pixel_2707/VDD pixel_2707/GND pixel_2707/VREF pixel_2707/ROW_SEL
+ pixel_2707/NB1 pixel_2707/VBIAS pixel_2707/NB2 pixel_2707/AMP_IN pixel_2707/SF_IB
+ pixel_2707/PIX_OUT pixel_2707/CSA_VREF pixel
Xpixel_6001 pixel_6001/gring pixel_6001/VDD pixel_6001/GND pixel_6001/VREF pixel_6001/ROW_SEL
+ pixel_6001/NB1 pixel_6001/VBIAS pixel_6001/NB2 pixel_6001/AMP_IN pixel_6001/SF_IB
+ pixel_6001/PIX_OUT pixel_6001/CSA_VREF pixel
Xpixel_6012 pixel_6012/gring pixel_6012/VDD pixel_6012/GND pixel_6012/VREF pixel_6012/ROW_SEL
+ pixel_6012/NB1 pixel_6012/VBIAS pixel_6012/NB2 pixel_6012/AMP_IN pixel_6012/SF_IB
+ pixel_6012/PIX_OUT pixel_6012/CSA_VREF pixel
Xpixel_6023 pixel_6023/gring pixel_6023/VDD pixel_6023/GND pixel_6023/VREF pixel_6023/ROW_SEL
+ pixel_6023/NB1 pixel_6023/VBIAS pixel_6023/NB2 pixel_6023/AMP_IN pixel_6023/SF_IB
+ pixel_6023/PIX_OUT pixel_6023/CSA_VREF pixel
Xpixel_6034 pixel_6034/gring pixel_6034/VDD pixel_6034/GND pixel_6034/VREF pixel_6034/ROW_SEL
+ pixel_6034/NB1 pixel_6034/VBIAS pixel_6034/NB2 pixel_6034/AMP_IN pixel_6034/SF_IB
+ pixel_6034/PIX_OUT pixel_6034/CSA_VREF pixel
Xpixel_6045 pixel_6045/gring pixel_6045/VDD pixel_6045/GND pixel_6045/VREF pixel_6045/ROW_SEL
+ pixel_6045/NB1 pixel_6045/VBIAS pixel_6045/NB2 pixel_6045/AMP_IN pixel_6045/SF_IB
+ pixel_6045/PIX_OUT pixel_6045/CSA_VREF pixel
Xpixel_6056 pixel_6056/gring pixel_6056/VDD pixel_6056/GND pixel_6056/VREF pixel_6056/ROW_SEL
+ pixel_6056/NB1 pixel_6056/VBIAS pixel_6056/NB2 pixel_6056/AMP_IN pixel_6056/SF_IB
+ pixel_6056/PIX_OUT pixel_6056/CSA_VREF pixel
Xpixel_6067 pixel_6067/gring pixel_6067/VDD pixel_6067/GND pixel_6067/VREF pixel_6067/ROW_SEL
+ pixel_6067/NB1 pixel_6067/VBIAS pixel_6067/NB2 pixel_6067/AMP_IN pixel_6067/SF_IB
+ pixel_6067/PIX_OUT pixel_6067/CSA_VREF pixel
Xpixel_5300 pixel_5300/gring pixel_5300/VDD pixel_5300/GND pixel_5300/VREF pixel_5300/ROW_SEL
+ pixel_5300/NB1 pixel_5300/VBIAS pixel_5300/NB2 pixel_5300/AMP_IN pixel_5300/SF_IB
+ pixel_5300/PIX_OUT pixel_5300/CSA_VREF pixel
Xpixel_5311 pixel_5311/gring pixel_5311/VDD pixel_5311/GND pixel_5311/VREF pixel_5311/ROW_SEL
+ pixel_5311/NB1 pixel_5311/VBIAS pixel_5311/NB2 pixel_5311/AMP_IN pixel_5311/SF_IB
+ pixel_5311/PIX_OUT pixel_5311/CSA_VREF pixel
Xpixel_5322 pixel_5322/gring pixel_5322/VDD pixel_5322/GND pixel_5322/VREF pixel_5322/ROW_SEL
+ pixel_5322/NB1 pixel_5322/VBIAS pixel_5322/NB2 pixel_5322/AMP_IN pixel_5322/SF_IB
+ pixel_5322/PIX_OUT pixel_5322/CSA_VREF pixel
Xpixel_6078 pixel_6078/gring pixel_6078/VDD pixel_6078/GND pixel_6078/VREF pixel_6078/ROW_SEL
+ pixel_6078/NB1 pixel_6078/VBIAS pixel_6078/NB2 pixel_6078/AMP_IN pixel_6078/SF_IB
+ pixel_6078/PIX_OUT pixel_6078/CSA_VREF pixel
Xpixel_6089 pixel_6089/gring pixel_6089/VDD pixel_6089/GND pixel_6089/VREF pixel_6089/ROW_SEL
+ pixel_6089/NB1 pixel_6089/VBIAS pixel_6089/NB2 pixel_6089/AMP_IN pixel_6089/SF_IB
+ pixel_6089/PIX_OUT pixel_6089/CSA_VREF pixel
Xpixel_5333 pixel_5333/gring pixel_5333/VDD pixel_5333/GND pixel_5333/VREF pixel_5333/ROW_SEL
+ pixel_5333/NB1 pixel_5333/VBIAS pixel_5333/NB2 pixel_5333/AMP_IN pixel_5333/SF_IB
+ pixel_5333/PIX_OUT pixel_5333/CSA_VREF pixel
Xpixel_5344 pixel_5344/gring pixel_5344/VDD pixel_5344/GND pixel_5344/VREF pixel_5344/ROW_SEL
+ pixel_5344/NB1 pixel_5344/VBIAS pixel_5344/NB2 pixel_5344/AMP_IN pixel_5344/SF_IB
+ pixel_5344/PIX_OUT pixel_5344/CSA_VREF pixel
Xpixel_5355 pixel_5355/gring pixel_5355/VDD pixel_5355/GND pixel_5355/VREF pixel_5355/ROW_SEL
+ pixel_5355/NB1 pixel_5355/VBIAS pixel_5355/NB2 pixel_5355/AMP_IN pixel_5355/SF_IB
+ pixel_5355/PIX_OUT pixel_5355/CSA_VREF pixel
Xpixel_5366 pixel_5366/gring pixel_5366/VDD pixel_5366/GND pixel_5366/VREF pixel_5366/ROW_SEL
+ pixel_5366/NB1 pixel_5366/VBIAS pixel_5366/NB2 pixel_5366/AMP_IN pixel_5366/SF_IB
+ pixel_5366/PIX_OUT pixel_5366/CSA_VREF pixel
Xpixel_4610 pixel_4610/gring pixel_4610/VDD pixel_4610/GND pixel_4610/VREF pixel_4610/ROW_SEL
+ pixel_4610/NB1 pixel_4610/VBIAS pixel_4610/NB2 pixel_4610/AMP_IN pixel_4610/SF_IB
+ pixel_4610/PIX_OUT pixel_4610/CSA_VREF pixel
Xpixel_4621 pixel_4621/gring pixel_4621/VDD pixel_4621/GND pixel_4621/VREF pixel_4621/ROW_SEL
+ pixel_4621/NB1 pixel_4621/VBIAS pixel_4621/NB2 pixel_4621/AMP_IN pixel_4621/SF_IB
+ pixel_4621/PIX_OUT pixel_4621/CSA_VREF pixel
Xpixel_5377 pixel_5377/gring pixel_5377/VDD pixel_5377/GND pixel_5377/VREF pixel_5377/ROW_SEL
+ pixel_5377/NB1 pixel_5377/VBIAS pixel_5377/NB2 pixel_5377/AMP_IN pixel_5377/SF_IB
+ pixel_5377/PIX_OUT pixel_5377/CSA_VREF pixel
Xpixel_5388 pixel_5388/gring pixel_5388/VDD pixel_5388/GND pixel_5388/VREF pixel_5388/ROW_SEL
+ pixel_5388/NB1 pixel_5388/VBIAS pixel_5388/NB2 pixel_5388/AMP_IN pixel_5388/SF_IB
+ pixel_5388/PIX_OUT pixel_5388/CSA_VREF pixel
Xpixel_5399 pixel_5399/gring pixel_5399/VDD pixel_5399/GND pixel_5399/VREF pixel_5399/ROW_SEL
+ pixel_5399/NB1 pixel_5399/VBIAS pixel_5399/NB2 pixel_5399/AMP_IN pixel_5399/SF_IB
+ pixel_5399/PIX_OUT pixel_5399/CSA_VREF pixel
Xpixel_4632 pixel_4632/gring pixel_4632/VDD pixel_4632/GND pixel_4632/VREF pixel_4632/ROW_SEL
+ pixel_4632/NB1 pixel_4632/VBIAS pixel_4632/NB2 pixel_4632/AMP_IN pixel_4632/SF_IB
+ pixel_4632/PIX_OUT pixel_4632/CSA_VREF pixel
Xpixel_4643 pixel_4643/gring pixel_4643/VDD pixel_4643/GND pixel_4643/VREF pixel_4643/ROW_SEL
+ pixel_4643/NB1 pixel_4643/VBIAS pixel_4643/NB2 pixel_4643/AMP_IN pixel_4643/SF_IB
+ pixel_4643/PIX_OUT pixel_4643/CSA_VREF pixel
Xpixel_4654 pixel_4654/gring pixel_4654/VDD pixel_4654/GND pixel_4654/VREF pixel_4654/ROW_SEL
+ pixel_4654/NB1 pixel_4654/VBIAS pixel_4654/NB2 pixel_4654/AMP_IN pixel_4654/SF_IB
+ pixel_4654/PIX_OUT pixel_4654/CSA_VREF pixel
Xpixel_693 pixel_693/gring pixel_693/VDD pixel_693/GND pixel_693/VREF pixel_693/ROW_SEL
+ pixel_693/NB1 pixel_693/VBIAS pixel_693/NB2 pixel_693/AMP_IN pixel_693/SF_IB pixel_693/PIX_OUT
+ pixel_693/CSA_VREF pixel
Xpixel_682 pixel_682/gring pixel_682/VDD pixel_682/GND pixel_682/VREF pixel_682/ROW_SEL
+ pixel_682/NB1 pixel_682/VBIAS pixel_682/NB2 pixel_682/AMP_IN pixel_682/SF_IB pixel_682/PIX_OUT
+ pixel_682/CSA_VREF pixel
Xpixel_671 pixel_671/gring pixel_671/VDD pixel_671/GND pixel_671/VREF pixel_671/ROW_SEL
+ pixel_671/NB1 pixel_671/VBIAS pixel_671/NB2 pixel_671/AMP_IN pixel_671/SF_IB pixel_671/PIX_OUT
+ pixel_671/CSA_VREF pixel
Xpixel_660 pixel_660/gring pixel_660/VDD pixel_660/GND pixel_660/VREF pixel_660/ROW_SEL
+ pixel_660/NB1 pixel_660/VBIAS pixel_660/NB2 pixel_660/AMP_IN pixel_660/SF_IB pixel_660/PIX_OUT
+ pixel_660/CSA_VREF pixel
Xpixel_4665 pixel_4665/gring pixel_4665/VDD pixel_4665/GND pixel_4665/VREF pixel_4665/ROW_SEL
+ pixel_4665/NB1 pixel_4665/VBIAS pixel_4665/NB2 pixel_4665/AMP_IN pixel_4665/SF_IB
+ pixel_4665/PIX_OUT pixel_4665/CSA_VREF pixel
Xpixel_4676 pixel_4676/gring pixel_4676/VDD pixel_4676/GND pixel_4676/VREF pixel_4676/ROW_SEL
+ pixel_4676/NB1 pixel_4676/VBIAS pixel_4676/NB2 pixel_4676/AMP_IN pixel_4676/SF_IB
+ pixel_4676/PIX_OUT pixel_4676/CSA_VREF pixel
Xpixel_4687 pixel_4687/gring pixel_4687/VDD pixel_4687/GND pixel_4687/VREF pixel_4687/ROW_SEL
+ pixel_4687/NB1 pixel_4687/VBIAS pixel_4687/NB2 pixel_4687/AMP_IN pixel_4687/SF_IB
+ pixel_4687/PIX_OUT pixel_4687/CSA_VREF pixel
Xpixel_4698 pixel_4698/gring pixel_4698/VDD pixel_4698/GND pixel_4698/VREF pixel_4698/ROW_SEL
+ pixel_4698/NB1 pixel_4698/VBIAS pixel_4698/NB2 pixel_4698/AMP_IN pixel_4698/SF_IB
+ pixel_4698/PIX_OUT pixel_4698/CSA_VREF pixel
Xpixel_3920 pixel_3920/gring pixel_3920/VDD pixel_3920/GND pixel_3920/VREF pixel_3920/ROW_SEL
+ pixel_3920/NB1 pixel_3920/VBIAS pixel_3920/NB2 pixel_3920/AMP_IN pixel_3920/SF_IB
+ pixel_3920/PIX_OUT pixel_3920/CSA_VREF pixel
Xpixel_3931 pixel_3931/gring pixel_3931/VDD pixel_3931/GND pixel_3931/VREF pixel_3931/ROW_SEL
+ pixel_3931/NB1 pixel_3931/VBIAS pixel_3931/NB2 pixel_3931/AMP_IN pixel_3931/SF_IB
+ pixel_3931/PIX_OUT pixel_3931/CSA_VREF pixel
Xpixel_3942 pixel_3942/gring pixel_3942/VDD pixel_3942/GND pixel_3942/VREF pixel_3942/ROW_SEL
+ pixel_3942/NB1 pixel_3942/VBIAS pixel_3942/NB2 pixel_3942/AMP_IN pixel_3942/SF_IB
+ pixel_3942/PIX_OUT pixel_3942/CSA_VREF pixel
Xpixel_3953 pixel_3953/gring pixel_3953/VDD pixel_3953/GND pixel_3953/VREF pixel_3953/ROW_SEL
+ pixel_3953/NB1 pixel_3953/VBIAS pixel_3953/NB2 pixel_3953/AMP_IN pixel_3953/SF_IB
+ pixel_3953/PIX_OUT pixel_3953/CSA_VREF pixel
Xpixel_3964 pixel_3964/gring pixel_3964/VDD pixel_3964/GND pixel_3964/VREF pixel_3964/ROW_SEL
+ pixel_3964/NB1 pixel_3964/VBIAS pixel_3964/NB2 pixel_3964/AMP_IN pixel_3964/SF_IB
+ pixel_3964/PIX_OUT pixel_3964/CSA_VREF pixel
Xpixel_3975 pixel_3975/gring pixel_3975/VDD pixel_3975/GND pixel_3975/VREF pixel_3975/ROW_SEL
+ pixel_3975/NB1 pixel_3975/VBIAS pixel_3975/NB2 pixel_3975/AMP_IN pixel_3975/SF_IB
+ pixel_3975/PIX_OUT pixel_3975/CSA_VREF pixel
Xpixel_3986 pixel_3986/gring pixel_3986/VDD pixel_3986/GND pixel_3986/VREF pixel_3986/ROW_SEL
+ pixel_3986/NB1 pixel_3986/VBIAS pixel_3986/NB2 pixel_3986/AMP_IN pixel_3986/SF_IB
+ pixel_3986/PIX_OUT pixel_3986/CSA_VREF pixel
Xpixel_3997 pixel_3997/gring pixel_3997/VDD pixel_3997/GND pixel_3997/VREF pixel_3997/ROW_SEL
+ pixel_3997/NB1 pixel_3997/VBIAS pixel_3997/NB2 pixel_3997/AMP_IN pixel_3997/SF_IB
+ pixel_3997/PIX_OUT pixel_3997/CSA_VREF pixel
Xpixel_7 pixel_7/gring pixel_7/VDD pixel_7/GND pixel_7/VREF pixel_7/ROW_SEL pixel_7/NB1
+ pixel_7/VBIAS pixel_7/NB2 pixel_7/AMP_IN pixel_7/SF_IB pixel_7/PIX_OUT pixel_7/CSA_VREF
+ pixel
Xpixel_7280 pixel_7280/gring pixel_7280/VDD pixel_7280/GND pixel_7280/VREF pixel_7280/ROW_SEL
+ pixel_7280/NB1 pixel_7280/VBIAS pixel_7280/NB2 pixel_7280/AMP_IN pixel_7280/SF_IB
+ pixel_7280/PIX_OUT pixel_7280/CSA_VREF pixel
Xpixel_7291 pixel_7291/gring pixel_7291/VDD pixel_7291/GND pixel_7291/VREF pixel_7291/ROW_SEL
+ pixel_7291/NB1 pixel_7291/VBIAS pixel_7291/NB2 pixel_7291/AMP_IN pixel_7291/SF_IB
+ pixel_7291/PIX_OUT pixel_7291/CSA_VREF pixel
Xpixel_6590 pixel_6590/gring pixel_6590/VDD pixel_6590/GND pixel_6590/VREF pixel_6590/ROW_SEL
+ pixel_6590/NB1 pixel_6590/VBIAS pixel_6590/NB2 pixel_6590/AMP_IN pixel_6590/SF_IB
+ pixel_6590/PIX_OUT pixel_6590/CSA_VREF pixel
Xpixel_8909 pixel_8909/gring pixel_8909/VDD pixel_8909/GND pixel_8909/VREF pixel_8909/ROW_SEL
+ pixel_8909/NB1 pixel_8909/VBIAS pixel_8909/NB2 pixel_8909/AMP_IN pixel_8909/SF_IB
+ pixel_8909/PIX_OUT pixel_8909/CSA_VREF pixel
Xpixel_3205 pixel_3205/gring pixel_3205/VDD pixel_3205/GND pixel_3205/VREF pixel_3205/ROW_SEL
+ pixel_3205/NB1 pixel_3205/VBIAS pixel_3205/NB2 pixel_3205/AMP_IN pixel_3205/SF_IB
+ pixel_3205/PIX_OUT pixel_3205/CSA_VREF pixel
Xpixel_3238 pixel_3238/gring pixel_3238/VDD pixel_3238/GND pixel_3238/VREF pixel_3238/ROW_SEL
+ pixel_3238/NB1 pixel_3238/VBIAS pixel_3238/NB2 pixel_3238/AMP_IN pixel_3238/SF_IB
+ pixel_3238/PIX_OUT pixel_3238/CSA_VREF pixel
Xpixel_3227 pixel_3227/gring pixel_3227/VDD pixel_3227/GND pixel_3227/VREF pixel_3227/ROW_SEL
+ pixel_3227/NB1 pixel_3227/VBIAS pixel_3227/NB2 pixel_3227/AMP_IN pixel_3227/SF_IB
+ pixel_3227/PIX_OUT pixel_3227/CSA_VREF pixel
Xpixel_3216 pixel_3216/gring pixel_3216/VDD pixel_3216/GND pixel_3216/VREF pixel_3216/ROW_SEL
+ pixel_3216/NB1 pixel_3216/VBIAS pixel_3216/NB2 pixel_3216/AMP_IN pixel_3216/SF_IB
+ pixel_3216/PIX_OUT pixel_3216/CSA_VREF pixel
Xpixel_2537 pixel_2537/gring pixel_2537/VDD pixel_2537/GND pixel_2537/VREF pixel_2537/ROW_SEL
+ pixel_2537/NB1 pixel_2537/VBIAS pixel_2537/NB2 pixel_2537/AMP_IN pixel_2537/SF_IB
+ pixel_2537/PIX_OUT pixel_2537/CSA_VREF pixel
Xpixel_2526 pixel_2526/gring pixel_2526/VDD pixel_2526/GND pixel_2526/VREF pixel_2526/ROW_SEL
+ pixel_2526/NB1 pixel_2526/VBIAS pixel_2526/NB2 pixel_2526/AMP_IN pixel_2526/SF_IB
+ pixel_2526/PIX_OUT pixel_2526/CSA_VREF pixel
Xpixel_2515 pixel_2515/gring pixel_2515/VDD pixel_2515/GND pixel_2515/VREF pixel_2515/ROW_SEL
+ pixel_2515/NB1 pixel_2515/VBIAS pixel_2515/NB2 pixel_2515/AMP_IN pixel_2515/SF_IB
+ pixel_2515/PIX_OUT pixel_2515/CSA_VREF pixel
Xpixel_2504 pixel_2504/gring pixel_2504/VDD pixel_2504/GND pixel_2504/VREF pixel_2504/ROW_SEL
+ pixel_2504/NB1 pixel_2504/VBIAS pixel_2504/NB2 pixel_2504/AMP_IN pixel_2504/SF_IB
+ pixel_2504/PIX_OUT pixel_2504/CSA_VREF pixel
Xpixel_3249 pixel_3249/gring pixel_3249/VDD pixel_3249/GND pixel_3249/VREF pixel_3249/ROW_SEL
+ pixel_3249/NB1 pixel_3249/VBIAS pixel_3249/NB2 pixel_3249/AMP_IN pixel_3249/SF_IB
+ pixel_3249/PIX_OUT pixel_3249/CSA_VREF pixel
Xpixel_1825 pixel_1825/gring pixel_1825/VDD pixel_1825/GND pixel_1825/VREF pixel_1825/ROW_SEL
+ pixel_1825/NB1 pixel_1825/VBIAS pixel_1825/NB2 pixel_1825/AMP_IN pixel_1825/SF_IB
+ pixel_1825/PIX_OUT pixel_1825/CSA_VREF pixel
Xpixel_1814 pixel_1814/gring pixel_1814/VDD pixel_1814/GND pixel_1814/VREF pixel_1814/ROW_SEL
+ pixel_1814/NB1 pixel_1814/VBIAS pixel_1814/NB2 pixel_1814/AMP_IN pixel_1814/SF_IB
+ pixel_1814/PIX_OUT pixel_1814/CSA_VREF pixel
Xpixel_1803 pixel_1803/gring pixel_1803/VDD pixel_1803/GND pixel_1803/VREF pixel_1803/ROW_SEL
+ pixel_1803/NB1 pixel_1803/VBIAS pixel_1803/NB2 pixel_1803/AMP_IN pixel_1803/SF_IB
+ pixel_1803/PIX_OUT pixel_1803/CSA_VREF pixel
Xpixel_2559 pixel_2559/gring pixel_2559/VDD pixel_2559/GND pixel_2559/VREF pixel_2559/ROW_SEL
+ pixel_2559/NB1 pixel_2559/VBIAS pixel_2559/NB2 pixel_2559/AMP_IN pixel_2559/SF_IB
+ pixel_2559/PIX_OUT pixel_2559/CSA_VREF pixel
Xpixel_2548 pixel_2548/gring pixel_2548/VDD pixel_2548/GND pixel_2548/VREF pixel_2548/ROW_SEL
+ pixel_2548/NB1 pixel_2548/VBIAS pixel_2548/NB2 pixel_2548/AMP_IN pixel_2548/SF_IB
+ pixel_2548/PIX_OUT pixel_2548/CSA_VREF pixel
Xpixel_1869 pixel_1869/gring pixel_1869/VDD pixel_1869/GND pixel_1869/VREF pixel_1869/ROW_SEL
+ pixel_1869/NB1 pixel_1869/VBIAS pixel_1869/NB2 pixel_1869/AMP_IN pixel_1869/SF_IB
+ pixel_1869/PIX_OUT pixel_1869/CSA_VREF pixel
Xpixel_1858 pixel_1858/gring pixel_1858/VDD pixel_1858/GND pixel_1858/VREF pixel_1858/ROW_SEL
+ pixel_1858/NB1 pixel_1858/VBIAS pixel_1858/NB2 pixel_1858/AMP_IN pixel_1858/SF_IB
+ pixel_1858/PIX_OUT pixel_1858/CSA_VREF pixel
Xpixel_1847 pixel_1847/gring pixel_1847/VDD pixel_1847/GND pixel_1847/VREF pixel_1847/ROW_SEL
+ pixel_1847/NB1 pixel_1847/VBIAS pixel_1847/NB2 pixel_1847/AMP_IN pixel_1847/SF_IB
+ pixel_1847/PIX_OUT pixel_1847/CSA_VREF pixel
Xpixel_1836 pixel_1836/gring pixel_1836/VDD pixel_1836/GND pixel_1836/VREF pixel_1836/ROW_SEL
+ pixel_1836/NB1 pixel_1836/VBIAS pixel_1836/NB2 pixel_1836/AMP_IN pixel_1836/SF_IB
+ pixel_1836/PIX_OUT pixel_1836/CSA_VREF pixel
Xpixel_5130 pixel_5130/gring pixel_5130/VDD pixel_5130/GND pixel_5130/VREF pixel_5130/ROW_SEL
+ pixel_5130/NB1 pixel_5130/VBIAS pixel_5130/NB2 pixel_5130/AMP_IN pixel_5130/SF_IB
+ pixel_5130/PIX_OUT pixel_5130/CSA_VREF pixel
Xpixel_5141 pixel_5141/gring pixel_5141/VDD pixel_5141/GND pixel_5141/VREF pixel_5141/ROW_SEL
+ pixel_5141/NB1 pixel_5141/VBIAS pixel_5141/NB2 pixel_5141/AMP_IN pixel_5141/SF_IB
+ pixel_5141/PIX_OUT pixel_5141/CSA_VREF pixel
Xpixel_5152 pixel_5152/gring pixel_5152/VDD pixel_5152/GND pixel_5152/VREF pixel_5152/ROW_SEL
+ pixel_5152/NB1 pixel_5152/VBIAS pixel_5152/NB2 pixel_5152/AMP_IN pixel_5152/SF_IB
+ pixel_5152/PIX_OUT pixel_5152/CSA_VREF pixel
Xpixel_5163 pixel_5163/gring pixel_5163/VDD pixel_5163/GND pixel_5163/VREF pixel_5163/ROW_SEL
+ pixel_5163/NB1 pixel_5163/VBIAS pixel_5163/NB2 pixel_5163/AMP_IN pixel_5163/SF_IB
+ pixel_5163/PIX_OUT pixel_5163/CSA_VREF pixel
Xpixel_5174 pixel_5174/gring pixel_5174/VDD pixel_5174/GND pixel_5174/VREF pixel_5174/ROW_SEL
+ pixel_5174/NB1 pixel_5174/VBIAS pixel_5174/NB2 pixel_5174/AMP_IN pixel_5174/SF_IB
+ pixel_5174/PIX_OUT pixel_5174/CSA_VREF pixel
Xpixel_5185 pixel_5185/gring pixel_5185/VDD pixel_5185/GND pixel_5185/VREF pixel_5185/ROW_SEL
+ pixel_5185/NB1 pixel_5185/VBIAS pixel_5185/NB2 pixel_5185/AMP_IN pixel_5185/SF_IB
+ pixel_5185/PIX_OUT pixel_5185/CSA_VREF pixel
Xpixel_5196 pixel_5196/gring pixel_5196/VDD pixel_5196/GND pixel_5196/VREF pixel_5196/ROW_SEL
+ pixel_5196/NB1 pixel_5196/VBIAS pixel_5196/NB2 pixel_5196/AMP_IN pixel_5196/SF_IB
+ pixel_5196/PIX_OUT pixel_5196/CSA_VREF pixel
Xpixel_4440 pixel_4440/gring pixel_4440/VDD pixel_4440/GND pixel_4440/VREF pixel_4440/ROW_SEL
+ pixel_4440/NB1 pixel_4440/VBIAS pixel_4440/NB2 pixel_4440/AMP_IN pixel_4440/SF_IB
+ pixel_4440/PIX_OUT pixel_4440/CSA_VREF pixel
Xpixel_4451 pixel_4451/gring pixel_4451/VDD pixel_4451/GND pixel_4451/VREF pixel_4451/ROW_SEL
+ pixel_4451/NB1 pixel_4451/VBIAS pixel_4451/NB2 pixel_4451/AMP_IN pixel_4451/SF_IB
+ pixel_4451/PIX_OUT pixel_4451/CSA_VREF pixel
Xpixel_4462 pixel_4462/gring pixel_4462/VDD pixel_4462/GND pixel_4462/VREF pixel_4462/ROW_SEL
+ pixel_4462/NB1 pixel_4462/VBIAS pixel_4462/NB2 pixel_4462/AMP_IN pixel_4462/SF_IB
+ pixel_4462/PIX_OUT pixel_4462/CSA_VREF pixel
Xpixel_490 pixel_490/gring pixel_490/VDD pixel_490/GND pixel_490/VREF pixel_490/ROW_SEL
+ pixel_490/NB1 pixel_490/VBIAS pixel_490/NB2 pixel_490/AMP_IN pixel_490/SF_IB pixel_490/PIX_OUT
+ pixel_490/CSA_VREF pixel
Xpixel_3761 pixel_3761/gring pixel_3761/VDD pixel_3761/GND pixel_3761/VREF pixel_3761/ROW_SEL
+ pixel_3761/NB1 pixel_3761/VBIAS pixel_3761/NB2 pixel_3761/AMP_IN pixel_3761/SF_IB
+ pixel_3761/PIX_OUT pixel_3761/CSA_VREF pixel
Xpixel_3750 pixel_3750/gring pixel_3750/VDD pixel_3750/GND pixel_3750/VREF pixel_3750/ROW_SEL
+ pixel_3750/NB1 pixel_3750/VBIAS pixel_3750/NB2 pixel_3750/AMP_IN pixel_3750/SF_IB
+ pixel_3750/PIX_OUT pixel_3750/CSA_VREF pixel
Xpixel_4473 pixel_4473/gring pixel_4473/VDD pixel_4473/GND pixel_4473/VREF pixel_4473/ROW_SEL
+ pixel_4473/NB1 pixel_4473/VBIAS pixel_4473/NB2 pixel_4473/AMP_IN pixel_4473/SF_IB
+ pixel_4473/PIX_OUT pixel_4473/CSA_VREF pixel
Xpixel_4484 pixel_4484/gring pixel_4484/VDD pixel_4484/GND pixel_4484/VREF pixel_4484/ROW_SEL
+ pixel_4484/NB1 pixel_4484/VBIAS pixel_4484/NB2 pixel_4484/AMP_IN pixel_4484/SF_IB
+ pixel_4484/PIX_OUT pixel_4484/CSA_VREF pixel
Xpixel_4495 pixel_4495/gring pixel_4495/VDD pixel_4495/GND pixel_4495/VREF pixel_4495/ROW_SEL
+ pixel_4495/NB1 pixel_4495/VBIAS pixel_4495/NB2 pixel_4495/AMP_IN pixel_4495/SF_IB
+ pixel_4495/PIX_OUT pixel_4495/CSA_VREF pixel
Xpixel_3794 pixel_3794/gring pixel_3794/VDD pixel_3794/GND pixel_3794/VREF pixel_3794/ROW_SEL
+ pixel_3794/NB1 pixel_3794/VBIAS pixel_3794/NB2 pixel_3794/AMP_IN pixel_3794/SF_IB
+ pixel_3794/PIX_OUT pixel_3794/CSA_VREF pixel
Xpixel_3783 pixel_3783/gring pixel_3783/VDD pixel_3783/GND pixel_3783/VREF pixel_3783/ROW_SEL
+ pixel_3783/NB1 pixel_3783/VBIAS pixel_3783/NB2 pixel_3783/AMP_IN pixel_3783/SF_IB
+ pixel_3783/PIX_OUT pixel_3783/CSA_VREF pixel
Xpixel_3772 pixel_3772/gring pixel_3772/VDD pixel_3772/GND pixel_3772/VREF pixel_3772/ROW_SEL
+ pixel_3772/NB1 pixel_3772/VBIAS pixel_3772/NB2 pixel_3772/AMP_IN pixel_3772/SF_IB
+ pixel_3772/PIX_OUT pixel_3772/CSA_VREF pixel
Xpixel_9429 pixel_9429/gring pixel_9429/VDD pixel_9429/GND pixel_9429/VREF pixel_9429/ROW_SEL
+ pixel_9429/NB1 pixel_9429/VBIAS pixel_9429/NB2 pixel_9429/AMP_IN pixel_9429/SF_IB
+ pixel_9429/PIX_OUT pixel_9429/CSA_VREF pixel
Xpixel_9418 pixel_9418/gring pixel_9418/VDD pixel_9418/GND pixel_9418/VREF pixel_9418/ROW_SEL
+ pixel_9418/NB1 pixel_9418/VBIAS pixel_9418/NB2 pixel_9418/AMP_IN pixel_9418/SF_IB
+ pixel_9418/PIX_OUT pixel_9418/CSA_VREF pixel
Xpixel_9407 pixel_9407/gring pixel_9407/VDD pixel_9407/GND pixel_9407/VREF pixel_9407/ROW_SEL
+ pixel_9407/NB1 pixel_9407/VBIAS pixel_9407/NB2 pixel_9407/AMP_IN pixel_9407/SF_IB
+ pixel_9407/PIX_OUT pixel_9407/CSA_VREF pixel
Xpixel_8717 pixel_8717/gring pixel_8717/VDD pixel_8717/GND pixel_8717/VREF pixel_8717/ROW_SEL
+ pixel_8717/NB1 pixel_8717/VBIAS pixel_8717/NB2 pixel_8717/AMP_IN pixel_8717/SF_IB
+ pixel_8717/PIX_OUT pixel_8717/CSA_VREF pixel
Xpixel_8706 pixel_8706/gring pixel_8706/VDD pixel_8706/GND pixel_8706/VREF pixel_8706/ROW_SEL
+ pixel_8706/NB1 pixel_8706/VBIAS pixel_8706/NB2 pixel_8706/AMP_IN pixel_8706/SF_IB
+ pixel_8706/PIX_OUT pixel_8706/CSA_VREF pixel
Xpixel_8739 pixel_8739/gring pixel_8739/VDD pixel_8739/GND pixel_8739/VREF pixel_8739/ROW_SEL
+ pixel_8739/NB1 pixel_8739/VBIAS pixel_8739/NB2 pixel_8739/AMP_IN pixel_8739/SF_IB
+ pixel_8739/PIX_OUT pixel_8739/CSA_VREF pixel
Xpixel_8728 pixel_8728/gring pixel_8728/VDD pixel_8728/GND pixel_8728/VREF pixel_8728/ROW_SEL
+ pixel_8728/NB1 pixel_8728/VBIAS pixel_8728/NB2 pixel_8728/AMP_IN pixel_8728/SF_IB
+ pixel_8728/PIX_OUT pixel_8728/CSA_VREF pixel
Xpixel_3013 pixel_3013/gring pixel_3013/VDD pixel_3013/GND pixel_3013/VREF pixel_3013/ROW_SEL
+ pixel_3013/NB1 pixel_3013/VBIAS pixel_3013/NB2 pixel_3013/AMP_IN pixel_3013/SF_IB
+ pixel_3013/PIX_OUT pixel_3013/CSA_VREF pixel
Xpixel_3002 pixel_3002/gring pixel_3002/VDD pixel_3002/GND pixel_3002/VREF pixel_3002/ROW_SEL
+ pixel_3002/NB1 pixel_3002/VBIAS pixel_3002/NB2 pixel_3002/AMP_IN pixel_3002/SF_IB
+ pixel_3002/PIX_OUT pixel_3002/CSA_VREF pixel
Xpixel_2312 pixel_2312/gring pixel_2312/VDD pixel_2312/GND pixel_2312/VREF pixel_2312/ROW_SEL
+ pixel_2312/NB1 pixel_2312/VBIAS pixel_2312/NB2 pixel_2312/AMP_IN pixel_2312/SF_IB
+ pixel_2312/PIX_OUT pixel_2312/CSA_VREF pixel
Xpixel_2301 pixel_2301/gring pixel_2301/VDD pixel_2301/GND pixel_2301/VREF pixel_2301/ROW_SEL
+ pixel_2301/NB1 pixel_2301/VBIAS pixel_2301/NB2 pixel_2301/AMP_IN pixel_2301/SF_IB
+ pixel_2301/PIX_OUT pixel_2301/CSA_VREF pixel
Xpixel_3057 pixel_3057/gring pixel_3057/VDD pixel_3057/GND pixel_3057/VREF pixel_3057/ROW_SEL
+ pixel_3057/NB1 pixel_3057/VBIAS pixel_3057/NB2 pixel_3057/AMP_IN pixel_3057/SF_IB
+ pixel_3057/PIX_OUT pixel_3057/CSA_VREF pixel
Xpixel_3046 pixel_3046/gring pixel_3046/VDD pixel_3046/GND pixel_3046/VREF pixel_3046/ROW_SEL
+ pixel_3046/NB1 pixel_3046/VBIAS pixel_3046/NB2 pixel_3046/AMP_IN pixel_3046/SF_IB
+ pixel_3046/PIX_OUT pixel_3046/CSA_VREF pixel
Xpixel_3035 pixel_3035/gring pixel_3035/VDD pixel_3035/GND pixel_3035/VREF pixel_3035/ROW_SEL
+ pixel_3035/NB1 pixel_3035/VBIAS pixel_3035/NB2 pixel_3035/AMP_IN pixel_3035/SF_IB
+ pixel_3035/PIX_OUT pixel_3035/CSA_VREF pixel
Xpixel_3024 pixel_3024/gring pixel_3024/VDD pixel_3024/GND pixel_3024/VREF pixel_3024/ROW_SEL
+ pixel_3024/NB1 pixel_3024/VBIAS pixel_3024/NB2 pixel_3024/AMP_IN pixel_3024/SF_IB
+ pixel_3024/PIX_OUT pixel_3024/CSA_VREF pixel
Xpixel_1600 pixel_1600/gring pixel_1600/VDD pixel_1600/GND pixel_1600/VREF pixel_1600/ROW_SEL
+ pixel_1600/NB1 pixel_1600/VBIAS pixel_1600/NB2 pixel_1600/AMP_IN pixel_1600/SF_IB
+ pixel_1600/PIX_OUT pixel_1600/CSA_VREF pixel
Xpixel_2345 pixel_2345/gring pixel_2345/VDD pixel_2345/GND pixel_2345/VREF pixel_2345/ROW_SEL
+ pixel_2345/NB1 pixel_2345/VBIAS pixel_2345/NB2 pixel_2345/AMP_IN pixel_2345/SF_IB
+ pixel_2345/PIX_OUT pixel_2345/CSA_VREF pixel
Xpixel_2334 pixel_2334/gring pixel_2334/VDD pixel_2334/GND pixel_2334/VREF pixel_2334/ROW_SEL
+ pixel_2334/NB1 pixel_2334/VBIAS pixel_2334/NB2 pixel_2334/AMP_IN pixel_2334/SF_IB
+ pixel_2334/PIX_OUT pixel_2334/CSA_VREF pixel
Xpixel_2323 pixel_2323/gring pixel_2323/VDD pixel_2323/GND pixel_2323/VREF pixel_2323/ROW_SEL
+ pixel_2323/NB1 pixel_2323/VBIAS pixel_2323/NB2 pixel_2323/AMP_IN pixel_2323/SF_IB
+ pixel_2323/PIX_OUT pixel_2323/CSA_VREF pixel
Xpixel_3079 pixel_3079/gring pixel_3079/VDD pixel_3079/GND pixel_3079/VREF pixel_3079/ROW_SEL
+ pixel_3079/NB1 pixel_3079/VBIAS pixel_3079/NB2 pixel_3079/AMP_IN pixel_3079/SF_IB
+ pixel_3079/PIX_OUT pixel_3079/CSA_VREF pixel
Xpixel_3068 pixel_3068/gring pixel_3068/VDD pixel_3068/GND pixel_3068/VREF pixel_3068/ROW_SEL
+ pixel_3068/NB1 pixel_3068/VBIAS pixel_3068/NB2 pixel_3068/AMP_IN pixel_3068/SF_IB
+ pixel_3068/PIX_OUT pixel_3068/CSA_VREF pixel
Xpixel_1633 pixel_1633/gring pixel_1633/VDD pixel_1633/GND pixel_1633/VREF pixel_1633/ROW_SEL
+ pixel_1633/NB1 pixel_1633/VBIAS pixel_1633/NB2 pixel_1633/AMP_IN pixel_1633/SF_IB
+ pixel_1633/PIX_OUT pixel_1633/CSA_VREF pixel
Xpixel_1622 pixel_1622/gring pixel_1622/VDD pixel_1622/GND pixel_1622/VREF pixel_1622/ROW_SEL
+ pixel_1622/NB1 pixel_1622/VBIAS pixel_1622/NB2 pixel_1622/AMP_IN pixel_1622/SF_IB
+ pixel_1622/PIX_OUT pixel_1622/CSA_VREF pixel
Xpixel_1611 pixel_1611/gring pixel_1611/VDD pixel_1611/GND pixel_1611/VREF pixel_1611/ROW_SEL
+ pixel_1611/NB1 pixel_1611/VBIAS pixel_1611/NB2 pixel_1611/AMP_IN pixel_1611/SF_IB
+ pixel_1611/PIX_OUT pixel_1611/CSA_VREF pixel
Xpixel_2378 pixel_2378/gring pixel_2378/VDD pixel_2378/GND pixel_2378/VREF pixel_2378/ROW_SEL
+ pixel_2378/NB1 pixel_2378/VBIAS pixel_2378/NB2 pixel_2378/AMP_IN pixel_2378/SF_IB
+ pixel_2378/PIX_OUT pixel_2378/CSA_VREF pixel
Xpixel_2367 pixel_2367/gring pixel_2367/VDD pixel_2367/GND pixel_2367/VREF pixel_2367/ROW_SEL
+ pixel_2367/NB1 pixel_2367/VBIAS pixel_2367/NB2 pixel_2367/AMP_IN pixel_2367/SF_IB
+ pixel_2367/PIX_OUT pixel_2367/CSA_VREF pixel
Xpixel_2356 pixel_2356/gring pixel_2356/VDD pixel_2356/GND pixel_2356/VREF pixel_2356/ROW_SEL
+ pixel_2356/NB1 pixel_2356/VBIAS pixel_2356/NB2 pixel_2356/AMP_IN pixel_2356/SF_IB
+ pixel_2356/PIX_OUT pixel_2356/CSA_VREF pixel
Xpixel_1677 pixel_1677/gring pixel_1677/VDD pixel_1677/GND pixel_1677/VREF pixel_1677/ROW_SEL
+ pixel_1677/NB1 pixel_1677/VBIAS pixel_1677/NB2 pixel_1677/AMP_IN pixel_1677/SF_IB
+ pixel_1677/PIX_OUT pixel_1677/CSA_VREF pixel
Xpixel_1666 pixel_1666/gring pixel_1666/VDD pixel_1666/GND pixel_1666/VREF pixel_1666/ROW_SEL
+ pixel_1666/NB1 pixel_1666/VBIAS pixel_1666/NB2 pixel_1666/AMP_IN pixel_1666/SF_IB
+ pixel_1666/PIX_OUT pixel_1666/CSA_VREF pixel
Xpixel_1655 pixel_1655/gring pixel_1655/VDD pixel_1655/GND pixel_1655/VREF pixel_1655/ROW_SEL
+ pixel_1655/NB1 pixel_1655/VBIAS pixel_1655/NB2 pixel_1655/AMP_IN pixel_1655/SF_IB
+ pixel_1655/PIX_OUT pixel_1655/CSA_VREF pixel
Xpixel_1644 pixel_1644/gring pixel_1644/VDD pixel_1644/GND pixel_1644/VREF pixel_1644/ROW_SEL
+ pixel_1644/NB1 pixel_1644/VBIAS pixel_1644/NB2 pixel_1644/AMP_IN pixel_1644/SF_IB
+ pixel_1644/PIX_OUT pixel_1644/CSA_VREF pixel
Xpixel_2389 pixel_2389/gring pixel_2389/VDD pixel_2389/GND pixel_2389/VREF pixel_2389/ROW_SEL
+ pixel_2389/NB1 pixel_2389/VBIAS pixel_2389/NB2 pixel_2389/AMP_IN pixel_2389/SF_IB
+ pixel_2389/PIX_OUT pixel_2389/CSA_VREF pixel
Xpixel_1699 pixel_1699/gring pixel_1699/VDD pixel_1699/GND pixel_1699/VREF pixel_1699/ROW_SEL
+ pixel_1699/NB1 pixel_1699/VBIAS pixel_1699/NB2 pixel_1699/AMP_IN pixel_1699/SF_IB
+ pixel_1699/PIX_OUT pixel_1699/CSA_VREF pixel
Xpixel_1688 pixel_1688/gring pixel_1688/VDD pixel_1688/GND pixel_1688/VREF pixel_1688/ROW_SEL
+ pixel_1688/NB1 pixel_1688/VBIAS pixel_1688/NB2 pixel_1688/AMP_IN pixel_1688/SF_IB
+ pixel_1688/PIX_OUT pixel_1688/CSA_VREF pixel
Xpixel_9941 pixel_9941/gring pixel_9941/VDD pixel_9941/GND pixel_9941/VREF pixel_9941/ROW_SEL
+ pixel_9941/NB1 pixel_9941/VBIAS pixel_9941/NB2 pixel_9941/AMP_IN pixel_9941/SF_IB
+ pixel_9941/PIX_OUT pixel_9941/CSA_VREF pixel
Xpixel_9930 pixel_9930/gring pixel_9930/VDD pixel_9930/GND pixel_9930/VREF pixel_9930/ROW_SEL
+ pixel_9930/NB1 pixel_9930/VBIAS pixel_9930/NB2 pixel_9930/AMP_IN pixel_9930/SF_IB
+ pixel_9930/PIX_OUT pixel_9930/CSA_VREF pixel
Xpixel_9952 pixel_9952/gring pixel_9952/VDD pixel_9952/GND pixel_9952/VREF pixel_9952/ROW_SEL
+ pixel_9952/NB1 pixel_9952/VBIAS pixel_9952/NB2 pixel_9952/AMP_IN pixel_9952/SF_IB
+ pixel_9952/PIX_OUT pixel_9952/CSA_VREF pixel
Xpixel_9963 pixel_9963/gring pixel_9963/VDD pixel_9963/GND pixel_9963/VREF pixel_9963/ROW_SEL
+ pixel_9963/NB1 pixel_9963/VBIAS pixel_9963/NB2 pixel_9963/AMP_IN pixel_9963/SF_IB
+ pixel_9963/PIX_OUT pixel_9963/CSA_VREF pixel
Xpixel_9974 pixel_9974/gring pixel_9974/VDD pixel_9974/GND pixel_9974/VREF pixel_9974/ROW_SEL
+ pixel_9974/NB1 pixel_9974/VBIAS pixel_9974/NB2 pixel_9974/AMP_IN pixel_9974/SF_IB
+ pixel_9974/PIX_OUT pixel_9974/CSA_VREF pixel
Xpixel_9985 pixel_9985/gring pixel_9985/VDD pixel_9985/GND pixel_9985/VREF pixel_9985/ROW_SEL
+ pixel_9985/NB1 pixel_9985/VBIAS pixel_9985/NB2 pixel_9985/AMP_IN pixel_9985/SF_IB
+ pixel_9985/PIX_OUT pixel_9985/CSA_VREF pixel
Xpixel_9996 pixel_9996/gring pixel_9996/VDD pixel_9996/GND pixel_9996/VREF pixel_9996/ROW_SEL
+ pixel_9996/NB1 pixel_9996/VBIAS pixel_9996/NB2 pixel_9996/AMP_IN pixel_9996/SF_IB
+ pixel_9996/PIX_OUT pixel_9996/CSA_VREF pixel
Xpixel_4270 pixel_4270/gring pixel_4270/VDD pixel_4270/GND pixel_4270/VREF pixel_4270/ROW_SEL
+ pixel_4270/NB1 pixel_4270/VBIAS pixel_4270/NB2 pixel_4270/AMP_IN pixel_4270/SF_IB
+ pixel_4270/PIX_OUT pixel_4270/CSA_VREF pixel
Xpixel_4281 pixel_4281/gring pixel_4281/VDD pixel_4281/GND pixel_4281/VREF pixel_4281/ROW_SEL
+ pixel_4281/NB1 pixel_4281/VBIAS pixel_4281/NB2 pixel_4281/AMP_IN pixel_4281/SF_IB
+ pixel_4281/PIX_OUT pixel_4281/CSA_VREF pixel
Xpixel_4292 pixel_4292/gring pixel_4292/VDD pixel_4292/GND pixel_4292/VREF pixel_4292/ROW_SEL
+ pixel_4292/NB1 pixel_4292/VBIAS pixel_4292/NB2 pixel_4292/AMP_IN pixel_4292/SF_IB
+ pixel_4292/PIX_OUT pixel_4292/CSA_VREF pixel
Xpixel_3591 pixel_3591/gring pixel_3591/VDD pixel_3591/GND pixel_3591/VREF pixel_3591/ROW_SEL
+ pixel_3591/NB1 pixel_3591/VBIAS pixel_3591/NB2 pixel_3591/AMP_IN pixel_3591/SF_IB
+ pixel_3591/PIX_OUT pixel_3591/CSA_VREF pixel
Xpixel_3580 pixel_3580/gring pixel_3580/VDD pixel_3580/GND pixel_3580/VREF pixel_3580/ROW_SEL
+ pixel_3580/NB1 pixel_3580/VBIAS pixel_3580/NB2 pixel_3580/AMP_IN pixel_3580/SF_IB
+ pixel_3580/PIX_OUT pixel_3580/CSA_VREF pixel
Xpixel_2890 pixel_2890/gring pixel_2890/VDD pixel_2890/GND pixel_2890/VREF pixel_2890/ROW_SEL
+ pixel_2890/NB1 pixel_2890/VBIAS pixel_2890/NB2 pixel_2890/AMP_IN pixel_2890/SF_IB
+ pixel_2890/PIX_OUT pixel_2890/CSA_VREF pixel
Xpixel_9204 pixel_9204/gring pixel_9204/VDD pixel_9204/GND pixel_9204/VREF pixel_9204/ROW_SEL
+ pixel_9204/NB1 pixel_9204/VBIAS pixel_9204/NB2 pixel_9204/AMP_IN pixel_9204/SF_IB
+ pixel_9204/PIX_OUT pixel_9204/CSA_VREF pixel
Xpixel_9237 pixel_9237/gring pixel_9237/VDD pixel_9237/GND pixel_9237/VREF pixel_9237/ROW_SEL
+ pixel_9237/NB1 pixel_9237/VBIAS pixel_9237/NB2 pixel_9237/AMP_IN pixel_9237/SF_IB
+ pixel_9237/PIX_OUT pixel_9237/CSA_VREF pixel
Xpixel_9226 pixel_9226/gring pixel_9226/VDD pixel_9226/GND pixel_9226/VREF pixel_9226/ROW_SEL
+ pixel_9226/NB1 pixel_9226/VBIAS pixel_9226/NB2 pixel_9226/AMP_IN pixel_9226/SF_IB
+ pixel_9226/PIX_OUT pixel_9226/CSA_VREF pixel
Xpixel_9215 pixel_9215/gring pixel_9215/VDD pixel_9215/GND pixel_9215/VREF pixel_9215/ROW_SEL
+ pixel_9215/NB1 pixel_9215/VBIAS pixel_9215/NB2 pixel_9215/AMP_IN pixel_9215/SF_IB
+ pixel_9215/PIX_OUT pixel_9215/CSA_VREF pixel
Xpixel_8536 pixel_8536/gring pixel_8536/VDD pixel_8536/GND pixel_8536/VREF pixel_8536/ROW_SEL
+ pixel_8536/NB1 pixel_8536/VBIAS pixel_8536/NB2 pixel_8536/AMP_IN pixel_8536/SF_IB
+ pixel_8536/PIX_OUT pixel_8536/CSA_VREF pixel
Xpixel_8525 pixel_8525/gring pixel_8525/VDD pixel_8525/GND pixel_8525/VREF pixel_8525/ROW_SEL
+ pixel_8525/NB1 pixel_8525/VBIAS pixel_8525/NB2 pixel_8525/AMP_IN pixel_8525/SF_IB
+ pixel_8525/PIX_OUT pixel_8525/CSA_VREF pixel
Xpixel_8514 pixel_8514/gring pixel_8514/VDD pixel_8514/GND pixel_8514/VREF pixel_8514/ROW_SEL
+ pixel_8514/NB1 pixel_8514/VBIAS pixel_8514/NB2 pixel_8514/AMP_IN pixel_8514/SF_IB
+ pixel_8514/PIX_OUT pixel_8514/CSA_VREF pixel
Xpixel_8503 pixel_8503/gring pixel_8503/VDD pixel_8503/GND pixel_8503/VREF pixel_8503/ROW_SEL
+ pixel_8503/NB1 pixel_8503/VBIAS pixel_8503/NB2 pixel_8503/AMP_IN pixel_8503/SF_IB
+ pixel_8503/PIX_OUT pixel_8503/CSA_VREF pixel
Xpixel_9259 pixel_9259/gring pixel_9259/VDD pixel_9259/GND pixel_9259/VREF pixel_9259/ROW_SEL
+ pixel_9259/NB1 pixel_9259/VBIAS pixel_9259/NB2 pixel_9259/AMP_IN pixel_9259/SF_IB
+ pixel_9259/PIX_OUT pixel_9259/CSA_VREF pixel
Xpixel_9248 pixel_9248/gring pixel_9248/VDD pixel_9248/GND pixel_9248/VREF pixel_9248/ROW_SEL
+ pixel_9248/NB1 pixel_9248/VBIAS pixel_9248/NB2 pixel_9248/AMP_IN pixel_9248/SF_IB
+ pixel_9248/PIX_OUT pixel_9248/CSA_VREF pixel
Xpixel_8569 pixel_8569/gring pixel_8569/VDD pixel_8569/GND pixel_8569/VREF pixel_8569/ROW_SEL
+ pixel_8569/NB1 pixel_8569/VBIAS pixel_8569/NB2 pixel_8569/AMP_IN pixel_8569/SF_IB
+ pixel_8569/PIX_OUT pixel_8569/CSA_VREF pixel
Xpixel_8558 pixel_8558/gring pixel_8558/VDD pixel_8558/GND pixel_8558/VREF pixel_8558/ROW_SEL
+ pixel_8558/NB1 pixel_8558/VBIAS pixel_8558/NB2 pixel_8558/AMP_IN pixel_8558/SF_IB
+ pixel_8558/PIX_OUT pixel_8558/CSA_VREF pixel
Xpixel_8547 pixel_8547/gring pixel_8547/VDD pixel_8547/GND pixel_8547/VREF pixel_8547/ROW_SEL
+ pixel_8547/NB1 pixel_8547/VBIAS pixel_8547/NB2 pixel_8547/AMP_IN pixel_8547/SF_IB
+ pixel_8547/PIX_OUT pixel_8547/CSA_VREF pixel
Xpixel_7802 pixel_7802/gring pixel_7802/VDD pixel_7802/GND pixel_7802/VREF pixel_7802/ROW_SEL
+ pixel_7802/NB1 pixel_7802/VBIAS pixel_7802/NB2 pixel_7802/AMP_IN pixel_7802/SF_IB
+ pixel_7802/PIX_OUT pixel_7802/CSA_VREF pixel
Xpixel_7813 pixel_7813/gring pixel_7813/VDD pixel_7813/GND pixel_7813/VREF pixel_7813/ROW_SEL
+ pixel_7813/NB1 pixel_7813/VBIAS pixel_7813/NB2 pixel_7813/AMP_IN pixel_7813/SF_IB
+ pixel_7813/PIX_OUT pixel_7813/CSA_VREF pixel
Xpixel_7824 pixel_7824/gring pixel_7824/VDD pixel_7824/GND pixel_7824/VREF pixel_7824/ROW_SEL
+ pixel_7824/NB1 pixel_7824/VBIAS pixel_7824/NB2 pixel_7824/AMP_IN pixel_7824/SF_IB
+ pixel_7824/PIX_OUT pixel_7824/CSA_VREF pixel
Xpixel_7835 pixel_7835/gring pixel_7835/VDD pixel_7835/GND pixel_7835/VREF pixel_7835/ROW_SEL
+ pixel_7835/NB1 pixel_7835/VBIAS pixel_7835/NB2 pixel_7835/AMP_IN pixel_7835/SF_IB
+ pixel_7835/PIX_OUT pixel_7835/CSA_VREF pixel
Xpixel_7846 pixel_7846/gring pixel_7846/VDD pixel_7846/GND pixel_7846/VREF pixel_7846/ROW_SEL
+ pixel_7846/NB1 pixel_7846/VBIAS pixel_7846/NB2 pixel_7846/AMP_IN pixel_7846/SF_IB
+ pixel_7846/PIX_OUT pixel_7846/CSA_VREF pixel
Xpixel_7857 pixel_7857/gring pixel_7857/VDD pixel_7857/GND pixel_7857/VREF pixel_7857/ROW_SEL
+ pixel_7857/NB1 pixel_7857/VBIAS pixel_7857/NB2 pixel_7857/AMP_IN pixel_7857/SF_IB
+ pixel_7857/PIX_OUT pixel_7857/CSA_VREF pixel
Xpixel_7868 pixel_7868/gring pixel_7868/VDD pixel_7868/GND pixel_7868/VREF pixel_7868/ROW_SEL
+ pixel_7868/NB1 pixel_7868/VBIAS pixel_7868/NB2 pixel_7868/AMP_IN pixel_7868/SF_IB
+ pixel_7868/PIX_OUT pixel_7868/CSA_VREF pixel
Xpixel_7879 pixel_7879/gring pixel_7879/VDD pixel_7879/GND pixel_7879/VREF pixel_7879/ROW_SEL
+ pixel_7879/NB1 pixel_7879/VBIAS pixel_7879/NB2 pixel_7879/AMP_IN pixel_7879/SF_IB
+ pixel_7879/PIX_OUT pixel_7879/CSA_VREF pixel
Xpixel_2120 pixel_2120/gring pixel_2120/VDD pixel_2120/GND pixel_2120/VREF pixel_2120/ROW_SEL
+ pixel_2120/NB1 pixel_2120/VBIAS pixel_2120/NB2 pixel_2120/AMP_IN pixel_2120/SF_IB
+ pixel_2120/PIX_OUT pixel_2120/CSA_VREF pixel
Xpixel_2153 pixel_2153/gring pixel_2153/VDD pixel_2153/GND pixel_2153/VREF pixel_2153/ROW_SEL
+ pixel_2153/NB1 pixel_2153/VBIAS pixel_2153/NB2 pixel_2153/AMP_IN pixel_2153/SF_IB
+ pixel_2153/PIX_OUT pixel_2153/CSA_VREF pixel
Xpixel_2142 pixel_2142/gring pixel_2142/VDD pixel_2142/GND pixel_2142/VREF pixel_2142/ROW_SEL
+ pixel_2142/NB1 pixel_2142/VBIAS pixel_2142/NB2 pixel_2142/AMP_IN pixel_2142/SF_IB
+ pixel_2142/PIX_OUT pixel_2142/CSA_VREF pixel
Xpixel_2131 pixel_2131/gring pixel_2131/VDD pixel_2131/GND pixel_2131/VREF pixel_2131/ROW_SEL
+ pixel_2131/NB1 pixel_2131/VBIAS pixel_2131/NB2 pixel_2131/AMP_IN pixel_2131/SF_IB
+ pixel_2131/PIX_OUT pixel_2131/CSA_VREF pixel
Xpixel_1452 pixel_1452/gring pixel_1452/VDD pixel_1452/GND pixel_1452/VREF pixel_1452/ROW_SEL
+ pixel_1452/NB1 pixel_1452/VBIAS pixel_1452/NB2 pixel_1452/AMP_IN pixel_1452/SF_IB
+ pixel_1452/PIX_OUT pixel_1452/CSA_VREF pixel
Xpixel_1441 pixel_1441/gring pixel_1441/VDD pixel_1441/GND pixel_1441/VREF pixel_1441/ROW_SEL
+ pixel_1441/NB1 pixel_1441/VBIAS pixel_1441/NB2 pixel_1441/AMP_IN pixel_1441/SF_IB
+ pixel_1441/PIX_OUT pixel_1441/CSA_VREF pixel
Xpixel_1430 pixel_1430/gring pixel_1430/VDD pixel_1430/GND pixel_1430/VREF pixel_1430/ROW_SEL
+ pixel_1430/NB1 pixel_1430/VBIAS pixel_1430/NB2 pixel_1430/AMP_IN pixel_1430/SF_IB
+ pixel_1430/PIX_OUT pixel_1430/CSA_VREF pixel
Xpixel_2197 pixel_2197/gring pixel_2197/VDD pixel_2197/GND pixel_2197/VREF pixel_2197/ROW_SEL
+ pixel_2197/NB1 pixel_2197/VBIAS pixel_2197/NB2 pixel_2197/AMP_IN pixel_2197/SF_IB
+ pixel_2197/PIX_OUT pixel_2197/CSA_VREF pixel
Xpixel_2186 pixel_2186/gring pixel_2186/VDD pixel_2186/GND pixel_2186/VREF pixel_2186/ROW_SEL
+ pixel_2186/NB1 pixel_2186/VBIAS pixel_2186/NB2 pixel_2186/AMP_IN pixel_2186/SF_IB
+ pixel_2186/PIX_OUT pixel_2186/CSA_VREF pixel
Xpixel_2175 pixel_2175/gring pixel_2175/VDD pixel_2175/GND pixel_2175/VREF pixel_2175/ROW_SEL
+ pixel_2175/NB1 pixel_2175/VBIAS pixel_2175/NB2 pixel_2175/AMP_IN pixel_2175/SF_IB
+ pixel_2175/PIX_OUT pixel_2175/CSA_VREF pixel
Xpixel_2164 pixel_2164/gring pixel_2164/VDD pixel_2164/GND pixel_2164/VREF pixel_2164/ROW_SEL
+ pixel_2164/NB1 pixel_2164/VBIAS pixel_2164/NB2 pixel_2164/AMP_IN pixel_2164/SF_IB
+ pixel_2164/PIX_OUT pixel_2164/CSA_VREF pixel
Xpixel_1485 pixel_1485/gring pixel_1485/VDD pixel_1485/GND pixel_1485/VREF pixel_1485/ROW_SEL
+ pixel_1485/NB1 pixel_1485/VBIAS pixel_1485/NB2 pixel_1485/AMP_IN pixel_1485/SF_IB
+ pixel_1485/PIX_OUT pixel_1485/CSA_VREF pixel
Xpixel_1474 pixel_1474/gring pixel_1474/VDD pixel_1474/GND pixel_1474/VREF pixel_1474/ROW_SEL
+ pixel_1474/NB1 pixel_1474/VBIAS pixel_1474/NB2 pixel_1474/AMP_IN pixel_1474/SF_IB
+ pixel_1474/PIX_OUT pixel_1474/CSA_VREF pixel
Xpixel_1463 pixel_1463/gring pixel_1463/VDD pixel_1463/GND pixel_1463/VREF pixel_1463/ROW_SEL
+ pixel_1463/NB1 pixel_1463/VBIAS pixel_1463/NB2 pixel_1463/AMP_IN pixel_1463/SF_IB
+ pixel_1463/PIX_OUT pixel_1463/CSA_VREF pixel
Xpixel_1496 pixel_1496/gring pixel_1496/VDD pixel_1496/GND pixel_1496/VREF pixel_1496/ROW_SEL
+ pixel_1496/NB1 pixel_1496/VBIAS pixel_1496/NB2 pixel_1496/AMP_IN pixel_1496/SF_IB
+ pixel_1496/PIX_OUT pixel_1496/CSA_VREF pixel
Xpixel_9760 pixel_9760/gring pixel_9760/VDD pixel_9760/GND pixel_9760/VREF pixel_9760/ROW_SEL
+ pixel_9760/NB1 pixel_9760/VBIAS pixel_9760/NB2 pixel_9760/AMP_IN pixel_9760/SF_IB
+ pixel_9760/PIX_OUT pixel_9760/CSA_VREF pixel
Xpixel_9771 pixel_9771/gring pixel_9771/VDD pixel_9771/GND pixel_9771/VREF pixel_9771/ROW_SEL
+ pixel_9771/NB1 pixel_9771/VBIAS pixel_9771/NB2 pixel_9771/AMP_IN pixel_9771/SF_IB
+ pixel_9771/PIX_OUT pixel_9771/CSA_VREF pixel
Xpixel_9782 pixel_9782/gring pixel_9782/VDD pixel_9782/GND pixel_9782/VREF pixel_9782/ROW_SEL
+ pixel_9782/NB1 pixel_9782/VBIAS pixel_9782/NB2 pixel_9782/AMP_IN pixel_9782/SF_IB
+ pixel_9782/PIX_OUT pixel_9782/CSA_VREF pixel
Xpixel_9793 pixel_9793/gring pixel_9793/VDD pixel_9793/GND pixel_9793/VREF pixel_9793/ROW_SEL
+ pixel_9793/NB1 pixel_9793/VBIAS pixel_9793/NB2 pixel_9793/AMP_IN pixel_9793/SF_IB
+ pixel_9793/PIX_OUT pixel_9793/CSA_VREF pixel
Xpixel_7109 pixel_7109/gring pixel_7109/VDD pixel_7109/GND pixel_7109/VREF pixel_7109/ROW_SEL
+ pixel_7109/NB1 pixel_7109/VBIAS pixel_7109/NB2 pixel_7109/AMP_IN pixel_7109/SF_IB
+ pixel_7109/PIX_OUT pixel_7109/CSA_VREF pixel
Xpixel_6408 pixel_6408/gring pixel_6408/VDD pixel_6408/GND pixel_6408/VREF pixel_6408/ROW_SEL
+ pixel_6408/NB1 pixel_6408/VBIAS pixel_6408/NB2 pixel_6408/AMP_IN pixel_6408/SF_IB
+ pixel_6408/PIX_OUT pixel_6408/CSA_VREF pixel
Xpixel_6419 pixel_6419/gring pixel_6419/VDD pixel_6419/GND pixel_6419/VREF pixel_6419/ROW_SEL
+ pixel_6419/NB1 pixel_6419/VBIAS pixel_6419/NB2 pixel_6419/AMP_IN pixel_6419/SF_IB
+ pixel_6419/PIX_OUT pixel_6419/CSA_VREF pixel
Xpixel_5707 pixel_5707/gring pixel_5707/VDD pixel_5707/GND pixel_5707/VREF pixel_5707/ROW_SEL
+ pixel_5707/NB1 pixel_5707/VBIAS pixel_5707/NB2 pixel_5707/AMP_IN pixel_5707/SF_IB
+ pixel_5707/PIX_OUT pixel_5707/CSA_VREF pixel
Xpixel_5718 pixel_5718/gring pixel_5718/VDD pixel_5718/GND pixel_5718/VREF pixel_5718/ROW_SEL
+ pixel_5718/NB1 pixel_5718/VBIAS pixel_5718/NB2 pixel_5718/AMP_IN pixel_5718/SF_IB
+ pixel_5718/PIX_OUT pixel_5718/CSA_VREF pixel
Xpixel_5729 pixel_5729/gring pixel_5729/VDD pixel_5729/GND pixel_5729/VREF pixel_5729/ROW_SEL
+ pixel_5729/NB1 pixel_5729/VBIAS pixel_5729/NB2 pixel_5729/AMP_IN pixel_5729/SF_IB
+ pixel_5729/PIX_OUT pixel_5729/CSA_VREF pixel
Xpixel_9012 pixel_9012/gring pixel_9012/VDD pixel_9012/GND pixel_9012/VREF pixel_9012/ROW_SEL
+ pixel_9012/NB1 pixel_9012/VBIAS pixel_9012/NB2 pixel_9012/AMP_IN pixel_9012/SF_IB
+ pixel_9012/PIX_OUT pixel_9012/CSA_VREF pixel
Xpixel_9001 pixel_9001/gring pixel_9001/VDD pixel_9001/GND pixel_9001/VREF pixel_9001/ROW_SEL
+ pixel_9001/NB1 pixel_9001/VBIAS pixel_9001/NB2 pixel_9001/AMP_IN pixel_9001/SF_IB
+ pixel_9001/PIX_OUT pixel_9001/CSA_VREF pixel
Xpixel_9045 pixel_9045/gring pixel_9045/VDD pixel_9045/GND pixel_9045/VREF pixel_9045/ROW_SEL
+ pixel_9045/NB1 pixel_9045/VBIAS pixel_9045/NB2 pixel_9045/AMP_IN pixel_9045/SF_IB
+ pixel_9045/PIX_OUT pixel_9045/CSA_VREF pixel
Xpixel_9034 pixel_9034/gring pixel_9034/VDD pixel_9034/GND pixel_9034/VREF pixel_9034/ROW_SEL
+ pixel_9034/NB1 pixel_9034/VBIAS pixel_9034/NB2 pixel_9034/AMP_IN pixel_9034/SF_IB
+ pixel_9034/PIX_OUT pixel_9034/CSA_VREF pixel
Xpixel_9023 pixel_9023/gring pixel_9023/VDD pixel_9023/GND pixel_9023/VREF pixel_9023/ROW_SEL
+ pixel_9023/NB1 pixel_9023/VBIAS pixel_9023/NB2 pixel_9023/AMP_IN pixel_9023/SF_IB
+ pixel_9023/PIX_OUT pixel_9023/CSA_VREF pixel
Xpixel_8300 pixel_8300/gring pixel_8300/VDD pixel_8300/GND pixel_8300/VREF pixel_8300/ROW_SEL
+ pixel_8300/NB1 pixel_8300/VBIAS pixel_8300/NB2 pixel_8300/AMP_IN pixel_8300/SF_IB
+ pixel_8300/PIX_OUT pixel_8300/CSA_VREF pixel
Xpixel_9089 pixel_9089/gring pixel_9089/VDD pixel_9089/GND pixel_9089/VREF pixel_9089/ROW_SEL
+ pixel_9089/NB1 pixel_9089/VBIAS pixel_9089/NB2 pixel_9089/AMP_IN pixel_9089/SF_IB
+ pixel_9089/PIX_OUT pixel_9089/CSA_VREF pixel
Xpixel_9078 pixel_9078/gring pixel_9078/VDD pixel_9078/GND pixel_9078/VREF pixel_9078/ROW_SEL
+ pixel_9078/NB1 pixel_9078/VBIAS pixel_9078/NB2 pixel_9078/AMP_IN pixel_9078/SF_IB
+ pixel_9078/PIX_OUT pixel_9078/CSA_VREF pixel
Xpixel_9067 pixel_9067/gring pixel_9067/VDD pixel_9067/GND pixel_9067/VREF pixel_9067/ROW_SEL
+ pixel_9067/NB1 pixel_9067/VBIAS pixel_9067/NB2 pixel_9067/AMP_IN pixel_9067/SF_IB
+ pixel_9067/PIX_OUT pixel_9067/CSA_VREF pixel
Xpixel_9056 pixel_9056/gring pixel_9056/VDD pixel_9056/GND pixel_9056/VREF pixel_9056/ROW_SEL
+ pixel_9056/NB1 pixel_9056/VBIAS pixel_9056/NB2 pixel_9056/AMP_IN pixel_9056/SF_IB
+ pixel_9056/PIX_OUT pixel_9056/CSA_VREF pixel
Xpixel_8311 pixel_8311/gring pixel_8311/VDD pixel_8311/GND pixel_8311/VREF pixel_8311/ROW_SEL
+ pixel_8311/NB1 pixel_8311/VBIAS pixel_8311/NB2 pixel_8311/AMP_IN pixel_8311/SF_IB
+ pixel_8311/PIX_OUT pixel_8311/CSA_VREF pixel
Xpixel_8322 pixel_8322/gring pixel_8322/VDD pixel_8322/GND pixel_8322/VREF pixel_8322/ROW_SEL
+ pixel_8322/NB1 pixel_8322/VBIAS pixel_8322/NB2 pixel_8322/AMP_IN pixel_8322/SF_IB
+ pixel_8322/PIX_OUT pixel_8322/CSA_VREF pixel
Xpixel_8333 pixel_8333/gring pixel_8333/VDD pixel_8333/GND pixel_8333/VREF pixel_8333/ROW_SEL
+ pixel_8333/NB1 pixel_8333/VBIAS pixel_8333/NB2 pixel_8333/AMP_IN pixel_8333/SF_IB
+ pixel_8333/PIX_OUT pixel_8333/CSA_VREF pixel
Xpixel_8344 pixel_8344/gring pixel_8344/VDD pixel_8344/GND pixel_8344/VREF pixel_8344/ROW_SEL
+ pixel_8344/NB1 pixel_8344/VBIAS pixel_8344/NB2 pixel_8344/AMP_IN pixel_8344/SF_IB
+ pixel_8344/PIX_OUT pixel_8344/CSA_VREF pixel
Xpixel_8355 pixel_8355/gring pixel_8355/VDD pixel_8355/GND pixel_8355/VREF pixel_8355/ROW_SEL
+ pixel_8355/NB1 pixel_8355/VBIAS pixel_8355/NB2 pixel_8355/AMP_IN pixel_8355/SF_IB
+ pixel_8355/PIX_OUT pixel_8355/CSA_VREF pixel
Xpixel_8366 pixel_8366/gring pixel_8366/VDD pixel_8366/GND pixel_8366/VREF pixel_8366/ROW_SEL
+ pixel_8366/NB1 pixel_8366/VBIAS pixel_8366/NB2 pixel_8366/AMP_IN pixel_8366/SF_IB
+ pixel_8366/PIX_OUT pixel_8366/CSA_VREF pixel
Xpixel_8377 pixel_8377/gring pixel_8377/VDD pixel_8377/GND pixel_8377/VREF pixel_8377/ROW_SEL
+ pixel_8377/NB1 pixel_8377/VBIAS pixel_8377/NB2 pixel_8377/AMP_IN pixel_8377/SF_IB
+ pixel_8377/PIX_OUT pixel_8377/CSA_VREF pixel
Xpixel_7610 pixel_7610/gring pixel_7610/VDD pixel_7610/GND pixel_7610/VREF pixel_7610/ROW_SEL
+ pixel_7610/NB1 pixel_7610/VBIAS pixel_7610/NB2 pixel_7610/AMP_IN pixel_7610/SF_IB
+ pixel_7610/PIX_OUT pixel_7610/CSA_VREF pixel
Xpixel_7621 pixel_7621/gring pixel_7621/VDD pixel_7621/GND pixel_7621/VREF pixel_7621/ROW_SEL
+ pixel_7621/NB1 pixel_7621/VBIAS pixel_7621/NB2 pixel_7621/AMP_IN pixel_7621/SF_IB
+ pixel_7621/PIX_OUT pixel_7621/CSA_VREF pixel
Xpixel_7632 pixel_7632/gring pixel_7632/VDD pixel_7632/GND pixel_7632/VREF pixel_7632/ROW_SEL
+ pixel_7632/NB1 pixel_7632/VBIAS pixel_7632/NB2 pixel_7632/AMP_IN pixel_7632/SF_IB
+ pixel_7632/PIX_OUT pixel_7632/CSA_VREF pixel
Xpixel_8388 pixel_8388/gring pixel_8388/VDD pixel_8388/GND pixel_8388/VREF pixel_8388/ROW_SEL
+ pixel_8388/NB1 pixel_8388/VBIAS pixel_8388/NB2 pixel_8388/AMP_IN pixel_8388/SF_IB
+ pixel_8388/PIX_OUT pixel_8388/CSA_VREF pixel
Xpixel_8399 pixel_8399/gring pixel_8399/VDD pixel_8399/GND pixel_8399/VREF pixel_8399/ROW_SEL
+ pixel_8399/NB1 pixel_8399/VBIAS pixel_8399/NB2 pixel_8399/AMP_IN pixel_8399/SF_IB
+ pixel_8399/PIX_OUT pixel_8399/CSA_VREF pixel
Xpixel_7643 pixel_7643/gring pixel_7643/VDD pixel_7643/GND pixel_7643/VREF pixel_7643/ROW_SEL
+ pixel_7643/NB1 pixel_7643/VBIAS pixel_7643/NB2 pixel_7643/AMP_IN pixel_7643/SF_IB
+ pixel_7643/PIX_OUT pixel_7643/CSA_VREF pixel
Xpixel_7654 pixel_7654/gring pixel_7654/VDD pixel_7654/GND pixel_7654/VREF pixel_7654/ROW_SEL
+ pixel_7654/NB1 pixel_7654/VBIAS pixel_7654/NB2 pixel_7654/AMP_IN pixel_7654/SF_IB
+ pixel_7654/PIX_OUT pixel_7654/CSA_VREF pixel
Xpixel_7665 pixel_7665/gring pixel_7665/VDD pixel_7665/GND pixel_7665/VREF pixel_7665/ROW_SEL
+ pixel_7665/NB1 pixel_7665/VBIAS pixel_7665/NB2 pixel_7665/AMP_IN pixel_7665/SF_IB
+ pixel_7665/PIX_OUT pixel_7665/CSA_VREF pixel
Xpixel_7676 pixel_7676/gring pixel_7676/VDD pixel_7676/GND pixel_7676/VREF pixel_7676/ROW_SEL
+ pixel_7676/NB1 pixel_7676/VBIAS pixel_7676/NB2 pixel_7676/AMP_IN pixel_7676/SF_IB
+ pixel_7676/PIX_OUT pixel_7676/CSA_VREF pixel
Xpixel_6920 pixel_6920/gring pixel_6920/VDD pixel_6920/GND pixel_6920/VREF pixel_6920/ROW_SEL
+ pixel_6920/NB1 pixel_6920/VBIAS pixel_6920/NB2 pixel_6920/AMP_IN pixel_6920/SF_IB
+ pixel_6920/PIX_OUT pixel_6920/CSA_VREF pixel
Xpixel_6931 pixel_6931/gring pixel_6931/VDD pixel_6931/GND pixel_6931/VREF pixel_6931/ROW_SEL
+ pixel_6931/NB1 pixel_6931/VBIAS pixel_6931/NB2 pixel_6931/AMP_IN pixel_6931/SF_IB
+ pixel_6931/PIX_OUT pixel_6931/CSA_VREF pixel
Xpixel_12 pixel_12/gring pixel_12/VDD pixel_12/GND pixel_12/VREF pixel_12/ROW_SEL
+ pixel_12/NB1 pixel_12/VBIAS pixel_12/NB2 pixel_12/AMP_IN pixel_12/SF_IB pixel_12/PIX_OUT
+ pixel_12/CSA_VREF pixel
Xpixel_7687 pixel_7687/gring pixel_7687/VDD pixel_7687/GND pixel_7687/VREF pixel_7687/ROW_SEL
+ pixel_7687/NB1 pixel_7687/VBIAS pixel_7687/NB2 pixel_7687/AMP_IN pixel_7687/SF_IB
+ pixel_7687/PIX_OUT pixel_7687/CSA_VREF pixel
Xpixel_7698 pixel_7698/gring pixel_7698/VDD pixel_7698/GND pixel_7698/VREF pixel_7698/ROW_SEL
+ pixel_7698/NB1 pixel_7698/VBIAS pixel_7698/NB2 pixel_7698/AMP_IN pixel_7698/SF_IB
+ pixel_7698/PIX_OUT pixel_7698/CSA_VREF pixel
Xpixel_6942 pixel_6942/gring pixel_6942/VDD pixel_6942/GND pixel_6942/VREF pixel_6942/ROW_SEL
+ pixel_6942/NB1 pixel_6942/VBIAS pixel_6942/NB2 pixel_6942/AMP_IN pixel_6942/SF_IB
+ pixel_6942/PIX_OUT pixel_6942/CSA_VREF pixel
Xpixel_6953 pixel_6953/gring pixel_6953/VDD pixel_6953/GND pixel_6953/VREF pixel_6953/ROW_SEL
+ pixel_6953/NB1 pixel_6953/VBIAS pixel_6953/NB2 pixel_6953/AMP_IN pixel_6953/SF_IB
+ pixel_6953/PIX_OUT pixel_6953/CSA_VREF pixel
Xpixel_6964 pixel_6964/gring pixel_6964/VDD pixel_6964/GND pixel_6964/VREF pixel_6964/ROW_SEL
+ pixel_6964/NB1 pixel_6964/VBIAS pixel_6964/NB2 pixel_6964/AMP_IN pixel_6964/SF_IB
+ pixel_6964/PIX_OUT pixel_6964/CSA_VREF pixel
Xpixel_45 pixel_45/gring pixel_45/VDD pixel_45/GND pixel_45/VREF pixel_45/ROW_SEL
+ pixel_45/NB1 pixel_45/VBIAS pixel_45/NB2 pixel_45/AMP_IN pixel_45/SF_IB pixel_45/PIX_OUT
+ pixel_45/CSA_VREF pixel
Xpixel_34 pixel_34/gring pixel_34/VDD pixel_34/GND pixel_34/VREF pixel_34/ROW_SEL
+ pixel_34/NB1 pixel_34/VBIAS pixel_34/NB2 pixel_34/AMP_IN pixel_34/SF_IB pixel_34/PIX_OUT
+ pixel_34/CSA_VREF pixel
Xpixel_23 pixel_23/gring pixel_23/VDD pixel_23/GND pixel_23/VREF pixel_23/ROW_SEL
+ pixel_23/NB1 pixel_23/VBIAS pixel_23/NB2 pixel_23/AMP_IN pixel_23/SF_IB pixel_23/PIX_OUT
+ pixel_23/CSA_VREF pixel
Xpixel_6975 pixel_6975/gring pixel_6975/VDD pixel_6975/GND pixel_6975/VREF pixel_6975/ROW_SEL
+ pixel_6975/NB1 pixel_6975/VBIAS pixel_6975/NB2 pixel_6975/AMP_IN pixel_6975/SF_IB
+ pixel_6975/PIX_OUT pixel_6975/CSA_VREF pixel
Xpixel_6986 pixel_6986/gring pixel_6986/VDD pixel_6986/GND pixel_6986/VREF pixel_6986/ROW_SEL
+ pixel_6986/NB1 pixel_6986/VBIAS pixel_6986/NB2 pixel_6986/AMP_IN pixel_6986/SF_IB
+ pixel_6986/PIX_OUT pixel_6986/CSA_VREF pixel
Xpixel_6997 pixel_6997/gring pixel_6997/VDD pixel_6997/GND pixel_6997/VREF pixel_6997/ROW_SEL
+ pixel_6997/NB1 pixel_6997/VBIAS pixel_6997/NB2 pixel_6997/AMP_IN pixel_6997/SF_IB
+ pixel_6997/PIX_OUT pixel_6997/CSA_VREF pixel
Xpixel_78 pixel_78/gring pixel_78/VDD pixel_78/GND pixel_78/VREF pixel_78/ROW_SEL
+ pixel_78/NB1 pixel_78/VBIAS pixel_78/NB2 pixel_78/AMP_IN pixel_78/SF_IB pixel_78/PIX_OUT
+ pixel_78/CSA_VREF pixel
Xpixel_67 pixel_67/gring pixel_67/VDD pixel_67/GND pixel_67/VREF pixel_67/ROW_SEL
+ pixel_67/NB1 pixel_67/VBIAS pixel_67/NB2 pixel_67/AMP_IN pixel_67/SF_IB pixel_67/PIX_OUT
+ pixel_67/CSA_VREF pixel
Xpixel_56 pixel_56/gring pixel_56/VDD pixel_56/GND pixel_56/VREF pixel_56/ROW_SEL
+ pixel_56/NB1 pixel_56/VBIAS pixel_56/NB2 pixel_56/AMP_IN pixel_56/SF_IB pixel_56/PIX_OUT
+ pixel_56/CSA_VREF pixel
Xpixel_89 pixel_89/gring pixel_89/VDD pixel_89/GND pixel_89/VREF pixel_89/ROW_SEL
+ pixel_89/NB1 pixel_89/VBIAS pixel_89/NB2 pixel_89/AMP_IN pixel_89/SF_IB pixel_89/PIX_OUT
+ pixel_89/CSA_VREF pixel
Xpixel_1260 pixel_1260/gring pixel_1260/VDD pixel_1260/GND pixel_1260/VREF pixel_1260/ROW_SEL
+ pixel_1260/NB1 pixel_1260/VBIAS pixel_1260/NB2 pixel_1260/AMP_IN pixel_1260/SF_IB
+ pixel_1260/PIX_OUT pixel_1260/CSA_VREF pixel
Xpixel_1293 pixel_1293/gring pixel_1293/VDD pixel_1293/GND pixel_1293/VREF pixel_1293/ROW_SEL
+ pixel_1293/NB1 pixel_1293/VBIAS pixel_1293/NB2 pixel_1293/AMP_IN pixel_1293/SF_IB
+ pixel_1293/PIX_OUT pixel_1293/CSA_VREF pixel
Xpixel_1282 pixel_1282/gring pixel_1282/VDD pixel_1282/GND pixel_1282/VREF pixel_1282/ROW_SEL
+ pixel_1282/NB1 pixel_1282/VBIAS pixel_1282/NB2 pixel_1282/AMP_IN pixel_1282/SF_IB
+ pixel_1282/PIX_OUT pixel_1282/CSA_VREF pixel
Xpixel_1271 pixel_1271/gring pixel_1271/VDD pixel_1271/GND pixel_1271/VREF pixel_1271/ROW_SEL
+ pixel_1271/NB1 pixel_1271/VBIAS pixel_1271/NB2 pixel_1271/AMP_IN pixel_1271/SF_IB
+ pixel_1271/PIX_OUT pixel_1271/CSA_VREF pixel
Xpixel_9590 pixel_9590/gring pixel_9590/VDD pixel_9590/GND pixel_9590/VREF pixel_9590/ROW_SEL
+ pixel_9590/NB1 pixel_9590/VBIAS pixel_9590/NB2 pixel_9590/AMP_IN pixel_9590/SF_IB
+ pixel_9590/PIX_OUT pixel_9590/CSA_VREF pixel
Xpixel_319 pixel_319/gring pixel_319/VDD pixel_319/GND pixel_319/VREF pixel_319/ROW_SEL
+ pixel_319/NB1 pixel_319/VBIAS pixel_319/NB2 pixel_319/AMP_IN pixel_319/SF_IB pixel_319/PIX_OUT
+ pixel_319/CSA_VREF pixel
Xpixel_308 pixel_308/gring pixel_308/VDD pixel_308/GND pixel_308/VREF pixel_308/ROW_SEL
+ pixel_308/NB1 pixel_308/VBIAS pixel_308/NB2 pixel_308/AMP_IN pixel_308/SF_IB pixel_308/PIX_OUT
+ pixel_308/CSA_VREF pixel
Xpixel_6205 pixel_6205/gring pixel_6205/VDD pixel_6205/GND pixel_6205/VREF pixel_6205/ROW_SEL
+ pixel_6205/NB1 pixel_6205/VBIAS pixel_6205/NB2 pixel_6205/AMP_IN pixel_6205/SF_IB
+ pixel_6205/PIX_OUT pixel_6205/CSA_VREF pixel
Xpixel_6216 pixel_6216/gring pixel_6216/VDD pixel_6216/GND pixel_6216/VREF pixel_6216/ROW_SEL
+ pixel_6216/NB1 pixel_6216/VBIAS pixel_6216/NB2 pixel_6216/AMP_IN pixel_6216/SF_IB
+ pixel_6216/PIX_OUT pixel_6216/CSA_VREF pixel
Xpixel_6227 pixel_6227/gring pixel_6227/VDD pixel_6227/GND pixel_6227/VREF pixel_6227/ROW_SEL
+ pixel_6227/NB1 pixel_6227/VBIAS pixel_6227/NB2 pixel_6227/AMP_IN pixel_6227/SF_IB
+ pixel_6227/PIX_OUT pixel_6227/CSA_VREF pixel
Xpixel_6238 pixel_6238/gring pixel_6238/VDD pixel_6238/GND pixel_6238/VREF pixel_6238/ROW_SEL
+ pixel_6238/NB1 pixel_6238/VBIAS pixel_6238/NB2 pixel_6238/AMP_IN pixel_6238/SF_IB
+ pixel_6238/PIX_OUT pixel_6238/CSA_VREF pixel
Xpixel_6249 pixel_6249/gring pixel_6249/VDD pixel_6249/GND pixel_6249/VREF pixel_6249/ROW_SEL
+ pixel_6249/NB1 pixel_6249/VBIAS pixel_6249/NB2 pixel_6249/AMP_IN pixel_6249/SF_IB
+ pixel_6249/PIX_OUT pixel_6249/CSA_VREF pixel
Xpixel_5504 pixel_5504/gring pixel_5504/VDD pixel_5504/GND pixel_5504/VREF pixel_5504/ROW_SEL
+ pixel_5504/NB1 pixel_5504/VBIAS pixel_5504/NB2 pixel_5504/AMP_IN pixel_5504/SF_IB
+ pixel_5504/PIX_OUT pixel_5504/CSA_VREF pixel
Xpixel_5515 pixel_5515/gring pixel_5515/VDD pixel_5515/GND pixel_5515/VREF pixel_5515/ROW_SEL
+ pixel_5515/NB1 pixel_5515/VBIAS pixel_5515/NB2 pixel_5515/AMP_IN pixel_5515/SF_IB
+ pixel_5515/PIX_OUT pixel_5515/CSA_VREF pixel
Xpixel_5526 pixel_5526/gring pixel_5526/VDD pixel_5526/GND pixel_5526/VREF pixel_5526/ROW_SEL
+ pixel_5526/NB1 pixel_5526/VBIAS pixel_5526/NB2 pixel_5526/AMP_IN pixel_5526/SF_IB
+ pixel_5526/PIX_OUT pixel_5526/CSA_VREF pixel
Xpixel_5537 pixel_5537/gring pixel_5537/VDD pixel_5537/GND pixel_5537/VREF pixel_5537/ROW_SEL
+ pixel_5537/NB1 pixel_5537/VBIAS pixel_5537/NB2 pixel_5537/AMP_IN pixel_5537/SF_IB
+ pixel_5537/PIX_OUT pixel_5537/CSA_VREF pixel
Xpixel_5548 pixel_5548/gring pixel_5548/VDD pixel_5548/GND pixel_5548/VREF pixel_5548/ROW_SEL
+ pixel_5548/NB1 pixel_5548/VBIAS pixel_5548/NB2 pixel_5548/AMP_IN pixel_5548/SF_IB
+ pixel_5548/PIX_OUT pixel_5548/CSA_VREF pixel
Xpixel_4803 pixel_4803/gring pixel_4803/VDD pixel_4803/GND pixel_4803/VREF pixel_4803/ROW_SEL
+ pixel_4803/NB1 pixel_4803/VBIAS pixel_4803/NB2 pixel_4803/AMP_IN pixel_4803/SF_IB
+ pixel_4803/PIX_OUT pixel_4803/CSA_VREF pixel
Xpixel_842 pixel_842/gring pixel_842/VDD pixel_842/GND pixel_842/VREF pixel_842/ROW_SEL
+ pixel_842/NB1 pixel_842/VBIAS pixel_842/NB2 pixel_842/AMP_IN pixel_842/SF_IB pixel_842/PIX_OUT
+ pixel_842/CSA_VREF pixel
Xpixel_831 pixel_831/gring pixel_831/VDD pixel_831/GND pixel_831/VREF pixel_831/ROW_SEL
+ pixel_831/NB1 pixel_831/VBIAS pixel_831/NB2 pixel_831/AMP_IN pixel_831/SF_IB pixel_831/PIX_OUT
+ pixel_831/CSA_VREF pixel
Xpixel_820 pixel_820/gring pixel_820/VDD pixel_820/GND pixel_820/VREF pixel_820/ROW_SEL
+ pixel_820/NB1 pixel_820/VBIAS pixel_820/NB2 pixel_820/AMP_IN pixel_820/SF_IB pixel_820/PIX_OUT
+ pixel_820/CSA_VREF pixel
Xpixel_5559 pixel_5559/gring pixel_5559/VDD pixel_5559/GND pixel_5559/VREF pixel_5559/ROW_SEL
+ pixel_5559/NB1 pixel_5559/VBIAS pixel_5559/NB2 pixel_5559/AMP_IN pixel_5559/SF_IB
+ pixel_5559/PIX_OUT pixel_5559/CSA_VREF pixel
Xpixel_4814 pixel_4814/gring pixel_4814/VDD pixel_4814/GND pixel_4814/VREF pixel_4814/ROW_SEL
+ pixel_4814/NB1 pixel_4814/VBIAS pixel_4814/NB2 pixel_4814/AMP_IN pixel_4814/SF_IB
+ pixel_4814/PIX_OUT pixel_4814/CSA_VREF pixel
Xpixel_4825 pixel_4825/gring pixel_4825/VDD pixel_4825/GND pixel_4825/VREF pixel_4825/ROW_SEL
+ pixel_4825/NB1 pixel_4825/VBIAS pixel_4825/NB2 pixel_4825/AMP_IN pixel_4825/SF_IB
+ pixel_4825/PIX_OUT pixel_4825/CSA_VREF pixel
Xpixel_4836 pixel_4836/gring pixel_4836/VDD pixel_4836/GND pixel_4836/VREF pixel_4836/ROW_SEL
+ pixel_4836/NB1 pixel_4836/VBIAS pixel_4836/NB2 pixel_4836/AMP_IN pixel_4836/SF_IB
+ pixel_4836/PIX_OUT pixel_4836/CSA_VREF pixel
Xpixel_4847 pixel_4847/gring pixel_4847/VDD pixel_4847/GND pixel_4847/VREF pixel_4847/ROW_SEL
+ pixel_4847/NB1 pixel_4847/VBIAS pixel_4847/NB2 pixel_4847/AMP_IN pixel_4847/SF_IB
+ pixel_4847/PIX_OUT pixel_4847/CSA_VREF pixel
Xpixel_875 pixel_875/gring pixel_875/VDD pixel_875/GND pixel_875/VREF pixel_875/ROW_SEL
+ pixel_875/NB1 pixel_875/VBIAS pixel_875/NB2 pixel_875/AMP_IN pixel_875/SF_IB pixel_875/PIX_OUT
+ pixel_875/CSA_VREF pixel
Xpixel_864 pixel_864/gring pixel_864/VDD pixel_864/GND pixel_864/VREF pixel_864/ROW_SEL
+ pixel_864/NB1 pixel_864/VBIAS pixel_864/NB2 pixel_864/AMP_IN pixel_864/SF_IB pixel_864/PIX_OUT
+ pixel_864/CSA_VREF pixel
Xpixel_853 pixel_853/gring pixel_853/VDD pixel_853/GND pixel_853/VREF pixel_853/ROW_SEL
+ pixel_853/NB1 pixel_853/VBIAS pixel_853/NB2 pixel_853/AMP_IN pixel_853/SF_IB pixel_853/PIX_OUT
+ pixel_853/CSA_VREF pixel
Xpixel_4858 pixel_4858/gring pixel_4858/VDD pixel_4858/GND pixel_4858/VREF pixel_4858/ROW_SEL
+ pixel_4858/NB1 pixel_4858/VBIAS pixel_4858/NB2 pixel_4858/AMP_IN pixel_4858/SF_IB
+ pixel_4858/PIX_OUT pixel_4858/CSA_VREF pixel
Xpixel_4869 pixel_4869/gring pixel_4869/VDD pixel_4869/GND pixel_4869/VREF pixel_4869/ROW_SEL
+ pixel_4869/NB1 pixel_4869/VBIAS pixel_4869/NB2 pixel_4869/AMP_IN pixel_4869/SF_IB
+ pixel_4869/PIX_OUT pixel_4869/CSA_VREF pixel
Xpixel_897 pixel_897/gring pixel_897/VDD pixel_897/GND pixel_897/VREF pixel_897/ROW_SEL
+ pixel_897/NB1 pixel_897/VBIAS pixel_897/NB2 pixel_897/AMP_IN pixel_897/SF_IB pixel_897/PIX_OUT
+ pixel_897/CSA_VREF pixel
Xpixel_886 pixel_886/gring pixel_886/VDD pixel_886/GND pixel_886/VREF pixel_886/ROW_SEL
+ pixel_886/NB1 pixel_886/VBIAS pixel_886/NB2 pixel_886/AMP_IN pixel_886/SF_IB pixel_886/PIX_OUT
+ pixel_886/CSA_VREF pixel
Xpixel_8130 pixel_8130/gring pixel_8130/VDD pixel_8130/GND pixel_8130/VREF pixel_8130/ROW_SEL
+ pixel_8130/NB1 pixel_8130/VBIAS pixel_8130/NB2 pixel_8130/AMP_IN pixel_8130/SF_IB
+ pixel_8130/PIX_OUT pixel_8130/CSA_VREF pixel
Xpixel_8141 pixel_8141/gring pixel_8141/VDD pixel_8141/GND pixel_8141/VREF pixel_8141/ROW_SEL
+ pixel_8141/NB1 pixel_8141/VBIAS pixel_8141/NB2 pixel_8141/AMP_IN pixel_8141/SF_IB
+ pixel_8141/PIX_OUT pixel_8141/CSA_VREF pixel
Xpixel_8152 pixel_8152/gring pixel_8152/VDD pixel_8152/GND pixel_8152/VREF pixel_8152/ROW_SEL
+ pixel_8152/NB1 pixel_8152/VBIAS pixel_8152/NB2 pixel_8152/AMP_IN pixel_8152/SF_IB
+ pixel_8152/PIX_OUT pixel_8152/CSA_VREF pixel
Xpixel_8163 pixel_8163/gring pixel_8163/VDD pixel_8163/GND pixel_8163/VREF pixel_8163/ROW_SEL
+ pixel_8163/NB1 pixel_8163/VBIAS pixel_8163/NB2 pixel_8163/AMP_IN pixel_8163/SF_IB
+ pixel_8163/PIX_OUT pixel_8163/CSA_VREF pixel
Xpixel_8174 pixel_8174/gring pixel_8174/VDD pixel_8174/GND pixel_8174/VREF pixel_8174/ROW_SEL
+ pixel_8174/NB1 pixel_8174/VBIAS pixel_8174/NB2 pixel_8174/AMP_IN pixel_8174/SF_IB
+ pixel_8174/PIX_OUT pixel_8174/CSA_VREF pixel
Xpixel_8185 pixel_8185/gring pixel_8185/VDD pixel_8185/GND pixel_8185/VREF pixel_8185/ROW_SEL
+ pixel_8185/NB1 pixel_8185/VBIAS pixel_8185/NB2 pixel_8185/AMP_IN pixel_8185/SF_IB
+ pixel_8185/PIX_OUT pixel_8185/CSA_VREF pixel
Xpixel_7440 pixel_7440/gring pixel_7440/VDD pixel_7440/GND pixel_7440/VREF pixel_7440/ROW_SEL
+ pixel_7440/NB1 pixel_7440/VBIAS pixel_7440/NB2 pixel_7440/AMP_IN pixel_7440/SF_IB
+ pixel_7440/PIX_OUT pixel_7440/CSA_VREF pixel
Xpixel_8196 pixel_8196/gring pixel_8196/VDD pixel_8196/GND pixel_8196/VREF pixel_8196/ROW_SEL
+ pixel_8196/NB1 pixel_8196/VBIAS pixel_8196/NB2 pixel_8196/AMP_IN pixel_8196/SF_IB
+ pixel_8196/PIX_OUT pixel_8196/CSA_VREF pixel
Xpixel_7451 pixel_7451/gring pixel_7451/VDD pixel_7451/GND pixel_7451/VREF pixel_7451/ROW_SEL
+ pixel_7451/NB1 pixel_7451/VBIAS pixel_7451/NB2 pixel_7451/AMP_IN pixel_7451/SF_IB
+ pixel_7451/PIX_OUT pixel_7451/CSA_VREF pixel
Xpixel_7462 pixel_7462/gring pixel_7462/VDD pixel_7462/GND pixel_7462/VREF pixel_7462/ROW_SEL
+ pixel_7462/NB1 pixel_7462/VBIAS pixel_7462/NB2 pixel_7462/AMP_IN pixel_7462/SF_IB
+ pixel_7462/PIX_OUT pixel_7462/CSA_VREF pixel
Xpixel_7473 pixel_7473/gring pixel_7473/VDD pixel_7473/GND pixel_7473/VREF pixel_7473/ROW_SEL
+ pixel_7473/NB1 pixel_7473/VBIAS pixel_7473/NB2 pixel_7473/AMP_IN pixel_7473/SF_IB
+ pixel_7473/PIX_OUT pixel_7473/CSA_VREF pixel
Xpixel_7484 pixel_7484/gring pixel_7484/VDD pixel_7484/GND pixel_7484/VREF pixel_7484/ROW_SEL
+ pixel_7484/NB1 pixel_7484/VBIAS pixel_7484/NB2 pixel_7484/AMP_IN pixel_7484/SF_IB
+ pixel_7484/PIX_OUT pixel_7484/CSA_VREF pixel
Xpixel_7495 pixel_7495/gring pixel_7495/VDD pixel_7495/GND pixel_7495/VREF pixel_7495/ROW_SEL
+ pixel_7495/NB1 pixel_7495/VBIAS pixel_7495/NB2 pixel_7495/AMP_IN pixel_7495/SF_IB
+ pixel_7495/PIX_OUT pixel_7495/CSA_VREF pixel
Xpixel_6750 pixel_6750/gring pixel_6750/VDD pixel_6750/GND pixel_6750/VREF pixel_6750/ROW_SEL
+ pixel_6750/NB1 pixel_6750/VBIAS pixel_6750/NB2 pixel_6750/AMP_IN pixel_6750/SF_IB
+ pixel_6750/PIX_OUT pixel_6750/CSA_VREF pixel
Xpixel_6761 pixel_6761/gring pixel_6761/VDD pixel_6761/GND pixel_6761/VREF pixel_6761/ROW_SEL
+ pixel_6761/NB1 pixel_6761/VBIAS pixel_6761/NB2 pixel_6761/AMP_IN pixel_6761/SF_IB
+ pixel_6761/PIX_OUT pixel_6761/CSA_VREF pixel
Xpixel_6772 pixel_6772/gring pixel_6772/VDD pixel_6772/GND pixel_6772/VREF pixel_6772/ROW_SEL
+ pixel_6772/NB1 pixel_6772/VBIAS pixel_6772/NB2 pixel_6772/AMP_IN pixel_6772/SF_IB
+ pixel_6772/PIX_OUT pixel_6772/CSA_VREF pixel
Xpixel_6783 pixel_6783/gring pixel_6783/VDD pixel_6783/GND pixel_6783/VREF pixel_6783/ROW_SEL
+ pixel_6783/NB1 pixel_6783/VBIAS pixel_6783/NB2 pixel_6783/AMP_IN pixel_6783/SF_IB
+ pixel_6783/PIX_OUT pixel_6783/CSA_VREF pixel
Xpixel_6794 pixel_6794/gring pixel_6794/VDD pixel_6794/GND pixel_6794/VREF pixel_6794/ROW_SEL
+ pixel_6794/NB1 pixel_6794/VBIAS pixel_6794/NB2 pixel_6794/AMP_IN pixel_6794/SF_IB
+ pixel_6794/PIX_OUT pixel_6794/CSA_VREF pixel
Xpixel_1090 pixel_1090/gring pixel_1090/VDD pixel_1090/GND pixel_1090/VREF pixel_1090/ROW_SEL
+ pixel_1090/NB1 pixel_1090/VBIAS pixel_1090/NB2 pixel_1090/AMP_IN pixel_1090/SF_IB
+ pixel_1090/PIX_OUT pixel_1090/CSA_VREF pixel
Xpixel_127 pixel_127/gring pixel_127/VDD pixel_127/GND pixel_127/VREF pixel_127/ROW_SEL
+ pixel_127/NB1 pixel_127/VBIAS pixel_127/NB2 pixel_127/AMP_IN pixel_127/SF_IB pixel_127/PIX_OUT
+ pixel_127/CSA_VREF pixel
Xpixel_116 pixel_116/gring pixel_116/VDD pixel_116/GND pixel_116/VREF pixel_116/ROW_SEL
+ pixel_116/NB1 pixel_116/VBIAS pixel_116/NB2 pixel_116/AMP_IN pixel_116/SF_IB pixel_116/PIX_OUT
+ pixel_116/CSA_VREF pixel
Xpixel_105 pixel_105/gring pixel_105/VDD pixel_105/GND pixel_105/VREF pixel_105/ROW_SEL
+ pixel_105/NB1 pixel_105/VBIAS pixel_105/NB2 pixel_105/AMP_IN pixel_105/SF_IB pixel_105/PIX_OUT
+ pixel_105/CSA_VREF pixel
Xpixel_149 pixel_149/gring pixel_149/VDD pixel_149/GND pixel_149/VREF pixel_149/ROW_SEL
+ pixel_149/NB1 pixel_149/VBIAS pixel_149/NB2 pixel_149/AMP_IN pixel_149/SF_IB pixel_149/PIX_OUT
+ pixel_149/CSA_VREF pixel
Xpixel_138 pixel_138/gring pixel_138/VDD pixel_138/GND pixel_138/VREF pixel_138/ROW_SEL
+ pixel_138/NB1 pixel_138/VBIAS pixel_138/NB2 pixel_138/AMP_IN pixel_138/SF_IB pixel_138/PIX_OUT
+ pixel_138/CSA_VREF pixel
Xpixel_3409 pixel_3409/gring pixel_3409/VDD pixel_3409/GND pixel_3409/VREF pixel_3409/ROW_SEL
+ pixel_3409/NB1 pixel_3409/VBIAS pixel_3409/NB2 pixel_3409/AMP_IN pixel_3409/SF_IB
+ pixel_3409/PIX_OUT pixel_3409/CSA_VREF pixel
Xpixel_2719 pixel_2719/gring pixel_2719/VDD pixel_2719/GND pixel_2719/VREF pixel_2719/ROW_SEL
+ pixel_2719/NB1 pixel_2719/VBIAS pixel_2719/NB2 pixel_2719/AMP_IN pixel_2719/SF_IB
+ pixel_2719/PIX_OUT pixel_2719/CSA_VREF pixel
Xpixel_2708 pixel_2708/gring pixel_2708/VDD pixel_2708/GND pixel_2708/VREF pixel_2708/ROW_SEL
+ pixel_2708/NB1 pixel_2708/VBIAS pixel_2708/NB2 pixel_2708/AMP_IN pixel_2708/SF_IB
+ pixel_2708/PIX_OUT pixel_2708/CSA_VREF pixel
Xpixel_6002 pixel_6002/gring pixel_6002/VDD pixel_6002/GND pixel_6002/VREF pixel_6002/ROW_SEL
+ pixel_6002/NB1 pixel_6002/VBIAS pixel_6002/NB2 pixel_6002/AMP_IN pixel_6002/SF_IB
+ pixel_6002/PIX_OUT pixel_6002/CSA_VREF pixel
Xpixel_6013 pixel_6013/gring pixel_6013/VDD pixel_6013/GND pixel_6013/VREF pixel_6013/ROW_SEL
+ pixel_6013/NB1 pixel_6013/VBIAS pixel_6013/NB2 pixel_6013/AMP_IN pixel_6013/SF_IB
+ pixel_6013/PIX_OUT pixel_6013/CSA_VREF pixel
Xpixel_6024 pixel_6024/gring pixel_6024/VDD pixel_6024/GND pixel_6024/VREF pixel_6024/ROW_SEL
+ pixel_6024/NB1 pixel_6024/VBIAS pixel_6024/NB2 pixel_6024/AMP_IN pixel_6024/SF_IB
+ pixel_6024/PIX_OUT pixel_6024/CSA_VREF pixel
Xpixel_6035 pixel_6035/gring pixel_6035/VDD pixel_6035/GND pixel_6035/VREF pixel_6035/ROW_SEL
+ pixel_6035/NB1 pixel_6035/VBIAS pixel_6035/NB2 pixel_6035/AMP_IN pixel_6035/SF_IB
+ pixel_6035/PIX_OUT pixel_6035/CSA_VREF pixel
Xpixel_6046 pixel_6046/gring pixel_6046/VDD pixel_6046/GND pixel_6046/VREF pixel_6046/ROW_SEL
+ pixel_6046/NB1 pixel_6046/VBIAS pixel_6046/NB2 pixel_6046/AMP_IN pixel_6046/SF_IB
+ pixel_6046/PIX_OUT pixel_6046/CSA_VREF pixel
Xpixel_6057 pixel_6057/gring pixel_6057/VDD pixel_6057/GND pixel_6057/VREF pixel_6057/ROW_SEL
+ pixel_6057/NB1 pixel_6057/VBIAS pixel_6057/NB2 pixel_6057/AMP_IN pixel_6057/SF_IB
+ pixel_6057/PIX_OUT pixel_6057/CSA_VREF pixel
Xpixel_6068 pixel_6068/gring pixel_6068/VDD pixel_6068/GND pixel_6068/VREF pixel_6068/ROW_SEL
+ pixel_6068/NB1 pixel_6068/VBIAS pixel_6068/NB2 pixel_6068/AMP_IN pixel_6068/SF_IB
+ pixel_6068/PIX_OUT pixel_6068/CSA_VREF pixel
Xpixel_5301 pixel_5301/gring pixel_5301/VDD pixel_5301/GND pixel_5301/VREF pixel_5301/ROW_SEL
+ pixel_5301/NB1 pixel_5301/VBIAS pixel_5301/NB2 pixel_5301/AMP_IN pixel_5301/SF_IB
+ pixel_5301/PIX_OUT pixel_5301/CSA_VREF pixel
Xpixel_5312 pixel_5312/gring pixel_5312/VDD pixel_5312/GND pixel_5312/VREF pixel_5312/ROW_SEL
+ pixel_5312/NB1 pixel_5312/VBIAS pixel_5312/NB2 pixel_5312/AMP_IN pixel_5312/SF_IB
+ pixel_5312/PIX_OUT pixel_5312/CSA_VREF pixel
Xpixel_5323 pixel_5323/gring pixel_5323/VDD pixel_5323/GND pixel_5323/VREF pixel_5323/ROW_SEL
+ pixel_5323/NB1 pixel_5323/VBIAS pixel_5323/NB2 pixel_5323/AMP_IN pixel_5323/SF_IB
+ pixel_5323/PIX_OUT pixel_5323/CSA_VREF pixel
Xpixel_6079 pixel_6079/gring pixel_6079/VDD pixel_6079/GND pixel_6079/VREF pixel_6079/ROW_SEL
+ pixel_6079/NB1 pixel_6079/VBIAS pixel_6079/NB2 pixel_6079/AMP_IN pixel_6079/SF_IB
+ pixel_6079/PIX_OUT pixel_6079/CSA_VREF pixel
Xpixel_5334 pixel_5334/gring pixel_5334/VDD pixel_5334/GND pixel_5334/VREF pixel_5334/ROW_SEL
+ pixel_5334/NB1 pixel_5334/VBIAS pixel_5334/NB2 pixel_5334/AMP_IN pixel_5334/SF_IB
+ pixel_5334/PIX_OUT pixel_5334/CSA_VREF pixel
Xpixel_5345 pixel_5345/gring pixel_5345/VDD pixel_5345/GND pixel_5345/VREF pixel_5345/ROW_SEL
+ pixel_5345/NB1 pixel_5345/VBIAS pixel_5345/NB2 pixel_5345/AMP_IN pixel_5345/SF_IB
+ pixel_5345/PIX_OUT pixel_5345/CSA_VREF pixel
Xpixel_5356 pixel_5356/gring pixel_5356/VDD pixel_5356/GND pixel_5356/VREF pixel_5356/ROW_SEL
+ pixel_5356/NB1 pixel_5356/VBIAS pixel_5356/NB2 pixel_5356/AMP_IN pixel_5356/SF_IB
+ pixel_5356/PIX_OUT pixel_5356/CSA_VREF pixel
Xpixel_4600 pixel_4600/gring pixel_4600/VDD pixel_4600/GND pixel_4600/VREF pixel_4600/ROW_SEL
+ pixel_4600/NB1 pixel_4600/VBIAS pixel_4600/NB2 pixel_4600/AMP_IN pixel_4600/SF_IB
+ pixel_4600/PIX_OUT pixel_4600/CSA_VREF pixel
Xpixel_4611 pixel_4611/gring pixel_4611/VDD pixel_4611/GND pixel_4611/VREF pixel_4611/ROW_SEL
+ pixel_4611/NB1 pixel_4611/VBIAS pixel_4611/NB2 pixel_4611/AMP_IN pixel_4611/SF_IB
+ pixel_4611/PIX_OUT pixel_4611/CSA_VREF pixel
Xpixel_650 pixel_650/gring pixel_650/VDD pixel_650/GND pixel_650/VREF pixel_650/ROW_SEL
+ pixel_650/NB1 pixel_650/VBIAS pixel_650/NB2 pixel_650/AMP_IN pixel_650/SF_IB pixel_650/PIX_OUT
+ pixel_650/CSA_VREF pixel
Xpixel_5367 pixel_5367/gring pixel_5367/VDD pixel_5367/GND pixel_5367/VREF pixel_5367/ROW_SEL
+ pixel_5367/NB1 pixel_5367/VBIAS pixel_5367/NB2 pixel_5367/AMP_IN pixel_5367/SF_IB
+ pixel_5367/PIX_OUT pixel_5367/CSA_VREF pixel
Xpixel_5378 pixel_5378/gring pixel_5378/VDD pixel_5378/GND pixel_5378/VREF pixel_5378/ROW_SEL
+ pixel_5378/NB1 pixel_5378/VBIAS pixel_5378/NB2 pixel_5378/AMP_IN pixel_5378/SF_IB
+ pixel_5378/PIX_OUT pixel_5378/CSA_VREF pixel
Xpixel_5389 pixel_5389/gring pixel_5389/VDD pixel_5389/GND pixel_5389/VREF pixel_5389/ROW_SEL
+ pixel_5389/NB1 pixel_5389/VBIAS pixel_5389/NB2 pixel_5389/AMP_IN pixel_5389/SF_IB
+ pixel_5389/PIX_OUT pixel_5389/CSA_VREF pixel
Xpixel_4622 pixel_4622/gring pixel_4622/VDD pixel_4622/GND pixel_4622/VREF pixel_4622/ROW_SEL
+ pixel_4622/NB1 pixel_4622/VBIAS pixel_4622/NB2 pixel_4622/AMP_IN pixel_4622/SF_IB
+ pixel_4622/PIX_OUT pixel_4622/CSA_VREF pixel
Xpixel_4633 pixel_4633/gring pixel_4633/VDD pixel_4633/GND pixel_4633/VREF pixel_4633/ROW_SEL
+ pixel_4633/NB1 pixel_4633/VBIAS pixel_4633/NB2 pixel_4633/AMP_IN pixel_4633/SF_IB
+ pixel_4633/PIX_OUT pixel_4633/CSA_VREF pixel
Xpixel_4644 pixel_4644/gring pixel_4644/VDD pixel_4644/GND pixel_4644/VREF pixel_4644/ROW_SEL
+ pixel_4644/NB1 pixel_4644/VBIAS pixel_4644/NB2 pixel_4644/AMP_IN pixel_4644/SF_IB
+ pixel_4644/PIX_OUT pixel_4644/CSA_VREF pixel
Xpixel_4655 pixel_4655/gring pixel_4655/VDD pixel_4655/GND pixel_4655/VREF pixel_4655/ROW_SEL
+ pixel_4655/NB1 pixel_4655/VBIAS pixel_4655/NB2 pixel_4655/AMP_IN pixel_4655/SF_IB
+ pixel_4655/PIX_OUT pixel_4655/CSA_VREF pixel
Xpixel_3910 pixel_3910/gring pixel_3910/VDD pixel_3910/GND pixel_3910/VREF pixel_3910/ROW_SEL
+ pixel_3910/NB1 pixel_3910/VBIAS pixel_3910/NB2 pixel_3910/AMP_IN pixel_3910/SF_IB
+ pixel_3910/PIX_OUT pixel_3910/CSA_VREF pixel
Xpixel_683 pixel_683/gring pixel_683/VDD pixel_683/GND pixel_683/VREF pixel_683/ROW_SEL
+ pixel_683/NB1 pixel_683/VBIAS pixel_683/NB2 pixel_683/AMP_IN pixel_683/SF_IB pixel_683/PIX_OUT
+ pixel_683/CSA_VREF pixel
Xpixel_672 pixel_672/gring pixel_672/VDD pixel_672/GND pixel_672/VREF pixel_672/ROW_SEL
+ pixel_672/NB1 pixel_672/VBIAS pixel_672/NB2 pixel_672/AMP_IN pixel_672/SF_IB pixel_672/PIX_OUT
+ pixel_672/CSA_VREF pixel
Xpixel_661 pixel_661/gring pixel_661/VDD pixel_661/GND pixel_661/VREF pixel_661/ROW_SEL
+ pixel_661/NB1 pixel_661/VBIAS pixel_661/NB2 pixel_661/AMP_IN pixel_661/SF_IB pixel_661/PIX_OUT
+ pixel_661/CSA_VREF pixel
Xpixel_4666 pixel_4666/gring pixel_4666/VDD pixel_4666/GND pixel_4666/VREF pixel_4666/ROW_SEL
+ pixel_4666/NB1 pixel_4666/VBIAS pixel_4666/NB2 pixel_4666/AMP_IN pixel_4666/SF_IB
+ pixel_4666/PIX_OUT pixel_4666/CSA_VREF pixel
Xpixel_4677 pixel_4677/gring pixel_4677/VDD pixel_4677/GND pixel_4677/VREF pixel_4677/ROW_SEL
+ pixel_4677/NB1 pixel_4677/VBIAS pixel_4677/NB2 pixel_4677/AMP_IN pixel_4677/SF_IB
+ pixel_4677/PIX_OUT pixel_4677/CSA_VREF pixel
Xpixel_4688 pixel_4688/gring pixel_4688/VDD pixel_4688/GND pixel_4688/VREF pixel_4688/ROW_SEL
+ pixel_4688/NB1 pixel_4688/VBIAS pixel_4688/NB2 pixel_4688/AMP_IN pixel_4688/SF_IB
+ pixel_4688/PIX_OUT pixel_4688/CSA_VREF pixel
Xpixel_3921 pixel_3921/gring pixel_3921/VDD pixel_3921/GND pixel_3921/VREF pixel_3921/ROW_SEL
+ pixel_3921/NB1 pixel_3921/VBIAS pixel_3921/NB2 pixel_3921/AMP_IN pixel_3921/SF_IB
+ pixel_3921/PIX_OUT pixel_3921/CSA_VREF pixel
Xpixel_3932 pixel_3932/gring pixel_3932/VDD pixel_3932/GND pixel_3932/VREF pixel_3932/ROW_SEL
+ pixel_3932/NB1 pixel_3932/VBIAS pixel_3932/NB2 pixel_3932/AMP_IN pixel_3932/SF_IB
+ pixel_3932/PIX_OUT pixel_3932/CSA_VREF pixel
Xpixel_3943 pixel_3943/gring pixel_3943/VDD pixel_3943/GND pixel_3943/VREF pixel_3943/ROW_SEL
+ pixel_3943/NB1 pixel_3943/VBIAS pixel_3943/NB2 pixel_3943/AMP_IN pixel_3943/SF_IB
+ pixel_3943/PIX_OUT pixel_3943/CSA_VREF pixel
Xpixel_694 pixel_694/gring pixel_694/VDD pixel_694/GND pixel_694/VREF pixel_694/ROW_SEL
+ pixel_694/NB1 pixel_694/VBIAS pixel_694/NB2 pixel_694/AMP_IN pixel_694/SF_IB pixel_694/PIX_OUT
+ pixel_694/CSA_VREF pixel
Xpixel_4699 pixel_4699/gring pixel_4699/VDD pixel_4699/GND pixel_4699/VREF pixel_4699/ROW_SEL
+ pixel_4699/NB1 pixel_4699/VBIAS pixel_4699/NB2 pixel_4699/AMP_IN pixel_4699/SF_IB
+ pixel_4699/PIX_OUT pixel_4699/CSA_VREF pixel
Xpixel_3954 pixel_3954/gring pixel_3954/VDD pixel_3954/GND pixel_3954/VREF pixel_3954/ROW_SEL
+ pixel_3954/NB1 pixel_3954/VBIAS pixel_3954/NB2 pixel_3954/AMP_IN pixel_3954/SF_IB
+ pixel_3954/PIX_OUT pixel_3954/CSA_VREF pixel
Xpixel_3965 pixel_3965/gring pixel_3965/VDD pixel_3965/GND pixel_3965/VREF pixel_3965/ROW_SEL
+ pixel_3965/NB1 pixel_3965/VBIAS pixel_3965/NB2 pixel_3965/AMP_IN pixel_3965/SF_IB
+ pixel_3965/PIX_OUT pixel_3965/CSA_VREF pixel
Xpixel_3976 pixel_3976/gring pixel_3976/VDD pixel_3976/GND pixel_3976/VREF pixel_3976/ROW_SEL
+ pixel_3976/NB1 pixel_3976/VBIAS pixel_3976/NB2 pixel_3976/AMP_IN pixel_3976/SF_IB
+ pixel_3976/PIX_OUT pixel_3976/CSA_VREF pixel
Xpixel_3987 pixel_3987/gring pixel_3987/VDD pixel_3987/GND pixel_3987/VREF pixel_3987/ROW_SEL
+ pixel_3987/NB1 pixel_3987/VBIAS pixel_3987/NB2 pixel_3987/AMP_IN pixel_3987/SF_IB
+ pixel_3987/PIX_OUT pixel_3987/CSA_VREF pixel
Xpixel_3998 pixel_3998/gring pixel_3998/VDD pixel_3998/GND pixel_3998/VREF pixel_3998/ROW_SEL
+ pixel_3998/NB1 pixel_3998/VBIAS pixel_3998/NB2 pixel_3998/AMP_IN pixel_3998/SF_IB
+ pixel_3998/PIX_OUT pixel_3998/CSA_VREF pixel
Xpixel_8 pixel_8/gring pixel_8/VDD pixel_8/GND pixel_8/VREF pixel_8/ROW_SEL pixel_8/NB1
+ pixel_8/VBIAS pixel_8/NB2 pixel_8/AMP_IN pixel_8/SF_IB pixel_8/PIX_OUT pixel_8/CSA_VREF
+ pixel
Xpixel_7270 pixel_7270/gring pixel_7270/VDD pixel_7270/GND pixel_7270/VREF pixel_7270/ROW_SEL
+ pixel_7270/NB1 pixel_7270/VBIAS pixel_7270/NB2 pixel_7270/AMP_IN pixel_7270/SF_IB
+ pixel_7270/PIX_OUT pixel_7270/CSA_VREF pixel
Xpixel_7281 pixel_7281/gring pixel_7281/VDD pixel_7281/GND pixel_7281/VREF pixel_7281/ROW_SEL
+ pixel_7281/NB1 pixel_7281/VBIAS pixel_7281/NB2 pixel_7281/AMP_IN pixel_7281/SF_IB
+ pixel_7281/PIX_OUT pixel_7281/CSA_VREF pixel
Xpixel_7292 pixel_7292/gring pixel_7292/VDD pixel_7292/GND pixel_7292/VREF pixel_7292/ROW_SEL
+ pixel_7292/NB1 pixel_7292/VBIAS pixel_7292/NB2 pixel_7292/AMP_IN pixel_7292/SF_IB
+ pixel_7292/PIX_OUT pixel_7292/CSA_VREF pixel
Xpixel_6580 pixel_6580/gring pixel_6580/VDD pixel_6580/GND pixel_6580/VREF pixel_6580/ROW_SEL
+ pixel_6580/NB1 pixel_6580/VBIAS pixel_6580/NB2 pixel_6580/AMP_IN pixel_6580/SF_IB
+ pixel_6580/PIX_OUT pixel_6580/CSA_VREF pixel
Xpixel_6591 pixel_6591/gring pixel_6591/VDD pixel_6591/GND pixel_6591/VREF pixel_6591/ROW_SEL
+ pixel_6591/NB1 pixel_6591/VBIAS pixel_6591/NB2 pixel_6591/AMP_IN pixel_6591/SF_IB
+ pixel_6591/PIX_OUT pixel_6591/CSA_VREF pixel
Xpixel_5890 pixel_5890/gring pixel_5890/VDD pixel_5890/GND pixel_5890/VREF pixel_5890/ROW_SEL
+ pixel_5890/NB1 pixel_5890/VBIAS pixel_5890/NB2 pixel_5890/AMP_IN pixel_5890/SF_IB
+ pixel_5890/PIX_OUT pixel_5890/CSA_VREF pixel
Xpixel_3206 pixel_3206/gring pixel_3206/VDD pixel_3206/GND pixel_3206/VREF pixel_3206/ROW_SEL
+ pixel_3206/NB1 pixel_3206/VBIAS pixel_3206/NB2 pixel_3206/AMP_IN pixel_3206/SF_IB
+ pixel_3206/PIX_OUT pixel_3206/CSA_VREF pixel
Xpixel_3239 pixel_3239/gring pixel_3239/VDD pixel_3239/GND pixel_3239/VREF pixel_3239/ROW_SEL
+ pixel_3239/NB1 pixel_3239/VBIAS pixel_3239/NB2 pixel_3239/AMP_IN pixel_3239/SF_IB
+ pixel_3239/PIX_OUT pixel_3239/CSA_VREF pixel
Xpixel_3228 pixel_3228/gring pixel_3228/VDD pixel_3228/GND pixel_3228/VREF pixel_3228/ROW_SEL
+ pixel_3228/NB1 pixel_3228/VBIAS pixel_3228/NB2 pixel_3228/AMP_IN pixel_3228/SF_IB
+ pixel_3228/PIX_OUT pixel_3228/CSA_VREF pixel
Xpixel_3217 pixel_3217/gring pixel_3217/VDD pixel_3217/GND pixel_3217/VREF pixel_3217/ROW_SEL
+ pixel_3217/NB1 pixel_3217/VBIAS pixel_3217/NB2 pixel_3217/AMP_IN pixel_3217/SF_IB
+ pixel_3217/PIX_OUT pixel_3217/CSA_VREF pixel
Xpixel_2527 pixel_2527/gring pixel_2527/VDD pixel_2527/GND pixel_2527/VREF pixel_2527/ROW_SEL
+ pixel_2527/NB1 pixel_2527/VBIAS pixel_2527/NB2 pixel_2527/AMP_IN pixel_2527/SF_IB
+ pixel_2527/PIX_OUT pixel_2527/CSA_VREF pixel
Xpixel_2516 pixel_2516/gring pixel_2516/VDD pixel_2516/GND pixel_2516/VREF pixel_2516/ROW_SEL
+ pixel_2516/NB1 pixel_2516/VBIAS pixel_2516/NB2 pixel_2516/AMP_IN pixel_2516/SF_IB
+ pixel_2516/PIX_OUT pixel_2516/CSA_VREF pixel
Xpixel_2505 pixel_2505/gring pixel_2505/VDD pixel_2505/GND pixel_2505/VREF pixel_2505/ROW_SEL
+ pixel_2505/NB1 pixel_2505/VBIAS pixel_2505/NB2 pixel_2505/AMP_IN pixel_2505/SF_IB
+ pixel_2505/PIX_OUT pixel_2505/CSA_VREF pixel
Xpixel_1826 pixel_1826/gring pixel_1826/VDD pixel_1826/GND pixel_1826/VREF pixel_1826/ROW_SEL
+ pixel_1826/NB1 pixel_1826/VBIAS pixel_1826/NB2 pixel_1826/AMP_IN pixel_1826/SF_IB
+ pixel_1826/PIX_OUT pixel_1826/CSA_VREF pixel
Xpixel_1815 pixel_1815/gring pixel_1815/VDD pixel_1815/GND pixel_1815/VREF pixel_1815/ROW_SEL
+ pixel_1815/NB1 pixel_1815/VBIAS pixel_1815/NB2 pixel_1815/AMP_IN pixel_1815/SF_IB
+ pixel_1815/PIX_OUT pixel_1815/CSA_VREF pixel
Xpixel_1804 pixel_1804/gring pixel_1804/VDD pixel_1804/GND pixel_1804/VREF pixel_1804/ROW_SEL
+ pixel_1804/NB1 pixel_1804/VBIAS pixel_1804/NB2 pixel_1804/AMP_IN pixel_1804/SF_IB
+ pixel_1804/PIX_OUT pixel_1804/CSA_VREF pixel
Xpixel_2549 pixel_2549/gring pixel_2549/VDD pixel_2549/GND pixel_2549/VREF pixel_2549/ROW_SEL
+ pixel_2549/NB1 pixel_2549/VBIAS pixel_2549/NB2 pixel_2549/AMP_IN pixel_2549/SF_IB
+ pixel_2549/PIX_OUT pixel_2549/CSA_VREF pixel
Xpixel_2538 pixel_2538/gring pixel_2538/VDD pixel_2538/GND pixel_2538/VREF pixel_2538/ROW_SEL
+ pixel_2538/NB1 pixel_2538/VBIAS pixel_2538/NB2 pixel_2538/AMP_IN pixel_2538/SF_IB
+ pixel_2538/PIX_OUT pixel_2538/CSA_VREF pixel
Xpixel_1859 pixel_1859/gring pixel_1859/VDD pixel_1859/GND pixel_1859/VREF pixel_1859/ROW_SEL
+ pixel_1859/NB1 pixel_1859/VBIAS pixel_1859/NB2 pixel_1859/AMP_IN pixel_1859/SF_IB
+ pixel_1859/PIX_OUT pixel_1859/CSA_VREF pixel
Xpixel_1848 pixel_1848/gring pixel_1848/VDD pixel_1848/GND pixel_1848/VREF pixel_1848/ROW_SEL
+ pixel_1848/NB1 pixel_1848/VBIAS pixel_1848/NB2 pixel_1848/AMP_IN pixel_1848/SF_IB
+ pixel_1848/PIX_OUT pixel_1848/CSA_VREF pixel
Xpixel_1837 pixel_1837/gring pixel_1837/VDD pixel_1837/GND pixel_1837/VREF pixel_1837/ROW_SEL
+ pixel_1837/NB1 pixel_1837/VBIAS pixel_1837/NB2 pixel_1837/AMP_IN pixel_1837/SF_IB
+ pixel_1837/PIX_OUT pixel_1837/CSA_VREF pixel
Xpixel_5120 pixel_5120/gring pixel_5120/VDD pixel_5120/GND pixel_5120/VREF pixel_5120/ROW_SEL
+ pixel_5120/NB1 pixel_5120/VBIAS pixel_5120/NB2 pixel_5120/AMP_IN pixel_5120/SF_IB
+ pixel_5120/PIX_OUT pixel_5120/CSA_VREF pixel
Xpixel_5131 pixel_5131/gring pixel_5131/VDD pixel_5131/GND pixel_5131/VREF pixel_5131/ROW_SEL
+ pixel_5131/NB1 pixel_5131/VBIAS pixel_5131/NB2 pixel_5131/AMP_IN pixel_5131/SF_IB
+ pixel_5131/PIX_OUT pixel_5131/CSA_VREF pixel
Xpixel_5142 pixel_5142/gring pixel_5142/VDD pixel_5142/GND pixel_5142/VREF pixel_5142/ROW_SEL
+ pixel_5142/NB1 pixel_5142/VBIAS pixel_5142/NB2 pixel_5142/AMP_IN pixel_5142/SF_IB
+ pixel_5142/PIX_OUT pixel_5142/CSA_VREF pixel
Xpixel_5153 pixel_5153/gring pixel_5153/VDD pixel_5153/GND pixel_5153/VREF pixel_5153/ROW_SEL
+ pixel_5153/NB1 pixel_5153/VBIAS pixel_5153/NB2 pixel_5153/AMP_IN pixel_5153/SF_IB
+ pixel_5153/PIX_OUT pixel_5153/CSA_VREF pixel
Xpixel_5164 pixel_5164/gring pixel_5164/VDD pixel_5164/GND pixel_5164/VREF pixel_5164/ROW_SEL
+ pixel_5164/NB1 pixel_5164/VBIAS pixel_5164/NB2 pixel_5164/AMP_IN pixel_5164/SF_IB
+ pixel_5164/PIX_OUT pixel_5164/CSA_VREF pixel
Xpixel_4430 pixel_4430/gring pixel_4430/VDD pixel_4430/GND pixel_4430/VREF pixel_4430/ROW_SEL
+ pixel_4430/NB1 pixel_4430/VBIAS pixel_4430/NB2 pixel_4430/AMP_IN pixel_4430/SF_IB
+ pixel_4430/PIX_OUT pixel_4430/CSA_VREF pixel
Xpixel_5175 pixel_5175/gring pixel_5175/VDD pixel_5175/GND pixel_5175/VREF pixel_5175/ROW_SEL
+ pixel_5175/NB1 pixel_5175/VBIAS pixel_5175/NB2 pixel_5175/AMP_IN pixel_5175/SF_IB
+ pixel_5175/PIX_OUT pixel_5175/CSA_VREF pixel
Xpixel_5186 pixel_5186/gring pixel_5186/VDD pixel_5186/GND pixel_5186/VREF pixel_5186/ROW_SEL
+ pixel_5186/NB1 pixel_5186/VBIAS pixel_5186/NB2 pixel_5186/AMP_IN pixel_5186/SF_IB
+ pixel_5186/PIX_OUT pixel_5186/CSA_VREF pixel
Xpixel_5197 pixel_5197/gring pixel_5197/VDD pixel_5197/GND pixel_5197/VREF pixel_5197/ROW_SEL
+ pixel_5197/NB1 pixel_5197/VBIAS pixel_5197/NB2 pixel_5197/AMP_IN pixel_5197/SF_IB
+ pixel_5197/PIX_OUT pixel_5197/CSA_VREF pixel
Xpixel_4441 pixel_4441/gring pixel_4441/VDD pixel_4441/GND pixel_4441/VREF pixel_4441/ROW_SEL
+ pixel_4441/NB1 pixel_4441/VBIAS pixel_4441/NB2 pixel_4441/AMP_IN pixel_4441/SF_IB
+ pixel_4441/PIX_OUT pixel_4441/CSA_VREF pixel
Xpixel_4452 pixel_4452/gring pixel_4452/VDD pixel_4452/GND pixel_4452/VREF pixel_4452/ROW_SEL
+ pixel_4452/NB1 pixel_4452/VBIAS pixel_4452/NB2 pixel_4452/AMP_IN pixel_4452/SF_IB
+ pixel_4452/PIX_OUT pixel_4452/CSA_VREF pixel
Xpixel_4463 pixel_4463/gring pixel_4463/VDD pixel_4463/GND pixel_4463/VREF pixel_4463/ROW_SEL
+ pixel_4463/NB1 pixel_4463/VBIAS pixel_4463/NB2 pixel_4463/AMP_IN pixel_4463/SF_IB
+ pixel_4463/PIX_OUT pixel_4463/CSA_VREF pixel
Xpixel_491 pixel_491/gring pixel_491/VDD pixel_491/GND pixel_491/VREF pixel_491/ROW_SEL
+ pixel_491/NB1 pixel_491/VBIAS pixel_491/NB2 pixel_491/AMP_IN pixel_491/SF_IB pixel_491/PIX_OUT
+ pixel_491/CSA_VREF pixel
Xpixel_480 pixel_480/gring pixel_480/VDD pixel_480/GND pixel_480/VREF pixel_480/ROW_SEL
+ pixel_480/NB1 pixel_480/VBIAS pixel_480/NB2 pixel_480/AMP_IN pixel_480/SF_IB pixel_480/PIX_OUT
+ pixel_480/CSA_VREF pixel
Xpixel_3751 pixel_3751/gring pixel_3751/VDD pixel_3751/GND pixel_3751/VREF pixel_3751/ROW_SEL
+ pixel_3751/NB1 pixel_3751/VBIAS pixel_3751/NB2 pixel_3751/AMP_IN pixel_3751/SF_IB
+ pixel_3751/PIX_OUT pixel_3751/CSA_VREF pixel
Xpixel_3740 pixel_3740/gring pixel_3740/VDD pixel_3740/GND pixel_3740/VREF pixel_3740/ROW_SEL
+ pixel_3740/NB1 pixel_3740/VBIAS pixel_3740/NB2 pixel_3740/AMP_IN pixel_3740/SF_IB
+ pixel_3740/PIX_OUT pixel_3740/CSA_VREF pixel
Xpixel_4474 pixel_4474/gring pixel_4474/VDD pixel_4474/GND pixel_4474/VREF pixel_4474/ROW_SEL
+ pixel_4474/NB1 pixel_4474/VBIAS pixel_4474/NB2 pixel_4474/AMP_IN pixel_4474/SF_IB
+ pixel_4474/PIX_OUT pixel_4474/CSA_VREF pixel
Xpixel_4485 pixel_4485/gring pixel_4485/VDD pixel_4485/GND pixel_4485/VREF pixel_4485/ROW_SEL
+ pixel_4485/NB1 pixel_4485/VBIAS pixel_4485/NB2 pixel_4485/AMP_IN pixel_4485/SF_IB
+ pixel_4485/PIX_OUT pixel_4485/CSA_VREF pixel
Xpixel_4496 pixel_4496/gring pixel_4496/VDD pixel_4496/GND pixel_4496/VREF pixel_4496/ROW_SEL
+ pixel_4496/NB1 pixel_4496/VBIAS pixel_4496/NB2 pixel_4496/AMP_IN pixel_4496/SF_IB
+ pixel_4496/PIX_OUT pixel_4496/CSA_VREF pixel
Xpixel_3795 pixel_3795/gring pixel_3795/VDD pixel_3795/GND pixel_3795/VREF pixel_3795/ROW_SEL
+ pixel_3795/NB1 pixel_3795/VBIAS pixel_3795/NB2 pixel_3795/AMP_IN pixel_3795/SF_IB
+ pixel_3795/PIX_OUT pixel_3795/CSA_VREF pixel
Xpixel_3784 pixel_3784/gring pixel_3784/VDD pixel_3784/GND pixel_3784/VREF pixel_3784/ROW_SEL
+ pixel_3784/NB1 pixel_3784/VBIAS pixel_3784/NB2 pixel_3784/AMP_IN pixel_3784/SF_IB
+ pixel_3784/PIX_OUT pixel_3784/CSA_VREF pixel
Xpixel_3773 pixel_3773/gring pixel_3773/VDD pixel_3773/GND pixel_3773/VREF pixel_3773/ROW_SEL
+ pixel_3773/NB1 pixel_3773/VBIAS pixel_3773/NB2 pixel_3773/AMP_IN pixel_3773/SF_IB
+ pixel_3773/PIX_OUT pixel_3773/CSA_VREF pixel
Xpixel_3762 pixel_3762/gring pixel_3762/VDD pixel_3762/GND pixel_3762/VREF pixel_3762/ROW_SEL
+ pixel_3762/NB1 pixel_3762/VBIAS pixel_3762/NB2 pixel_3762/AMP_IN pixel_3762/SF_IB
+ pixel_3762/PIX_OUT pixel_3762/CSA_VREF pixel
Xpixel_9419 pixel_9419/gring pixel_9419/VDD pixel_9419/GND pixel_9419/VREF pixel_9419/ROW_SEL
+ pixel_9419/NB1 pixel_9419/VBIAS pixel_9419/NB2 pixel_9419/AMP_IN pixel_9419/SF_IB
+ pixel_9419/PIX_OUT pixel_9419/CSA_VREF pixel
Xpixel_9408 pixel_9408/gring pixel_9408/VDD pixel_9408/GND pixel_9408/VREF pixel_9408/ROW_SEL
+ pixel_9408/NB1 pixel_9408/VBIAS pixel_9408/NB2 pixel_9408/AMP_IN pixel_9408/SF_IB
+ pixel_9408/PIX_OUT pixel_9408/CSA_VREF pixel
Xpixel_8718 pixel_8718/gring pixel_8718/VDD pixel_8718/GND pixel_8718/VREF pixel_8718/ROW_SEL
+ pixel_8718/NB1 pixel_8718/VBIAS pixel_8718/NB2 pixel_8718/AMP_IN pixel_8718/SF_IB
+ pixel_8718/PIX_OUT pixel_8718/CSA_VREF pixel
Xpixel_8707 pixel_8707/gring pixel_8707/VDD pixel_8707/GND pixel_8707/VREF pixel_8707/ROW_SEL
+ pixel_8707/NB1 pixel_8707/VBIAS pixel_8707/NB2 pixel_8707/AMP_IN pixel_8707/SF_IB
+ pixel_8707/PIX_OUT pixel_8707/CSA_VREF pixel
Xpixel_8729 pixel_8729/gring pixel_8729/VDD pixel_8729/GND pixel_8729/VREF pixel_8729/ROW_SEL
+ pixel_8729/NB1 pixel_8729/VBIAS pixel_8729/NB2 pixel_8729/AMP_IN pixel_8729/SF_IB
+ pixel_8729/PIX_OUT pixel_8729/CSA_VREF pixel
Xpixel_3014 pixel_3014/gring pixel_3014/VDD pixel_3014/GND pixel_3014/VREF pixel_3014/ROW_SEL
+ pixel_3014/NB1 pixel_3014/VBIAS pixel_3014/NB2 pixel_3014/AMP_IN pixel_3014/SF_IB
+ pixel_3014/PIX_OUT pixel_3014/CSA_VREF pixel
Xpixel_3003 pixel_3003/gring pixel_3003/VDD pixel_3003/GND pixel_3003/VREF pixel_3003/ROW_SEL
+ pixel_3003/NB1 pixel_3003/VBIAS pixel_3003/NB2 pixel_3003/AMP_IN pixel_3003/SF_IB
+ pixel_3003/PIX_OUT pixel_3003/CSA_VREF pixel
Xpixel_2302 pixel_2302/gring pixel_2302/VDD pixel_2302/GND pixel_2302/VREF pixel_2302/ROW_SEL
+ pixel_2302/NB1 pixel_2302/VBIAS pixel_2302/NB2 pixel_2302/AMP_IN pixel_2302/SF_IB
+ pixel_2302/PIX_OUT pixel_2302/CSA_VREF pixel
Xpixel_3047 pixel_3047/gring pixel_3047/VDD pixel_3047/GND pixel_3047/VREF pixel_3047/ROW_SEL
+ pixel_3047/NB1 pixel_3047/VBIAS pixel_3047/NB2 pixel_3047/AMP_IN pixel_3047/SF_IB
+ pixel_3047/PIX_OUT pixel_3047/CSA_VREF pixel
Xpixel_3036 pixel_3036/gring pixel_3036/VDD pixel_3036/GND pixel_3036/VREF pixel_3036/ROW_SEL
+ pixel_3036/NB1 pixel_3036/VBIAS pixel_3036/NB2 pixel_3036/AMP_IN pixel_3036/SF_IB
+ pixel_3036/PIX_OUT pixel_3036/CSA_VREF pixel
Xpixel_3025 pixel_3025/gring pixel_3025/VDD pixel_3025/GND pixel_3025/VREF pixel_3025/ROW_SEL
+ pixel_3025/NB1 pixel_3025/VBIAS pixel_3025/NB2 pixel_3025/AMP_IN pixel_3025/SF_IB
+ pixel_3025/PIX_OUT pixel_3025/CSA_VREF pixel
Xpixel_1601 pixel_1601/gring pixel_1601/VDD pixel_1601/GND pixel_1601/VREF pixel_1601/ROW_SEL
+ pixel_1601/NB1 pixel_1601/VBIAS pixel_1601/NB2 pixel_1601/AMP_IN pixel_1601/SF_IB
+ pixel_1601/PIX_OUT pixel_1601/CSA_VREF pixel
Xpixel_2335 pixel_2335/gring pixel_2335/VDD pixel_2335/GND pixel_2335/VREF pixel_2335/ROW_SEL
+ pixel_2335/NB1 pixel_2335/VBIAS pixel_2335/NB2 pixel_2335/AMP_IN pixel_2335/SF_IB
+ pixel_2335/PIX_OUT pixel_2335/CSA_VREF pixel
Xpixel_2324 pixel_2324/gring pixel_2324/VDD pixel_2324/GND pixel_2324/VREF pixel_2324/ROW_SEL
+ pixel_2324/NB1 pixel_2324/VBIAS pixel_2324/NB2 pixel_2324/AMP_IN pixel_2324/SF_IB
+ pixel_2324/PIX_OUT pixel_2324/CSA_VREF pixel
Xpixel_2313 pixel_2313/gring pixel_2313/VDD pixel_2313/GND pixel_2313/VREF pixel_2313/ROW_SEL
+ pixel_2313/NB1 pixel_2313/VBIAS pixel_2313/NB2 pixel_2313/AMP_IN pixel_2313/SF_IB
+ pixel_2313/PIX_OUT pixel_2313/CSA_VREF pixel
Xpixel_3069 pixel_3069/gring pixel_3069/VDD pixel_3069/GND pixel_3069/VREF pixel_3069/ROW_SEL
+ pixel_3069/NB1 pixel_3069/VBIAS pixel_3069/NB2 pixel_3069/AMP_IN pixel_3069/SF_IB
+ pixel_3069/PIX_OUT pixel_3069/CSA_VREF pixel
Xpixel_3058 pixel_3058/gring pixel_3058/VDD pixel_3058/GND pixel_3058/VREF pixel_3058/ROW_SEL
+ pixel_3058/NB1 pixel_3058/VBIAS pixel_3058/NB2 pixel_3058/AMP_IN pixel_3058/SF_IB
+ pixel_3058/PIX_OUT pixel_3058/CSA_VREF pixel
Xpixel_1634 pixel_1634/gring pixel_1634/VDD pixel_1634/GND pixel_1634/VREF pixel_1634/ROW_SEL
+ pixel_1634/NB1 pixel_1634/VBIAS pixel_1634/NB2 pixel_1634/AMP_IN pixel_1634/SF_IB
+ pixel_1634/PIX_OUT pixel_1634/CSA_VREF pixel
Xpixel_1623 pixel_1623/gring pixel_1623/VDD pixel_1623/GND pixel_1623/VREF pixel_1623/ROW_SEL
+ pixel_1623/NB1 pixel_1623/VBIAS pixel_1623/NB2 pixel_1623/AMP_IN pixel_1623/SF_IB
+ pixel_1623/PIX_OUT pixel_1623/CSA_VREF pixel
Xpixel_1612 pixel_1612/gring pixel_1612/VDD pixel_1612/GND pixel_1612/VREF pixel_1612/ROW_SEL
+ pixel_1612/NB1 pixel_1612/VBIAS pixel_1612/NB2 pixel_1612/AMP_IN pixel_1612/SF_IB
+ pixel_1612/PIX_OUT pixel_1612/CSA_VREF pixel
Xpixel_2379 pixel_2379/gring pixel_2379/VDD pixel_2379/GND pixel_2379/VREF pixel_2379/ROW_SEL
+ pixel_2379/NB1 pixel_2379/VBIAS pixel_2379/NB2 pixel_2379/AMP_IN pixel_2379/SF_IB
+ pixel_2379/PIX_OUT pixel_2379/CSA_VREF pixel
Xpixel_2368 pixel_2368/gring pixel_2368/VDD pixel_2368/GND pixel_2368/VREF pixel_2368/ROW_SEL
+ pixel_2368/NB1 pixel_2368/VBIAS pixel_2368/NB2 pixel_2368/AMP_IN pixel_2368/SF_IB
+ pixel_2368/PIX_OUT pixel_2368/CSA_VREF pixel
Xpixel_2357 pixel_2357/gring pixel_2357/VDD pixel_2357/GND pixel_2357/VREF pixel_2357/ROW_SEL
+ pixel_2357/NB1 pixel_2357/VBIAS pixel_2357/NB2 pixel_2357/AMP_IN pixel_2357/SF_IB
+ pixel_2357/PIX_OUT pixel_2357/CSA_VREF pixel
Xpixel_2346 pixel_2346/gring pixel_2346/VDD pixel_2346/GND pixel_2346/VREF pixel_2346/ROW_SEL
+ pixel_2346/NB1 pixel_2346/VBIAS pixel_2346/NB2 pixel_2346/AMP_IN pixel_2346/SF_IB
+ pixel_2346/PIX_OUT pixel_2346/CSA_VREF pixel
Xpixel_1667 pixel_1667/gring pixel_1667/VDD pixel_1667/GND pixel_1667/VREF pixel_1667/ROW_SEL
+ pixel_1667/NB1 pixel_1667/VBIAS pixel_1667/NB2 pixel_1667/AMP_IN pixel_1667/SF_IB
+ pixel_1667/PIX_OUT pixel_1667/CSA_VREF pixel
Xpixel_1656 pixel_1656/gring pixel_1656/VDD pixel_1656/GND pixel_1656/VREF pixel_1656/ROW_SEL
+ pixel_1656/NB1 pixel_1656/VBIAS pixel_1656/NB2 pixel_1656/AMP_IN pixel_1656/SF_IB
+ pixel_1656/PIX_OUT pixel_1656/CSA_VREF pixel
Xpixel_1645 pixel_1645/gring pixel_1645/VDD pixel_1645/GND pixel_1645/VREF pixel_1645/ROW_SEL
+ pixel_1645/NB1 pixel_1645/VBIAS pixel_1645/NB2 pixel_1645/AMP_IN pixel_1645/SF_IB
+ pixel_1645/PIX_OUT pixel_1645/CSA_VREF pixel
Xpixel_1689 pixel_1689/gring pixel_1689/VDD pixel_1689/GND pixel_1689/VREF pixel_1689/ROW_SEL
+ pixel_1689/NB1 pixel_1689/VBIAS pixel_1689/NB2 pixel_1689/AMP_IN pixel_1689/SF_IB
+ pixel_1689/PIX_OUT pixel_1689/CSA_VREF pixel
Xpixel_1678 pixel_1678/gring pixel_1678/VDD pixel_1678/GND pixel_1678/VREF pixel_1678/ROW_SEL
+ pixel_1678/NB1 pixel_1678/VBIAS pixel_1678/NB2 pixel_1678/AMP_IN pixel_1678/SF_IB
+ pixel_1678/PIX_OUT pixel_1678/CSA_VREF pixel
Xpixel_9942 pixel_9942/gring pixel_9942/VDD pixel_9942/GND pixel_9942/VREF pixel_9942/ROW_SEL
+ pixel_9942/NB1 pixel_9942/VBIAS pixel_9942/NB2 pixel_9942/AMP_IN pixel_9942/SF_IB
+ pixel_9942/PIX_OUT pixel_9942/CSA_VREF pixel
Xpixel_9931 pixel_9931/gring pixel_9931/VDD pixel_9931/GND pixel_9931/VREF pixel_9931/ROW_SEL
+ pixel_9931/NB1 pixel_9931/VBIAS pixel_9931/NB2 pixel_9931/AMP_IN pixel_9931/SF_IB
+ pixel_9931/PIX_OUT pixel_9931/CSA_VREF pixel
Xpixel_9920 pixel_9920/gring pixel_9920/VDD pixel_9920/GND pixel_9920/VREF pixel_9920/ROW_SEL
+ pixel_9920/NB1 pixel_9920/VBIAS pixel_9920/NB2 pixel_9920/AMP_IN pixel_9920/SF_IB
+ pixel_9920/PIX_OUT pixel_9920/CSA_VREF pixel
Xpixel_9953 pixel_9953/gring pixel_9953/VDD pixel_9953/GND pixel_9953/VREF pixel_9953/ROW_SEL
+ pixel_9953/NB1 pixel_9953/VBIAS pixel_9953/NB2 pixel_9953/AMP_IN pixel_9953/SF_IB
+ pixel_9953/PIX_OUT pixel_9953/CSA_VREF pixel
Xpixel_9964 pixel_9964/gring pixel_9964/VDD pixel_9964/GND pixel_9964/VREF pixel_9964/ROW_SEL
+ pixel_9964/NB1 pixel_9964/VBIAS pixel_9964/NB2 pixel_9964/AMP_IN pixel_9964/SF_IB
+ pixel_9964/PIX_OUT pixel_9964/CSA_VREF pixel
Xpixel_9975 pixel_9975/gring pixel_9975/VDD pixel_9975/GND pixel_9975/VREF pixel_9975/ROW_SEL
+ pixel_9975/NB1 pixel_9975/VBIAS pixel_9975/NB2 pixel_9975/AMP_IN pixel_9975/SF_IB
+ pixel_9975/PIX_OUT pixel_9975/CSA_VREF pixel
Xpixel_9986 pixel_9986/gring pixel_9986/VDD pixel_9986/GND pixel_9986/VREF pixel_9986/ROW_SEL
+ pixel_9986/NB1 pixel_9986/VBIAS pixel_9986/NB2 pixel_9986/AMP_IN pixel_9986/SF_IB
+ pixel_9986/PIX_OUT pixel_9986/CSA_VREF pixel
Xpixel_9997 pixel_9997/gring pixel_9997/VDD pixel_9997/GND pixel_9997/VREF pixel_9997/ROW_SEL
+ pixel_9997/NB1 pixel_9997/VBIAS pixel_9997/NB2 pixel_9997/AMP_IN pixel_9997/SF_IB
+ pixel_9997/PIX_OUT pixel_9997/CSA_VREF pixel
Xpixel_4260 pixel_4260/gring pixel_4260/VDD pixel_4260/GND pixel_4260/VREF pixel_4260/ROW_SEL
+ pixel_4260/NB1 pixel_4260/VBIAS pixel_4260/NB2 pixel_4260/AMP_IN pixel_4260/SF_IB
+ pixel_4260/PIX_OUT pixel_4260/CSA_VREF pixel
Xpixel_4271 pixel_4271/gring pixel_4271/VDD pixel_4271/GND pixel_4271/VREF pixel_4271/ROW_SEL
+ pixel_4271/NB1 pixel_4271/VBIAS pixel_4271/NB2 pixel_4271/AMP_IN pixel_4271/SF_IB
+ pixel_4271/PIX_OUT pixel_4271/CSA_VREF pixel
Xpixel_3570 pixel_3570/gring pixel_3570/VDD pixel_3570/GND pixel_3570/VREF pixel_3570/ROW_SEL
+ pixel_3570/NB1 pixel_3570/VBIAS pixel_3570/NB2 pixel_3570/AMP_IN pixel_3570/SF_IB
+ pixel_3570/PIX_OUT pixel_3570/CSA_VREF pixel
Xpixel_4282 pixel_4282/gring pixel_4282/VDD pixel_4282/GND pixel_4282/VREF pixel_4282/ROW_SEL
+ pixel_4282/NB1 pixel_4282/VBIAS pixel_4282/NB2 pixel_4282/AMP_IN pixel_4282/SF_IB
+ pixel_4282/PIX_OUT pixel_4282/CSA_VREF pixel
Xpixel_4293 pixel_4293/gring pixel_4293/VDD pixel_4293/GND pixel_4293/VREF pixel_4293/ROW_SEL
+ pixel_4293/NB1 pixel_4293/VBIAS pixel_4293/NB2 pixel_4293/AMP_IN pixel_4293/SF_IB
+ pixel_4293/PIX_OUT pixel_4293/CSA_VREF pixel
Xpixel_3592 pixel_3592/gring pixel_3592/VDD pixel_3592/GND pixel_3592/VREF pixel_3592/ROW_SEL
+ pixel_3592/NB1 pixel_3592/VBIAS pixel_3592/NB2 pixel_3592/AMP_IN pixel_3592/SF_IB
+ pixel_3592/PIX_OUT pixel_3592/CSA_VREF pixel
Xpixel_3581 pixel_3581/gring pixel_3581/VDD pixel_3581/GND pixel_3581/VREF pixel_3581/ROW_SEL
+ pixel_3581/NB1 pixel_3581/VBIAS pixel_3581/NB2 pixel_3581/AMP_IN pixel_3581/SF_IB
+ pixel_3581/PIX_OUT pixel_3581/CSA_VREF pixel
Xpixel_2891 pixel_2891/gring pixel_2891/VDD pixel_2891/GND pixel_2891/VREF pixel_2891/ROW_SEL
+ pixel_2891/NB1 pixel_2891/VBIAS pixel_2891/NB2 pixel_2891/AMP_IN pixel_2891/SF_IB
+ pixel_2891/PIX_OUT pixel_2891/CSA_VREF pixel
Xpixel_2880 pixel_2880/gring pixel_2880/VDD pixel_2880/GND pixel_2880/VREF pixel_2880/ROW_SEL
+ pixel_2880/NB1 pixel_2880/VBIAS pixel_2880/NB2 pixel_2880/AMP_IN pixel_2880/SF_IB
+ pixel_2880/PIX_OUT pixel_2880/CSA_VREF pixel
Xpixel_9238 pixel_9238/gring pixel_9238/VDD pixel_9238/GND pixel_9238/VREF pixel_9238/ROW_SEL
+ pixel_9238/NB1 pixel_9238/VBIAS pixel_9238/NB2 pixel_9238/AMP_IN pixel_9238/SF_IB
+ pixel_9238/PIX_OUT pixel_9238/CSA_VREF pixel
Xpixel_9227 pixel_9227/gring pixel_9227/VDD pixel_9227/GND pixel_9227/VREF pixel_9227/ROW_SEL
+ pixel_9227/NB1 pixel_9227/VBIAS pixel_9227/NB2 pixel_9227/AMP_IN pixel_9227/SF_IB
+ pixel_9227/PIX_OUT pixel_9227/CSA_VREF pixel
Xpixel_9216 pixel_9216/gring pixel_9216/VDD pixel_9216/GND pixel_9216/VREF pixel_9216/ROW_SEL
+ pixel_9216/NB1 pixel_9216/VBIAS pixel_9216/NB2 pixel_9216/AMP_IN pixel_9216/SF_IB
+ pixel_9216/PIX_OUT pixel_9216/CSA_VREF pixel
Xpixel_9205 pixel_9205/gring pixel_9205/VDD pixel_9205/GND pixel_9205/VREF pixel_9205/ROW_SEL
+ pixel_9205/NB1 pixel_9205/VBIAS pixel_9205/NB2 pixel_9205/AMP_IN pixel_9205/SF_IB
+ pixel_9205/PIX_OUT pixel_9205/CSA_VREF pixel
Xpixel_8526 pixel_8526/gring pixel_8526/VDD pixel_8526/GND pixel_8526/VREF pixel_8526/ROW_SEL
+ pixel_8526/NB1 pixel_8526/VBIAS pixel_8526/NB2 pixel_8526/AMP_IN pixel_8526/SF_IB
+ pixel_8526/PIX_OUT pixel_8526/CSA_VREF pixel
Xpixel_8515 pixel_8515/gring pixel_8515/VDD pixel_8515/GND pixel_8515/VREF pixel_8515/ROW_SEL
+ pixel_8515/NB1 pixel_8515/VBIAS pixel_8515/NB2 pixel_8515/AMP_IN pixel_8515/SF_IB
+ pixel_8515/PIX_OUT pixel_8515/CSA_VREF pixel
Xpixel_8504 pixel_8504/gring pixel_8504/VDD pixel_8504/GND pixel_8504/VREF pixel_8504/ROW_SEL
+ pixel_8504/NB1 pixel_8504/VBIAS pixel_8504/NB2 pixel_8504/AMP_IN pixel_8504/SF_IB
+ pixel_8504/PIX_OUT pixel_8504/CSA_VREF pixel
Xpixel_9249 pixel_9249/gring pixel_9249/VDD pixel_9249/GND pixel_9249/VREF pixel_9249/ROW_SEL
+ pixel_9249/NB1 pixel_9249/VBIAS pixel_9249/NB2 pixel_9249/AMP_IN pixel_9249/SF_IB
+ pixel_9249/PIX_OUT pixel_9249/CSA_VREF pixel
Xpixel_8559 pixel_8559/gring pixel_8559/VDD pixel_8559/GND pixel_8559/VREF pixel_8559/ROW_SEL
+ pixel_8559/NB1 pixel_8559/VBIAS pixel_8559/NB2 pixel_8559/AMP_IN pixel_8559/SF_IB
+ pixel_8559/PIX_OUT pixel_8559/CSA_VREF pixel
Xpixel_8548 pixel_8548/gring pixel_8548/VDD pixel_8548/GND pixel_8548/VREF pixel_8548/ROW_SEL
+ pixel_8548/NB1 pixel_8548/VBIAS pixel_8548/NB2 pixel_8548/AMP_IN pixel_8548/SF_IB
+ pixel_8548/PIX_OUT pixel_8548/CSA_VREF pixel
Xpixel_8537 pixel_8537/gring pixel_8537/VDD pixel_8537/GND pixel_8537/VREF pixel_8537/ROW_SEL
+ pixel_8537/NB1 pixel_8537/VBIAS pixel_8537/NB2 pixel_8537/AMP_IN pixel_8537/SF_IB
+ pixel_8537/PIX_OUT pixel_8537/CSA_VREF pixel
Xpixel_7803 pixel_7803/gring pixel_7803/VDD pixel_7803/GND pixel_7803/VREF pixel_7803/ROW_SEL
+ pixel_7803/NB1 pixel_7803/VBIAS pixel_7803/NB2 pixel_7803/AMP_IN pixel_7803/SF_IB
+ pixel_7803/PIX_OUT pixel_7803/CSA_VREF pixel
Xpixel_7814 pixel_7814/gring pixel_7814/VDD pixel_7814/GND pixel_7814/VREF pixel_7814/ROW_SEL
+ pixel_7814/NB1 pixel_7814/VBIAS pixel_7814/NB2 pixel_7814/AMP_IN pixel_7814/SF_IB
+ pixel_7814/PIX_OUT pixel_7814/CSA_VREF pixel
Xpixel_7825 pixel_7825/gring pixel_7825/VDD pixel_7825/GND pixel_7825/VREF pixel_7825/ROW_SEL
+ pixel_7825/NB1 pixel_7825/VBIAS pixel_7825/NB2 pixel_7825/AMP_IN pixel_7825/SF_IB
+ pixel_7825/PIX_OUT pixel_7825/CSA_VREF pixel
Xpixel_7836 pixel_7836/gring pixel_7836/VDD pixel_7836/GND pixel_7836/VREF pixel_7836/ROW_SEL
+ pixel_7836/NB1 pixel_7836/VBIAS pixel_7836/NB2 pixel_7836/AMP_IN pixel_7836/SF_IB
+ pixel_7836/PIX_OUT pixel_7836/CSA_VREF pixel
Xpixel_7847 pixel_7847/gring pixel_7847/VDD pixel_7847/GND pixel_7847/VREF pixel_7847/ROW_SEL
+ pixel_7847/NB1 pixel_7847/VBIAS pixel_7847/NB2 pixel_7847/AMP_IN pixel_7847/SF_IB
+ pixel_7847/PIX_OUT pixel_7847/CSA_VREF pixel
Xpixel_7858 pixel_7858/gring pixel_7858/VDD pixel_7858/GND pixel_7858/VREF pixel_7858/ROW_SEL
+ pixel_7858/NB1 pixel_7858/VBIAS pixel_7858/NB2 pixel_7858/AMP_IN pixel_7858/SF_IB
+ pixel_7858/PIX_OUT pixel_7858/CSA_VREF pixel
Xpixel_7869 pixel_7869/gring pixel_7869/VDD pixel_7869/GND pixel_7869/VREF pixel_7869/ROW_SEL
+ pixel_7869/NB1 pixel_7869/VBIAS pixel_7869/NB2 pixel_7869/AMP_IN pixel_7869/SF_IB
+ pixel_7869/PIX_OUT pixel_7869/CSA_VREF pixel
Xpixel_2110 pixel_2110/gring pixel_2110/VDD pixel_2110/GND pixel_2110/VREF pixel_2110/ROW_SEL
+ pixel_2110/NB1 pixel_2110/VBIAS pixel_2110/NB2 pixel_2110/AMP_IN pixel_2110/SF_IB
+ pixel_2110/PIX_OUT pixel_2110/CSA_VREF pixel
Xpixel_2154 pixel_2154/gring pixel_2154/VDD pixel_2154/GND pixel_2154/VREF pixel_2154/ROW_SEL
+ pixel_2154/NB1 pixel_2154/VBIAS pixel_2154/NB2 pixel_2154/AMP_IN pixel_2154/SF_IB
+ pixel_2154/PIX_OUT pixel_2154/CSA_VREF pixel
Xpixel_2143 pixel_2143/gring pixel_2143/VDD pixel_2143/GND pixel_2143/VREF pixel_2143/ROW_SEL
+ pixel_2143/NB1 pixel_2143/VBIAS pixel_2143/NB2 pixel_2143/AMP_IN pixel_2143/SF_IB
+ pixel_2143/PIX_OUT pixel_2143/CSA_VREF pixel
Xpixel_2132 pixel_2132/gring pixel_2132/VDD pixel_2132/GND pixel_2132/VREF pixel_2132/ROW_SEL
+ pixel_2132/NB1 pixel_2132/VBIAS pixel_2132/NB2 pixel_2132/AMP_IN pixel_2132/SF_IB
+ pixel_2132/PIX_OUT pixel_2132/CSA_VREF pixel
Xpixel_2121 pixel_2121/gring pixel_2121/VDD pixel_2121/GND pixel_2121/VREF pixel_2121/ROW_SEL
+ pixel_2121/NB1 pixel_2121/VBIAS pixel_2121/NB2 pixel_2121/AMP_IN pixel_2121/SF_IB
+ pixel_2121/PIX_OUT pixel_2121/CSA_VREF pixel
Xpixel_1442 pixel_1442/gring pixel_1442/VDD pixel_1442/GND pixel_1442/VREF pixel_1442/ROW_SEL
+ pixel_1442/NB1 pixel_1442/VBIAS pixel_1442/NB2 pixel_1442/AMP_IN pixel_1442/SF_IB
+ pixel_1442/PIX_OUT pixel_1442/CSA_VREF pixel
Xpixel_1431 pixel_1431/gring pixel_1431/VDD pixel_1431/GND pixel_1431/VREF pixel_1431/ROW_SEL
+ pixel_1431/NB1 pixel_1431/VBIAS pixel_1431/NB2 pixel_1431/AMP_IN pixel_1431/SF_IB
+ pixel_1431/PIX_OUT pixel_1431/CSA_VREF pixel
Xpixel_1420 pixel_1420/gring pixel_1420/VDD pixel_1420/GND pixel_1420/VREF pixel_1420/ROW_SEL
+ pixel_1420/NB1 pixel_1420/VBIAS pixel_1420/NB2 pixel_1420/AMP_IN pixel_1420/SF_IB
+ pixel_1420/PIX_OUT pixel_1420/CSA_VREF pixel
Xpixel_2187 pixel_2187/gring pixel_2187/VDD pixel_2187/GND pixel_2187/VREF pixel_2187/ROW_SEL
+ pixel_2187/NB1 pixel_2187/VBIAS pixel_2187/NB2 pixel_2187/AMP_IN pixel_2187/SF_IB
+ pixel_2187/PIX_OUT pixel_2187/CSA_VREF pixel
Xpixel_2176 pixel_2176/gring pixel_2176/VDD pixel_2176/GND pixel_2176/VREF pixel_2176/ROW_SEL
+ pixel_2176/NB1 pixel_2176/VBIAS pixel_2176/NB2 pixel_2176/AMP_IN pixel_2176/SF_IB
+ pixel_2176/PIX_OUT pixel_2176/CSA_VREF pixel
Xpixel_2165 pixel_2165/gring pixel_2165/VDD pixel_2165/GND pixel_2165/VREF pixel_2165/ROW_SEL
+ pixel_2165/NB1 pixel_2165/VBIAS pixel_2165/NB2 pixel_2165/AMP_IN pixel_2165/SF_IB
+ pixel_2165/PIX_OUT pixel_2165/CSA_VREF pixel
Xpixel_1475 pixel_1475/gring pixel_1475/VDD pixel_1475/GND pixel_1475/VREF pixel_1475/ROW_SEL
+ pixel_1475/NB1 pixel_1475/VBIAS pixel_1475/NB2 pixel_1475/AMP_IN pixel_1475/SF_IB
+ pixel_1475/PIX_OUT pixel_1475/CSA_VREF pixel
Xpixel_1464 pixel_1464/gring pixel_1464/VDD pixel_1464/GND pixel_1464/VREF pixel_1464/ROW_SEL
+ pixel_1464/NB1 pixel_1464/VBIAS pixel_1464/NB2 pixel_1464/AMP_IN pixel_1464/SF_IB
+ pixel_1464/PIX_OUT pixel_1464/CSA_VREF pixel
Xpixel_1453 pixel_1453/gring pixel_1453/VDD pixel_1453/GND pixel_1453/VREF pixel_1453/ROW_SEL
+ pixel_1453/NB1 pixel_1453/VBIAS pixel_1453/NB2 pixel_1453/AMP_IN pixel_1453/SF_IB
+ pixel_1453/PIX_OUT pixel_1453/CSA_VREF pixel
Xpixel_2198 pixel_2198/gring pixel_2198/VDD pixel_2198/GND pixel_2198/VREF pixel_2198/ROW_SEL
+ pixel_2198/NB1 pixel_2198/VBIAS pixel_2198/NB2 pixel_2198/AMP_IN pixel_2198/SF_IB
+ pixel_2198/PIX_OUT pixel_2198/CSA_VREF pixel
Xpixel_1497 pixel_1497/gring pixel_1497/VDD pixel_1497/GND pixel_1497/VREF pixel_1497/ROW_SEL
+ pixel_1497/NB1 pixel_1497/VBIAS pixel_1497/NB2 pixel_1497/AMP_IN pixel_1497/SF_IB
+ pixel_1497/PIX_OUT pixel_1497/CSA_VREF pixel
Xpixel_1486 pixel_1486/gring pixel_1486/VDD pixel_1486/GND pixel_1486/VREF pixel_1486/ROW_SEL
+ pixel_1486/NB1 pixel_1486/VBIAS pixel_1486/NB2 pixel_1486/AMP_IN pixel_1486/SF_IB
+ pixel_1486/PIX_OUT pixel_1486/CSA_VREF pixel
Xpixel_9750 pixel_9750/gring pixel_9750/VDD pixel_9750/GND pixel_9750/VREF pixel_9750/ROW_SEL
+ pixel_9750/NB1 pixel_9750/VBIAS pixel_9750/NB2 pixel_9750/AMP_IN pixel_9750/SF_IB
+ pixel_9750/PIX_OUT pixel_9750/CSA_VREF pixel
Xpixel_9761 pixel_9761/gring pixel_9761/VDD pixel_9761/GND pixel_9761/VREF pixel_9761/ROW_SEL
+ pixel_9761/NB1 pixel_9761/VBIAS pixel_9761/NB2 pixel_9761/AMP_IN pixel_9761/SF_IB
+ pixel_9761/PIX_OUT pixel_9761/CSA_VREF pixel
Xpixel_9772 pixel_9772/gring pixel_9772/VDD pixel_9772/GND pixel_9772/VREF pixel_9772/ROW_SEL
+ pixel_9772/NB1 pixel_9772/VBIAS pixel_9772/NB2 pixel_9772/AMP_IN pixel_9772/SF_IB
+ pixel_9772/PIX_OUT pixel_9772/CSA_VREF pixel
Xpixel_9783 pixel_9783/gring pixel_9783/VDD pixel_9783/GND pixel_9783/VREF pixel_9783/ROW_SEL
+ pixel_9783/NB1 pixel_9783/VBIAS pixel_9783/NB2 pixel_9783/AMP_IN pixel_9783/SF_IB
+ pixel_9783/PIX_OUT pixel_9783/CSA_VREF pixel
Xpixel_9794 pixel_9794/gring pixel_9794/VDD pixel_9794/GND pixel_9794/VREF pixel_9794/ROW_SEL
+ pixel_9794/NB1 pixel_9794/VBIAS pixel_9794/NB2 pixel_9794/AMP_IN pixel_9794/SF_IB
+ pixel_9794/PIX_OUT pixel_9794/CSA_VREF pixel
Xpixel_4090 pixel_4090/gring pixel_4090/VDD pixel_4090/GND pixel_4090/VREF pixel_4090/ROW_SEL
+ pixel_4090/NB1 pixel_4090/VBIAS pixel_4090/NB2 pixel_4090/AMP_IN pixel_4090/SF_IB
+ pixel_4090/PIX_OUT pixel_4090/CSA_VREF pixel
Xpixel_6409 pixel_6409/gring pixel_6409/VDD pixel_6409/GND pixel_6409/VREF pixel_6409/ROW_SEL
+ pixel_6409/NB1 pixel_6409/VBIAS pixel_6409/NB2 pixel_6409/AMP_IN pixel_6409/SF_IB
+ pixel_6409/PIX_OUT pixel_6409/CSA_VREF pixel
Xpixel_5708 pixel_5708/gring pixel_5708/VDD pixel_5708/GND pixel_5708/VREF pixel_5708/ROW_SEL
+ pixel_5708/NB1 pixel_5708/VBIAS pixel_5708/NB2 pixel_5708/AMP_IN pixel_5708/SF_IB
+ pixel_5708/PIX_OUT pixel_5708/CSA_VREF pixel
Xpixel_5719 pixel_5719/gring pixel_5719/VDD pixel_5719/GND pixel_5719/VREF pixel_5719/ROW_SEL
+ pixel_5719/NB1 pixel_5719/VBIAS pixel_5719/NB2 pixel_5719/AMP_IN pixel_5719/SF_IB
+ pixel_5719/PIX_OUT pixel_5719/CSA_VREF pixel
Xpixel_9013 pixel_9013/gring pixel_9013/VDD pixel_9013/GND pixel_9013/VREF pixel_9013/ROW_SEL
+ pixel_9013/NB1 pixel_9013/VBIAS pixel_9013/NB2 pixel_9013/AMP_IN pixel_9013/SF_IB
+ pixel_9013/PIX_OUT pixel_9013/CSA_VREF pixel
Xpixel_9002 pixel_9002/gring pixel_9002/VDD pixel_9002/GND pixel_9002/VREF pixel_9002/ROW_SEL
+ pixel_9002/NB1 pixel_9002/VBIAS pixel_9002/NB2 pixel_9002/AMP_IN pixel_9002/SF_IB
+ pixel_9002/PIX_OUT pixel_9002/CSA_VREF pixel
Xpixel_9046 pixel_9046/gring pixel_9046/VDD pixel_9046/GND pixel_9046/VREF pixel_9046/ROW_SEL
+ pixel_9046/NB1 pixel_9046/VBIAS pixel_9046/NB2 pixel_9046/AMP_IN pixel_9046/SF_IB
+ pixel_9046/PIX_OUT pixel_9046/CSA_VREF pixel
Xpixel_9035 pixel_9035/gring pixel_9035/VDD pixel_9035/GND pixel_9035/VREF pixel_9035/ROW_SEL
+ pixel_9035/NB1 pixel_9035/VBIAS pixel_9035/NB2 pixel_9035/AMP_IN pixel_9035/SF_IB
+ pixel_9035/PIX_OUT pixel_9035/CSA_VREF pixel
Xpixel_9024 pixel_9024/gring pixel_9024/VDD pixel_9024/GND pixel_9024/VREF pixel_9024/ROW_SEL
+ pixel_9024/NB1 pixel_9024/VBIAS pixel_9024/NB2 pixel_9024/AMP_IN pixel_9024/SF_IB
+ pixel_9024/PIX_OUT pixel_9024/CSA_VREF pixel
Xpixel_8301 pixel_8301/gring pixel_8301/VDD pixel_8301/GND pixel_8301/VREF pixel_8301/ROW_SEL
+ pixel_8301/NB1 pixel_8301/VBIAS pixel_8301/NB2 pixel_8301/AMP_IN pixel_8301/SF_IB
+ pixel_8301/PIX_OUT pixel_8301/CSA_VREF pixel
Xpixel_9079 pixel_9079/gring pixel_9079/VDD pixel_9079/GND pixel_9079/VREF pixel_9079/ROW_SEL
+ pixel_9079/NB1 pixel_9079/VBIAS pixel_9079/NB2 pixel_9079/AMP_IN pixel_9079/SF_IB
+ pixel_9079/PIX_OUT pixel_9079/CSA_VREF pixel
Xpixel_9068 pixel_9068/gring pixel_9068/VDD pixel_9068/GND pixel_9068/VREF pixel_9068/ROW_SEL
+ pixel_9068/NB1 pixel_9068/VBIAS pixel_9068/NB2 pixel_9068/AMP_IN pixel_9068/SF_IB
+ pixel_9068/PIX_OUT pixel_9068/CSA_VREF pixel
Xpixel_9057 pixel_9057/gring pixel_9057/VDD pixel_9057/GND pixel_9057/VREF pixel_9057/ROW_SEL
+ pixel_9057/NB1 pixel_9057/VBIAS pixel_9057/NB2 pixel_9057/AMP_IN pixel_9057/SF_IB
+ pixel_9057/PIX_OUT pixel_9057/CSA_VREF pixel
Xpixel_8312 pixel_8312/gring pixel_8312/VDD pixel_8312/GND pixel_8312/VREF pixel_8312/ROW_SEL
+ pixel_8312/NB1 pixel_8312/VBIAS pixel_8312/NB2 pixel_8312/AMP_IN pixel_8312/SF_IB
+ pixel_8312/PIX_OUT pixel_8312/CSA_VREF pixel
Xpixel_8323 pixel_8323/gring pixel_8323/VDD pixel_8323/GND pixel_8323/VREF pixel_8323/ROW_SEL
+ pixel_8323/NB1 pixel_8323/VBIAS pixel_8323/NB2 pixel_8323/AMP_IN pixel_8323/SF_IB
+ pixel_8323/PIX_OUT pixel_8323/CSA_VREF pixel
Xpixel_8334 pixel_8334/gring pixel_8334/VDD pixel_8334/GND pixel_8334/VREF pixel_8334/ROW_SEL
+ pixel_8334/NB1 pixel_8334/VBIAS pixel_8334/NB2 pixel_8334/AMP_IN pixel_8334/SF_IB
+ pixel_8334/PIX_OUT pixel_8334/CSA_VREF pixel
Xpixel_8345 pixel_8345/gring pixel_8345/VDD pixel_8345/GND pixel_8345/VREF pixel_8345/ROW_SEL
+ pixel_8345/NB1 pixel_8345/VBIAS pixel_8345/NB2 pixel_8345/AMP_IN pixel_8345/SF_IB
+ pixel_8345/PIX_OUT pixel_8345/CSA_VREF pixel
Xpixel_8356 pixel_8356/gring pixel_8356/VDD pixel_8356/GND pixel_8356/VREF pixel_8356/ROW_SEL
+ pixel_8356/NB1 pixel_8356/VBIAS pixel_8356/NB2 pixel_8356/AMP_IN pixel_8356/SF_IB
+ pixel_8356/PIX_OUT pixel_8356/CSA_VREF pixel
Xpixel_8367 pixel_8367/gring pixel_8367/VDD pixel_8367/GND pixel_8367/VREF pixel_8367/ROW_SEL
+ pixel_8367/NB1 pixel_8367/VBIAS pixel_8367/NB2 pixel_8367/AMP_IN pixel_8367/SF_IB
+ pixel_8367/PIX_OUT pixel_8367/CSA_VREF pixel
Xpixel_8378 pixel_8378/gring pixel_8378/VDD pixel_8378/GND pixel_8378/VREF pixel_8378/ROW_SEL
+ pixel_8378/NB1 pixel_8378/VBIAS pixel_8378/NB2 pixel_8378/AMP_IN pixel_8378/SF_IB
+ pixel_8378/PIX_OUT pixel_8378/CSA_VREF pixel
Xpixel_7600 pixel_7600/gring pixel_7600/VDD pixel_7600/GND pixel_7600/VREF pixel_7600/ROW_SEL
+ pixel_7600/NB1 pixel_7600/VBIAS pixel_7600/NB2 pixel_7600/AMP_IN pixel_7600/SF_IB
+ pixel_7600/PIX_OUT pixel_7600/CSA_VREF pixel
Xpixel_7611 pixel_7611/gring pixel_7611/VDD pixel_7611/GND pixel_7611/VREF pixel_7611/ROW_SEL
+ pixel_7611/NB1 pixel_7611/VBIAS pixel_7611/NB2 pixel_7611/AMP_IN pixel_7611/SF_IB
+ pixel_7611/PIX_OUT pixel_7611/CSA_VREF pixel
Xpixel_7622 pixel_7622/gring pixel_7622/VDD pixel_7622/GND pixel_7622/VREF pixel_7622/ROW_SEL
+ pixel_7622/NB1 pixel_7622/VBIAS pixel_7622/NB2 pixel_7622/AMP_IN pixel_7622/SF_IB
+ pixel_7622/PIX_OUT pixel_7622/CSA_VREF pixel
Xpixel_7633 pixel_7633/gring pixel_7633/VDD pixel_7633/GND pixel_7633/VREF pixel_7633/ROW_SEL
+ pixel_7633/NB1 pixel_7633/VBIAS pixel_7633/NB2 pixel_7633/AMP_IN pixel_7633/SF_IB
+ pixel_7633/PIX_OUT pixel_7633/CSA_VREF pixel
Xpixel_8389 pixel_8389/gring pixel_8389/VDD pixel_8389/GND pixel_8389/VREF pixel_8389/ROW_SEL
+ pixel_8389/NB1 pixel_8389/VBIAS pixel_8389/NB2 pixel_8389/AMP_IN pixel_8389/SF_IB
+ pixel_8389/PIX_OUT pixel_8389/CSA_VREF pixel
Xpixel_7644 pixel_7644/gring pixel_7644/VDD pixel_7644/GND pixel_7644/VREF pixel_7644/ROW_SEL
+ pixel_7644/NB1 pixel_7644/VBIAS pixel_7644/NB2 pixel_7644/AMP_IN pixel_7644/SF_IB
+ pixel_7644/PIX_OUT pixel_7644/CSA_VREF pixel
Xpixel_7655 pixel_7655/gring pixel_7655/VDD pixel_7655/GND pixel_7655/VREF pixel_7655/ROW_SEL
+ pixel_7655/NB1 pixel_7655/VBIAS pixel_7655/NB2 pixel_7655/AMP_IN pixel_7655/SF_IB
+ pixel_7655/PIX_OUT pixel_7655/CSA_VREF pixel
Xpixel_7666 pixel_7666/gring pixel_7666/VDD pixel_7666/GND pixel_7666/VREF pixel_7666/ROW_SEL
+ pixel_7666/NB1 pixel_7666/VBIAS pixel_7666/NB2 pixel_7666/AMP_IN pixel_7666/SF_IB
+ pixel_7666/PIX_OUT pixel_7666/CSA_VREF pixel
Xpixel_6910 pixel_6910/gring pixel_6910/VDD pixel_6910/GND pixel_6910/VREF pixel_6910/ROW_SEL
+ pixel_6910/NB1 pixel_6910/VBIAS pixel_6910/NB2 pixel_6910/AMP_IN pixel_6910/SF_IB
+ pixel_6910/PIX_OUT pixel_6910/CSA_VREF pixel
Xpixel_6921 pixel_6921/gring pixel_6921/VDD pixel_6921/GND pixel_6921/VREF pixel_6921/ROW_SEL
+ pixel_6921/NB1 pixel_6921/VBIAS pixel_6921/NB2 pixel_6921/AMP_IN pixel_6921/SF_IB
+ pixel_6921/PIX_OUT pixel_6921/CSA_VREF pixel
Xpixel_7677 pixel_7677/gring pixel_7677/VDD pixel_7677/GND pixel_7677/VREF pixel_7677/ROW_SEL
+ pixel_7677/NB1 pixel_7677/VBIAS pixel_7677/NB2 pixel_7677/AMP_IN pixel_7677/SF_IB
+ pixel_7677/PIX_OUT pixel_7677/CSA_VREF pixel
Xpixel_7688 pixel_7688/gring pixel_7688/VDD pixel_7688/GND pixel_7688/VREF pixel_7688/ROW_SEL
+ pixel_7688/NB1 pixel_7688/VBIAS pixel_7688/NB2 pixel_7688/AMP_IN pixel_7688/SF_IB
+ pixel_7688/PIX_OUT pixel_7688/CSA_VREF pixel
Xpixel_7699 pixel_7699/gring pixel_7699/VDD pixel_7699/GND pixel_7699/VREF pixel_7699/ROW_SEL
+ pixel_7699/NB1 pixel_7699/VBIAS pixel_7699/NB2 pixel_7699/AMP_IN pixel_7699/SF_IB
+ pixel_7699/PIX_OUT pixel_7699/CSA_VREF pixel
Xpixel_6932 pixel_6932/gring pixel_6932/VDD pixel_6932/GND pixel_6932/VREF pixel_6932/ROW_SEL
+ pixel_6932/NB1 pixel_6932/VBIAS pixel_6932/NB2 pixel_6932/AMP_IN pixel_6932/SF_IB
+ pixel_6932/PIX_OUT pixel_6932/CSA_VREF pixel
Xpixel_6943 pixel_6943/gring pixel_6943/VDD pixel_6943/GND pixel_6943/VREF pixel_6943/ROW_SEL
+ pixel_6943/NB1 pixel_6943/VBIAS pixel_6943/NB2 pixel_6943/AMP_IN pixel_6943/SF_IB
+ pixel_6943/PIX_OUT pixel_6943/CSA_VREF pixel
Xpixel_6954 pixel_6954/gring pixel_6954/VDD pixel_6954/GND pixel_6954/VREF pixel_6954/ROW_SEL
+ pixel_6954/NB1 pixel_6954/VBIAS pixel_6954/NB2 pixel_6954/AMP_IN pixel_6954/SF_IB
+ pixel_6954/PIX_OUT pixel_6954/CSA_VREF pixel
Xpixel_46 pixel_46/gring pixel_46/VDD pixel_46/GND pixel_46/VREF pixel_46/ROW_SEL
+ pixel_46/NB1 pixel_46/VBIAS pixel_46/NB2 pixel_46/AMP_IN pixel_46/SF_IB pixel_46/PIX_OUT
+ pixel_46/CSA_VREF pixel
Xpixel_35 pixel_35/gring pixel_35/VDD pixel_35/GND pixel_35/VREF pixel_35/ROW_SEL
+ pixel_35/NB1 pixel_35/VBIAS pixel_35/NB2 pixel_35/AMP_IN pixel_35/SF_IB pixel_35/PIX_OUT
+ pixel_35/CSA_VREF pixel
Xpixel_24 pixel_24/gring pixel_24/VDD pixel_24/GND pixel_24/VREF pixel_24/ROW_SEL
+ pixel_24/NB1 pixel_24/VBIAS pixel_24/NB2 pixel_24/AMP_IN pixel_24/SF_IB pixel_24/PIX_OUT
+ pixel_24/CSA_VREF pixel
Xpixel_13 pixel_13/gring pixel_13/VDD pixel_13/GND pixel_13/VREF pixel_13/ROW_SEL
+ pixel_13/NB1 pixel_13/VBIAS pixel_13/NB2 pixel_13/AMP_IN pixel_13/SF_IB pixel_13/PIX_OUT
+ pixel_13/CSA_VREF pixel
Xpixel_6965 pixel_6965/gring pixel_6965/VDD pixel_6965/GND pixel_6965/VREF pixel_6965/ROW_SEL
+ pixel_6965/NB1 pixel_6965/VBIAS pixel_6965/NB2 pixel_6965/AMP_IN pixel_6965/SF_IB
+ pixel_6965/PIX_OUT pixel_6965/CSA_VREF pixel
Xpixel_6976 pixel_6976/gring pixel_6976/VDD pixel_6976/GND pixel_6976/VREF pixel_6976/ROW_SEL
+ pixel_6976/NB1 pixel_6976/VBIAS pixel_6976/NB2 pixel_6976/AMP_IN pixel_6976/SF_IB
+ pixel_6976/PIX_OUT pixel_6976/CSA_VREF pixel
Xpixel_6987 pixel_6987/gring pixel_6987/VDD pixel_6987/GND pixel_6987/VREF pixel_6987/ROW_SEL
+ pixel_6987/NB1 pixel_6987/VBIAS pixel_6987/NB2 pixel_6987/AMP_IN pixel_6987/SF_IB
+ pixel_6987/PIX_OUT pixel_6987/CSA_VREF pixel
Xpixel_6998 pixel_6998/gring pixel_6998/VDD pixel_6998/GND pixel_6998/VREF pixel_6998/ROW_SEL
+ pixel_6998/NB1 pixel_6998/VBIAS pixel_6998/NB2 pixel_6998/AMP_IN pixel_6998/SF_IB
+ pixel_6998/PIX_OUT pixel_6998/CSA_VREF pixel
Xpixel_79 pixel_79/gring pixel_79/VDD pixel_79/GND pixel_79/VREF pixel_79/ROW_SEL
+ pixel_79/NB1 pixel_79/VBIAS pixel_79/NB2 pixel_79/AMP_IN pixel_79/SF_IB pixel_79/PIX_OUT
+ pixel_79/CSA_VREF pixel
Xpixel_68 pixel_68/gring pixel_68/VDD pixel_68/GND pixel_68/VREF pixel_68/ROW_SEL
+ pixel_68/NB1 pixel_68/VBIAS pixel_68/NB2 pixel_68/AMP_IN pixel_68/SF_IB pixel_68/PIX_OUT
+ pixel_68/CSA_VREF pixel
Xpixel_57 pixel_57/gring pixel_57/VDD pixel_57/GND pixel_57/VREF pixel_57/ROW_SEL
+ pixel_57/NB1 pixel_57/VBIAS pixel_57/NB2 pixel_57/AMP_IN pixel_57/SF_IB pixel_57/PIX_OUT
+ pixel_57/CSA_VREF pixel
Xpixel_1250 pixel_1250/gring pixel_1250/VDD pixel_1250/GND pixel_1250/VREF pixel_1250/ROW_SEL
+ pixel_1250/NB1 pixel_1250/VBIAS pixel_1250/NB2 pixel_1250/AMP_IN pixel_1250/SF_IB
+ pixel_1250/PIX_OUT pixel_1250/CSA_VREF pixel
Xpixel_1294 pixel_1294/gring pixel_1294/VDD pixel_1294/GND pixel_1294/VREF pixel_1294/ROW_SEL
+ pixel_1294/NB1 pixel_1294/VBIAS pixel_1294/NB2 pixel_1294/AMP_IN pixel_1294/SF_IB
+ pixel_1294/PIX_OUT pixel_1294/CSA_VREF pixel
Xpixel_1283 pixel_1283/gring pixel_1283/VDD pixel_1283/GND pixel_1283/VREF pixel_1283/ROW_SEL
+ pixel_1283/NB1 pixel_1283/VBIAS pixel_1283/NB2 pixel_1283/AMP_IN pixel_1283/SF_IB
+ pixel_1283/PIX_OUT pixel_1283/CSA_VREF pixel
Xpixel_1272 pixel_1272/gring pixel_1272/VDD pixel_1272/GND pixel_1272/VREF pixel_1272/ROW_SEL
+ pixel_1272/NB1 pixel_1272/VBIAS pixel_1272/NB2 pixel_1272/AMP_IN pixel_1272/SF_IB
+ pixel_1272/PIX_OUT pixel_1272/CSA_VREF pixel
Xpixel_1261 pixel_1261/gring pixel_1261/VDD pixel_1261/GND pixel_1261/VREF pixel_1261/ROW_SEL
+ pixel_1261/NB1 pixel_1261/VBIAS pixel_1261/NB2 pixel_1261/AMP_IN pixel_1261/SF_IB
+ pixel_1261/PIX_OUT pixel_1261/CSA_VREF pixel
Xpixel_9591 pixel_9591/gring pixel_9591/VDD pixel_9591/GND pixel_9591/VREF pixel_9591/ROW_SEL
+ pixel_9591/NB1 pixel_9591/VBIAS pixel_9591/NB2 pixel_9591/AMP_IN pixel_9591/SF_IB
+ pixel_9591/PIX_OUT pixel_9591/CSA_VREF pixel
Xpixel_9580 pixel_9580/gring pixel_9580/VDD pixel_9580/GND pixel_9580/VREF pixel_9580/ROW_SEL
+ pixel_9580/NB1 pixel_9580/VBIAS pixel_9580/NB2 pixel_9580/AMP_IN pixel_9580/SF_IB
+ pixel_9580/PIX_OUT pixel_9580/CSA_VREF pixel
Xpixel_8890 pixel_8890/gring pixel_8890/VDD pixel_8890/GND pixel_8890/VREF pixel_8890/ROW_SEL
+ pixel_8890/NB1 pixel_8890/VBIAS pixel_8890/NB2 pixel_8890/AMP_IN pixel_8890/SF_IB
+ pixel_8890/PIX_OUT pixel_8890/CSA_VREF pixel
Xpixel_309 pixel_309/gring pixel_309/VDD pixel_309/GND pixel_309/VREF pixel_309/ROW_SEL
+ pixel_309/NB1 pixel_309/VBIAS pixel_309/NB2 pixel_309/AMP_IN pixel_309/SF_IB pixel_309/PIX_OUT
+ pixel_309/CSA_VREF pixel
Xpixel_6206 pixel_6206/gring pixel_6206/VDD pixel_6206/GND pixel_6206/VREF pixel_6206/ROW_SEL
+ pixel_6206/NB1 pixel_6206/VBIAS pixel_6206/NB2 pixel_6206/AMP_IN pixel_6206/SF_IB
+ pixel_6206/PIX_OUT pixel_6206/CSA_VREF pixel
Xpixel_6217 pixel_6217/gring pixel_6217/VDD pixel_6217/GND pixel_6217/VREF pixel_6217/ROW_SEL
+ pixel_6217/NB1 pixel_6217/VBIAS pixel_6217/NB2 pixel_6217/AMP_IN pixel_6217/SF_IB
+ pixel_6217/PIX_OUT pixel_6217/CSA_VREF pixel
Xpixel_6228 pixel_6228/gring pixel_6228/VDD pixel_6228/GND pixel_6228/VREF pixel_6228/ROW_SEL
+ pixel_6228/NB1 pixel_6228/VBIAS pixel_6228/NB2 pixel_6228/AMP_IN pixel_6228/SF_IB
+ pixel_6228/PIX_OUT pixel_6228/CSA_VREF pixel
Xpixel_6239 pixel_6239/gring pixel_6239/VDD pixel_6239/GND pixel_6239/VREF pixel_6239/ROW_SEL
+ pixel_6239/NB1 pixel_6239/VBIAS pixel_6239/NB2 pixel_6239/AMP_IN pixel_6239/SF_IB
+ pixel_6239/PIX_OUT pixel_6239/CSA_VREF pixel
Xpixel_5505 pixel_5505/gring pixel_5505/VDD pixel_5505/GND pixel_5505/VREF pixel_5505/ROW_SEL
+ pixel_5505/NB1 pixel_5505/VBIAS pixel_5505/NB2 pixel_5505/AMP_IN pixel_5505/SF_IB
+ pixel_5505/PIX_OUT pixel_5505/CSA_VREF pixel
Xpixel_5516 pixel_5516/gring pixel_5516/VDD pixel_5516/GND pixel_5516/VREF pixel_5516/ROW_SEL
+ pixel_5516/NB1 pixel_5516/VBIAS pixel_5516/NB2 pixel_5516/AMP_IN pixel_5516/SF_IB
+ pixel_5516/PIX_OUT pixel_5516/CSA_VREF pixel
Xpixel_5527 pixel_5527/gring pixel_5527/VDD pixel_5527/GND pixel_5527/VREF pixel_5527/ROW_SEL
+ pixel_5527/NB1 pixel_5527/VBIAS pixel_5527/NB2 pixel_5527/AMP_IN pixel_5527/SF_IB
+ pixel_5527/PIX_OUT pixel_5527/CSA_VREF pixel
Xpixel_5538 pixel_5538/gring pixel_5538/VDD pixel_5538/GND pixel_5538/VREF pixel_5538/ROW_SEL
+ pixel_5538/NB1 pixel_5538/VBIAS pixel_5538/NB2 pixel_5538/AMP_IN pixel_5538/SF_IB
+ pixel_5538/PIX_OUT pixel_5538/CSA_VREF pixel
Xpixel_5549 pixel_5549/gring pixel_5549/VDD pixel_5549/GND pixel_5549/VREF pixel_5549/ROW_SEL
+ pixel_5549/NB1 pixel_5549/VBIAS pixel_5549/NB2 pixel_5549/AMP_IN pixel_5549/SF_IB
+ pixel_5549/PIX_OUT pixel_5549/CSA_VREF pixel
Xpixel_4804 pixel_4804/gring pixel_4804/VDD pixel_4804/GND pixel_4804/VREF pixel_4804/ROW_SEL
+ pixel_4804/NB1 pixel_4804/VBIAS pixel_4804/NB2 pixel_4804/AMP_IN pixel_4804/SF_IB
+ pixel_4804/PIX_OUT pixel_4804/CSA_VREF pixel
Xpixel_832 pixel_832/gring pixel_832/VDD pixel_832/GND pixel_832/VREF pixel_832/ROW_SEL
+ pixel_832/NB1 pixel_832/VBIAS pixel_832/NB2 pixel_832/AMP_IN pixel_832/SF_IB pixel_832/PIX_OUT
+ pixel_832/CSA_VREF pixel
Xpixel_821 pixel_821/gring pixel_821/VDD pixel_821/GND pixel_821/VREF pixel_821/ROW_SEL
+ pixel_821/NB1 pixel_821/VBIAS pixel_821/NB2 pixel_821/AMP_IN pixel_821/SF_IB pixel_821/PIX_OUT
+ pixel_821/CSA_VREF pixel
Xpixel_810 pixel_810/gring pixel_810/VDD pixel_810/GND pixel_810/VREF pixel_810/ROW_SEL
+ pixel_810/NB1 pixel_810/VBIAS pixel_810/NB2 pixel_810/AMP_IN pixel_810/SF_IB pixel_810/PIX_OUT
+ pixel_810/CSA_VREF pixel
Xpixel_4815 pixel_4815/gring pixel_4815/VDD pixel_4815/GND pixel_4815/VREF pixel_4815/ROW_SEL
+ pixel_4815/NB1 pixel_4815/VBIAS pixel_4815/NB2 pixel_4815/AMP_IN pixel_4815/SF_IB
+ pixel_4815/PIX_OUT pixel_4815/CSA_VREF pixel
Xpixel_4826 pixel_4826/gring pixel_4826/VDD pixel_4826/GND pixel_4826/VREF pixel_4826/ROW_SEL
+ pixel_4826/NB1 pixel_4826/VBIAS pixel_4826/NB2 pixel_4826/AMP_IN pixel_4826/SF_IB
+ pixel_4826/PIX_OUT pixel_4826/CSA_VREF pixel
Xpixel_4837 pixel_4837/gring pixel_4837/VDD pixel_4837/GND pixel_4837/VREF pixel_4837/ROW_SEL
+ pixel_4837/NB1 pixel_4837/VBIAS pixel_4837/NB2 pixel_4837/AMP_IN pixel_4837/SF_IB
+ pixel_4837/PIX_OUT pixel_4837/CSA_VREF pixel
Xpixel_876 pixel_876/gring pixel_876/VDD pixel_876/GND pixel_876/VREF pixel_876/ROW_SEL
+ pixel_876/NB1 pixel_876/VBIAS pixel_876/NB2 pixel_876/AMP_IN pixel_876/SF_IB pixel_876/PIX_OUT
+ pixel_876/CSA_VREF pixel
Xpixel_865 pixel_865/gring pixel_865/VDD pixel_865/GND pixel_865/VREF pixel_865/ROW_SEL
+ pixel_865/NB1 pixel_865/VBIAS pixel_865/NB2 pixel_865/AMP_IN pixel_865/SF_IB pixel_865/PIX_OUT
+ pixel_865/CSA_VREF pixel
Xpixel_854 pixel_854/gring pixel_854/VDD pixel_854/GND pixel_854/VREF pixel_854/ROW_SEL
+ pixel_854/NB1 pixel_854/VBIAS pixel_854/NB2 pixel_854/AMP_IN pixel_854/SF_IB pixel_854/PIX_OUT
+ pixel_854/CSA_VREF pixel
Xpixel_843 pixel_843/gring pixel_843/VDD pixel_843/GND pixel_843/VREF pixel_843/ROW_SEL
+ pixel_843/NB1 pixel_843/VBIAS pixel_843/NB2 pixel_843/AMP_IN pixel_843/SF_IB pixel_843/PIX_OUT
+ pixel_843/CSA_VREF pixel
Xpixel_4848 pixel_4848/gring pixel_4848/VDD pixel_4848/GND pixel_4848/VREF pixel_4848/ROW_SEL
+ pixel_4848/NB1 pixel_4848/VBIAS pixel_4848/NB2 pixel_4848/AMP_IN pixel_4848/SF_IB
+ pixel_4848/PIX_OUT pixel_4848/CSA_VREF pixel
Xpixel_4859 pixel_4859/gring pixel_4859/VDD pixel_4859/GND pixel_4859/VREF pixel_4859/ROW_SEL
+ pixel_4859/NB1 pixel_4859/VBIAS pixel_4859/NB2 pixel_4859/AMP_IN pixel_4859/SF_IB
+ pixel_4859/PIX_OUT pixel_4859/CSA_VREF pixel
Xpixel_898 pixel_898/gring pixel_898/VDD pixel_898/GND pixel_898/VREF pixel_898/ROW_SEL
+ pixel_898/NB1 pixel_898/VBIAS pixel_898/NB2 pixel_898/AMP_IN pixel_898/SF_IB pixel_898/PIX_OUT
+ pixel_898/CSA_VREF pixel
Xpixel_887 pixel_887/gring pixel_887/VDD pixel_887/GND pixel_887/VREF pixel_887/ROW_SEL
+ pixel_887/NB1 pixel_887/VBIAS pixel_887/NB2 pixel_887/AMP_IN pixel_887/SF_IB pixel_887/PIX_OUT
+ pixel_887/CSA_VREF pixel
Xpixel_8120 pixel_8120/gring pixel_8120/VDD pixel_8120/GND pixel_8120/VREF pixel_8120/ROW_SEL
+ pixel_8120/NB1 pixel_8120/VBIAS pixel_8120/NB2 pixel_8120/AMP_IN pixel_8120/SF_IB
+ pixel_8120/PIX_OUT pixel_8120/CSA_VREF pixel
Xpixel_8131 pixel_8131/gring pixel_8131/VDD pixel_8131/GND pixel_8131/VREF pixel_8131/ROW_SEL
+ pixel_8131/NB1 pixel_8131/VBIAS pixel_8131/NB2 pixel_8131/AMP_IN pixel_8131/SF_IB
+ pixel_8131/PIX_OUT pixel_8131/CSA_VREF pixel
Xpixel_8142 pixel_8142/gring pixel_8142/VDD pixel_8142/GND pixel_8142/VREF pixel_8142/ROW_SEL
+ pixel_8142/NB1 pixel_8142/VBIAS pixel_8142/NB2 pixel_8142/AMP_IN pixel_8142/SF_IB
+ pixel_8142/PIX_OUT pixel_8142/CSA_VREF pixel
Xpixel_8153 pixel_8153/gring pixel_8153/VDD pixel_8153/GND pixel_8153/VREF pixel_8153/ROW_SEL
+ pixel_8153/NB1 pixel_8153/VBIAS pixel_8153/NB2 pixel_8153/AMP_IN pixel_8153/SF_IB
+ pixel_8153/PIX_OUT pixel_8153/CSA_VREF pixel
Xpixel_8164 pixel_8164/gring pixel_8164/VDD pixel_8164/GND pixel_8164/VREF pixel_8164/ROW_SEL
+ pixel_8164/NB1 pixel_8164/VBIAS pixel_8164/NB2 pixel_8164/AMP_IN pixel_8164/SF_IB
+ pixel_8164/PIX_OUT pixel_8164/CSA_VREF pixel
Xpixel_8175 pixel_8175/gring pixel_8175/VDD pixel_8175/GND pixel_8175/VREF pixel_8175/ROW_SEL
+ pixel_8175/NB1 pixel_8175/VBIAS pixel_8175/NB2 pixel_8175/AMP_IN pixel_8175/SF_IB
+ pixel_8175/PIX_OUT pixel_8175/CSA_VREF pixel
Xpixel_8186 pixel_8186/gring pixel_8186/VDD pixel_8186/GND pixel_8186/VREF pixel_8186/ROW_SEL
+ pixel_8186/NB1 pixel_8186/VBIAS pixel_8186/NB2 pixel_8186/AMP_IN pixel_8186/SF_IB
+ pixel_8186/PIX_OUT pixel_8186/CSA_VREF pixel
Xpixel_7430 pixel_7430/gring pixel_7430/VDD pixel_7430/GND pixel_7430/VREF pixel_7430/ROW_SEL
+ pixel_7430/NB1 pixel_7430/VBIAS pixel_7430/NB2 pixel_7430/AMP_IN pixel_7430/SF_IB
+ pixel_7430/PIX_OUT pixel_7430/CSA_VREF pixel
Xpixel_7441 pixel_7441/gring pixel_7441/VDD pixel_7441/GND pixel_7441/VREF pixel_7441/ROW_SEL
+ pixel_7441/NB1 pixel_7441/VBIAS pixel_7441/NB2 pixel_7441/AMP_IN pixel_7441/SF_IB
+ pixel_7441/PIX_OUT pixel_7441/CSA_VREF pixel
Xpixel_8197 pixel_8197/gring pixel_8197/VDD pixel_8197/GND pixel_8197/VREF pixel_8197/ROW_SEL
+ pixel_8197/NB1 pixel_8197/VBIAS pixel_8197/NB2 pixel_8197/AMP_IN pixel_8197/SF_IB
+ pixel_8197/PIX_OUT pixel_8197/CSA_VREF pixel
Xpixel_7452 pixel_7452/gring pixel_7452/VDD pixel_7452/GND pixel_7452/VREF pixel_7452/ROW_SEL
+ pixel_7452/NB1 pixel_7452/VBIAS pixel_7452/NB2 pixel_7452/AMP_IN pixel_7452/SF_IB
+ pixel_7452/PIX_OUT pixel_7452/CSA_VREF pixel
Xpixel_7463 pixel_7463/gring pixel_7463/VDD pixel_7463/GND pixel_7463/VREF pixel_7463/ROW_SEL
+ pixel_7463/NB1 pixel_7463/VBIAS pixel_7463/NB2 pixel_7463/AMP_IN pixel_7463/SF_IB
+ pixel_7463/PIX_OUT pixel_7463/CSA_VREF pixel
Xpixel_7474 pixel_7474/gring pixel_7474/VDD pixel_7474/GND pixel_7474/VREF pixel_7474/ROW_SEL
+ pixel_7474/NB1 pixel_7474/VBIAS pixel_7474/NB2 pixel_7474/AMP_IN pixel_7474/SF_IB
+ pixel_7474/PIX_OUT pixel_7474/CSA_VREF pixel
Xpixel_7485 pixel_7485/gring pixel_7485/VDD pixel_7485/GND pixel_7485/VREF pixel_7485/ROW_SEL
+ pixel_7485/NB1 pixel_7485/VBIAS pixel_7485/NB2 pixel_7485/AMP_IN pixel_7485/SF_IB
+ pixel_7485/PIX_OUT pixel_7485/CSA_VREF pixel
Xpixel_7496 pixel_7496/gring pixel_7496/VDD pixel_7496/GND pixel_7496/VREF pixel_7496/ROW_SEL
+ pixel_7496/NB1 pixel_7496/VBIAS pixel_7496/NB2 pixel_7496/AMP_IN pixel_7496/SF_IB
+ pixel_7496/PIX_OUT pixel_7496/CSA_VREF pixel
Xpixel_6740 pixel_6740/gring pixel_6740/VDD pixel_6740/GND pixel_6740/VREF pixel_6740/ROW_SEL
+ pixel_6740/NB1 pixel_6740/VBIAS pixel_6740/NB2 pixel_6740/AMP_IN pixel_6740/SF_IB
+ pixel_6740/PIX_OUT pixel_6740/CSA_VREF pixel
Xpixel_6751 pixel_6751/gring pixel_6751/VDD pixel_6751/GND pixel_6751/VREF pixel_6751/ROW_SEL
+ pixel_6751/NB1 pixel_6751/VBIAS pixel_6751/NB2 pixel_6751/AMP_IN pixel_6751/SF_IB
+ pixel_6751/PIX_OUT pixel_6751/CSA_VREF pixel
Xpixel_6762 pixel_6762/gring pixel_6762/VDD pixel_6762/GND pixel_6762/VREF pixel_6762/ROW_SEL
+ pixel_6762/NB1 pixel_6762/VBIAS pixel_6762/NB2 pixel_6762/AMP_IN pixel_6762/SF_IB
+ pixel_6762/PIX_OUT pixel_6762/CSA_VREF pixel
Xpixel_6773 pixel_6773/gring pixel_6773/VDD pixel_6773/GND pixel_6773/VREF pixel_6773/ROW_SEL
+ pixel_6773/NB1 pixel_6773/VBIAS pixel_6773/NB2 pixel_6773/AMP_IN pixel_6773/SF_IB
+ pixel_6773/PIX_OUT pixel_6773/CSA_VREF pixel
Xpixel_6784 pixel_6784/gring pixel_6784/VDD pixel_6784/GND pixel_6784/VREF pixel_6784/ROW_SEL
+ pixel_6784/NB1 pixel_6784/VBIAS pixel_6784/NB2 pixel_6784/AMP_IN pixel_6784/SF_IB
+ pixel_6784/PIX_OUT pixel_6784/CSA_VREF pixel
Xpixel_6795 pixel_6795/gring pixel_6795/VDD pixel_6795/GND pixel_6795/VREF pixel_6795/ROW_SEL
+ pixel_6795/NB1 pixel_6795/VBIAS pixel_6795/NB2 pixel_6795/AMP_IN pixel_6795/SF_IB
+ pixel_6795/PIX_OUT pixel_6795/CSA_VREF pixel
Xpixel_1091 pixel_1091/gring pixel_1091/VDD pixel_1091/GND pixel_1091/VREF pixel_1091/ROW_SEL
+ pixel_1091/NB1 pixel_1091/VBIAS pixel_1091/NB2 pixel_1091/AMP_IN pixel_1091/SF_IB
+ pixel_1091/PIX_OUT pixel_1091/CSA_VREF pixel
Xpixel_1080 pixel_1080/gring pixel_1080/VDD pixel_1080/GND pixel_1080/VREF pixel_1080/ROW_SEL
+ pixel_1080/NB1 pixel_1080/VBIAS pixel_1080/NB2 pixel_1080/AMP_IN pixel_1080/SF_IB
+ pixel_1080/PIX_OUT pixel_1080/CSA_VREF pixel
Xpixel_128 pixel_128/gring pixel_128/VDD pixel_128/GND pixel_128/VREF pixel_128/ROW_SEL
+ pixel_128/NB1 pixel_128/VBIAS pixel_128/NB2 pixel_128/AMP_IN pixel_128/SF_IB pixel_128/PIX_OUT
+ pixel_128/CSA_VREF pixel
Xpixel_117 pixel_117/gring pixel_117/VDD pixel_117/GND pixel_117/VREF pixel_117/ROW_SEL
+ pixel_117/NB1 pixel_117/VBIAS pixel_117/NB2 pixel_117/AMP_IN pixel_117/SF_IB pixel_117/PIX_OUT
+ pixel_117/CSA_VREF pixel
Xpixel_106 pixel_106/gring pixel_106/VDD pixel_106/GND pixel_106/VREF pixel_106/ROW_SEL
+ pixel_106/NB1 pixel_106/VBIAS pixel_106/NB2 pixel_106/AMP_IN pixel_106/SF_IB pixel_106/PIX_OUT
+ pixel_106/CSA_VREF pixel
Xpixel_139 pixel_139/gring pixel_139/VDD pixel_139/GND pixel_139/VREF pixel_139/ROW_SEL
+ pixel_139/NB1 pixel_139/VBIAS pixel_139/NB2 pixel_139/AMP_IN pixel_139/SF_IB pixel_139/PIX_OUT
+ pixel_139/CSA_VREF pixel
Xpixel_2709 pixel_2709/gring pixel_2709/VDD pixel_2709/GND pixel_2709/VREF pixel_2709/ROW_SEL
+ pixel_2709/NB1 pixel_2709/VBIAS pixel_2709/NB2 pixel_2709/AMP_IN pixel_2709/SF_IB
+ pixel_2709/PIX_OUT pixel_2709/CSA_VREF pixel
Xpixel_6003 pixel_6003/gring pixel_6003/VDD pixel_6003/GND pixel_6003/VREF pixel_6003/ROW_SEL
+ pixel_6003/NB1 pixel_6003/VBIAS pixel_6003/NB2 pixel_6003/AMP_IN pixel_6003/SF_IB
+ pixel_6003/PIX_OUT pixel_6003/CSA_VREF pixel
Xpixel_6014 pixel_6014/gring pixel_6014/VDD pixel_6014/GND pixel_6014/VREF pixel_6014/ROW_SEL
+ pixel_6014/NB1 pixel_6014/VBIAS pixel_6014/NB2 pixel_6014/AMP_IN pixel_6014/SF_IB
+ pixel_6014/PIX_OUT pixel_6014/CSA_VREF pixel
Xpixel_6025 pixel_6025/gring pixel_6025/VDD pixel_6025/GND pixel_6025/VREF pixel_6025/ROW_SEL
+ pixel_6025/NB1 pixel_6025/VBIAS pixel_6025/NB2 pixel_6025/AMP_IN pixel_6025/SF_IB
+ pixel_6025/PIX_OUT pixel_6025/CSA_VREF pixel
Xpixel_6036 pixel_6036/gring pixel_6036/VDD pixel_6036/GND pixel_6036/VREF pixel_6036/ROW_SEL
+ pixel_6036/NB1 pixel_6036/VBIAS pixel_6036/NB2 pixel_6036/AMP_IN pixel_6036/SF_IB
+ pixel_6036/PIX_OUT pixel_6036/CSA_VREF pixel
Xpixel_6047 pixel_6047/gring pixel_6047/VDD pixel_6047/GND pixel_6047/VREF pixel_6047/ROW_SEL
+ pixel_6047/NB1 pixel_6047/VBIAS pixel_6047/NB2 pixel_6047/AMP_IN pixel_6047/SF_IB
+ pixel_6047/PIX_OUT pixel_6047/CSA_VREF pixel
Xpixel_6058 pixel_6058/gring pixel_6058/VDD pixel_6058/GND pixel_6058/VREF pixel_6058/ROW_SEL
+ pixel_6058/NB1 pixel_6058/VBIAS pixel_6058/NB2 pixel_6058/AMP_IN pixel_6058/SF_IB
+ pixel_6058/PIX_OUT pixel_6058/CSA_VREF pixel
Xpixel_5302 pixel_5302/gring pixel_5302/VDD pixel_5302/GND pixel_5302/VREF pixel_5302/ROW_SEL
+ pixel_5302/NB1 pixel_5302/VBIAS pixel_5302/NB2 pixel_5302/AMP_IN pixel_5302/SF_IB
+ pixel_5302/PIX_OUT pixel_5302/CSA_VREF pixel
Xpixel_5313 pixel_5313/gring pixel_5313/VDD pixel_5313/GND pixel_5313/VREF pixel_5313/ROW_SEL
+ pixel_5313/NB1 pixel_5313/VBIAS pixel_5313/NB2 pixel_5313/AMP_IN pixel_5313/SF_IB
+ pixel_5313/PIX_OUT pixel_5313/CSA_VREF pixel
Xpixel_6069 pixel_6069/gring pixel_6069/VDD pixel_6069/GND pixel_6069/VREF pixel_6069/ROW_SEL
+ pixel_6069/NB1 pixel_6069/VBIAS pixel_6069/NB2 pixel_6069/AMP_IN pixel_6069/SF_IB
+ pixel_6069/PIX_OUT pixel_6069/CSA_VREF pixel
Xpixel_5324 pixel_5324/gring pixel_5324/VDD pixel_5324/GND pixel_5324/VREF pixel_5324/ROW_SEL
+ pixel_5324/NB1 pixel_5324/VBIAS pixel_5324/NB2 pixel_5324/AMP_IN pixel_5324/SF_IB
+ pixel_5324/PIX_OUT pixel_5324/CSA_VREF pixel
Xpixel_5335 pixel_5335/gring pixel_5335/VDD pixel_5335/GND pixel_5335/VREF pixel_5335/ROW_SEL
+ pixel_5335/NB1 pixel_5335/VBIAS pixel_5335/NB2 pixel_5335/AMP_IN pixel_5335/SF_IB
+ pixel_5335/PIX_OUT pixel_5335/CSA_VREF pixel
Xpixel_5346 pixel_5346/gring pixel_5346/VDD pixel_5346/GND pixel_5346/VREF pixel_5346/ROW_SEL
+ pixel_5346/NB1 pixel_5346/VBIAS pixel_5346/NB2 pixel_5346/AMP_IN pixel_5346/SF_IB
+ pixel_5346/PIX_OUT pixel_5346/CSA_VREF pixel
Xpixel_5357 pixel_5357/gring pixel_5357/VDD pixel_5357/GND pixel_5357/VREF pixel_5357/ROW_SEL
+ pixel_5357/NB1 pixel_5357/VBIAS pixel_5357/NB2 pixel_5357/AMP_IN pixel_5357/SF_IB
+ pixel_5357/PIX_OUT pixel_5357/CSA_VREF pixel
Xpixel_4601 pixel_4601/gring pixel_4601/VDD pixel_4601/GND pixel_4601/VREF pixel_4601/ROW_SEL
+ pixel_4601/NB1 pixel_4601/VBIAS pixel_4601/NB2 pixel_4601/AMP_IN pixel_4601/SF_IB
+ pixel_4601/PIX_OUT pixel_4601/CSA_VREF pixel
Xpixel_4612 pixel_4612/gring pixel_4612/VDD pixel_4612/GND pixel_4612/VREF pixel_4612/ROW_SEL
+ pixel_4612/NB1 pixel_4612/VBIAS pixel_4612/NB2 pixel_4612/AMP_IN pixel_4612/SF_IB
+ pixel_4612/PIX_OUT pixel_4612/CSA_VREF pixel
Xpixel_640 pixel_640/gring pixel_640/VDD pixel_640/GND pixel_640/VREF pixel_640/ROW_SEL
+ pixel_640/NB1 pixel_640/VBIAS pixel_640/NB2 pixel_640/AMP_IN pixel_640/SF_IB pixel_640/PIX_OUT
+ pixel_640/CSA_VREF pixel
Xpixel_5368 pixel_5368/gring pixel_5368/VDD pixel_5368/GND pixel_5368/VREF pixel_5368/ROW_SEL
+ pixel_5368/NB1 pixel_5368/VBIAS pixel_5368/NB2 pixel_5368/AMP_IN pixel_5368/SF_IB
+ pixel_5368/PIX_OUT pixel_5368/CSA_VREF pixel
Xpixel_5379 pixel_5379/gring pixel_5379/VDD pixel_5379/GND pixel_5379/VREF pixel_5379/ROW_SEL
+ pixel_5379/NB1 pixel_5379/VBIAS pixel_5379/NB2 pixel_5379/AMP_IN pixel_5379/SF_IB
+ pixel_5379/PIX_OUT pixel_5379/CSA_VREF pixel
Xpixel_4623 pixel_4623/gring pixel_4623/VDD pixel_4623/GND pixel_4623/VREF pixel_4623/ROW_SEL
+ pixel_4623/NB1 pixel_4623/VBIAS pixel_4623/NB2 pixel_4623/AMP_IN pixel_4623/SF_IB
+ pixel_4623/PIX_OUT pixel_4623/CSA_VREF pixel
Xpixel_4634 pixel_4634/gring pixel_4634/VDD pixel_4634/GND pixel_4634/VREF pixel_4634/ROW_SEL
+ pixel_4634/NB1 pixel_4634/VBIAS pixel_4634/NB2 pixel_4634/AMP_IN pixel_4634/SF_IB
+ pixel_4634/PIX_OUT pixel_4634/CSA_VREF pixel
Xpixel_4645 pixel_4645/gring pixel_4645/VDD pixel_4645/GND pixel_4645/VREF pixel_4645/ROW_SEL
+ pixel_4645/NB1 pixel_4645/VBIAS pixel_4645/NB2 pixel_4645/AMP_IN pixel_4645/SF_IB
+ pixel_4645/PIX_OUT pixel_4645/CSA_VREF pixel
Xpixel_3900 pixel_3900/gring pixel_3900/VDD pixel_3900/GND pixel_3900/VREF pixel_3900/ROW_SEL
+ pixel_3900/NB1 pixel_3900/VBIAS pixel_3900/NB2 pixel_3900/AMP_IN pixel_3900/SF_IB
+ pixel_3900/PIX_OUT pixel_3900/CSA_VREF pixel
Xpixel_684 pixel_684/gring pixel_684/VDD pixel_684/GND pixel_684/VREF pixel_684/ROW_SEL
+ pixel_684/NB1 pixel_684/VBIAS pixel_684/NB2 pixel_684/AMP_IN pixel_684/SF_IB pixel_684/PIX_OUT
+ pixel_684/CSA_VREF pixel
Xpixel_673 pixel_673/gring pixel_673/VDD pixel_673/GND pixel_673/VREF pixel_673/ROW_SEL
+ pixel_673/NB1 pixel_673/VBIAS pixel_673/NB2 pixel_673/AMP_IN pixel_673/SF_IB pixel_673/PIX_OUT
+ pixel_673/CSA_VREF pixel
Xpixel_662 pixel_662/gring pixel_662/VDD pixel_662/GND pixel_662/VREF pixel_662/ROW_SEL
+ pixel_662/NB1 pixel_662/VBIAS pixel_662/NB2 pixel_662/AMP_IN pixel_662/SF_IB pixel_662/PIX_OUT
+ pixel_662/CSA_VREF pixel
Xpixel_651 pixel_651/gring pixel_651/VDD pixel_651/GND pixel_651/VREF pixel_651/ROW_SEL
+ pixel_651/NB1 pixel_651/VBIAS pixel_651/NB2 pixel_651/AMP_IN pixel_651/SF_IB pixel_651/PIX_OUT
+ pixel_651/CSA_VREF pixel
Xpixel_4656 pixel_4656/gring pixel_4656/VDD pixel_4656/GND pixel_4656/VREF pixel_4656/ROW_SEL
+ pixel_4656/NB1 pixel_4656/VBIAS pixel_4656/NB2 pixel_4656/AMP_IN pixel_4656/SF_IB
+ pixel_4656/PIX_OUT pixel_4656/CSA_VREF pixel
Xpixel_4667 pixel_4667/gring pixel_4667/VDD pixel_4667/GND pixel_4667/VREF pixel_4667/ROW_SEL
+ pixel_4667/NB1 pixel_4667/VBIAS pixel_4667/NB2 pixel_4667/AMP_IN pixel_4667/SF_IB
+ pixel_4667/PIX_OUT pixel_4667/CSA_VREF pixel
Xpixel_4678 pixel_4678/gring pixel_4678/VDD pixel_4678/GND pixel_4678/VREF pixel_4678/ROW_SEL
+ pixel_4678/NB1 pixel_4678/VBIAS pixel_4678/NB2 pixel_4678/AMP_IN pixel_4678/SF_IB
+ pixel_4678/PIX_OUT pixel_4678/CSA_VREF pixel
Xpixel_4689 pixel_4689/gring pixel_4689/VDD pixel_4689/GND pixel_4689/VREF pixel_4689/ROW_SEL
+ pixel_4689/NB1 pixel_4689/VBIAS pixel_4689/NB2 pixel_4689/AMP_IN pixel_4689/SF_IB
+ pixel_4689/PIX_OUT pixel_4689/CSA_VREF pixel
Xpixel_3911 pixel_3911/gring pixel_3911/VDD pixel_3911/GND pixel_3911/VREF pixel_3911/ROW_SEL
+ pixel_3911/NB1 pixel_3911/VBIAS pixel_3911/NB2 pixel_3911/AMP_IN pixel_3911/SF_IB
+ pixel_3911/PIX_OUT pixel_3911/CSA_VREF pixel
Xpixel_3922 pixel_3922/gring pixel_3922/VDD pixel_3922/GND pixel_3922/VREF pixel_3922/ROW_SEL
+ pixel_3922/NB1 pixel_3922/VBIAS pixel_3922/NB2 pixel_3922/AMP_IN pixel_3922/SF_IB
+ pixel_3922/PIX_OUT pixel_3922/CSA_VREF pixel
Xpixel_3933 pixel_3933/gring pixel_3933/VDD pixel_3933/GND pixel_3933/VREF pixel_3933/ROW_SEL
+ pixel_3933/NB1 pixel_3933/VBIAS pixel_3933/NB2 pixel_3933/AMP_IN pixel_3933/SF_IB
+ pixel_3933/PIX_OUT pixel_3933/CSA_VREF pixel
Xpixel_3944 pixel_3944/gring pixel_3944/VDD pixel_3944/GND pixel_3944/VREF pixel_3944/ROW_SEL
+ pixel_3944/NB1 pixel_3944/VBIAS pixel_3944/NB2 pixel_3944/AMP_IN pixel_3944/SF_IB
+ pixel_3944/PIX_OUT pixel_3944/CSA_VREF pixel
Xpixel_695 pixel_695/gring pixel_695/VDD pixel_695/GND pixel_695/VREF pixel_695/ROW_SEL
+ pixel_695/NB1 pixel_695/VBIAS pixel_695/NB2 pixel_695/AMP_IN pixel_695/SF_IB pixel_695/PIX_OUT
+ pixel_695/CSA_VREF pixel
Xpixel_3955 pixel_3955/gring pixel_3955/VDD pixel_3955/GND pixel_3955/VREF pixel_3955/ROW_SEL
+ pixel_3955/NB1 pixel_3955/VBIAS pixel_3955/NB2 pixel_3955/AMP_IN pixel_3955/SF_IB
+ pixel_3955/PIX_OUT pixel_3955/CSA_VREF pixel
Xpixel_3966 pixel_3966/gring pixel_3966/VDD pixel_3966/GND pixel_3966/VREF pixel_3966/ROW_SEL
+ pixel_3966/NB1 pixel_3966/VBIAS pixel_3966/NB2 pixel_3966/AMP_IN pixel_3966/SF_IB
+ pixel_3966/PIX_OUT pixel_3966/CSA_VREF pixel
Xpixel_3977 pixel_3977/gring pixel_3977/VDD pixel_3977/GND pixel_3977/VREF pixel_3977/ROW_SEL
+ pixel_3977/NB1 pixel_3977/VBIAS pixel_3977/NB2 pixel_3977/AMP_IN pixel_3977/SF_IB
+ pixel_3977/PIX_OUT pixel_3977/CSA_VREF pixel
Xpixel_3988 pixel_3988/gring pixel_3988/VDD pixel_3988/GND pixel_3988/VREF pixel_3988/ROW_SEL
+ pixel_3988/NB1 pixel_3988/VBIAS pixel_3988/NB2 pixel_3988/AMP_IN pixel_3988/SF_IB
+ pixel_3988/PIX_OUT pixel_3988/CSA_VREF pixel
Xpixel_3999 pixel_3999/gring pixel_3999/VDD pixel_3999/GND pixel_3999/VREF pixel_3999/ROW_SEL
+ pixel_3999/NB1 pixel_3999/VBIAS pixel_3999/NB2 pixel_3999/AMP_IN pixel_3999/SF_IB
+ pixel_3999/PIX_OUT pixel_3999/CSA_VREF pixel
Xpixel_9 pixel_9/gring pixel_9/VDD pixel_9/GND pixel_9/VREF pixel_9/ROW_SEL pixel_9/NB1
+ pixel_9/VBIAS pixel_9/NB2 pixel_9/AMP_IN pixel_9/SF_IB pixel_9/PIX_OUT pixel_9/CSA_VREF
+ pixel
Xpixel_7260 pixel_7260/gring pixel_7260/VDD pixel_7260/GND pixel_7260/VREF pixel_7260/ROW_SEL
+ pixel_7260/NB1 pixel_7260/VBIAS pixel_7260/NB2 pixel_7260/AMP_IN pixel_7260/SF_IB
+ pixel_7260/PIX_OUT pixel_7260/CSA_VREF pixel
Xpixel_7271 pixel_7271/gring pixel_7271/VDD pixel_7271/GND pixel_7271/VREF pixel_7271/ROW_SEL
+ pixel_7271/NB1 pixel_7271/VBIAS pixel_7271/NB2 pixel_7271/AMP_IN pixel_7271/SF_IB
+ pixel_7271/PIX_OUT pixel_7271/CSA_VREF pixel
Xpixel_7282 pixel_7282/gring pixel_7282/VDD pixel_7282/GND pixel_7282/VREF pixel_7282/ROW_SEL
+ pixel_7282/NB1 pixel_7282/VBIAS pixel_7282/NB2 pixel_7282/AMP_IN pixel_7282/SF_IB
+ pixel_7282/PIX_OUT pixel_7282/CSA_VREF pixel
Xpixel_7293 pixel_7293/gring pixel_7293/VDD pixel_7293/GND pixel_7293/VREF pixel_7293/ROW_SEL
+ pixel_7293/NB1 pixel_7293/VBIAS pixel_7293/NB2 pixel_7293/AMP_IN pixel_7293/SF_IB
+ pixel_7293/PIX_OUT pixel_7293/CSA_VREF pixel
Xpixel_6570 pixel_6570/gring pixel_6570/VDD pixel_6570/GND pixel_6570/VREF pixel_6570/ROW_SEL
+ pixel_6570/NB1 pixel_6570/VBIAS pixel_6570/NB2 pixel_6570/AMP_IN pixel_6570/SF_IB
+ pixel_6570/PIX_OUT pixel_6570/CSA_VREF pixel
Xpixel_6581 pixel_6581/gring pixel_6581/VDD pixel_6581/GND pixel_6581/VREF pixel_6581/ROW_SEL
+ pixel_6581/NB1 pixel_6581/VBIAS pixel_6581/NB2 pixel_6581/AMP_IN pixel_6581/SF_IB
+ pixel_6581/PIX_OUT pixel_6581/CSA_VREF pixel
Xpixel_6592 pixel_6592/gring pixel_6592/VDD pixel_6592/GND pixel_6592/VREF pixel_6592/ROW_SEL
+ pixel_6592/NB1 pixel_6592/VBIAS pixel_6592/NB2 pixel_6592/AMP_IN pixel_6592/SF_IB
+ pixel_6592/PIX_OUT pixel_6592/CSA_VREF pixel
Xpixel_5880 pixel_5880/gring pixel_5880/VDD pixel_5880/GND pixel_5880/VREF pixel_5880/ROW_SEL
+ pixel_5880/NB1 pixel_5880/VBIAS pixel_5880/NB2 pixel_5880/AMP_IN pixel_5880/SF_IB
+ pixel_5880/PIX_OUT pixel_5880/CSA_VREF pixel
Xpixel_5891 pixel_5891/gring pixel_5891/VDD pixel_5891/GND pixel_5891/VREF pixel_5891/ROW_SEL
+ pixel_5891/NB1 pixel_5891/VBIAS pixel_5891/NB2 pixel_5891/AMP_IN pixel_5891/SF_IB
+ pixel_5891/PIX_OUT pixel_5891/CSA_VREF pixel
Xpixel_3229 pixel_3229/gring pixel_3229/VDD pixel_3229/GND pixel_3229/VREF pixel_3229/ROW_SEL
+ pixel_3229/NB1 pixel_3229/VBIAS pixel_3229/NB2 pixel_3229/AMP_IN pixel_3229/SF_IB
+ pixel_3229/PIX_OUT pixel_3229/CSA_VREF pixel
Xpixel_3218 pixel_3218/gring pixel_3218/VDD pixel_3218/GND pixel_3218/VREF pixel_3218/ROW_SEL
+ pixel_3218/NB1 pixel_3218/VBIAS pixel_3218/NB2 pixel_3218/AMP_IN pixel_3218/SF_IB
+ pixel_3218/PIX_OUT pixel_3218/CSA_VREF pixel
Xpixel_3207 pixel_3207/gring pixel_3207/VDD pixel_3207/GND pixel_3207/VREF pixel_3207/ROW_SEL
+ pixel_3207/NB1 pixel_3207/VBIAS pixel_3207/NB2 pixel_3207/AMP_IN pixel_3207/SF_IB
+ pixel_3207/PIX_OUT pixel_3207/CSA_VREF pixel
Xpixel_2528 pixel_2528/gring pixel_2528/VDD pixel_2528/GND pixel_2528/VREF pixel_2528/ROW_SEL
+ pixel_2528/NB1 pixel_2528/VBIAS pixel_2528/NB2 pixel_2528/AMP_IN pixel_2528/SF_IB
+ pixel_2528/PIX_OUT pixel_2528/CSA_VREF pixel
Xpixel_2517 pixel_2517/gring pixel_2517/VDD pixel_2517/GND pixel_2517/VREF pixel_2517/ROW_SEL
+ pixel_2517/NB1 pixel_2517/VBIAS pixel_2517/NB2 pixel_2517/AMP_IN pixel_2517/SF_IB
+ pixel_2517/PIX_OUT pixel_2517/CSA_VREF pixel
Xpixel_2506 pixel_2506/gring pixel_2506/VDD pixel_2506/GND pixel_2506/VREF pixel_2506/ROW_SEL
+ pixel_2506/NB1 pixel_2506/VBIAS pixel_2506/NB2 pixel_2506/AMP_IN pixel_2506/SF_IB
+ pixel_2506/PIX_OUT pixel_2506/CSA_VREF pixel
Xpixel_1816 pixel_1816/gring pixel_1816/VDD pixel_1816/GND pixel_1816/VREF pixel_1816/ROW_SEL
+ pixel_1816/NB1 pixel_1816/VBIAS pixel_1816/NB2 pixel_1816/AMP_IN pixel_1816/SF_IB
+ pixel_1816/PIX_OUT pixel_1816/CSA_VREF pixel
Xpixel_1805 pixel_1805/gring pixel_1805/VDD pixel_1805/GND pixel_1805/VREF pixel_1805/ROW_SEL
+ pixel_1805/NB1 pixel_1805/VBIAS pixel_1805/NB2 pixel_1805/AMP_IN pixel_1805/SF_IB
+ pixel_1805/PIX_OUT pixel_1805/CSA_VREF pixel
Xpixel_2539 pixel_2539/gring pixel_2539/VDD pixel_2539/GND pixel_2539/VREF pixel_2539/ROW_SEL
+ pixel_2539/NB1 pixel_2539/VBIAS pixel_2539/NB2 pixel_2539/AMP_IN pixel_2539/SF_IB
+ pixel_2539/PIX_OUT pixel_2539/CSA_VREF pixel
Xpixel_1849 pixel_1849/gring pixel_1849/VDD pixel_1849/GND pixel_1849/VREF pixel_1849/ROW_SEL
+ pixel_1849/NB1 pixel_1849/VBIAS pixel_1849/NB2 pixel_1849/AMP_IN pixel_1849/SF_IB
+ pixel_1849/PIX_OUT pixel_1849/CSA_VREF pixel
Xpixel_1838 pixel_1838/gring pixel_1838/VDD pixel_1838/GND pixel_1838/VREF pixel_1838/ROW_SEL
+ pixel_1838/NB1 pixel_1838/VBIAS pixel_1838/NB2 pixel_1838/AMP_IN pixel_1838/SF_IB
+ pixel_1838/PIX_OUT pixel_1838/CSA_VREF pixel
Xpixel_1827 pixel_1827/gring pixel_1827/VDD pixel_1827/GND pixel_1827/VREF pixel_1827/ROW_SEL
+ pixel_1827/NB1 pixel_1827/VBIAS pixel_1827/NB2 pixel_1827/AMP_IN pixel_1827/SF_IB
+ pixel_1827/PIX_OUT pixel_1827/CSA_VREF pixel
Xpixel_5110 pixel_5110/gring pixel_5110/VDD pixel_5110/GND pixel_5110/VREF pixel_5110/ROW_SEL
+ pixel_5110/NB1 pixel_5110/VBIAS pixel_5110/NB2 pixel_5110/AMP_IN pixel_5110/SF_IB
+ pixel_5110/PIX_OUT pixel_5110/CSA_VREF pixel
Xpixel_5121 pixel_5121/gring pixel_5121/VDD pixel_5121/GND pixel_5121/VREF pixel_5121/ROW_SEL
+ pixel_5121/NB1 pixel_5121/VBIAS pixel_5121/NB2 pixel_5121/AMP_IN pixel_5121/SF_IB
+ pixel_5121/PIX_OUT pixel_5121/CSA_VREF pixel
Xpixel_5132 pixel_5132/gring pixel_5132/VDD pixel_5132/GND pixel_5132/VREF pixel_5132/ROW_SEL
+ pixel_5132/NB1 pixel_5132/VBIAS pixel_5132/NB2 pixel_5132/AMP_IN pixel_5132/SF_IB
+ pixel_5132/PIX_OUT pixel_5132/CSA_VREF pixel
Xpixel_5143 pixel_5143/gring pixel_5143/VDD pixel_5143/GND pixel_5143/VREF pixel_5143/ROW_SEL
+ pixel_5143/NB1 pixel_5143/VBIAS pixel_5143/NB2 pixel_5143/AMP_IN pixel_5143/SF_IB
+ pixel_5143/PIX_OUT pixel_5143/CSA_VREF pixel
Xpixel_5154 pixel_5154/gring pixel_5154/VDD pixel_5154/GND pixel_5154/VREF pixel_5154/ROW_SEL
+ pixel_5154/NB1 pixel_5154/VBIAS pixel_5154/NB2 pixel_5154/AMP_IN pixel_5154/SF_IB
+ pixel_5154/PIX_OUT pixel_5154/CSA_VREF pixel
Xpixel_5165 pixel_5165/gring pixel_5165/VDD pixel_5165/GND pixel_5165/VREF pixel_5165/ROW_SEL
+ pixel_5165/NB1 pixel_5165/VBIAS pixel_5165/NB2 pixel_5165/AMP_IN pixel_5165/SF_IB
+ pixel_5165/PIX_OUT pixel_5165/CSA_VREF pixel
Xpixel_4420 pixel_4420/gring pixel_4420/VDD pixel_4420/GND pixel_4420/VREF pixel_4420/ROW_SEL
+ pixel_4420/NB1 pixel_4420/VBIAS pixel_4420/NB2 pixel_4420/AMP_IN pixel_4420/SF_IB
+ pixel_4420/PIX_OUT pixel_4420/CSA_VREF pixel
Xpixel_5176 pixel_5176/gring pixel_5176/VDD pixel_5176/GND pixel_5176/VREF pixel_5176/ROW_SEL
+ pixel_5176/NB1 pixel_5176/VBIAS pixel_5176/NB2 pixel_5176/AMP_IN pixel_5176/SF_IB
+ pixel_5176/PIX_OUT pixel_5176/CSA_VREF pixel
Xpixel_5187 pixel_5187/gring pixel_5187/VDD pixel_5187/GND pixel_5187/VREF pixel_5187/ROW_SEL
+ pixel_5187/NB1 pixel_5187/VBIAS pixel_5187/NB2 pixel_5187/AMP_IN pixel_5187/SF_IB
+ pixel_5187/PIX_OUT pixel_5187/CSA_VREF pixel
Xpixel_5198 pixel_5198/gring pixel_5198/VDD pixel_5198/GND pixel_5198/VREF pixel_5198/ROW_SEL
+ pixel_5198/NB1 pixel_5198/VBIAS pixel_5198/NB2 pixel_5198/AMP_IN pixel_5198/SF_IB
+ pixel_5198/PIX_OUT pixel_5198/CSA_VREF pixel
Xpixel_4431 pixel_4431/gring pixel_4431/VDD pixel_4431/GND pixel_4431/VREF pixel_4431/ROW_SEL
+ pixel_4431/NB1 pixel_4431/VBIAS pixel_4431/NB2 pixel_4431/AMP_IN pixel_4431/SF_IB
+ pixel_4431/PIX_OUT pixel_4431/CSA_VREF pixel
Xpixel_4442 pixel_4442/gring pixel_4442/VDD pixel_4442/GND pixel_4442/VREF pixel_4442/ROW_SEL
+ pixel_4442/NB1 pixel_4442/VBIAS pixel_4442/NB2 pixel_4442/AMP_IN pixel_4442/SF_IB
+ pixel_4442/PIX_OUT pixel_4442/CSA_VREF pixel
Xpixel_4453 pixel_4453/gring pixel_4453/VDD pixel_4453/GND pixel_4453/VREF pixel_4453/ROW_SEL
+ pixel_4453/NB1 pixel_4453/VBIAS pixel_4453/NB2 pixel_4453/AMP_IN pixel_4453/SF_IB
+ pixel_4453/PIX_OUT pixel_4453/CSA_VREF pixel
Xpixel_492 pixel_492/gring pixel_492/VDD pixel_492/GND pixel_492/VREF pixel_492/ROW_SEL
+ pixel_492/NB1 pixel_492/VBIAS pixel_492/NB2 pixel_492/AMP_IN pixel_492/SF_IB pixel_492/PIX_OUT
+ pixel_492/CSA_VREF pixel
Xpixel_481 pixel_481/gring pixel_481/VDD pixel_481/GND pixel_481/VREF pixel_481/ROW_SEL
+ pixel_481/NB1 pixel_481/VBIAS pixel_481/NB2 pixel_481/AMP_IN pixel_481/SF_IB pixel_481/PIX_OUT
+ pixel_481/CSA_VREF pixel
Xpixel_470 pixel_470/gring pixel_470/VDD pixel_470/GND pixel_470/VREF pixel_470/ROW_SEL
+ pixel_470/NB1 pixel_470/VBIAS pixel_470/NB2 pixel_470/AMP_IN pixel_470/SF_IB pixel_470/PIX_OUT
+ pixel_470/CSA_VREF pixel
Xpixel_3752 pixel_3752/gring pixel_3752/VDD pixel_3752/GND pixel_3752/VREF pixel_3752/ROW_SEL
+ pixel_3752/NB1 pixel_3752/VBIAS pixel_3752/NB2 pixel_3752/AMP_IN pixel_3752/SF_IB
+ pixel_3752/PIX_OUT pixel_3752/CSA_VREF pixel
Xpixel_3741 pixel_3741/gring pixel_3741/VDD pixel_3741/GND pixel_3741/VREF pixel_3741/ROW_SEL
+ pixel_3741/NB1 pixel_3741/VBIAS pixel_3741/NB2 pixel_3741/AMP_IN pixel_3741/SF_IB
+ pixel_3741/PIX_OUT pixel_3741/CSA_VREF pixel
Xpixel_3730 pixel_3730/gring pixel_3730/VDD pixel_3730/GND pixel_3730/VREF pixel_3730/ROW_SEL
+ pixel_3730/NB1 pixel_3730/VBIAS pixel_3730/NB2 pixel_3730/AMP_IN pixel_3730/SF_IB
+ pixel_3730/PIX_OUT pixel_3730/CSA_VREF pixel
Xpixel_4464 pixel_4464/gring pixel_4464/VDD pixel_4464/GND pixel_4464/VREF pixel_4464/ROW_SEL
+ pixel_4464/NB1 pixel_4464/VBIAS pixel_4464/NB2 pixel_4464/AMP_IN pixel_4464/SF_IB
+ pixel_4464/PIX_OUT pixel_4464/CSA_VREF pixel
Xpixel_4475 pixel_4475/gring pixel_4475/VDD pixel_4475/GND pixel_4475/VREF pixel_4475/ROW_SEL
+ pixel_4475/NB1 pixel_4475/VBIAS pixel_4475/NB2 pixel_4475/AMP_IN pixel_4475/SF_IB
+ pixel_4475/PIX_OUT pixel_4475/CSA_VREF pixel
Xpixel_4486 pixel_4486/gring pixel_4486/VDD pixel_4486/GND pixel_4486/VREF pixel_4486/ROW_SEL
+ pixel_4486/NB1 pixel_4486/VBIAS pixel_4486/NB2 pixel_4486/AMP_IN pixel_4486/SF_IB
+ pixel_4486/PIX_OUT pixel_4486/CSA_VREF pixel
Xpixel_4497 pixel_4497/gring pixel_4497/VDD pixel_4497/GND pixel_4497/VREF pixel_4497/ROW_SEL
+ pixel_4497/NB1 pixel_4497/VBIAS pixel_4497/NB2 pixel_4497/AMP_IN pixel_4497/SF_IB
+ pixel_4497/PIX_OUT pixel_4497/CSA_VREF pixel
Xpixel_3785 pixel_3785/gring pixel_3785/VDD pixel_3785/GND pixel_3785/VREF pixel_3785/ROW_SEL
+ pixel_3785/NB1 pixel_3785/VBIAS pixel_3785/NB2 pixel_3785/AMP_IN pixel_3785/SF_IB
+ pixel_3785/PIX_OUT pixel_3785/CSA_VREF pixel
Xpixel_3774 pixel_3774/gring pixel_3774/VDD pixel_3774/GND pixel_3774/VREF pixel_3774/ROW_SEL
+ pixel_3774/NB1 pixel_3774/VBIAS pixel_3774/NB2 pixel_3774/AMP_IN pixel_3774/SF_IB
+ pixel_3774/PIX_OUT pixel_3774/CSA_VREF pixel
Xpixel_3763 pixel_3763/gring pixel_3763/VDD pixel_3763/GND pixel_3763/VREF pixel_3763/ROW_SEL
+ pixel_3763/NB1 pixel_3763/VBIAS pixel_3763/NB2 pixel_3763/AMP_IN pixel_3763/SF_IB
+ pixel_3763/PIX_OUT pixel_3763/CSA_VREF pixel
Xpixel_3796 pixel_3796/gring pixel_3796/VDD pixel_3796/GND pixel_3796/VREF pixel_3796/ROW_SEL
+ pixel_3796/NB1 pixel_3796/VBIAS pixel_3796/NB2 pixel_3796/AMP_IN pixel_3796/SF_IB
+ pixel_3796/PIX_OUT pixel_3796/CSA_VREF pixel
Xpixel_7090 pixel_7090/gring pixel_7090/VDD pixel_7090/GND pixel_7090/VREF pixel_7090/ROW_SEL
+ pixel_7090/NB1 pixel_7090/VBIAS pixel_7090/NB2 pixel_7090/AMP_IN pixel_7090/SF_IB
+ pixel_7090/PIX_OUT pixel_7090/CSA_VREF pixel
Xpixel_9409 pixel_9409/gring pixel_9409/VDD pixel_9409/GND pixel_9409/VREF pixel_9409/ROW_SEL
+ pixel_9409/NB1 pixel_9409/VBIAS pixel_9409/NB2 pixel_9409/AMP_IN pixel_9409/SF_IB
+ pixel_9409/PIX_OUT pixel_9409/CSA_VREF pixel
Xpixel_8708 pixel_8708/gring pixel_8708/VDD pixel_8708/GND pixel_8708/VREF pixel_8708/ROW_SEL
+ pixel_8708/NB1 pixel_8708/VBIAS pixel_8708/NB2 pixel_8708/AMP_IN pixel_8708/SF_IB
+ pixel_8708/PIX_OUT pixel_8708/CSA_VREF pixel
Xpixel_8719 pixel_8719/gring pixel_8719/VDD pixel_8719/GND pixel_8719/VREF pixel_8719/ROW_SEL
+ pixel_8719/NB1 pixel_8719/VBIAS pixel_8719/NB2 pixel_8719/AMP_IN pixel_8719/SF_IB
+ pixel_8719/PIX_OUT pixel_8719/CSA_VREF pixel
Xpixel_3004 pixel_3004/gring pixel_3004/VDD pixel_3004/GND pixel_3004/VREF pixel_3004/ROW_SEL
+ pixel_3004/NB1 pixel_3004/VBIAS pixel_3004/NB2 pixel_3004/AMP_IN pixel_3004/SF_IB
+ pixel_3004/PIX_OUT pixel_3004/CSA_VREF pixel
Xpixel_2303 pixel_2303/gring pixel_2303/VDD pixel_2303/GND pixel_2303/VREF pixel_2303/ROW_SEL
+ pixel_2303/NB1 pixel_2303/VBIAS pixel_2303/NB2 pixel_2303/AMP_IN pixel_2303/SF_IB
+ pixel_2303/PIX_OUT pixel_2303/CSA_VREF pixel
Xpixel_3048 pixel_3048/gring pixel_3048/VDD pixel_3048/GND pixel_3048/VREF pixel_3048/ROW_SEL
+ pixel_3048/NB1 pixel_3048/VBIAS pixel_3048/NB2 pixel_3048/AMP_IN pixel_3048/SF_IB
+ pixel_3048/PIX_OUT pixel_3048/CSA_VREF pixel
Xpixel_3037 pixel_3037/gring pixel_3037/VDD pixel_3037/GND pixel_3037/VREF pixel_3037/ROW_SEL
+ pixel_3037/NB1 pixel_3037/VBIAS pixel_3037/NB2 pixel_3037/AMP_IN pixel_3037/SF_IB
+ pixel_3037/PIX_OUT pixel_3037/CSA_VREF pixel
Xpixel_3026 pixel_3026/gring pixel_3026/VDD pixel_3026/GND pixel_3026/VREF pixel_3026/ROW_SEL
+ pixel_3026/NB1 pixel_3026/VBIAS pixel_3026/NB2 pixel_3026/AMP_IN pixel_3026/SF_IB
+ pixel_3026/PIX_OUT pixel_3026/CSA_VREF pixel
Xpixel_3015 pixel_3015/gring pixel_3015/VDD pixel_3015/GND pixel_3015/VREF pixel_3015/ROW_SEL
+ pixel_3015/NB1 pixel_3015/VBIAS pixel_3015/NB2 pixel_3015/AMP_IN pixel_3015/SF_IB
+ pixel_3015/PIX_OUT pixel_3015/CSA_VREF pixel
Xpixel_2336 pixel_2336/gring pixel_2336/VDD pixel_2336/GND pixel_2336/VREF pixel_2336/ROW_SEL
+ pixel_2336/NB1 pixel_2336/VBIAS pixel_2336/NB2 pixel_2336/AMP_IN pixel_2336/SF_IB
+ pixel_2336/PIX_OUT pixel_2336/CSA_VREF pixel
Xpixel_2325 pixel_2325/gring pixel_2325/VDD pixel_2325/GND pixel_2325/VREF pixel_2325/ROW_SEL
+ pixel_2325/NB1 pixel_2325/VBIAS pixel_2325/NB2 pixel_2325/AMP_IN pixel_2325/SF_IB
+ pixel_2325/PIX_OUT pixel_2325/CSA_VREF pixel
Xpixel_2314 pixel_2314/gring pixel_2314/VDD pixel_2314/GND pixel_2314/VREF pixel_2314/ROW_SEL
+ pixel_2314/NB1 pixel_2314/VBIAS pixel_2314/NB2 pixel_2314/AMP_IN pixel_2314/SF_IB
+ pixel_2314/PIX_OUT pixel_2314/CSA_VREF pixel
Xpixel_3059 pixel_3059/gring pixel_3059/VDD pixel_3059/GND pixel_3059/VREF pixel_3059/ROW_SEL
+ pixel_3059/NB1 pixel_3059/VBIAS pixel_3059/NB2 pixel_3059/AMP_IN pixel_3059/SF_IB
+ pixel_3059/PIX_OUT pixel_3059/CSA_VREF pixel
Xpixel_1624 pixel_1624/gring pixel_1624/VDD pixel_1624/GND pixel_1624/VREF pixel_1624/ROW_SEL
+ pixel_1624/NB1 pixel_1624/VBIAS pixel_1624/NB2 pixel_1624/AMP_IN pixel_1624/SF_IB
+ pixel_1624/PIX_OUT pixel_1624/CSA_VREF pixel
Xpixel_1613 pixel_1613/gring pixel_1613/VDD pixel_1613/GND pixel_1613/VREF pixel_1613/ROW_SEL
+ pixel_1613/NB1 pixel_1613/VBIAS pixel_1613/NB2 pixel_1613/AMP_IN pixel_1613/SF_IB
+ pixel_1613/PIX_OUT pixel_1613/CSA_VREF pixel
Xpixel_1602 pixel_1602/gring pixel_1602/VDD pixel_1602/GND pixel_1602/VREF pixel_1602/ROW_SEL
+ pixel_1602/NB1 pixel_1602/VBIAS pixel_1602/NB2 pixel_1602/AMP_IN pixel_1602/SF_IB
+ pixel_1602/PIX_OUT pixel_1602/CSA_VREF pixel
Xpixel_2369 pixel_2369/gring pixel_2369/VDD pixel_2369/GND pixel_2369/VREF pixel_2369/ROW_SEL
+ pixel_2369/NB1 pixel_2369/VBIAS pixel_2369/NB2 pixel_2369/AMP_IN pixel_2369/SF_IB
+ pixel_2369/PIX_OUT pixel_2369/CSA_VREF pixel
Xpixel_2358 pixel_2358/gring pixel_2358/VDD pixel_2358/GND pixel_2358/VREF pixel_2358/ROW_SEL
+ pixel_2358/NB1 pixel_2358/VBIAS pixel_2358/NB2 pixel_2358/AMP_IN pixel_2358/SF_IB
+ pixel_2358/PIX_OUT pixel_2358/CSA_VREF pixel
Xpixel_2347 pixel_2347/gring pixel_2347/VDD pixel_2347/GND pixel_2347/VREF pixel_2347/ROW_SEL
+ pixel_2347/NB1 pixel_2347/VBIAS pixel_2347/NB2 pixel_2347/AMP_IN pixel_2347/SF_IB
+ pixel_2347/PIX_OUT pixel_2347/CSA_VREF pixel
Xpixel_1668 pixel_1668/gring pixel_1668/VDD pixel_1668/GND pixel_1668/VREF pixel_1668/ROW_SEL
+ pixel_1668/NB1 pixel_1668/VBIAS pixel_1668/NB2 pixel_1668/AMP_IN pixel_1668/SF_IB
+ pixel_1668/PIX_OUT pixel_1668/CSA_VREF pixel
Xpixel_1657 pixel_1657/gring pixel_1657/VDD pixel_1657/GND pixel_1657/VREF pixel_1657/ROW_SEL
+ pixel_1657/NB1 pixel_1657/VBIAS pixel_1657/NB2 pixel_1657/AMP_IN pixel_1657/SF_IB
+ pixel_1657/PIX_OUT pixel_1657/CSA_VREF pixel
Xpixel_1646 pixel_1646/gring pixel_1646/VDD pixel_1646/GND pixel_1646/VREF pixel_1646/ROW_SEL
+ pixel_1646/NB1 pixel_1646/VBIAS pixel_1646/NB2 pixel_1646/AMP_IN pixel_1646/SF_IB
+ pixel_1646/PIX_OUT pixel_1646/CSA_VREF pixel
Xpixel_1635 pixel_1635/gring pixel_1635/VDD pixel_1635/GND pixel_1635/VREF pixel_1635/ROW_SEL
+ pixel_1635/NB1 pixel_1635/VBIAS pixel_1635/NB2 pixel_1635/AMP_IN pixel_1635/SF_IB
+ pixel_1635/PIX_OUT pixel_1635/CSA_VREF pixel
Xpixel_1679 pixel_1679/gring pixel_1679/VDD pixel_1679/GND pixel_1679/VREF pixel_1679/ROW_SEL
+ pixel_1679/NB1 pixel_1679/VBIAS pixel_1679/NB2 pixel_1679/AMP_IN pixel_1679/SF_IB
+ pixel_1679/PIX_OUT pixel_1679/CSA_VREF pixel
Xpixel_9932 pixel_9932/gring pixel_9932/VDD pixel_9932/GND pixel_9932/VREF pixel_9932/ROW_SEL
+ pixel_9932/NB1 pixel_9932/VBIAS pixel_9932/NB2 pixel_9932/AMP_IN pixel_9932/SF_IB
+ pixel_9932/PIX_OUT pixel_9932/CSA_VREF pixel
Xpixel_9921 pixel_9921/gring pixel_9921/VDD pixel_9921/GND pixel_9921/VREF pixel_9921/ROW_SEL
+ pixel_9921/NB1 pixel_9921/VBIAS pixel_9921/NB2 pixel_9921/AMP_IN pixel_9921/SF_IB
+ pixel_9921/PIX_OUT pixel_9921/CSA_VREF pixel
Xpixel_9910 pixel_9910/gring pixel_9910/VDD pixel_9910/GND pixel_9910/VREF pixel_9910/ROW_SEL
+ pixel_9910/NB1 pixel_9910/VBIAS pixel_9910/NB2 pixel_9910/AMP_IN pixel_9910/SF_IB
+ pixel_9910/PIX_OUT pixel_9910/CSA_VREF pixel
Xpixel_9943 pixel_9943/gring pixel_9943/VDD pixel_9943/GND pixel_9943/VREF pixel_9943/ROW_SEL
+ pixel_9943/NB1 pixel_9943/VBIAS pixel_9943/NB2 pixel_9943/AMP_IN pixel_9943/SF_IB
+ pixel_9943/PIX_OUT pixel_9943/CSA_VREF pixel
Xpixel_9954 pixel_9954/gring pixel_9954/VDD pixel_9954/GND pixel_9954/VREF pixel_9954/ROW_SEL
+ pixel_9954/NB1 pixel_9954/VBIAS pixel_9954/NB2 pixel_9954/AMP_IN pixel_9954/SF_IB
+ pixel_9954/PIX_OUT pixel_9954/CSA_VREF pixel
Xpixel_9965 pixel_9965/gring pixel_9965/VDD pixel_9965/GND pixel_9965/VREF pixel_9965/ROW_SEL
+ pixel_9965/NB1 pixel_9965/VBIAS pixel_9965/NB2 pixel_9965/AMP_IN pixel_9965/SF_IB
+ pixel_9965/PIX_OUT pixel_9965/CSA_VREF pixel
Xpixel_9976 pixel_9976/gring pixel_9976/VDD pixel_9976/GND pixel_9976/VREF pixel_9976/ROW_SEL
+ pixel_9976/NB1 pixel_9976/VBIAS pixel_9976/NB2 pixel_9976/AMP_IN pixel_9976/SF_IB
+ pixel_9976/PIX_OUT pixel_9976/CSA_VREF pixel
Xpixel_9987 pixel_9987/gring pixel_9987/VDD pixel_9987/GND pixel_9987/VREF pixel_9987/ROW_SEL
+ pixel_9987/NB1 pixel_9987/VBIAS pixel_9987/NB2 pixel_9987/AMP_IN pixel_9987/SF_IB
+ pixel_9987/PIX_OUT pixel_9987/CSA_VREF pixel
Xpixel_9998 pixel_9998/gring pixel_9998/VDD pixel_9998/GND pixel_9998/VREF pixel_9998/ROW_SEL
+ pixel_9998/NB1 pixel_9998/VBIAS pixel_9998/NB2 pixel_9998/AMP_IN pixel_9998/SF_IB
+ pixel_9998/PIX_OUT pixel_9998/CSA_VREF pixel
Xpixel_4250 pixel_4250/gring pixel_4250/VDD pixel_4250/GND pixel_4250/VREF pixel_4250/ROW_SEL
+ pixel_4250/NB1 pixel_4250/VBIAS pixel_4250/NB2 pixel_4250/AMP_IN pixel_4250/SF_IB
+ pixel_4250/PIX_OUT pixel_4250/CSA_VREF pixel
Xpixel_4261 pixel_4261/gring pixel_4261/VDD pixel_4261/GND pixel_4261/VREF pixel_4261/ROW_SEL
+ pixel_4261/NB1 pixel_4261/VBIAS pixel_4261/NB2 pixel_4261/AMP_IN pixel_4261/SF_IB
+ pixel_4261/PIX_OUT pixel_4261/CSA_VREF pixel
Xpixel_4272 pixel_4272/gring pixel_4272/VDD pixel_4272/GND pixel_4272/VREF pixel_4272/ROW_SEL
+ pixel_4272/NB1 pixel_4272/VBIAS pixel_4272/NB2 pixel_4272/AMP_IN pixel_4272/SF_IB
+ pixel_4272/PIX_OUT pixel_4272/CSA_VREF pixel
Xpixel_3560 pixel_3560/gring pixel_3560/VDD pixel_3560/GND pixel_3560/VREF pixel_3560/ROW_SEL
+ pixel_3560/NB1 pixel_3560/VBIAS pixel_3560/NB2 pixel_3560/AMP_IN pixel_3560/SF_IB
+ pixel_3560/PIX_OUT pixel_3560/CSA_VREF pixel
Xpixel_4283 pixel_4283/gring pixel_4283/VDD pixel_4283/GND pixel_4283/VREF pixel_4283/ROW_SEL
+ pixel_4283/NB1 pixel_4283/VBIAS pixel_4283/NB2 pixel_4283/AMP_IN pixel_4283/SF_IB
+ pixel_4283/PIX_OUT pixel_4283/CSA_VREF pixel
Xpixel_4294 pixel_4294/gring pixel_4294/VDD pixel_4294/GND pixel_4294/VREF pixel_4294/ROW_SEL
+ pixel_4294/NB1 pixel_4294/VBIAS pixel_4294/NB2 pixel_4294/AMP_IN pixel_4294/SF_IB
+ pixel_4294/PIX_OUT pixel_4294/CSA_VREF pixel
Xpixel_3593 pixel_3593/gring pixel_3593/VDD pixel_3593/GND pixel_3593/VREF pixel_3593/ROW_SEL
+ pixel_3593/NB1 pixel_3593/VBIAS pixel_3593/NB2 pixel_3593/AMP_IN pixel_3593/SF_IB
+ pixel_3593/PIX_OUT pixel_3593/CSA_VREF pixel
Xpixel_3582 pixel_3582/gring pixel_3582/VDD pixel_3582/GND pixel_3582/VREF pixel_3582/ROW_SEL
+ pixel_3582/NB1 pixel_3582/VBIAS pixel_3582/NB2 pixel_3582/AMP_IN pixel_3582/SF_IB
+ pixel_3582/PIX_OUT pixel_3582/CSA_VREF pixel
Xpixel_3571 pixel_3571/gring pixel_3571/VDD pixel_3571/GND pixel_3571/VREF pixel_3571/ROW_SEL
+ pixel_3571/NB1 pixel_3571/VBIAS pixel_3571/NB2 pixel_3571/AMP_IN pixel_3571/SF_IB
+ pixel_3571/PIX_OUT pixel_3571/CSA_VREF pixel
Xpixel_2892 pixel_2892/gring pixel_2892/VDD pixel_2892/GND pixel_2892/VREF pixel_2892/ROW_SEL
+ pixel_2892/NB1 pixel_2892/VBIAS pixel_2892/NB2 pixel_2892/AMP_IN pixel_2892/SF_IB
+ pixel_2892/PIX_OUT pixel_2892/CSA_VREF pixel
Xpixel_2881 pixel_2881/gring pixel_2881/VDD pixel_2881/GND pixel_2881/VREF pixel_2881/ROW_SEL
+ pixel_2881/NB1 pixel_2881/VBIAS pixel_2881/NB2 pixel_2881/AMP_IN pixel_2881/SF_IB
+ pixel_2881/PIX_OUT pixel_2881/CSA_VREF pixel
Xpixel_2870 pixel_2870/gring pixel_2870/VDD pixel_2870/GND pixel_2870/VREF pixel_2870/ROW_SEL
+ pixel_2870/NB1 pixel_2870/VBIAS pixel_2870/NB2 pixel_2870/AMP_IN pixel_2870/SF_IB
+ pixel_2870/PIX_OUT pixel_2870/CSA_VREF pixel
Xpixel_9228 pixel_9228/gring pixel_9228/VDD pixel_9228/GND pixel_9228/VREF pixel_9228/ROW_SEL
+ pixel_9228/NB1 pixel_9228/VBIAS pixel_9228/NB2 pixel_9228/AMP_IN pixel_9228/SF_IB
+ pixel_9228/PIX_OUT pixel_9228/CSA_VREF pixel
Xpixel_9217 pixel_9217/gring pixel_9217/VDD pixel_9217/GND pixel_9217/VREF pixel_9217/ROW_SEL
+ pixel_9217/NB1 pixel_9217/VBIAS pixel_9217/NB2 pixel_9217/AMP_IN pixel_9217/SF_IB
+ pixel_9217/PIX_OUT pixel_9217/CSA_VREF pixel
Xpixel_9206 pixel_9206/gring pixel_9206/VDD pixel_9206/GND pixel_9206/VREF pixel_9206/ROW_SEL
+ pixel_9206/NB1 pixel_9206/VBIAS pixel_9206/NB2 pixel_9206/AMP_IN pixel_9206/SF_IB
+ pixel_9206/PIX_OUT pixel_9206/CSA_VREF pixel
Xpixel_8527 pixel_8527/gring pixel_8527/VDD pixel_8527/GND pixel_8527/VREF pixel_8527/ROW_SEL
+ pixel_8527/NB1 pixel_8527/VBIAS pixel_8527/NB2 pixel_8527/AMP_IN pixel_8527/SF_IB
+ pixel_8527/PIX_OUT pixel_8527/CSA_VREF pixel
Xpixel_8516 pixel_8516/gring pixel_8516/VDD pixel_8516/GND pixel_8516/VREF pixel_8516/ROW_SEL
+ pixel_8516/NB1 pixel_8516/VBIAS pixel_8516/NB2 pixel_8516/AMP_IN pixel_8516/SF_IB
+ pixel_8516/PIX_OUT pixel_8516/CSA_VREF pixel
Xpixel_8505 pixel_8505/gring pixel_8505/VDD pixel_8505/GND pixel_8505/VREF pixel_8505/ROW_SEL
+ pixel_8505/NB1 pixel_8505/VBIAS pixel_8505/NB2 pixel_8505/AMP_IN pixel_8505/SF_IB
+ pixel_8505/PIX_OUT pixel_8505/CSA_VREF pixel
Xpixel_9239 pixel_9239/gring pixel_9239/VDD pixel_9239/GND pixel_9239/VREF pixel_9239/ROW_SEL
+ pixel_9239/NB1 pixel_9239/VBIAS pixel_9239/NB2 pixel_9239/AMP_IN pixel_9239/SF_IB
+ pixel_9239/PIX_OUT pixel_9239/CSA_VREF pixel
Xpixel_8549 pixel_8549/gring pixel_8549/VDD pixel_8549/GND pixel_8549/VREF pixel_8549/ROW_SEL
+ pixel_8549/NB1 pixel_8549/VBIAS pixel_8549/NB2 pixel_8549/AMP_IN pixel_8549/SF_IB
+ pixel_8549/PIX_OUT pixel_8549/CSA_VREF pixel
Xpixel_8538 pixel_8538/gring pixel_8538/VDD pixel_8538/GND pixel_8538/VREF pixel_8538/ROW_SEL
+ pixel_8538/NB1 pixel_8538/VBIAS pixel_8538/NB2 pixel_8538/AMP_IN pixel_8538/SF_IB
+ pixel_8538/PIX_OUT pixel_8538/CSA_VREF pixel
Xpixel_7804 pixel_7804/gring pixel_7804/VDD pixel_7804/GND pixel_7804/VREF pixel_7804/ROW_SEL
+ pixel_7804/NB1 pixel_7804/VBIAS pixel_7804/NB2 pixel_7804/AMP_IN pixel_7804/SF_IB
+ pixel_7804/PIX_OUT pixel_7804/CSA_VREF pixel
Xpixel_7815 pixel_7815/gring pixel_7815/VDD pixel_7815/GND pixel_7815/VREF pixel_7815/ROW_SEL
+ pixel_7815/NB1 pixel_7815/VBIAS pixel_7815/NB2 pixel_7815/AMP_IN pixel_7815/SF_IB
+ pixel_7815/PIX_OUT pixel_7815/CSA_VREF pixel
Xpixel_7826 pixel_7826/gring pixel_7826/VDD pixel_7826/GND pixel_7826/VREF pixel_7826/ROW_SEL
+ pixel_7826/NB1 pixel_7826/VBIAS pixel_7826/NB2 pixel_7826/AMP_IN pixel_7826/SF_IB
+ pixel_7826/PIX_OUT pixel_7826/CSA_VREF pixel
Xpixel_7837 pixel_7837/gring pixel_7837/VDD pixel_7837/GND pixel_7837/VREF pixel_7837/ROW_SEL
+ pixel_7837/NB1 pixel_7837/VBIAS pixel_7837/NB2 pixel_7837/AMP_IN pixel_7837/SF_IB
+ pixel_7837/PIX_OUT pixel_7837/CSA_VREF pixel
Xpixel_7848 pixel_7848/gring pixel_7848/VDD pixel_7848/GND pixel_7848/VREF pixel_7848/ROW_SEL
+ pixel_7848/NB1 pixel_7848/VBIAS pixel_7848/NB2 pixel_7848/AMP_IN pixel_7848/SF_IB
+ pixel_7848/PIX_OUT pixel_7848/CSA_VREF pixel
Xpixel_7859 pixel_7859/gring pixel_7859/VDD pixel_7859/GND pixel_7859/VREF pixel_7859/ROW_SEL
+ pixel_7859/NB1 pixel_7859/VBIAS pixel_7859/NB2 pixel_7859/AMP_IN pixel_7859/SF_IB
+ pixel_7859/PIX_OUT pixel_7859/CSA_VREF pixel
Xpixel_2111 pixel_2111/gring pixel_2111/VDD pixel_2111/GND pixel_2111/VREF pixel_2111/ROW_SEL
+ pixel_2111/NB1 pixel_2111/VBIAS pixel_2111/NB2 pixel_2111/AMP_IN pixel_2111/SF_IB
+ pixel_2111/PIX_OUT pixel_2111/CSA_VREF pixel
Xpixel_2100 pixel_2100/gring pixel_2100/VDD pixel_2100/GND pixel_2100/VREF pixel_2100/ROW_SEL
+ pixel_2100/NB1 pixel_2100/VBIAS pixel_2100/NB2 pixel_2100/AMP_IN pixel_2100/SF_IB
+ pixel_2100/PIX_OUT pixel_2100/CSA_VREF pixel
Xpixel_2144 pixel_2144/gring pixel_2144/VDD pixel_2144/GND pixel_2144/VREF pixel_2144/ROW_SEL
+ pixel_2144/NB1 pixel_2144/VBIAS pixel_2144/NB2 pixel_2144/AMP_IN pixel_2144/SF_IB
+ pixel_2144/PIX_OUT pixel_2144/CSA_VREF pixel
Xpixel_2133 pixel_2133/gring pixel_2133/VDD pixel_2133/GND pixel_2133/VREF pixel_2133/ROW_SEL
+ pixel_2133/NB1 pixel_2133/VBIAS pixel_2133/NB2 pixel_2133/AMP_IN pixel_2133/SF_IB
+ pixel_2133/PIX_OUT pixel_2133/CSA_VREF pixel
Xpixel_2122 pixel_2122/gring pixel_2122/VDD pixel_2122/GND pixel_2122/VREF pixel_2122/ROW_SEL
+ pixel_2122/NB1 pixel_2122/VBIAS pixel_2122/NB2 pixel_2122/AMP_IN pixel_2122/SF_IB
+ pixel_2122/PIX_OUT pixel_2122/CSA_VREF pixel
Xpixel_1443 pixel_1443/gring pixel_1443/VDD pixel_1443/GND pixel_1443/VREF pixel_1443/ROW_SEL
+ pixel_1443/NB1 pixel_1443/VBIAS pixel_1443/NB2 pixel_1443/AMP_IN pixel_1443/SF_IB
+ pixel_1443/PIX_OUT pixel_1443/CSA_VREF pixel
Xpixel_1432 pixel_1432/gring pixel_1432/VDD pixel_1432/GND pixel_1432/VREF pixel_1432/ROW_SEL
+ pixel_1432/NB1 pixel_1432/VBIAS pixel_1432/NB2 pixel_1432/AMP_IN pixel_1432/SF_IB
+ pixel_1432/PIX_OUT pixel_1432/CSA_VREF pixel
Xpixel_1421 pixel_1421/gring pixel_1421/VDD pixel_1421/GND pixel_1421/VREF pixel_1421/ROW_SEL
+ pixel_1421/NB1 pixel_1421/VBIAS pixel_1421/NB2 pixel_1421/AMP_IN pixel_1421/SF_IB
+ pixel_1421/PIX_OUT pixel_1421/CSA_VREF pixel
Xpixel_1410 pixel_1410/gring pixel_1410/VDD pixel_1410/GND pixel_1410/VREF pixel_1410/ROW_SEL
+ pixel_1410/NB1 pixel_1410/VBIAS pixel_1410/NB2 pixel_1410/AMP_IN pixel_1410/SF_IB
+ pixel_1410/PIX_OUT pixel_1410/CSA_VREF pixel
Xpixel_2177 pixel_2177/gring pixel_2177/VDD pixel_2177/GND pixel_2177/VREF pixel_2177/ROW_SEL
+ pixel_2177/NB1 pixel_2177/VBIAS pixel_2177/NB2 pixel_2177/AMP_IN pixel_2177/SF_IB
+ pixel_2177/PIX_OUT pixel_2177/CSA_VREF pixel
Xpixel_2166 pixel_2166/gring pixel_2166/VDD pixel_2166/GND pixel_2166/VREF pixel_2166/ROW_SEL
+ pixel_2166/NB1 pixel_2166/VBIAS pixel_2166/NB2 pixel_2166/AMP_IN pixel_2166/SF_IB
+ pixel_2166/PIX_OUT pixel_2166/CSA_VREF pixel
Xpixel_2155 pixel_2155/gring pixel_2155/VDD pixel_2155/GND pixel_2155/VREF pixel_2155/ROW_SEL
+ pixel_2155/NB1 pixel_2155/VBIAS pixel_2155/NB2 pixel_2155/AMP_IN pixel_2155/SF_IB
+ pixel_2155/PIX_OUT pixel_2155/CSA_VREF pixel
Xpixel_1476 pixel_1476/gring pixel_1476/VDD pixel_1476/GND pixel_1476/VREF pixel_1476/ROW_SEL
+ pixel_1476/NB1 pixel_1476/VBIAS pixel_1476/NB2 pixel_1476/AMP_IN pixel_1476/SF_IB
+ pixel_1476/PIX_OUT pixel_1476/CSA_VREF pixel
Xpixel_1465 pixel_1465/gring pixel_1465/VDD pixel_1465/GND pixel_1465/VREF pixel_1465/ROW_SEL
+ pixel_1465/NB1 pixel_1465/VBIAS pixel_1465/NB2 pixel_1465/AMP_IN pixel_1465/SF_IB
+ pixel_1465/PIX_OUT pixel_1465/CSA_VREF pixel
Xpixel_1454 pixel_1454/gring pixel_1454/VDD pixel_1454/GND pixel_1454/VREF pixel_1454/ROW_SEL
+ pixel_1454/NB1 pixel_1454/VBIAS pixel_1454/NB2 pixel_1454/AMP_IN pixel_1454/SF_IB
+ pixel_1454/PIX_OUT pixel_1454/CSA_VREF pixel
Xpixel_2199 pixel_2199/gring pixel_2199/VDD pixel_2199/GND pixel_2199/VREF pixel_2199/ROW_SEL
+ pixel_2199/NB1 pixel_2199/VBIAS pixel_2199/NB2 pixel_2199/AMP_IN pixel_2199/SF_IB
+ pixel_2199/PIX_OUT pixel_2199/CSA_VREF pixel
Xpixel_2188 pixel_2188/gring pixel_2188/VDD pixel_2188/GND pixel_2188/VREF pixel_2188/ROW_SEL
+ pixel_2188/NB1 pixel_2188/VBIAS pixel_2188/NB2 pixel_2188/AMP_IN pixel_2188/SF_IB
+ pixel_2188/PIX_OUT pixel_2188/CSA_VREF pixel
Xpixel_1498 pixel_1498/gring pixel_1498/VDD pixel_1498/GND pixel_1498/VREF pixel_1498/ROW_SEL
+ pixel_1498/NB1 pixel_1498/VBIAS pixel_1498/NB2 pixel_1498/AMP_IN pixel_1498/SF_IB
+ pixel_1498/PIX_OUT pixel_1498/CSA_VREF pixel
Xpixel_1487 pixel_1487/gring pixel_1487/VDD pixel_1487/GND pixel_1487/VREF pixel_1487/ROW_SEL
+ pixel_1487/NB1 pixel_1487/VBIAS pixel_1487/NB2 pixel_1487/AMP_IN pixel_1487/SF_IB
+ pixel_1487/PIX_OUT pixel_1487/CSA_VREF pixel
Xpixel_9740 pixel_9740/gring pixel_9740/VDD pixel_9740/GND pixel_9740/VREF pixel_9740/ROW_SEL
+ pixel_9740/NB1 pixel_9740/VBIAS pixel_9740/NB2 pixel_9740/AMP_IN pixel_9740/SF_IB
+ pixel_9740/PIX_OUT pixel_9740/CSA_VREF pixel
Xpixel_9751 pixel_9751/gring pixel_9751/VDD pixel_9751/GND pixel_9751/VREF pixel_9751/ROW_SEL
+ pixel_9751/NB1 pixel_9751/VBIAS pixel_9751/NB2 pixel_9751/AMP_IN pixel_9751/SF_IB
+ pixel_9751/PIX_OUT pixel_9751/CSA_VREF pixel
Xpixel_9762 pixel_9762/gring pixel_9762/VDD pixel_9762/GND pixel_9762/VREF pixel_9762/ROW_SEL
+ pixel_9762/NB1 pixel_9762/VBIAS pixel_9762/NB2 pixel_9762/AMP_IN pixel_9762/SF_IB
+ pixel_9762/PIX_OUT pixel_9762/CSA_VREF pixel
Xpixel_9773 pixel_9773/gring pixel_9773/VDD pixel_9773/GND pixel_9773/VREF pixel_9773/ROW_SEL
+ pixel_9773/NB1 pixel_9773/VBIAS pixel_9773/NB2 pixel_9773/AMP_IN pixel_9773/SF_IB
+ pixel_9773/PIX_OUT pixel_9773/CSA_VREF pixel
Xpixel_9784 pixel_9784/gring pixel_9784/VDD pixel_9784/GND pixel_9784/VREF pixel_9784/ROW_SEL
+ pixel_9784/NB1 pixel_9784/VBIAS pixel_9784/NB2 pixel_9784/AMP_IN pixel_9784/SF_IB
+ pixel_9784/PIX_OUT pixel_9784/CSA_VREF pixel
Xpixel_9795 pixel_9795/gring pixel_9795/VDD pixel_9795/GND pixel_9795/VREF pixel_9795/ROW_SEL
+ pixel_9795/NB1 pixel_9795/VBIAS pixel_9795/NB2 pixel_9795/AMP_IN pixel_9795/SF_IB
+ pixel_9795/PIX_OUT pixel_9795/CSA_VREF pixel
Xpixel_4080 pixel_4080/gring pixel_4080/VDD pixel_4080/GND pixel_4080/VREF pixel_4080/ROW_SEL
+ pixel_4080/NB1 pixel_4080/VBIAS pixel_4080/NB2 pixel_4080/AMP_IN pixel_4080/SF_IB
+ pixel_4080/PIX_OUT pixel_4080/CSA_VREF pixel
Xpixel_4091 pixel_4091/gring pixel_4091/VDD pixel_4091/GND pixel_4091/VREF pixel_4091/ROW_SEL
+ pixel_4091/NB1 pixel_4091/VBIAS pixel_4091/NB2 pixel_4091/AMP_IN pixel_4091/SF_IB
+ pixel_4091/PIX_OUT pixel_4091/CSA_VREF pixel
Xpixel_3390 pixel_3390/gring pixel_3390/VDD pixel_3390/GND pixel_3390/VREF pixel_3390/ROW_SEL
+ pixel_3390/NB1 pixel_3390/VBIAS pixel_3390/NB2 pixel_3390/AMP_IN pixel_3390/SF_IB
+ pixel_3390/PIX_OUT pixel_3390/CSA_VREF pixel
Xpixel_5709 pixel_5709/gring pixel_5709/VDD pixel_5709/GND pixel_5709/VREF pixel_5709/ROW_SEL
+ pixel_5709/NB1 pixel_5709/VBIAS pixel_5709/NB2 pixel_5709/AMP_IN pixel_5709/SF_IB
+ pixel_5709/PIX_OUT pixel_5709/CSA_VREF pixel
Xpixel_9003 pixel_9003/gring pixel_9003/VDD pixel_9003/GND pixel_9003/VREF pixel_9003/ROW_SEL
+ pixel_9003/NB1 pixel_9003/VBIAS pixel_9003/NB2 pixel_9003/AMP_IN pixel_9003/SF_IB
+ pixel_9003/PIX_OUT pixel_9003/CSA_VREF pixel
Xpixel_9036 pixel_9036/gring pixel_9036/VDD pixel_9036/GND pixel_9036/VREF pixel_9036/ROW_SEL
+ pixel_9036/NB1 pixel_9036/VBIAS pixel_9036/NB2 pixel_9036/AMP_IN pixel_9036/SF_IB
+ pixel_9036/PIX_OUT pixel_9036/CSA_VREF pixel
Xpixel_9025 pixel_9025/gring pixel_9025/VDD pixel_9025/GND pixel_9025/VREF pixel_9025/ROW_SEL
+ pixel_9025/NB1 pixel_9025/VBIAS pixel_9025/NB2 pixel_9025/AMP_IN pixel_9025/SF_IB
+ pixel_9025/PIX_OUT pixel_9025/CSA_VREF pixel
Xpixel_9014 pixel_9014/gring pixel_9014/VDD pixel_9014/GND pixel_9014/VREF pixel_9014/ROW_SEL
+ pixel_9014/NB1 pixel_9014/VBIAS pixel_9014/NB2 pixel_9014/AMP_IN pixel_9014/SF_IB
+ pixel_9014/PIX_OUT pixel_9014/CSA_VREF pixel
Xpixel_9069 pixel_9069/gring pixel_9069/VDD pixel_9069/GND pixel_9069/VREF pixel_9069/ROW_SEL
+ pixel_9069/NB1 pixel_9069/VBIAS pixel_9069/NB2 pixel_9069/AMP_IN pixel_9069/SF_IB
+ pixel_9069/PIX_OUT pixel_9069/CSA_VREF pixel
Xpixel_9058 pixel_9058/gring pixel_9058/VDD pixel_9058/GND pixel_9058/VREF pixel_9058/ROW_SEL
+ pixel_9058/NB1 pixel_9058/VBIAS pixel_9058/NB2 pixel_9058/AMP_IN pixel_9058/SF_IB
+ pixel_9058/PIX_OUT pixel_9058/CSA_VREF pixel
Xpixel_9047 pixel_9047/gring pixel_9047/VDD pixel_9047/GND pixel_9047/VREF pixel_9047/ROW_SEL
+ pixel_9047/NB1 pixel_9047/VBIAS pixel_9047/NB2 pixel_9047/AMP_IN pixel_9047/SF_IB
+ pixel_9047/PIX_OUT pixel_9047/CSA_VREF pixel
Xpixel_8302 pixel_8302/gring pixel_8302/VDD pixel_8302/GND pixel_8302/VREF pixel_8302/ROW_SEL
+ pixel_8302/NB1 pixel_8302/VBIAS pixel_8302/NB2 pixel_8302/AMP_IN pixel_8302/SF_IB
+ pixel_8302/PIX_OUT pixel_8302/CSA_VREF pixel
Xpixel_8313 pixel_8313/gring pixel_8313/VDD pixel_8313/GND pixel_8313/VREF pixel_8313/ROW_SEL
+ pixel_8313/NB1 pixel_8313/VBIAS pixel_8313/NB2 pixel_8313/AMP_IN pixel_8313/SF_IB
+ pixel_8313/PIX_OUT pixel_8313/CSA_VREF pixel
Xpixel_8324 pixel_8324/gring pixel_8324/VDD pixel_8324/GND pixel_8324/VREF pixel_8324/ROW_SEL
+ pixel_8324/NB1 pixel_8324/VBIAS pixel_8324/NB2 pixel_8324/AMP_IN pixel_8324/SF_IB
+ pixel_8324/PIX_OUT pixel_8324/CSA_VREF pixel
Xpixel_8335 pixel_8335/gring pixel_8335/VDD pixel_8335/GND pixel_8335/VREF pixel_8335/ROW_SEL
+ pixel_8335/NB1 pixel_8335/VBIAS pixel_8335/NB2 pixel_8335/AMP_IN pixel_8335/SF_IB
+ pixel_8335/PIX_OUT pixel_8335/CSA_VREF pixel
Xpixel_8346 pixel_8346/gring pixel_8346/VDD pixel_8346/GND pixel_8346/VREF pixel_8346/ROW_SEL
+ pixel_8346/NB1 pixel_8346/VBIAS pixel_8346/NB2 pixel_8346/AMP_IN pixel_8346/SF_IB
+ pixel_8346/PIX_OUT pixel_8346/CSA_VREF pixel
Xpixel_8357 pixel_8357/gring pixel_8357/VDD pixel_8357/GND pixel_8357/VREF pixel_8357/ROW_SEL
+ pixel_8357/NB1 pixel_8357/VBIAS pixel_8357/NB2 pixel_8357/AMP_IN pixel_8357/SF_IB
+ pixel_8357/PIX_OUT pixel_8357/CSA_VREF pixel
Xpixel_8368 pixel_8368/gring pixel_8368/VDD pixel_8368/GND pixel_8368/VREF pixel_8368/ROW_SEL
+ pixel_8368/NB1 pixel_8368/VBIAS pixel_8368/NB2 pixel_8368/AMP_IN pixel_8368/SF_IB
+ pixel_8368/PIX_OUT pixel_8368/CSA_VREF pixel
Xpixel_7601 pixel_7601/gring pixel_7601/VDD pixel_7601/GND pixel_7601/VREF pixel_7601/ROW_SEL
+ pixel_7601/NB1 pixel_7601/VBIAS pixel_7601/NB2 pixel_7601/AMP_IN pixel_7601/SF_IB
+ pixel_7601/PIX_OUT pixel_7601/CSA_VREF pixel
Xpixel_7612 pixel_7612/gring pixel_7612/VDD pixel_7612/GND pixel_7612/VREF pixel_7612/ROW_SEL
+ pixel_7612/NB1 pixel_7612/VBIAS pixel_7612/NB2 pixel_7612/AMP_IN pixel_7612/SF_IB
+ pixel_7612/PIX_OUT pixel_7612/CSA_VREF pixel
Xpixel_7623 pixel_7623/gring pixel_7623/VDD pixel_7623/GND pixel_7623/VREF pixel_7623/ROW_SEL
+ pixel_7623/NB1 pixel_7623/VBIAS pixel_7623/NB2 pixel_7623/AMP_IN pixel_7623/SF_IB
+ pixel_7623/PIX_OUT pixel_7623/CSA_VREF pixel
Xpixel_8379 pixel_8379/gring pixel_8379/VDD pixel_8379/GND pixel_8379/VREF pixel_8379/ROW_SEL
+ pixel_8379/NB1 pixel_8379/VBIAS pixel_8379/NB2 pixel_8379/AMP_IN pixel_8379/SF_IB
+ pixel_8379/PIX_OUT pixel_8379/CSA_VREF pixel
Xpixel_7634 pixel_7634/gring pixel_7634/VDD pixel_7634/GND pixel_7634/VREF pixel_7634/ROW_SEL
+ pixel_7634/NB1 pixel_7634/VBIAS pixel_7634/NB2 pixel_7634/AMP_IN pixel_7634/SF_IB
+ pixel_7634/PIX_OUT pixel_7634/CSA_VREF pixel
Xpixel_7645 pixel_7645/gring pixel_7645/VDD pixel_7645/GND pixel_7645/VREF pixel_7645/ROW_SEL
+ pixel_7645/NB1 pixel_7645/VBIAS pixel_7645/NB2 pixel_7645/AMP_IN pixel_7645/SF_IB
+ pixel_7645/PIX_OUT pixel_7645/CSA_VREF pixel
Xpixel_7656 pixel_7656/gring pixel_7656/VDD pixel_7656/GND pixel_7656/VREF pixel_7656/ROW_SEL
+ pixel_7656/NB1 pixel_7656/VBIAS pixel_7656/NB2 pixel_7656/AMP_IN pixel_7656/SF_IB
+ pixel_7656/PIX_OUT pixel_7656/CSA_VREF pixel
Xpixel_6900 pixel_6900/gring pixel_6900/VDD pixel_6900/GND pixel_6900/VREF pixel_6900/ROW_SEL
+ pixel_6900/NB1 pixel_6900/VBIAS pixel_6900/NB2 pixel_6900/AMP_IN pixel_6900/SF_IB
+ pixel_6900/PIX_OUT pixel_6900/CSA_VREF pixel
Xpixel_6911 pixel_6911/gring pixel_6911/VDD pixel_6911/GND pixel_6911/VREF pixel_6911/ROW_SEL
+ pixel_6911/NB1 pixel_6911/VBIAS pixel_6911/NB2 pixel_6911/AMP_IN pixel_6911/SF_IB
+ pixel_6911/PIX_OUT pixel_6911/CSA_VREF pixel
Xpixel_6922 pixel_6922/gring pixel_6922/VDD pixel_6922/GND pixel_6922/VREF pixel_6922/ROW_SEL
+ pixel_6922/NB1 pixel_6922/VBIAS pixel_6922/NB2 pixel_6922/AMP_IN pixel_6922/SF_IB
+ pixel_6922/PIX_OUT pixel_6922/CSA_VREF pixel
Xpixel_7667 pixel_7667/gring pixel_7667/VDD pixel_7667/GND pixel_7667/VREF pixel_7667/ROW_SEL
+ pixel_7667/NB1 pixel_7667/VBIAS pixel_7667/NB2 pixel_7667/AMP_IN pixel_7667/SF_IB
+ pixel_7667/PIX_OUT pixel_7667/CSA_VREF pixel
Xpixel_7678 pixel_7678/gring pixel_7678/VDD pixel_7678/GND pixel_7678/VREF pixel_7678/ROW_SEL
+ pixel_7678/NB1 pixel_7678/VBIAS pixel_7678/NB2 pixel_7678/AMP_IN pixel_7678/SF_IB
+ pixel_7678/PIX_OUT pixel_7678/CSA_VREF pixel
Xpixel_7689 pixel_7689/gring pixel_7689/VDD pixel_7689/GND pixel_7689/VREF pixel_7689/ROW_SEL
+ pixel_7689/NB1 pixel_7689/VBIAS pixel_7689/NB2 pixel_7689/AMP_IN pixel_7689/SF_IB
+ pixel_7689/PIX_OUT pixel_7689/CSA_VREF pixel
Xpixel_6933 pixel_6933/gring pixel_6933/VDD pixel_6933/GND pixel_6933/VREF pixel_6933/ROW_SEL
+ pixel_6933/NB1 pixel_6933/VBIAS pixel_6933/NB2 pixel_6933/AMP_IN pixel_6933/SF_IB
+ pixel_6933/PIX_OUT pixel_6933/CSA_VREF pixel
Xpixel_6944 pixel_6944/gring pixel_6944/VDD pixel_6944/GND pixel_6944/VREF pixel_6944/ROW_SEL
+ pixel_6944/NB1 pixel_6944/VBIAS pixel_6944/NB2 pixel_6944/AMP_IN pixel_6944/SF_IB
+ pixel_6944/PIX_OUT pixel_6944/CSA_VREF pixel
Xpixel_6955 pixel_6955/gring pixel_6955/VDD pixel_6955/GND pixel_6955/VREF pixel_6955/ROW_SEL
+ pixel_6955/NB1 pixel_6955/VBIAS pixel_6955/NB2 pixel_6955/AMP_IN pixel_6955/SF_IB
+ pixel_6955/PIX_OUT pixel_6955/CSA_VREF pixel
Xpixel_36 pixel_36/gring pixel_36/VDD pixel_36/GND pixel_36/VREF pixel_36/ROW_SEL
+ pixel_36/NB1 pixel_36/VBIAS pixel_36/NB2 pixel_36/AMP_IN pixel_36/SF_IB pixel_36/PIX_OUT
+ pixel_36/CSA_VREF pixel
Xpixel_25 pixel_25/gring pixel_25/VDD pixel_25/GND pixel_25/VREF pixel_25/ROW_SEL
+ pixel_25/NB1 pixel_25/VBIAS pixel_25/NB2 pixel_25/AMP_IN pixel_25/SF_IB pixel_25/PIX_OUT
+ pixel_25/CSA_VREF pixel
Xpixel_14 pixel_14/gring pixel_14/VDD pixel_14/GND pixel_14/VREF pixel_14/ROW_SEL
+ pixel_14/NB1 pixel_14/VBIAS pixel_14/NB2 pixel_14/AMP_IN pixel_14/SF_IB pixel_14/PIX_OUT
+ pixel_14/CSA_VREF pixel
Xpixel_6966 pixel_6966/gring pixel_6966/VDD pixel_6966/GND pixel_6966/VREF pixel_6966/ROW_SEL
+ pixel_6966/NB1 pixel_6966/VBIAS pixel_6966/NB2 pixel_6966/AMP_IN pixel_6966/SF_IB
+ pixel_6966/PIX_OUT pixel_6966/CSA_VREF pixel
Xpixel_6977 pixel_6977/gring pixel_6977/VDD pixel_6977/GND pixel_6977/VREF pixel_6977/ROW_SEL
+ pixel_6977/NB1 pixel_6977/VBIAS pixel_6977/NB2 pixel_6977/AMP_IN pixel_6977/SF_IB
+ pixel_6977/PIX_OUT pixel_6977/CSA_VREF pixel
Xpixel_6988 pixel_6988/gring pixel_6988/VDD pixel_6988/GND pixel_6988/VREF pixel_6988/ROW_SEL
+ pixel_6988/NB1 pixel_6988/VBIAS pixel_6988/NB2 pixel_6988/AMP_IN pixel_6988/SF_IB
+ pixel_6988/PIX_OUT pixel_6988/CSA_VREF pixel
Xpixel_69 pixel_69/gring pixel_69/VDD pixel_69/GND pixel_69/VREF pixel_69/ROW_SEL
+ pixel_69/NB1 pixel_69/VBIAS pixel_69/NB2 pixel_69/AMP_IN pixel_69/SF_IB pixel_69/PIX_OUT
+ pixel_69/CSA_VREF pixel
Xpixel_58 pixel_58/gring pixel_58/VDD pixel_58/GND pixel_58/VREF pixel_58/ROW_SEL
+ pixel_58/NB1 pixel_58/VBIAS pixel_58/NB2 pixel_58/AMP_IN pixel_58/SF_IB pixel_58/PIX_OUT
+ pixel_58/CSA_VREF pixel
Xpixel_47 pixel_47/gring pixel_47/VDD pixel_47/GND pixel_47/VREF pixel_47/ROW_SEL
+ pixel_47/NB1 pixel_47/VBIAS pixel_47/NB2 pixel_47/AMP_IN pixel_47/SF_IB pixel_47/PIX_OUT
+ pixel_47/CSA_VREF pixel
Xpixel_6999 pixel_6999/gring pixel_6999/VDD pixel_6999/GND pixel_6999/VREF pixel_6999/ROW_SEL
+ pixel_6999/NB1 pixel_6999/VBIAS pixel_6999/NB2 pixel_6999/AMP_IN pixel_6999/SF_IB
+ pixel_6999/PIX_OUT pixel_6999/CSA_VREF pixel
Xpixel_1251 pixel_1251/gring pixel_1251/VDD pixel_1251/GND pixel_1251/VREF pixel_1251/ROW_SEL
+ pixel_1251/NB1 pixel_1251/VBIAS pixel_1251/NB2 pixel_1251/AMP_IN pixel_1251/SF_IB
+ pixel_1251/PIX_OUT pixel_1251/CSA_VREF pixel
Xpixel_1240 pixel_1240/gring pixel_1240/VDD pixel_1240/GND pixel_1240/VREF pixel_1240/ROW_SEL
+ pixel_1240/NB1 pixel_1240/VBIAS pixel_1240/NB2 pixel_1240/AMP_IN pixel_1240/SF_IB
+ pixel_1240/PIX_OUT pixel_1240/CSA_VREF pixel
Xpixel_1284 pixel_1284/gring pixel_1284/VDD pixel_1284/GND pixel_1284/VREF pixel_1284/ROW_SEL
+ pixel_1284/NB1 pixel_1284/VBIAS pixel_1284/NB2 pixel_1284/AMP_IN pixel_1284/SF_IB
+ pixel_1284/PIX_OUT pixel_1284/CSA_VREF pixel
Xpixel_1273 pixel_1273/gring pixel_1273/VDD pixel_1273/GND pixel_1273/VREF pixel_1273/ROW_SEL
+ pixel_1273/NB1 pixel_1273/VBIAS pixel_1273/NB2 pixel_1273/AMP_IN pixel_1273/SF_IB
+ pixel_1273/PIX_OUT pixel_1273/CSA_VREF pixel
Xpixel_1262 pixel_1262/gring pixel_1262/VDD pixel_1262/GND pixel_1262/VREF pixel_1262/ROW_SEL
+ pixel_1262/NB1 pixel_1262/VBIAS pixel_1262/NB2 pixel_1262/AMP_IN pixel_1262/SF_IB
+ pixel_1262/PIX_OUT pixel_1262/CSA_VREF pixel
Xpixel_1295 pixel_1295/gring pixel_1295/VDD pixel_1295/GND pixel_1295/VREF pixel_1295/ROW_SEL
+ pixel_1295/NB1 pixel_1295/VBIAS pixel_1295/NB2 pixel_1295/AMP_IN pixel_1295/SF_IB
+ pixel_1295/PIX_OUT pixel_1295/CSA_VREF pixel
Xpixel_9592 pixel_9592/gring pixel_9592/VDD pixel_9592/GND pixel_9592/VREF pixel_9592/ROW_SEL
+ pixel_9592/NB1 pixel_9592/VBIAS pixel_9592/NB2 pixel_9592/AMP_IN pixel_9592/SF_IB
+ pixel_9592/PIX_OUT pixel_9592/CSA_VREF pixel
Xpixel_9581 pixel_9581/gring pixel_9581/VDD pixel_9581/GND pixel_9581/VREF pixel_9581/ROW_SEL
+ pixel_9581/NB1 pixel_9581/VBIAS pixel_9581/NB2 pixel_9581/AMP_IN pixel_9581/SF_IB
+ pixel_9581/PIX_OUT pixel_9581/CSA_VREF pixel
Xpixel_9570 pixel_9570/gring pixel_9570/VDD pixel_9570/GND pixel_9570/VREF pixel_9570/ROW_SEL
+ pixel_9570/NB1 pixel_9570/VBIAS pixel_9570/NB2 pixel_9570/AMP_IN pixel_9570/SF_IB
+ pixel_9570/PIX_OUT pixel_9570/CSA_VREF pixel
Xpixel_8891 pixel_8891/gring pixel_8891/VDD pixel_8891/GND pixel_8891/VREF pixel_8891/ROW_SEL
+ pixel_8891/NB1 pixel_8891/VBIAS pixel_8891/NB2 pixel_8891/AMP_IN pixel_8891/SF_IB
+ pixel_8891/PIX_OUT pixel_8891/CSA_VREF pixel
Xpixel_8880 pixel_8880/gring pixel_8880/VDD pixel_8880/GND pixel_8880/VREF pixel_8880/ROW_SEL
+ pixel_8880/NB1 pixel_8880/VBIAS pixel_8880/NB2 pixel_8880/AMP_IN pixel_8880/SF_IB
+ pixel_8880/PIX_OUT pixel_8880/CSA_VREF pixel
Xpixel_6207 pixel_6207/gring pixel_6207/VDD pixel_6207/GND pixel_6207/VREF pixel_6207/ROW_SEL
+ pixel_6207/NB1 pixel_6207/VBIAS pixel_6207/NB2 pixel_6207/AMP_IN pixel_6207/SF_IB
+ pixel_6207/PIX_OUT pixel_6207/CSA_VREF pixel
Xpixel_6218 pixel_6218/gring pixel_6218/VDD pixel_6218/GND pixel_6218/VREF pixel_6218/ROW_SEL
+ pixel_6218/NB1 pixel_6218/VBIAS pixel_6218/NB2 pixel_6218/AMP_IN pixel_6218/SF_IB
+ pixel_6218/PIX_OUT pixel_6218/CSA_VREF pixel
Xpixel_6229 pixel_6229/gring pixel_6229/VDD pixel_6229/GND pixel_6229/VREF pixel_6229/ROW_SEL
+ pixel_6229/NB1 pixel_6229/VBIAS pixel_6229/NB2 pixel_6229/AMP_IN pixel_6229/SF_IB
+ pixel_6229/PIX_OUT pixel_6229/CSA_VREF pixel
Xpixel_5506 pixel_5506/gring pixel_5506/VDD pixel_5506/GND pixel_5506/VREF pixel_5506/ROW_SEL
+ pixel_5506/NB1 pixel_5506/VBIAS pixel_5506/NB2 pixel_5506/AMP_IN pixel_5506/SF_IB
+ pixel_5506/PIX_OUT pixel_5506/CSA_VREF pixel
Xpixel_5517 pixel_5517/gring pixel_5517/VDD pixel_5517/GND pixel_5517/VREF pixel_5517/ROW_SEL
+ pixel_5517/NB1 pixel_5517/VBIAS pixel_5517/NB2 pixel_5517/AMP_IN pixel_5517/SF_IB
+ pixel_5517/PIX_OUT pixel_5517/CSA_VREF pixel
Xpixel_5528 pixel_5528/gring pixel_5528/VDD pixel_5528/GND pixel_5528/VREF pixel_5528/ROW_SEL
+ pixel_5528/NB1 pixel_5528/VBIAS pixel_5528/NB2 pixel_5528/AMP_IN pixel_5528/SF_IB
+ pixel_5528/PIX_OUT pixel_5528/CSA_VREF pixel
Xpixel_5539 pixel_5539/gring pixel_5539/VDD pixel_5539/GND pixel_5539/VREF pixel_5539/ROW_SEL
+ pixel_5539/NB1 pixel_5539/VBIAS pixel_5539/NB2 pixel_5539/AMP_IN pixel_5539/SF_IB
+ pixel_5539/PIX_OUT pixel_5539/CSA_VREF pixel
Xpixel_833 pixel_833/gring pixel_833/VDD pixel_833/GND pixel_833/VREF pixel_833/ROW_SEL
+ pixel_833/NB1 pixel_833/VBIAS pixel_833/NB2 pixel_833/AMP_IN pixel_833/SF_IB pixel_833/PIX_OUT
+ pixel_833/CSA_VREF pixel
Xpixel_822 pixel_822/gring pixel_822/VDD pixel_822/GND pixel_822/VREF pixel_822/ROW_SEL
+ pixel_822/NB1 pixel_822/VBIAS pixel_822/NB2 pixel_822/AMP_IN pixel_822/SF_IB pixel_822/PIX_OUT
+ pixel_822/CSA_VREF pixel
Xpixel_811 pixel_811/gring pixel_811/VDD pixel_811/GND pixel_811/VREF pixel_811/ROW_SEL
+ pixel_811/NB1 pixel_811/VBIAS pixel_811/NB2 pixel_811/AMP_IN pixel_811/SF_IB pixel_811/PIX_OUT
+ pixel_811/CSA_VREF pixel
Xpixel_800 pixel_800/gring pixel_800/VDD pixel_800/GND pixel_800/VREF pixel_800/ROW_SEL
+ pixel_800/NB1 pixel_800/VBIAS pixel_800/NB2 pixel_800/AMP_IN pixel_800/SF_IB pixel_800/PIX_OUT
+ pixel_800/CSA_VREF pixel
Xpixel_4805 pixel_4805/gring pixel_4805/VDD pixel_4805/GND pixel_4805/VREF pixel_4805/ROW_SEL
+ pixel_4805/NB1 pixel_4805/VBIAS pixel_4805/NB2 pixel_4805/AMP_IN pixel_4805/SF_IB
+ pixel_4805/PIX_OUT pixel_4805/CSA_VREF pixel
Xpixel_4816 pixel_4816/gring pixel_4816/VDD pixel_4816/GND pixel_4816/VREF pixel_4816/ROW_SEL
+ pixel_4816/NB1 pixel_4816/VBIAS pixel_4816/NB2 pixel_4816/AMP_IN pixel_4816/SF_IB
+ pixel_4816/PIX_OUT pixel_4816/CSA_VREF pixel
Xpixel_4827 pixel_4827/gring pixel_4827/VDD pixel_4827/GND pixel_4827/VREF pixel_4827/ROW_SEL
+ pixel_4827/NB1 pixel_4827/VBIAS pixel_4827/NB2 pixel_4827/AMP_IN pixel_4827/SF_IB
+ pixel_4827/PIX_OUT pixel_4827/CSA_VREF pixel
Xpixel_4838 pixel_4838/gring pixel_4838/VDD pixel_4838/GND pixel_4838/VREF pixel_4838/ROW_SEL
+ pixel_4838/NB1 pixel_4838/VBIAS pixel_4838/NB2 pixel_4838/AMP_IN pixel_4838/SF_IB
+ pixel_4838/PIX_OUT pixel_4838/CSA_VREF pixel
Xpixel_866 pixel_866/gring pixel_866/VDD pixel_866/GND pixel_866/VREF pixel_866/ROW_SEL
+ pixel_866/NB1 pixel_866/VBIAS pixel_866/NB2 pixel_866/AMP_IN pixel_866/SF_IB pixel_866/PIX_OUT
+ pixel_866/CSA_VREF pixel
Xpixel_855 pixel_855/gring pixel_855/VDD pixel_855/GND pixel_855/VREF pixel_855/ROW_SEL
+ pixel_855/NB1 pixel_855/VBIAS pixel_855/NB2 pixel_855/AMP_IN pixel_855/SF_IB pixel_855/PIX_OUT
+ pixel_855/CSA_VREF pixel
Xpixel_844 pixel_844/gring pixel_844/VDD pixel_844/GND pixel_844/VREF pixel_844/ROW_SEL
+ pixel_844/NB1 pixel_844/VBIAS pixel_844/NB2 pixel_844/AMP_IN pixel_844/SF_IB pixel_844/PIX_OUT
+ pixel_844/CSA_VREF pixel
Xpixel_4849 pixel_4849/gring pixel_4849/VDD pixel_4849/GND pixel_4849/VREF pixel_4849/ROW_SEL
+ pixel_4849/NB1 pixel_4849/VBIAS pixel_4849/NB2 pixel_4849/AMP_IN pixel_4849/SF_IB
+ pixel_4849/PIX_OUT pixel_4849/CSA_VREF pixel
Xpixel_899 pixel_899/gring pixel_899/VDD pixel_899/GND pixel_899/VREF pixel_899/ROW_SEL
+ pixel_899/NB1 pixel_899/VBIAS pixel_899/NB2 pixel_899/AMP_IN pixel_899/SF_IB pixel_899/PIX_OUT
+ pixel_899/CSA_VREF pixel
Xpixel_888 pixel_888/gring pixel_888/VDD pixel_888/GND pixel_888/VREF pixel_888/ROW_SEL
+ pixel_888/NB1 pixel_888/VBIAS pixel_888/NB2 pixel_888/AMP_IN pixel_888/SF_IB pixel_888/PIX_OUT
+ pixel_888/CSA_VREF pixel
Xpixel_877 pixel_877/gring pixel_877/VDD pixel_877/GND pixel_877/VREF pixel_877/ROW_SEL
+ pixel_877/NB1 pixel_877/VBIAS pixel_877/NB2 pixel_877/AMP_IN pixel_877/SF_IB pixel_877/PIX_OUT
+ pixel_877/CSA_VREF pixel
Xpixel_8110 pixel_8110/gring pixel_8110/VDD pixel_8110/GND pixel_8110/VREF pixel_8110/ROW_SEL
+ pixel_8110/NB1 pixel_8110/VBIAS pixel_8110/NB2 pixel_8110/AMP_IN pixel_8110/SF_IB
+ pixel_8110/PIX_OUT pixel_8110/CSA_VREF pixel
Xpixel_8121 pixel_8121/gring pixel_8121/VDD pixel_8121/GND pixel_8121/VREF pixel_8121/ROW_SEL
+ pixel_8121/NB1 pixel_8121/VBIAS pixel_8121/NB2 pixel_8121/AMP_IN pixel_8121/SF_IB
+ pixel_8121/PIX_OUT pixel_8121/CSA_VREF pixel
Xpixel_8132 pixel_8132/gring pixel_8132/VDD pixel_8132/GND pixel_8132/VREF pixel_8132/ROW_SEL
+ pixel_8132/NB1 pixel_8132/VBIAS pixel_8132/NB2 pixel_8132/AMP_IN pixel_8132/SF_IB
+ pixel_8132/PIX_OUT pixel_8132/CSA_VREF pixel
Xpixel_8143 pixel_8143/gring pixel_8143/VDD pixel_8143/GND pixel_8143/VREF pixel_8143/ROW_SEL
+ pixel_8143/NB1 pixel_8143/VBIAS pixel_8143/NB2 pixel_8143/AMP_IN pixel_8143/SF_IB
+ pixel_8143/PIX_OUT pixel_8143/CSA_VREF pixel
Xpixel_8154 pixel_8154/gring pixel_8154/VDD pixel_8154/GND pixel_8154/VREF pixel_8154/ROW_SEL
+ pixel_8154/NB1 pixel_8154/VBIAS pixel_8154/NB2 pixel_8154/AMP_IN pixel_8154/SF_IB
+ pixel_8154/PIX_OUT pixel_8154/CSA_VREF pixel
Xpixel_8165 pixel_8165/gring pixel_8165/VDD pixel_8165/GND pixel_8165/VREF pixel_8165/ROW_SEL
+ pixel_8165/NB1 pixel_8165/VBIAS pixel_8165/NB2 pixel_8165/AMP_IN pixel_8165/SF_IB
+ pixel_8165/PIX_OUT pixel_8165/CSA_VREF pixel
Xpixel_8176 pixel_8176/gring pixel_8176/VDD pixel_8176/GND pixel_8176/VREF pixel_8176/ROW_SEL
+ pixel_8176/NB1 pixel_8176/VBIAS pixel_8176/NB2 pixel_8176/AMP_IN pixel_8176/SF_IB
+ pixel_8176/PIX_OUT pixel_8176/CSA_VREF pixel
Xpixel_7420 pixel_7420/gring pixel_7420/VDD pixel_7420/GND pixel_7420/VREF pixel_7420/ROW_SEL
+ pixel_7420/NB1 pixel_7420/VBIAS pixel_7420/NB2 pixel_7420/AMP_IN pixel_7420/SF_IB
+ pixel_7420/PIX_OUT pixel_7420/CSA_VREF pixel
Xpixel_7431 pixel_7431/gring pixel_7431/VDD pixel_7431/GND pixel_7431/VREF pixel_7431/ROW_SEL
+ pixel_7431/NB1 pixel_7431/VBIAS pixel_7431/NB2 pixel_7431/AMP_IN pixel_7431/SF_IB
+ pixel_7431/PIX_OUT pixel_7431/CSA_VREF pixel
Xpixel_8187 pixel_8187/gring pixel_8187/VDD pixel_8187/GND pixel_8187/VREF pixel_8187/ROW_SEL
+ pixel_8187/NB1 pixel_8187/VBIAS pixel_8187/NB2 pixel_8187/AMP_IN pixel_8187/SF_IB
+ pixel_8187/PIX_OUT pixel_8187/CSA_VREF pixel
Xpixel_8198 pixel_8198/gring pixel_8198/VDD pixel_8198/GND pixel_8198/VREF pixel_8198/ROW_SEL
+ pixel_8198/NB1 pixel_8198/VBIAS pixel_8198/NB2 pixel_8198/AMP_IN pixel_8198/SF_IB
+ pixel_8198/PIX_OUT pixel_8198/CSA_VREF pixel
Xpixel_7442 pixel_7442/gring pixel_7442/VDD pixel_7442/GND pixel_7442/VREF pixel_7442/ROW_SEL
+ pixel_7442/NB1 pixel_7442/VBIAS pixel_7442/NB2 pixel_7442/AMP_IN pixel_7442/SF_IB
+ pixel_7442/PIX_OUT pixel_7442/CSA_VREF pixel
Xpixel_7453 pixel_7453/gring pixel_7453/VDD pixel_7453/GND pixel_7453/VREF pixel_7453/ROW_SEL
+ pixel_7453/NB1 pixel_7453/VBIAS pixel_7453/NB2 pixel_7453/AMP_IN pixel_7453/SF_IB
+ pixel_7453/PIX_OUT pixel_7453/CSA_VREF pixel
Xpixel_7464 pixel_7464/gring pixel_7464/VDD pixel_7464/GND pixel_7464/VREF pixel_7464/ROW_SEL
+ pixel_7464/NB1 pixel_7464/VBIAS pixel_7464/NB2 pixel_7464/AMP_IN pixel_7464/SF_IB
+ pixel_7464/PIX_OUT pixel_7464/CSA_VREF pixel
Xpixel_7475 pixel_7475/gring pixel_7475/VDD pixel_7475/GND pixel_7475/VREF pixel_7475/ROW_SEL
+ pixel_7475/NB1 pixel_7475/VBIAS pixel_7475/NB2 pixel_7475/AMP_IN pixel_7475/SF_IB
+ pixel_7475/PIX_OUT pixel_7475/CSA_VREF pixel
Xpixel_6730 pixel_6730/gring pixel_6730/VDD pixel_6730/GND pixel_6730/VREF pixel_6730/ROW_SEL
+ pixel_6730/NB1 pixel_6730/VBIAS pixel_6730/NB2 pixel_6730/AMP_IN pixel_6730/SF_IB
+ pixel_6730/PIX_OUT pixel_6730/CSA_VREF pixel
Xpixel_7486 pixel_7486/gring pixel_7486/VDD pixel_7486/GND pixel_7486/VREF pixel_7486/ROW_SEL
+ pixel_7486/NB1 pixel_7486/VBIAS pixel_7486/NB2 pixel_7486/AMP_IN pixel_7486/SF_IB
+ pixel_7486/PIX_OUT pixel_7486/CSA_VREF pixel
Xpixel_7497 pixel_7497/gring pixel_7497/VDD pixel_7497/GND pixel_7497/VREF pixel_7497/ROW_SEL
+ pixel_7497/NB1 pixel_7497/VBIAS pixel_7497/NB2 pixel_7497/AMP_IN pixel_7497/SF_IB
+ pixel_7497/PIX_OUT pixel_7497/CSA_VREF pixel
Xpixel_6741 pixel_6741/gring pixel_6741/VDD pixel_6741/GND pixel_6741/VREF pixel_6741/ROW_SEL
+ pixel_6741/NB1 pixel_6741/VBIAS pixel_6741/NB2 pixel_6741/AMP_IN pixel_6741/SF_IB
+ pixel_6741/PIX_OUT pixel_6741/CSA_VREF pixel
Xpixel_6752 pixel_6752/gring pixel_6752/VDD pixel_6752/GND pixel_6752/VREF pixel_6752/ROW_SEL
+ pixel_6752/NB1 pixel_6752/VBIAS pixel_6752/NB2 pixel_6752/AMP_IN pixel_6752/SF_IB
+ pixel_6752/PIX_OUT pixel_6752/CSA_VREF pixel
Xpixel_6763 pixel_6763/gring pixel_6763/VDD pixel_6763/GND pixel_6763/VREF pixel_6763/ROW_SEL
+ pixel_6763/NB1 pixel_6763/VBIAS pixel_6763/NB2 pixel_6763/AMP_IN pixel_6763/SF_IB
+ pixel_6763/PIX_OUT pixel_6763/CSA_VREF pixel
Xpixel_6774 pixel_6774/gring pixel_6774/VDD pixel_6774/GND pixel_6774/VREF pixel_6774/ROW_SEL
+ pixel_6774/NB1 pixel_6774/VBIAS pixel_6774/NB2 pixel_6774/AMP_IN pixel_6774/SF_IB
+ pixel_6774/PIX_OUT pixel_6774/CSA_VREF pixel
Xpixel_6785 pixel_6785/gring pixel_6785/VDD pixel_6785/GND pixel_6785/VREF pixel_6785/ROW_SEL
+ pixel_6785/NB1 pixel_6785/VBIAS pixel_6785/NB2 pixel_6785/AMP_IN pixel_6785/SF_IB
+ pixel_6785/PIX_OUT pixel_6785/CSA_VREF pixel
Xpixel_6796 pixel_6796/gring pixel_6796/VDD pixel_6796/GND pixel_6796/VREF pixel_6796/ROW_SEL
+ pixel_6796/NB1 pixel_6796/VBIAS pixel_6796/NB2 pixel_6796/AMP_IN pixel_6796/SF_IB
+ pixel_6796/PIX_OUT pixel_6796/CSA_VREF pixel
Xpixel_1092 pixel_1092/gring pixel_1092/VDD pixel_1092/GND pixel_1092/VREF pixel_1092/ROW_SEL
+ pixel_1092/NB1 pixel_1092/VBIAS pixel_1092/NB2 pixel_1092/AMP_IN pixel_1092/SF_IB
+ pixel_1092/PIX_OUT pixel_1092/CSA_VREF pixel
Xpixel_1081 pixel_1081/gring pixel_1081/VDD pixel_1081/GND pixel_1081/VREF pixel_1081/ROW_SEL
+ pixel_1081/NB1 pixel_1081/VBIAS pixel_1081/NB2 pixel_1081/AMP_IN pixel_1081/SF_IB
+ pixel_1081/PIX_OUT pixel_1081/CSA_VREF pixel
Xpixel_1070 pixel_1070/gring pixel_1070/VDD pixel_1070/GND pixel_1070/VREF pixel_1070/ROW_SEL
+ pixel_1070/NB1 pixel_1070/VBIAS pixel_1070/NB2 pixel_1070/AMP_IN pixel_1070/SF_IB
+ pixel_1070/PIX_OUT pixel_1070/CSA_VREF pixel
Xpixel_118 pixel_118/gring pixel_118/VDD pixel_118/GND pixel_118/VREF pixel_118/ROW_SEL
+ pixel_118/NB1 pixel_118/VBIAS pixel_118/NB2 pixel_118/AMP_IN pixel_118/SF_IB pixel_118/PIX_OUT
+ pixel_118/CSA_VREF pixel
Xpixel_107 pixel_107/gring pixel_107/VDD pixel_107/GND pixel_107/VREF pixel_107/ROW_SEL
+ pixel_107/NB1 pixel_107/VBIAS pixel_107/NB2 pixel_107/AMP_IN pixel_107/SF_IB pixel_107/PIX_OUT
+ pixel_107/CSA_VREF pixel
Xpixel_129 pixel_129/gring pixel_129/VDD pixel_129/GND pixel_129/VREF pixel_129/ROW_SEL
+ pixel_129/NB1 pixel_129/VBIAS pixel_129/NB2 pixel_129/AMP_IN pixel_129/SF_IB pixel_129/PIX_OUT
+ pixel_129/CSA_VREF pixel
Xpixel_6004 pixel_6004/gring pixel_6004/VDD pixel_6004/GND pixel_6004/VREF pixel_6004/ROW_SEL
+ pixel_6004/NB1 pixel_6004/VBIAS pixel_6004/NB2 pixel_6004/AMP_IN pixel_6004/SF_IB
+ pixel_6004/PIX_OUT pixel_6004/CSA_VREF pixel
Xpixel_6015 pixel_6015/gring pixel_6015/VDD pixel_6015/GND pixel_6015/VREF pixel_6015/ROW_SEL
+ pixel_6015/NB1 pixel_6015/VBIAS pixel_6015/NB2 pixel_6015/AMP_IN pixel_6015/SF_IB
+ pixel_6015/PIX_OUT pixel_6015/CSA_VREF pixel
Xpixel_6026 pixel_6026/gring pixel_6026/VDD pixel_6026/GND pixel_6026/VREF pixel_6026/ROW_SEL
+ pixel_6026/NB1 pixel_6026/VBIAS pixel_6026/NB2 pixel_6026/AMP_IN pixel_6026/SF_IB
+ pixel_6026/PIX_OUT pixel_6026/CSA_VREF pixel
Xpixel_6037 pixel_6037/gring pixel_6037/VDD pixel_6037/GND pixel_6037/VREF pixel_6037/ROW_SEL
+ pixel_6037/NB1 pixel_6037/VBIAS pixel_6037/NB2 pixel_6037/AMP_IN pixel_6037/SF_IB
+ pixel_6037/PIX_OUT pixel_6037/CSA_VREF pixel
Xpixel_6048 pixel_6048/gring pixel_6048/VDD pixel_6048/GND pixel_6048/VREF pixel_6048/ROW_SEL
+ pixel_6048/NB1 pixel_6048/VBIAS pixel_6048/NB2 pixel_6048/AMP_IN pixel_6048/SF_IB
+ pixel_6048/PIX_OUT pixel_6048/CSA_VREF pixel
Xpixel_6059 pixel_6059/gring pixel_6059/VDD pixel_6059/GND pixel_6059/VREF pixel_6059/ROW_SEL
+ pixel_6059/NB1 pixel_6059/VBIAS pixel_6059/NB2 pixel_6059/AMP_IN pixel_6059/SF_IB
+ pixel_6059/PIX_OUT pixel_6059/CSA_VREF pixel
Xpixel_5303 pixel_5303/gring pixel_5303/VDD pixel_5303/GND pixel_5303/VREF pixel_5303/ROW_SEL
+ pixel_5303/NB1 pixel_5303/VBIAS pixel_5303/NB2 pixel_5303/AMP_IN pixel_5303/SF_IB
+ pixel_5303/PIX_OUT pixel_5303/CSA_VREF pixel
Xpixel_5314 pixel_5314/gring pixel_5314/VDD pixel_5314/GND pixel_5314/VREF pixel_5314/ROW_SEL
+ pixel_5314/NB1 pixel_5314/VBIAS pixel_5314/NB2 pixel_5314/AMP_IN pixel_5314/SF_IB
+ pixel_5314/PIX_OUT pixel_5314/CSA_VREF pixel
Xpixel_5325 pixel_5325/gring pixel_5325/VDD pixel_5325/GND pixel_5325/VREF pixel_5325/ROW_SEL
+ pixel_5325/NB1 pixel_5325/VBIAS pixel_5325/NB2 pixel_5325/AMP_IN pixel_5325/SF_IB
+ pixel_5325/PIX_OUT pixel_5325/CSA_VREF pixel
Xpixel_5336 pixel_5336/gring pixel_5336/VDD pixel_5336/GND pixel_5336/VREF pixel_5336/ROW_SEL
+ pixel_5336/NB1 pixel_5336/VBIAS pixel_5336/NB2 pixel_5336/AMP_IN pixel_5336/SF_IB
+ pixel_5336/PIX_OUT pixel_5336/CSA_VREF pixel
Xpixel_5347 pixel_5347/gring pixel_5347/VDD pixel_5347/GND pixel_5347/VREF pixel_5347/ROW_SEL
+ pixel_5347/NB1 pixel_5347/VBIAS pixel_5347/NB2 pixel_5347/AMP_IN pixel_5347/SF_IB
+ pixel_5347/PIX_OUT pixel_5347/CSA_VREF pixel
Xpixel_4602 pixel_4602/gring pixel_4602/VDD pixel_4602/GND pixel_4602/VREF pixel_4602/ROW_SEL
+ pixel_4602/NB1 pixel_4602/VBIAS pixel_4602/NB2 pixel_4602/AMP_IN pixel_4602/SF_IB
+ pixel_4602/PIX_OUT pixel_4602/CSA_VREF pixel
Xpixel_641 pixel_641/gring pixel_641/VDD pixel_641/GND pixel_641/VREF pixel_641/ROW_SEL
+ pixel_641/NB1 pixel_641/VBIAS pixel_641/NB2 pixel_641/AMP_IN pixel_641/SF_IB pixel_641/PIX_OUT
+ pixel_641/CSA_VREF pixel
Xpixel_630 pixel_630/gring pixel_630/VDD pixel_630/GND pixel_630/VREF pixel_630/ROW_SEL
+ pixel_630/NB1 pixel_630/VBIAS pixel_630/NB2 pixel_630/AMP_IN pixel_630/SF_IB pixel_630/PIX_OUT
+ pixel_630/CSA_VREF pixel
Xpixel_5358 pixel_5358/gring pixel_5358/VDD pixel_5358/GND pixel_5358/VREF pixel_5358/ROW_SEL
+ pixel_5358/NB1 pixel_5358/VBIAS pixel_5358/NB2 pixel_5358/AMP_IN pixel_5358/SF_IB
+ pixel_5358/PIX_OUT pixel_5358/CSA_VREF pixel
Xpixel_5369 pixel_5369/gring pixel_5369/VDD pixel_5369/GND pixel_5369/VREF pixel_5369/ROW_SEL
+ pixel_5369/NB1 pixel_5369/VBIAS pixel_5369/NB2 pixel_5369/AMP_IN pixel_5369/SF_IB
+ pixel_5369/PIX_OUT pixel_5369/CSA_VREF pixel
Xpixel_4613 pixel_4613/gring pixel_4613/VDD pixel_4613/GND pixel_4613/VREF pixel_4613/ROW_SEL
+ pixel_4613/NB1 pixel_4613/VBIAS pixel_4613/NB2 pixel_4613/AMP_IN pixel_4613/SF_IB
+ pixel_4613/PIX_OUT pixel_4613/CSA_VREF pixel
Xpixel_4624 pixel_4624/gring pixel_4624/VDD pixel_4624/GND pixel_4624/VREF pixel_4624/ROW_SEL
+ pixel_4624/NB1 pixel_4624/VBIAS pixel_4624/NB2 pixel_4624/AMP_IN pixel_4624/SF_IB
+ pixel_4624/PIX_OUT pixel_4624/CSA_VREF pixel
Xpixel_4635 pixel_4635/gring pixel_4635/VDD pixel_4635/GND pixel_4635/VREF pixel_4635/ROW_SEL
+ pixel_4635/NB1 pixel_4635/VBIAS pixel_4635/NB2 pixel_4635/AMP_IN pixel_4635/SF_IB
+ pixel_4635/PIX_OUT pixel_4635/CSA_VREF pixel
Xpixel_4646 pixel_4646/gring pixel_4646/VDD pixel_4646/GND pixel_4646/VREF pixel_4646/ROW_SEL
+ pixel_4646/NB1 pixel_4646/VBIAS pixel_4646/NB2 pixel_4646/AMP_IN pixel_4646/SF_IB
+ pixel_4646/PIX_OUT pixel_4646/CSA_VREF pixel
Xpixel_3901 pixel_3901/gring pixel_3901/VDD pixel_3901/GND pixel_3901/VREF pixel_3901/ROW_SEL
+ pixel_3901/NB1 pixel_3901/VBIAS pixel_3901/NB2 pixel_3901/AMP_IN pixel_3901/SF_IB
+ pixel_3901/PIX_OUT pixel_3901/CSA_VREF pixel
Xpixel_674 pixel_674/gring pixel_674/VDD pixel_674/GND pixel_674/VREF pixel_674/ROW_SEL
+ pixel_674/NB1 pixel_674/VBIAS pixel_674/NB2 pixel_674/AMP_IN pixel_674/SF_IB pixel_674/PIX_OUT
+ pixel_674/CSA_VREF pixel
Xpixel_663 pixel_663/gring pixel_663/VDD pixel_663/GND pixel_663/VREF pixel_663/ROW_SEL
+ pixel_663/NB1 pixel_663/VBIAS pixel_663/NB2 pixel_663/AMP_IN pixel_663/SF_IB pixel_663/PIX_OUT
+ pixel_663/CSA_VREF pixel
Xpixel_652 pixel_652/gring pixel_652/VDD pixel_652/GND pixel_652/VREF pixel_652/ROW_SEL
+ pixel_652/NB1 pixel_652/VBIAS pixel_652/NB2 pixel_652/AMP_IN pixel_652/SF_IB pixel_652/PIX_OUT
+ pixel_652/CSA_VREF pixel
Xpixel_4657 pixel_4657/gring pixel_4657/VDD pixel_4657/GND pixel_4657/VREF pixel_4657/ROW_SEL
+ pixel_4657/NB1 pixel_4657/VBIAS pixel_4657/NB2 pixel_4657/AMP_IN pixel_4657/SF_IB
+ pixel_4657/PIX_OUT pixel_4657/CSA_VREF pixel
Xpixel_4668 pixel_4668/gring pixel_4668/VDD pixel_4668/GND pixel_4668/VREF pixel_4668/ROW_SEL
+ pixel_4668/NB1 pixel_4668/VBIAS pixel_4668/NB2 pixel_4668/AMP_IN pixel_4668/SF_IB
+ pixel_4668/PIX_OUT pixel_4668/CSA_VREF pixel
Xpixel_4679 pixel_4679/gring pixel_4679/VDD pixel_4679/GND pixel_4679/VREF pixel_4679/ROW_SEL
+ pixel_4679/NB1 pixel_4679/VBIAS pixel_4679/NB2 pixel_4679/AMP_IN pixel_4679/SF_IB
+ pixel_4679/PIX_OUT pixel_4679/CSA_VREF pixel
Xpixel_3912 pixel_3912/gring pixel_3912/VDD pixel_3912/GND pixel_3912/VREF pixel_3912/ROW_SEL
+ pixel_3912/NB1 pixel_3912/VBIAS pixel_3912/NB2 pixel_3912/AMP_IN pixel_3912/SF_IB
+ pixel_3912/PIX_OUT pixel_3912/CSA_VREF pixel
Xpixel_3923 pixel_3923/gring pixel_3923/VDD pixel_3923/GND pixel_3923/VREF pixel_3923/ROW_SEL
+ pixel_3923/NB1 pixel_3923/VBIAS pixel_3923/NB2 pixel_3923/AMP_IN pixel_3923/SF_IB
+ pixel_3923/PIX_OUT pixel_3923/CSA_VREF pixel
Xpixel_3934 pixel_3934/gring pixel_3934/VDD pixel_3934/GND pixel_3934/VREF pixel_3934/ROW_SEL
+ pixel_3934/NB1 pixel_3934/VBIAS pixel_3934/NB2 pixel_3934/AMP_IN pixel_3934/SF_IB
+ pixel_3934/PIX_OUT pixel_3934/CSA_VREF pixel
Xpixel_696 pixel_696/gring pixel_696/VDD pixel_696/GND pixel_696/VREF pixel_696/ROW_SEL
+ pixel_696/NB1 pixel_696/VBIAS pixel_696/NB2 pixel_696/AMP_IN pixel_696/SF_IB pixel_696/PIX_OUT
+ pixel_696/CSA_VREF pixel
Xpixel_685 pixel_685/gring pixel_685/VDD pixel_685/GND pixel_685/VREF pixel_685/ROW_SEL
+ pixel_685/NB1 pixel_685/VBIAS pixel_685/NB2 pixel_685/AMP_IN pixel_685/SF_IB pixel_685/PIX_OUT
+ pixel_685/CSA_VREF pixel
Xpixel_3945 pixel_3945/gring pixel_3945/VDD pixel_3945/GND pixel_3945/VREF pixel_3945/ROW_SEL
+ pixel_3945/NB1 pixel_3945/VBIAS pixel_3945/NB2 pixel_3945/AMP_IN pixel_3945/SF_IB
+ pixel_3945/PIX_OUT pixel_3945/CSA_VREF pixel
Xpixel_3956 pixel_3956/gring pixel_3956/VDD pixel_3956/GND pixel_3956/VREF pixel_3956/ROW_SEL
+ pixel_3956/NB1 pixel_3956/VBIAS pixel_3956/NB2 pixel_3956/AMP_IN pixel_3956/SF_IB
+ pixel_3956/PIX_OUT pixel_3956/CSA_VREF pixel
Xpixel_3967 pixel_3967/gring pixel_3967/VDD pixel_3967/GND pixel_3967/VREF pixel_3967/ROW_SEL
+ pixel_3967/NB1 pixel_3967/VBIAS pixel_3967/NB2 pixel_3967/AMP_IN pixel_3967/SF_IB
+ pixel_3967/PIX_OUT pixel_3967/CSA_VREF pixel
Xpixel_3978 pixel_3978/gring pixel_3978/VDD pixel_3978/GND pixel_3978/VREF pixel_3978/ROW_SEL
+ pixel_3978/NB1 pixel_3978/VBIAS pixel_3978/NB2 pixel_3978/AMP_IN pixel_3978/SF_IB
+ pixel_3978/PIX_OUT pixel_3978/CSA_VREF pixel
Xpixel_3989 pixel_3989/gring pixel_3989/VDD pixel_3989/GND pixel_3989/VREF pixel_3989/ROW_SEL
+ pixel_3989/NB1 pixel_3989/VBIAS pixel_3989/NB2 pixel_3989/AMP_IN pixel_3989/SF_IB
+ pixel_3989/PIX_OUT pixel_3989/CSA_VREF pixel
Xpixel_7250 pixel_7250/gring pixel_7250/VDD pixel_7250/GND pixel_7250/VREF pixel_7250/ROW_SEL
+ pixel_7250/NB1 pixel_7250/VBIAS pixel_7250/NB2 pixel_7250/AMP_IN pixel_7250/SF_IB
+ pixel_7250/PIX_OUT pixel_7250/CSA_VREF pixel
Xpixel_7261 pixel_7261/gring pixel_7261/VDD pixel_7261/GND pixel_7261/VREF pixel_7261/ROW_SEL
+ pixel_7261/NB1 pixel_7261/VBIAS pixel_7261/NB2 pixel_7261/AMP_IN pixel_7261/SF_IB
+ pixel_7261/PIX_OUT pixel_7261/CSA_VREF pixel
Xpixel_7272 pixel_7272/gring pixel_7272/VDD pixel_7272/GND pixel_7272/VREF pixel_7272/ROW_SEL
+ pixel_7272/NB1 pixel_7272/VBIAS pixel_7272/NB2 pixel_7272/AMP_IN pixel_7272/SF_IB
+ pixel_7272/PIX_OUT pixel_7272/CSA_VREF pixel
Xpixel_7283 pixel_7283/gring pixel_7283/VDD pixel_7283/GND pixel_7283/VREF pixel_7283/ROW_SEL
+ pixel_7283/NB1 pixel_7283/VBIAS pixel_7283/NB2 pixel_7283/AMP_IN pixel_7283/SF_IB
+ pixel_7283/PIX_OUT pixel_7283/CSA_VREF pixel
Xpixel_7294 pixel_7294/gring pixel_7294/VDD pixel_7294/GND pixel_7294/VREF pixel_7294/ROW_SEL
+ pixel_7294/NB1 pixel_7294/VBIAS pixel_7294/NB2 pixel_7294/AMP_IN pixel_7294/SF_IB
+ pixel_7294/PIX_OUT pixel_7294/CSA_VREF pixel
Xpixel_6560 pixel_6560/gring pixel_6560/VDD pixel_6560/GND pixel_6560/VREF pixel_6560/ROW_SEL
+ pixel_6560/NB1 pixel_6560/VBIAS pixel_6560/NB2 pixel_6560/AMP_IN pixel_6560/SF_IB
+ pixel_6560/PIX_OUT pixel_6560/CSA_VREF pixel
Xpixel_6571 pixel_6571/gring pixel_6571/VDD pixel_6571/GND pixel_6571/VREF pixel_6571/ROW_SEL
+ pixel_6571/NB1 pixel_6571/VBIAS pixel_6571/NB2 pixel_6571/AMP_IN pixel_6571/SF_IB
+ pixel_6571/PIX_OUT pixel_6571/CSA_VREF pixel
Xpixel_6582 pixel_6582/gring pixel_6582/VDD pixel_6582/GND pixel_6582/VREF pixel_6582/ROW_SEL
+ pixel_6582/NB1 pixel_6582/VBIAS pixel_6582/NB2 pixel_6582/AMP_IN pixel_6582/SF_IB
+ pixel_6582/PIX_OUT pixel_6582/CSA_VREF pixel
Xpixel_6593 pixel_6593/gring pixel_6593/VDD pixel_6593/GND pixel_6593/VREF pixel_6593/ROW_SEL
+ pixel_6593/NB1 pixel_6593/VBIAS pixel_6593/NB2 pixel_6593/AMP_IN pixel_6593/SF_IB
+ pixel_6593/PIX_OUT pixel_6593/CSA_VREF pixel
Xpixel_5870 pixel_5870/gring pixel_5870/VDD pixel_5870/GND pixel_5870/VREF pixel_5870/ROW_SEL
+ pixel_5870/NB1 pixel_5870/VBIAS pixel_5870/NB2 pixel_5870/AMP_IN pixel_5870/SF_IB
+ pixel_5870/PIX_OUT pixel_5870/CSA_VREF pixel
Xpixel_5881 pixel_5881/gring pixel_5881/VDD pixel_5881/GND pixel_5881/VREF pixel_5881/ROW_SEL
+ pixel_5881/NB1 pixel_5881/VBIAS pixel_5881/NB2 pixel_5881/AMP_IN pixel_5881/SF_IB
+ pixel_5881/PIX_OUT pixel_5881/CSA_VREF pixel
Xpixel_5892 pixel_5892/gring pixel_5892/VDD pixel_5892/GND pixel_5892/VREF pixel_5892/ROW_SEL
+ pixel_5892/NB1 pixel_5892/VBIAS pixel_5892/NB2 pixel_5892/AMP_IN pixel_5892/SF_IB
+ pixel_5892/PIX_OUT pixel_5892/CSA_VREF pixel
Xpixel_3219 pixel_3219/gring pixel_3219/VDD pixel_3219/GND pixel_3219/VREF pixel_3219/ROW_SEL
+ pixel_3219/NB1 pixel_3219/VBIAS pixel_3219/NB2 pixel_3219/AMP_IN pixel_3219/SF_IB
+ pixel_3219/PIX_OUT pixel_3219/CSA_VREF pixel
Xpixel_3208 pixel_3208/gring pixel_3208/VDD pixel_3208/GND pixel_3208/VREF pixel_3208/ROW_SEL
+ pixel_3208/NB1 pixel_3208/VBIAS pixel_3208/NB2 pixel_3208/AMP_IN pixel_3208/SF_IB
+ pixel_3208/PIX_OUT pixel_3208/CSA_VREF pixel
Xpixel_2518 pixel_2518/gring pixel_2518/VDD pixel_2518/GND pixel_2518/VREF pixel_2518/ROW_SEL
+ pixel_2518/NB1 pixel_2518/VBIAS pixel_2518/NB2 pixel_2518/AMP_IN pixel_2518/SF_IB
+ pixel_2518/PIX_OUT pixel_2518/CSA_VREF pixel
Xpixel_2507 pixel_2507/gring pixel_2507/VDD pixel_2507/GND pixel_2507/VREF pixel_2507/ROW_SEL
+ pixel_2507/NB1 pixel_2507/VBIAS pixel_2507/NB2 pixel_2507/AMP_IN pixel_2507/SF_IB
+ pixel_2507/PIX_OUT pixel_2507/CSA_VREF pixel
Xpixel_1817 pixel_1817/gring pixel_1817/VDD pixel_1817/GND pixel_1817/VREF pixel_1817/ROW_SEL
+ pixel_1817/NB1 pixel_1817/VBIAS pixel_1817/NB2 pixel_1817/AMP_IN pixel_1817/SF_IB
+ pixel_1817/PIX_OUT pixel_1817/CSA_VREF pixel
Xpixel_1806 pixel_1806/gring pixel_1806/VDD pixel_1806/GND pixel_1806/VREF pixel_1806/ROW_SEL
+ pixel_1806/NB1 pixel_1806/VBIAS pixel_1806/NB2 pixel_1806/AMP_IN pixel_1806/SF_IB
+ pixel_1806/PIX_OUT pixel_1806/CSA_VREF pixel
Xpixel_2529 pixel_2529/gring pixel_2529/VDD pixel_2529/GND pixel_2529/VREF pixel_2529/ROW_SEL
+ pixel_2529/NB1 pixel_2529/VBIAS pixel_2529/NB2 pixel_2529/AMP_IN pixel_2529/SF_IB
+ pixel_2529/PIX_OUT pixel_2529/CSA_VREF pixel
Xpixel_1839 pixel_1839/gring pixel_1839/VDD pixel_1839/GND pixel_1839/VREF pixel_1839/ROW_SEL
+ pixel_1839/NB1 pixel_1839/VBIAS pixel_1839/NB2 pixel_1839/AMP_IN pixel_1839/SF_IB
+ pixel_1839/PIX_OUT pixel_1839/CSA_VREF pixel
Xpixel_1828 pixel_1828/gring pixel_1828/VDD pixel_1828/GND pixel_1828/VREF pixel_1828/ROW_SEL
+ pixel_1828/NB1 pixel_1828/VBIAS pixel_1828/NB2 pixel_1828/AMP_IN pixel_1828/SF_IB
+ pixel_1828/PIX_OUT pixel_1828/CSA_VREF pixel
Xpixel_5100 pixel_5100/gring pixel_5100/VDD pixel_5100/GND pixel_5100/VREF pixel_5100/ROW_SEL
+ pixel_5100/NB1 pixel_5100/VBIAS pixel_5100/NB2 pixel_5100/AMP_IN pixel_5100/SF_IB
+ pixel_5100/PIX_OUT pixel_5100/CSA_VREF pixel
Xpixel_5111 pixel_5111/gring pixel_5111/VDD pixel_5111/GND pixel_5111/VREF pixel_5111/ROW_SEL
+ pixel_5111/NB1 pixel_5111/VBIAS pixel_5111/NB2 pixel_5111/AMP_IN pixel_5111/SF_IB
+ pixel_5111/PIX_OUT pixel_5111/CSA_VREF pixel
Xpixel_5122 pixel_5122/gring pixel_5122/VDD pixel_5122/GND pixel_5122/VREF pixel_5122/ROW_SEL
+ pixel_5122/NB1 pixel_5122/VBIAS pixel_5122/NB2 pixel_5122/AMP_IN pixel_5122/SF_IB
+ pixel_5122/PIX_OUT pixel_5122/CSA_VREF pixel
Xpixel_5133 pixel_5133/gring pixel_5133/VDD pixel_5133/GND pixel_5133/VREF pixel_5133/ROW_SEL
+ pixel_5133/NB1 pixel_5133/VBIAS pixel_5133/NB2 pixel_5133/AMP_IN pixel_5133/SF_IB
+ pixel_5133/PIX_OUT pixel_5133/CSA_VREF pixel
Xpixel_5144 pixel_5144/gring pixel_5144/VDD pixel_5144/GND pixel_5144/VREF pixel_5144/ROW_SEL
+ pixel_5144/NB1 pixel_5144/VBIAS pixel_5144/NB2 pixel_5144/AMP_IN pixel_5144/SF_IB
+ pixel_5144/PIX_OUT pixel_5144/CSA_VREF pixel
Xpixel_5155 pixel_5155/gring pixel_5155/VDD pixel_5155/GND pixel_5155/VREF pixel_5155/ROW_SEL
+ pixel_5155/NB1 pixel_5155/VBIAS pixel_5155/NB2 pixel_5155/AMP_IN pixel_5155/SF_IB
+ pixel_5155/PIX_OUT pixel_5155/CSA_VREF pixel
Xpixel_4410 pixel_4410/gring pixel_4410/VDD pixel_4410/GND pixel_4410/VREF pixel_4410/ROW_SEL
+ pixel_4410/NB1 pixel_4410/VBIAS pixel_4410/NB2 pixel_4410/AMP_IN pixel_4410/SF_IB
+ pixel_4410/PIX_OUT pixel_4410/CSA_VREF pixel
Xpixel_4421 pixel_4421/gring pixel_4421/VDD pixel_4421/GND pixel_4421/VREF pixel_4421/ROW_SEL
+ pixel_4421/NB1 pixel_4421/VBIAS pixel_4421/NB2 pixel_4421/AMP_IN pixel_4421/SF_IB
+ pixel_4421/PIX_OUT pixel_4421/CSA_VREF pixel
Xpixel_5166 pixel_5166/gring pixel_5166/VDD pixel_5166/GND pixel_5166/VREF pixel_5166/ROW_SEL
+ pixel_5166/NB1 pixel_5166/VBIAS pixel_5166/NB2 pixel_5166/AMP_IN pixel_5166/SF_IB
+ pixel_5166/PIX_OUT pixel_5166/CSA_VREF pixel
Xpixel_5177 pixel_5177/gring pixel_5177/VDD pixel_5177/GND pixel_5177/VREF pixel_5177/ROW_SEL
+ pixel_5177/NB1 pixel_5177/VBIAS pixel_5177/NB2 pixel_5177/AMP_IN pixel_5177/SF_IB
+ pixel_5177/PIX_OUT pixel_5177/CSA_VREF pixel
Xpixel_5188 pixel_5188/gring pixel_5188/VDD pixel_5188/GND pixel_5188/VREF pixel_5188/ROW_SEL
+ pixel_5188/NB1 pixel_5188/VBIAS pixel_5188/NB2 pixel_5188/AMP_IN pixel_5188/SF_IB
+ pixel_5188/PIX_OUT pixel_5188/CSA_VREF pixel
Xpixel_5199 pixel_5199/gring pixel_5199/VDD pixel_5199/GND pixel_5199/VREF pixel_5199/ROW_SEL
+ pixel_5199/NB1 pixel_5199/VBIAS pixel_5199/NB2 pixel_5199/AMP_IN pixel_5199/SF_IB
+ pixel_5199/PIX_OUT pixel_5199/CSA_VREF pixel
Xpixel_4432 pixel_4432/gring pixel_4432/VDD pixel_4432/GND pixel_4432/VREF pixel_4432/ROW_SEL
+ pixel_4432/NB1 pixel_4432/VBIAS pixel_4432/NB2 pixel_4432/AMP_IN pixel_4432/SF_IB
+ pixel_4432/PIX_OUT pixel_4432/CSA_VREF pixel
Xpixel_4443 pixel_4443/gring pixel_4443/VDD pixel_4443/GND pixel_4443/VREF pixel_4443/ROW_SEL
+ pixel_4443/NB1 pixel_4443/VBIAS pixel_4443/NB2 pixel_4443/AMP_IN pixel_4443/SF_IB
+ pixel_4443/PIX_OUT pixel_4443/CSA_VREF pixel
Xpixel_4454 pixel_4454/gring pixel_4454/VDD pixel_4454/GND pixel_4454/VREF pixel_4454/ROW_SEL
+ pixel_4454/NB1 pixel_4454/VBIAS pixel_4454/NB2 pixel_4454/AMP_IN pixel_4454/SF_IB
+ pixel_4454/PIX_OUT pixel_4454/CSA_VREF pixel
Xpixel_482 pixel_482/gring pixel_482/VDD pixel_482/GND pixel_482/VREF pixel_482/ROW_SEL
+ pixel_482/NB1 pixel_482/VBIAS pixel_482/NB2 pixel_482/AMP_IN pixel_482/SF_IB pixel_482/PIX_OUT
+ pixel_482/CSA_VREF pixel
Xpixel_471 pixel_471/gring pixel_471/VDD pixel_471/GND pixel_471/VREF pixel_471/ROW_SEL
+ pixel_471/NB1 pixel_471/VBIAS pixel_471/NB2 pixel_471/AMP_IN pixel_471/SF_IB pixel_471/PIX_OUT
+ pixel_471/CSA_VREF pixel
Xpixel_460 pixel_460/gring pixel_460/VDD pixel_460/GND pixel_460/VREF pixel_460/ROW_SEL
+ pixel_460/NB1 pixel_460/VBIAS pixel_460/NB2 pixel_460/AMP_IN pixel_460/SF_IB pixel_460/PIX_OUT
+ pixel_460/CSA_VREF pixel
Xpixel_3742 pixel_3742/gring pixel_3742/VDD pixel_3742/GND pixel_3742/VREF pixel_3742/ROW_SEL
+ pixel_3742/NB1 pixel_3742/VBIAS pixel_3742/NB2 pixel_3742/AMP_IN pixel_3742/SF_IB
+ pixel_3742/PIX_OUT pixel_3742/CSA_VREF pixel
Xpixel_3731 pixel_3731/gring pixel_3731/VDD pixel_3731/GND pixel_3731/VREF pixel_3731/ROW_SEL
+ pixel_3731/NB1 pixel_3731/VBIAS pixel_3731/NB2 pixel_3731/AMP_IN pixel_3731/SF_IB
+ pixel_3731/PIX_OUT pixel_3731/CSA_VREF pixel
Xpixel_3720 pixel_3720/gring pixel_3720/VDD pixel_3720/GND pixel_3720/VREF pixel_3720/ROW_SEL
+ pixel_3720/NB1 pixel_3720/VBIAS pixel_3720/NB2 pixel_3720/AMP_IN pixel_3720/SF_IB
+ pixel_3720/PIX_OUT pixel_3720/CSA_VREF pixel
Xpixel_4465 pixel_4465/gring pixel_4465/VDD pixel_4465/GND pixel_4465/VREF pixel_4465/ROW_SEL
+ pixel_4465/NB1 pixel_4465/VBIAS pixel_4465/NB2 pixel_4465/AMP_IN pixel_4465/SF_IB
+ pixel_4465/PIX_OUT pixel_4465/CSA_VREF pixel
Xpixel_4476 pixel_4476/gring pixel_4476/VDD pixel_4476/GND pixel_4476/VREF pixel_4476/ROW_SEL
+ pixel_4476/NB1 pixel_4476/VBIAS pixel_4476/NB2 pixel_4476/AMP_IN pixel_4476/SF_IB
+ pixel_4476/PIX_OUT pixel_4476/CSA_VREF pixel
Xpixel_4487 pixel_4487/gring pixel_4487/VDD pixel_4487/GND pixel_4487/VREF pixel_4487/ROW_SEL
+ pixel_4487/NB1 pixel_4487/VBIAS pixel_4487/NB2 pixel_4487/AMP_IN pixel_4487/SF_IB
+ pixel_4487/PIX_OUT pixel_4487/CSA_VREF pixel
Xpixel_493 pixel_493/gring pixel_493/VDD pixel_493/GND pixel_493/VREF pixel_493/ROW_SEL
+ pixel_493/NB1 pixel_493/VBIAS pixel_493/NB2 pixel_493/AMP_IN pixel_493/SF_IB pixel_493/PIX_OUT
+ pixel_493/CSA_VREF pixel
Xpixel_3786 pixel_3786/gring pixel_3786/VDD pixel_3786/GND pixel_3786/VREF pixel_3786/ROW_SEL
+ pixel_3786/NB1 pixel_3786/VBIAS pixel_3786/NB2 pixel_3786/AMP_IN pixel_3786/SF_IB
+ pixel_3786/PIX_OUT pixel_3786/CSA_VREF pixel
Xpixel_3775 pixel_3775/gring pixel_3775/VDD pixel_3775/GND pixel_3775/VREF pixel_3775/ROW_SEL
+ pixel_3775/NB1 pixel_3775/VBIAS pixel_3775/NB2 pixel_3775/AMP_IN pixel_3775/SF_IB
+ pixel_3775/PIX_OUT pixel_3775/CSA_VREF pixel
Xpixel_3764 pixel_3764/gring pixel_3764/VDD pixel_3764/GND pixel_3764/VREF pixel_3764/ROW_SEL
+ pixel_3764/NB1 pixel_3764/VBIAS pixel_3764/NB2 pixel_3764/AMP_IN pixel_3764/SF_IB
+ pixel_3764/PIX_OUT pixel_3764/CSA_VREF pixel
Xpixel_3753 pixel_3753/gring pixel_3753/VDD pixel_3753/GND pixel_3753/VREF pixel_3753/ROW_SEL
+ pixel_3753/NB1 pixel_3753/VBIAS pixel_3753/NB2 pixel_3753/AMP_IN pixel_3753/SF_IB
+ pixel_3753/PIX_OUT pixel_3753/CSA_VREF pixel
Xpixel_4498 pixel_4498/gring pixel_4498/VDD pixel_4498/GND pixel_4498/VREF pixel_4498/ROW_SEL
+ pixel_4498/NB1 pixel_4498/VBIAS pixel_4498/NB2 pixel_4498/AMP_IN pixel_4498/SF_IB
+ pixel_4498/PIX_OUT pixel_4498/CSA_VREF pixel
Xpixel_3797 pixel_3797/gring pixel_3797/VDD pixel_3797/GND pixel_3797/VREF pixel_3797/ROW_SEL
+ pixel_3797/NB1 pixel_3797/VBIAS pixel_3797/NB2 pixel_3797/AMP_IN pixel_3797/SF_IB
+ pixel_3797/PIX_OUT pixel_3797/CSA_VREF pixel
Xpixel_7080 pixel_7080/gring pixel_7080/VDD pixel_7080/GND pixel_7080/VREF pixel_7080/ROW_SEL
+ pixel_7080/NB1 pixel_7080/VBIAS pixel_7080/NB2 pixel_7080/AMP_IN pixel_7080/SF_IB
+ pixel_7080/PIX_OUT pixel_7080/CSA_VREF pixel
Xpixel_7091 pixel_7091/gring pixel_7091/VDD pixel_7091/GND pixel_7091/VREF pixel_7091/ROW_SEL
+ pixel_7091/NB1 pixel_7091/VBIAS pixel_7091/NB2 pixel_7091/AMP_IN pixel_7091/SF_IB
+ pixel_7091/PIX_OUT pixel_7091/CSA_VREF pixel
Xpixel_6390 pixel_6390/gring pixel_6390/VDD pixel_6390/GND pixel_6390/VREF pixel_6390/ROW_SEL
+ pixel_6390/NB1 pixel_6390/VBIAS pixel_6390/NB2 pixel_6390/AMP_IN pixel_6390/SF_IB
+ pixel_6390/PIX_OUT pixel_6390/CSA_VREF pixel
Xpixel_8709 pixel_8709/gring pixel_8709/VDD pixel_8709/GND pixel_8709/VREF pixel_8709/ROW_SEL
+ pixel_8709/NB1 pixel_8709/VBIAS pixel_8709/NB2 pixel_8709/AMP_IN pixel_8709/SF_IB
+ pixel_8709/PIX_OUT pixel_8709/CSA_VREF pixel
Xpixel_3005 pixel_3005/gring pixel_3005/VDD pixel_3005/GND pixel_3005/VREF pixel_3005/ROW_SEL
+ pixel_3005/NB1 pixel_3005/VBIAS pixel_3005/NB2 pixel_3005/AMP_IN pixel_3005/SF_IB
+ pixel_3005/PIX_OUT pixel_3005/CSA_VREF pixel
Xpixel_3038 pixel_3038/gring pixel_3038/VDD pixel_3038/GND pixel_3038/VREF pixel_3038/ROW_SEL
+ pixel_3038/NB1 pixel_3038/VBIAS pixel_3038/NB2 pixel_3038/AMP_IN pixel_3038/SF_IB
+ pixel_3038/PIX_OUT pixel_3038/CSA_VREF pixel
Xpixel_3027 pixel_3027/gring pixel_3027/VDD pixel_3027/GND pixel_3027/VREF pixel_3027/ROW_SEL
+ pixel_3027/NB1 pixel_3027/VBIAS pixel_3027/NB2 pixel_3027/AMP_IN pixel_3027/SF_IB
+ pixel_3027/PIX_OUT pixel_3027/CSA_VREF pixel
Xpixel_3016 pixel_3016/gring pixel_3016/VDD pixel_3016/GND pixel_3016/VREF pixel_3016/ROW_SEL
+ pixel_3016/NB1 pixel_3016/VBIAS pixel_3016/NB2 pixel_3016/AMP_IN pixel_3016/SF_IB
+ pixel_3016/PIX_OUT pixel_3016/CSA_VREF pixel
Xpixel_2326 pixel_2326/gring pixel_2326/VDD pixel_2326/GND pixel_2326/VREF pixel_2326/ROW_SEL
+ pixel_2326/NB1 pixel_2326/VBIAS pixel_2326/NB2 pixel_2326/AMP_IN pixel_2326/SF_IB
+ pixel_2326/PIX_OUT pixel_2326/CSA_VREF pixel
Xpixel_2315 pixel_2315/gring pixel_2315/VDD pixel_2315/GND pixel_2315/VREF pixel_2315/ROW_SEL
+ pixel_2315/NB1 pixel_2315/VBIAS pixel_2315/NB2 pixel_2315/AMP_IN pixel_2315/SF_IB
+ pixel_2315/PIX_OUT pixel_2315/CSA_VREF pixel
Xpixel_2304 pixel_2304/gring pixel_2304/VDD pixel_2304/GND pixel_2304/VREF pixel_2304/ROW_SEL
+ pixel_2304/NB1 pixel_2304/VBIAS pixel_2304/NB2 pixel_2304/AMP_IN pixel_2304/SF_IB
+ pixel_2304/PIX_OUT pixel_2304/CSA_VREF pixel
Xpixel_3049 pixel_3049/gring pixel_3049/VDD pixel_3049/GND pixel_3049/VREF pixel_3049/ROW_SEL
+ pixel_3049/NB1 pixel_3049/VBIAS pixel_3049/NB2 pixel_3049/AMP_IN pixel_3049/SF_IB
+ pixel_3049/PIX_OUT pixel_3049/CSA_VREF pixel
Xpixel_1625 pixel_1625/gring pixel_1625/VDD pixel_1625/GND pixel_1625/VREF pixel_1625/ROW_SEL
+ pixel_1625/NB1 pixel_1625/VBIAS pixel_1625/NB2 pixel_1625/AMP_IN pixel_1625/SF_IB
+ pixel_1625/PIX_OUT pixel_1625/CSA_VREF pixel
Xpixel_1614 pixel_1614/gring pixel_1614/VDD pixel_1614/GND pixel_1614/VREF pixel_1614/ROW_SEL
+ pixel_1614/NB1 pixel_1614/VBIAS pixel_1614/NB2 pixel_1614/AMP_IN pixel_1614/SF_IB
+ pixel_1614/PIX_OUT pixel_1614/CSA_VREF pixel
Xpixel_1603 pixel_1603/gring pixel_1603/VDD pixel_1603/GND pixel_1603/VREF pixel_1603/ROW_SEL
+ pixel_1603/NB1 pixel_1603/VBIAS pixel_1603/NB2 pixel_1603/AMP_IN pixel_1603/SF_IB
+ pixel_1603/PIX_OUT pixel_1603/CSA_VREF pixel
Xpixel_2359 pixel_2359/gring pixel_2359/VDD pixel_2359/GND pixel_2359/VREF pixel_2359/ROW_SEL
+ pixel_2359/NB1 pixel_2359/VBIAS pixel_2359/NB2 pixel_2359/AMP_IN pixel_2359/SF_IB
+ pixel_2359/PIX_OUT pixel_2359/CSA_VREF pixel
Xpixel_2348 pixel_2348/gring pixel_2348/VDD pixel_2348/GND pixel_2348/VREF pixel_2348/ROW_SEL
+ pixel_2348/NB1 pixel_2348/VBIAS pixel_2348/NB2 pixel_2348/AMP_IN pixel_2348/SF_IB
+ pixel_2348/PIX_OUT pixel_2348/CSA_VREF pixel
Xpixel_2337 pixel_2337/gring pixel_2337/VDD pixel_2337/GND pixel_2337/VREF pixel_2337/ROW_SEL
+ pixel_2337/NB1 pixel_2337/VBIAS pixel_2337/NB2 pixel_2337/AMP_IN pixel_2337/SF_IB
+ pixel_2337/PIX_OUT pixel_2337/CSA_VREF pixel
Xpixel_1658 pixel_1658/gring pixel_1658/VDD pixel_1658/GND pixel_1658/VREF pixel_1658/ROW_SEL
+ pixel_1658/NB1 pixel_1658/VBIAS pixel_1658/NB2 pixel_1658/AMP_IN pixel_1658/SF_IB
+ pixel_1658/PIX_OUT pixel_1658/CSA_VREF pixel
Xpixel_1647 pixel_1647/gring pixel_1647/VDD pixel_1647/GND pixel_1647/VREF pixel_1647/ROW_SEL
+ pixel_1647/NB1 pixel_1647/VBIAS pixel_1647/NB2 pixel_1647/AMP_IN pixel_1647/SF_IB
+ pixel_1647/PIX_OUT pixel_1647/CSA_VREF pixel
Xpixel_1636 pixel_1636/gring pixel_1636/VDD pixel_1636/GND pixel_1636/VREF pixel_1636/ROW_SEL
+ pixel_1636/NB1 pixel_1636/VBIAS pixel_1636/NB2 pixel_1636/AMP_IN pixel_1636/SF_IB
+ pixel_1636/PIX_OUT pixel_1636/CSA_VREF pixel
Xpixel_1669 pixel_1669/gring pixel_1669/VDD pixel_1669/GND pixel_1669/VREF pixel_1669/ROW_SEL
+ pixel_1669/NB1 pixel_1669/VBIAS pixel_1669/NB2 pixel_1669/AMP_IN pixel_1669/SF_IB
+ pixel_1669/PIX_OUT pixel_1669/CSA_VREF pixel
Xpixel_9900 pixel_9900/gring pixel_9900/VDD pixel_9900/GND pixel_9900/VREF pixel_9900/ROW_SEL
+ pixel_9900/NB1 pixel_9900/VBIAS pixel_9900/NB2 pixel_9900/AMP_IN pixel_9900/SF_IB
+ pixel_9900/PIX_OUT pixel_9900/CSA_VREF pixel
Xpixel_9933 pixel_9933/gring pixel_9933/VDD pixel_9933/GND pixel_9933/VREF pixel_9933/ROW_SEL
+ pixel_9933/NB1 pixel_9933/VBIAS pixel_9933/NB2 pixel_9933/AMP_IN pixel_9933/SF_IB
+ pixel_9933/PIX_OUT pixel_9933/CSA_VREF pixel
Xpixel_9922 pixel_9922/gring pixel_9922/VDD pixel_9922/GND pixel_9922/VREF pixel_9922/ROW_SEL
+ pixel_9922/NB1 pixel_9922/VBIAS pixel_9922/NB2 pixel_9922/AMP_IN pixel_9922/SF_IB
+ pixel_9922/PIX_OUT pixel_9922/CSA_VREF pixel
Xpixel_9911 pixel_9911/gring pixel_9911/VDD pixel_9911/GND pixel_9911/VREF pixel_9911/ROW_SEL
+ pixel_9911/NB1 pixel_9911/VBIAS pixel_9911/NB2 pixel_9911/AMP_IN pixel_9911/SF_IB
+ pixel_9911/PIX_OUT pixel_9911/CSA_VREF pixel
Xpixel_9944 pixel_9944/gring pixel_9944/VDD pixel_9944/GND pixel_9944/VREF pixel_9944/ROW_SEL
+ pixel_9944/NB1 pixel_9944/VBIAS pixel_9944/NB2 pixel_9944/AMP_IN pixel_9944/SF_IB
+ pixel_9944/PIX_OUT pixel_9944/CSA_VREF pixel
Xpixel_9955 pixel_9955/gring pixel_9955/VDD pixel_9955/GND pixel_9955/VREF pixel_9955/ROW_SEL
+ pixel_9955/NB1 pixel_9955/VBIAS pixel_9955/NB2 pixel_9955/AMP_IN pixel_9955/SF_IB
+ pixel_9955/PIX_OUT pixel_9955/CSA_VREF pixel
Xpixel_9966 pixel_9966/gring pixel_9966/VDD pixel_9966/GND pixel_9966/VREF pixel_9966/ROW_SEL
+ pixel_9966/NB1 pixel_9966/VBIAS pixel_9966/NB2 pixel_9966/AMP_IN pixel_9966/SF_IB
+ pixel_9966/PIX_OUT pixel_9966/CSA_VREF pixel
Xpixel_9977 pixel_9977/gring pixel_9977/VDD pixel_9977/GND pixel_9977/VREF pixel_9977/ROW_SEL
+ pixel_9977/NB1 pixel_9977/VBIAS pixel_9977/NB2 pixel_9977/AMP_IN pixel_9977/SF_IB
+ pixel_9977/PIX_OUT pixel_9977/CSA_VREF pixel
Xpixel_9988 pixel_9988/gring pixel_9988/VDD pixel_9988/GND pixel_9988/VREF pixel_9988/ROW_SEL
+ pixel_9988/NB1 pixel_9988/VBIAS pixel_9988/NB2 pixel_9988/AMP_IN pixel_9988/SF_IB
+ pixel_9988/PIX_OUT pixel_9988/CSA_VREF pixel
Xpixel_9999 pixel_9999/gring pixel_9999/VDD pixel_9999/GND pixel_9999/VREF pixel_9999/ROW_SEL
+ pixel_9999/NB1 pixel_9999/VBIAS pixel_9999/NB2 pixel_9999/AMP_IN pixel_9999/SF_IB
+ pixel_9999/PIX_OUT pixel_9999/CSA_VREF pixel
Xpixel_4240 pixel_4240/gring pixel_4240/VDD pixel_4240/GND pixel_4240/VREF pixel_4240/ROW_SEL
+ pixel_4240/NB1 pixel_4240/VBIAS pixel_4240/NB2 pixel_4240/AMP_IN pixel_4240/SF_IB
+ pixel_4240/PIX_OUT pixel_4240/CSA_VREF pixel
Xpixel_4251 pixel_4251/gring pixel_4251/VDD pixel_4251/GND pixel_4251/VREF pixel_4251/ROW_SEL
+ pixel_4251/NB1 pixel_4251/VBIAS pixel_4251/NB2 pixel_4251/AMP_IN pixel_4251/SF_IB
+ pixel_4251/PIX_OUT pixel_4251/CSA_VREF pixel
Xpixel_4262 pixel_4262/gring pixel_4262/VDD pixel_4262/GND pixel_4262/VREF pixel_4262/ROW_SEL
+ pixel_4262/NB1 pixel_4262/VBIAS pixel_4262/NB2 pixel_4262/AMP_IN pixel_4262/SF_IB
+ pixel_4262/PIX_OUT pixel_4262/CSA_VREF pixel
Xpixel_290 pixel_290/gring pixel_290/VDD pixel_290/GND pixel_290/VREF pixel_290/ROW_SEL
+ pixel_290/NB1 pixel_290/VBIAS pixel_290/NB2 pixel_290/AMP_IN pixel_290/SF_IB pixel_290/PIX_OUT
+ pixel_290/CSA_VREF pixel
Xpixel_3561 pixel_3561/gring pixel_3561/VDD pixel_3561/GND pixel_3561/VREF pixel_3561/ROW_SEL
+ pixel_3561/NB1 pixel_3561/VBIAS pixel_3561/NB2 pixel_3561/AMP_IN pixel_3561/SF_IB
+ pixel_3561/PIX_OUT pixel_3561/CSA_VREF pixel
Xpixel_3550 pixel_3550/gring pixel_3550/VDD pixel_3550/GND pixel_3550/VREF pixel_3550/ROW_SEL
+ pixel_3550/NB1 pixel_3550/VBIAS pixel_3550/NB2 pixel_3550/AMP_IN pixel_3550/SF_IB
+ pixel_3550/PIX_OUT pixel_3550/CSA_VREF pixel
Xpixel_4273 pixel_4273/gring pixel_4273/VDD pixel_4273/GND pixel_4273/VREF pixel_4273/ROW_SEL
+ pixel_4273/NB1 pixel_4273/VBIAS pixel_4273/NB2 pixel_4273/AMP_IN pixel_4273/SF_IB
+ pixel_4273/PIX_OUT pixel_4273/CSA_VREF pixel
Xpixel_4284 pixel_4284/gring pixel_4284/VDD pixel_4284/GND pixel_4284/VREF pixel_4284/ROW_SEL
+ pixel_4284/NB1 pixel_4284/VBIAS pixel_4284/NB2 pixel_4284/AMP_IN pixel_4284/SF_IB
+ pixel_4284/PIX_OUT pixel_4284/CSA_VREF pixel
Xpixel_4295 pixel_4295/gring pixel_4295/VDD pixel_4295/GND pixel_4295/VREF pixel_4295/ROW_SEL
+ pixel_4295/NB1 pixel_4295/VBIAS pixel_4295/NB2 pixel_4295/AMP_IN pixel_4295/SF_IB
+ pixel_4295/PIX_OUT pixel_4295/CSA_VREF pixel
Xpixel_3594 pixel_3594/gring pixel_3594/VDD pixel_3594/GND pixel_3594/VREF pixel_3594/ROW_SEL
+ pixel_3594/NB1 pixel_3594/VBIAS pixel_3594/NB2 pixel_3594/AMP_IN pixel_3594/SF_IB
+ pixel_3594/PIX_OUT pixel_3594/CSA_VREF pixel
Xpixel_3583 pixel_3583/gring pixel_3583/VDD pixel_3583/GND pixel_3583/VREF pixel_3583/ROW_SEL
+ pixel_3583/NB1 pixel_3583/VBIAS pixel_3583/NB2 pixel_3583/AMP_IN pixel_3583/SF_IB
+ pixel_3583/PIX_OUT pixel_3583/CSA_VREF pixel
Xpixel_3572 pixel_3572/gring pixel_3572/VDD pixel_3572/GND pixel_3572/VREF pixel_3572/ROW_SEL
+ pixel_3572/NB1 pixel_3572/VBIAS pixel_3572/NB2 pixel_3572/AMP_IN pixel_3572/SF_IB
+ pixel_3572/PIX_OUT pixel_3572/CSA_VREF pixel
Xpixel_2882 pixel_2882/gring pixel_2882/VDD pixel_2882/GND pixel_2882/VREF pixel_2882/ROW_SEL
+ pixel_2882/NB1 pixel_2882/VBIAS pixel_2882/NB2 pixel_2882/AMP_IN pixel_2882/SF_IB
+ pixel_2882/PIX_OUT pixel_2882/CSA_VREF pixel
Xpixel_2871 pixel_2871/gring pixel_2871/VDD pixel_2871/GND pixel_2871/VREF pixel_2871/ROW_SEL
+ pixel_2871/NB1 pixel_2871/VBIAS pixel_2871/NB2 pixel_2871/AMP_IN pixel_2871/SF_IB
+ pixel_2871/PIX_OUT pixel_2871/CSA_VREF pixel
Xpixel_2860 pixel_2860/gring pixel_2860/VDD pixel_2860/GND pixel_2860/VREF pixel_2860/ROW_SEL
+ pixel_2860/NB1 pixel_2860/VBIAS pixel_2860/NB2 pixel_2860/AMP_IN pixel_2860/SF_IB
+ pixel_2860/PIX_OUT pixel_2860/CSA_VREF pixel
Xpixel_2893 pixel_2893/gring pixel_2893/VDD pixel_2893/GND pixel_2893/VREF pixel_2893/ROW_SEL
+ pixel_2893/NB1 pixel_2893/VBIAS pixel_2893/NB2 pixel_2893/AMP_IN pixel_2893/SF_IB
+ pixel_2893/PIX_OUT pixel_2893/CSA_VREF pixel
Xpixel_9229 pixel_9229/gring pixel_9229/VDD pixel_9229/GND pixel_9229/VREF pixel_9229/ROW_SEL
+ pixel_9229/NB1 pixel_9229/VBIAS pixel_9229/NB2 pixel_9229/AMP_IN pixel_9229/SF_IB
+ pixel_9229/PIX_OUT pixel_9229/CSA_VREF pixel
Xpixel_9218 pixel_9218/gring pixel_9218/VDD pixel_9218/GND pixel_9218/VREF pixel_9218/ROW_SEL
+ pixel_9218/NB1 pixel_9218/VBIAS pixel_9218/NB2 pixel_9218/AMP_IN pixel_9218/SF_IB
+ pixel_9218/PIX_OUT pixel_9218/CSA_VREF pixel
Xpixel_9207 pixel_9207/gring pixel_9207/VDD pixel_9207/GND pixel_9207/VREF pixel_9207/ROW_SEL
+ pixel_9207/NB1 pixel_9207/VBIAS pixel_9207/NB2 pixel_9207/AMP_IN pixel_9207/SF_IB
+ pixel_9207/PIX_OUT pixel_9207/CSA_VREF pixel
Xpixel_8517 pixel_8517/gring pixel_8517/VDD pixel_8517/GND pixel_8517/VREF pixel_8517/ROW_SEL
+ pixel_8517/NB1 pixel_8517/VBIAS pixel_8517/NB2 pixel_8517/AMP_IN pixel_8517/SF_IB
+ pixel_8517/PIX_OUT pixel_8517/CSA_VREF pixel
Xpixel_8506 pixel_8506/gring pixel_8506/VDD pixel_8506/GND pixel_8506/VREF pixel_8506/ROW_SEL
+ pixel_8506/NB1 pixel_8506/VBIAS pixel_8506/NB2 pixel_8506/AMP_IN pixel_8506/SF_IB
+ pixel_8506/PIX_OUT pixel_8506/CSA_VREF pixel
Xpixel_8539 pixel_8539/gring pixel_8539/VDD pixel_8539/GND pixel_8539/VREF pixel_8539/ROW_SEL
+ pixel_8539/NB1 pixel_8539/VBIAS pixel_8539/NB2 pixel_8539/AMP_IN pixel_8539/SF_IB
+ pixel_8539/PIX_OUT pixel_8539/CSA_VREF pixel
Xpixel_8528 pixel_8528/gring pixel_8528/VDD pixel_8528/GND pixel_8528/VREF pixel_8528/ROW_SEL
+ pixel_8528/NB1 pixel_8528/VBIAS pixel_8528/NB2 pixel_8528/AMP_IN pixel_8528/SF_IB
+ pixel_8528/PIX_OUT pixel_8528/CSA_VREF pixel
Xpixel_7805 pixel_7805/gring pixel_7805/VDD pixel_7805/GND pixel_7805/VREF pixel_7805/ROW_SEL
+ pixel_7805/NB1 pixel_7805/VBIAS pixel_7805/NB2 pixel_7805/AMP_IN pixel_7805/SF_IB
+ pixel_7805/PIX_OUT pixel_7805/CSA_VREF pixel
Xpixel_7816 pixel_7816/gring pixel_7816/VDD pixel_7816/GND pixel_7816/VREF pixel_7816/ROW_SEL
+ pixel_7816/NB1 pixel_7816/VBIAS pixel_7816/NB2 pixel_7816/AMP_IN pixel_7816/SF_IB
+ pixel_7816/PIX_OUT pixel_7816/CSA_VREF pixel
Xpixel_7827 pixel_7827/gring pixel_7827/VDD pixel_7827/GND pixel_7827/VREF pixel_7827/ROW_SEL
+ pixel_7827/NB1 pixel_7827/VBIAS pixel_7827/NB2 pixel_7827/AMP_IN pixel_7827/SF_IB
+ pixel_7827/PIX_OUT pixel_7827/CSA_VREF pixel
Xpixel_7838 pixel_7838/gring pixel_7838/VDD pixel_7838/GND pixel_7838/VREF pixel_7838/ROW_SEL
+ pixel_7838/NB1 pixel_7838/VBIAS pixel_7838/NB2 pixel_7838/AMP_IN pixel_7838/SF_IB
+ pixel_7838/PIX_OUT pixel_7838/CSA_VREF pixel
Xpixel_7849 pixel_7849/gring pixel_7849/VDD pixel_7849/GND pixel_7849/VREF pixel_7849/ROW_SEL
+ pixel_7849/NB1 pixel_7849/VBIAS pixel_7849/NB2 pixel_7849/AMP_IN pixel_7849/SF_IB
+ pixel_7849/PIX_OUT pixel_7849/CSA_VREF pixel
Xpixel_2101 pixel_2101/gring pixel_2101/VDD pixel_2101/GND pixel_2101/VREF pixel_2101/ROW_SEL
+ pixel_2101/NB1 pixel_2101/VBIAS pixel_2101/NB2 pixel_2101/AMP_IN pixel_2101/SF_IB
+ pixel_2101/PIX_OUT pixel_2101/CSA_VREF pixel
Xpixel_1400 pixel_1400/gring pixel_1400/VDD pixel_1400/GND pixel_1400/VREF pixel_1400/ROW_SEL
+ pixel_1400/NB1 pixel_1400/VBIAS pixel_1400/NB2 pixel_1400/AMP_IN pixel_1400/SF_IB
+ pixel_1400/PIX_OUT pixel_1400/CSA_VREF pixel
Xpixel_2145 pixel_2145/gring pixel_2145/VDD pixel_2145/GND pixel_2145/VREF pixel_2145/ROW_SEL
+ pixel_2145/NB1 pixel_2145/VBIAS pixel_2145/NB2 pixel_2145/AMP_IN pixel_2145/SF_IB
+ pixel_2145/PIX_OUT pixel_2145/CSA_VREF pixel
Xpixel_2134 pixel_2134/gring pixel_2134/VDD pixel_2134/GND pixel_2134/VREF pixel_2134/ROW_SEL
+ pixel_2134/NB1 pixel_2134/VBIAS pixel_2134/NB2 pixel_2134/AMP_IN pixel_2134/SF_IB
+ pixel_2134/PIX_OUT pixel_2134/CSA_VREF pixel
Xpixel_2123 pixel_2123/gring pixel_2123/VDD pixel_2123/GND pixel_2123/VREF pixel_2123/ROW_SEL
+ pixel_2123/NB1 pixel_2123/VBIAS pixel_2123/NB2 pixel_2123/AMP_IN pixel_2123/SF_IB
+ pixel_2123/PIX_OUT pixel_2123/CSA_VREF pixel
Xpixel_2112 pixel_2112/gring pixel_2112/VDD pixel_2112/GND pixel_2112/VREF pixel_2112/ROW_SEL
+ pixel_2112/NB1 pixel_2112/VBIAS pixel_2112/NB2 pixel_2112/AMP_IN pixel_2112/SF_IB
+ pixel_2112/PIX_OUT pixel_2112/CSA_VREF pixel
Xpixel_1433 pixel_1433/gring pixel_1433/VDD pixel_1433/GND pixel_1433/VREF pixel_1433/ROW_SEL
+ pixel_1433/NB1 pixel_1433/VBIAS pixel_1433/NB2 pixel_1433/AMP_IN pixel_1433/SF_IB
+ pixel_1433/PIX_OUT pixel_1433/CSA_VREF pixel
Xpixel_1422 pixel_1422/gring pixel_1422/VDD pixel_1422/GND pixel_1422/VREF pixel_1422/ROW_SEL
+ pixel_1422/NB1 pixel_1422/VBIAS pixel_1422/NB2 pixel_1422/AMP_IN pixel_1422/SF_IB
+ pixel_1422/PIX_OUT pixel_1422/CSA_VREF pixel
Xpixel_1411 pixel_1411/gring pixel_1411/VDD pixel_1411/GND pixel_1411/VREF pixel_1411/ROW_SEL
+ pixel_1411/NB1 pixel_1411/VBIAS pixel_1411/NB2 pixel_1411/AMP_IN pixel_1411/SF_IB
+ pixel_1411/PIX_OUT pixel_1411/CSA_VREF pixel
Xpixel_2178 pixel_2178/gring pixel_2178/VDD pixel_2178/GND pixel_2178/VREF pixel_2178/ROW_SEL
+ pixel_2178/NB1 pixel_2178/VBIAS pixel_2178/NB2 pixel_2178/AMP_IN pixel_2178/SF_IB
+ pixel_2178/PIX_OUT pixel_2178/CSA_VREF pixel
Xpixel_2167 pixel_2167/gring pixel_2167/VDD pixel_2167/GND pixel_2167/VREF pixel_2167/ROW_SEL
+ pixel_2167/NB1 pixel_2167/VBIAS pixel_2167/NB2 pixel_2167/AMP_IN pixel_2167/SF_IB
+ pixel_2167/PIX_OUT pixel_2167/CSA_VREF pixel
Xpixel_2156 pixel_2156/gring pixel_2156/VDD pixel_2156/GND pixel_2156/VREF pixel_2156/ROW_SEL
+ pixel_2156/NB1 pixel_2156/VBIAS pixel_2156/NB2 pixel_2156/AMP_IN pixel_2156/SF_IB
+ pixel_2156/PIX_OUT pixel_2156/CSA_VREF pixel
Xpixel_1466 pixel_1466/gring pixel_1466/VDD pixel_1466/GND pixel_1466/VREF pixel_1466/ROW_SEL
+ pixel_1466/NB1 pixel_1466/VBIAS pixel_1466/NB2 pixel_1466/AMP_IN pixel_1466/SF_IB
+ pixel_1466/PIX_OUT pixel_1466/CSA_VREF pixel
Xpixel_1455 pixel_1455/gring pixel_1455/VDD pixel_1455/GND pixel_1455/VREF pixel_1455/ROW_SEL
+ pixel_1455/NB1 pixel_1455/VBIAS pixel_1455/NB2 pixel_1455/AMP_IN pixel_1455/SF_IB
+ pixel_1455/PIX_OUT pixel_1455/CSA_VREF pixel
Xpixel_1444 pixel_1444/gring pixel_1444/VDD pixel_1444/GND pixel_1444/VREF pixel_1444/ROW_SEL
+ pixel_1444/NB1 pixel_1444/VBIAS pixel_1444/NB2 pixel_1444/AMP_IN pixel_1444/SF_IB
+ pixel_1444/PIX_OUT pixel_1444/CSA_VREF pixel
Xpixel_2189 pixel_2189/gring pixel_2189/VDD pixel_2189/GND pixel_2189/VREF pixel_2189/ROW_SEL
+ pixel_2189/NB1 pixel_2189/VBIAS pixel_2189/NB2 pixel_2189/AMP_IN pixel_2189/SF_IB
+ pixel_2189/PIX_OUT pixel_2189/CSA_VREF pixel
Xpixel_1499 pixel_1499/gring pixel_1499/VDD pixel_1499/GND pixel_1499/VREF pixel_1499/ROW_SEL
+ pixel_1499/NB1 pixel_1499/VBIAS pixel_1499/NB2 pixel_1499/AMP_IN pixel_1499/SF_IB
+ pixel_1499/PIX_OUT pixel_1499/CSA_VREF pixel
Xpixel_1488 pixel_1488/gring pixel_1488/VDD pixel_1488/GND pixel_1488/VREF pixel_1488/ROW_SEL
+ pixel_1488/NB1 pixel_1488/VBIAS pixel_1488/NB2 pixel_1488/AMP_IN pixel_1488/SF_IB
+ pixel_1488/PIX_OUT pixel_1488/CSA_VREF pixel
Xpixel_1477 pixel_1477/gring pixel_1477/VDD pixel_1477/GND pixel_1477/VREF pixel_1477/ROW_SEL
+ pixel_1477/NB1 pixel_1477/VBIAS pixel_1477/NB2 pixel_1477/AMP_IN pixel_1477/SF_IB
+ pixel_1477/PIX_OUT pixel_1477/CSA_VREF pixel
Xpixel_9730 pixel_9730/gring pixel_9730/VDD pixel_9730/GND pixel_9730/VREF pixel_9730/ROW_SEL
+ pixel_9730/NB1 pixel_9730/VBIAS pixel_9730/NB2 pixel_9730/AMP_IN pixel_9730/SF_IB
+ pixel_9730/PIX_OUT pixel_9730/CSA_VREF pixel
Xpixel_9741 pixel_9741/gring pixel_9741/VDD pixel_9741/GND pixel_9741/VREF pixel_9741/ROW_SEL
+ pixel_9741/NB1 pixel_9741/VBIAS pixel_9741/NB2 pixel_9741/AMP_IN pixel_9741/SF_IB
+ pixel_9741/PIX_OUT pixel_9741/CSA_VREF pixel
Xpixel_9752 pixel_9752/gring pixel_9752/VDD pixel_9752/GND pixel_9752/VREF pixel_9752/ROW_SEL
+ pixel_9752/NB1 pixel_9752/VBIAS pixel_9752/NB2 pixel_9752/AMP_IN pixel_9752/SF_IB
+ pixel_9752/PIX_OUT pixel_9752/CSA_VREF pixel
Xpixel_9763 pixel_9763/gring pixel_9763/VDD pixel_9763/GND pixel_9763/VREF pixel_9763/ROW_SEL
+ pixel_9763/NB1 pixel_9763/VBIAS pixel_9763/NB2 pixel_9763/AMP_IN pixel_9763/SF_IB
+ pixel_9763/PIX_OUT pixel_9763/CSA_VREF pixel
Xpixel_9774 pixel_9774/gring pixel_9774/VDD pixel_9774/GND pixel_9774/VREF pixel_9774/ROW_SEL
+ pixel_9774/NB1 pixel_9774/VBIAS pixel_9774/NB2 pixel_9774/AMP_IN pixel_9774/SF_IB
+ pixel_9774/PIX_OUT pixel_9774/CSA_VREF pixel
Xpixel_9785 pixel_9785/gring pixel_9785/VDD pixel_9785/GND pixel_9785/VREF pixel_9785/ROW_SEL
+ pixel_9785/NB1 pixel_9785/VBIAS pixel_9785/NB2 pixel_9785/AMP_IN pixel_9785/SF_IB
+ pixel_9785/PIX_OUT pixel_9785/CSA_VREF pixel
Xpixel_9796 pixel_9796/gring pixel_9796/VDD pixel_9796/GND pixel_9796/VREF pixel_9796/ROW_SEL
+ pixel_9796/NB1 pixel_9796/VBIAS pixel_9796/NB2 pixel_9796/AMP_IN pixel_9796/SF_IB
+ pixel_9796/PIX_OUT pixel_9796/CSA_VREF pixel
Xpixel_4070 pixel_4070/gring pixel_4070/VDD pixel_4070/GND pixel_4070/VREF pixel_4070/ROW_SEL
+ pixel_4070/NB1 pixel_4070/VBIAS pixel_4070/NB2 pixel_4070/AMP_IN pixel_4070/SF_IB
+ pixel_4070/PIX_OUT pixel_4070/CSA_VREF pixel
Xpixel_4081 pixel_4081/gring pixel_4081/VDD pixel_4081/GND pixel_4081/VREF pixel_4081/ROW_SEL
+ pixel_4081/NB1 pixel_4081/VBIAS pixel_4081/NB2 pixel_4081/AMP_IN pixel_4081/SF_IB
+ pixel_4081/PIX_OUT pixel_4081/CSA_VREF pixel
Xpixel_4092 pixel_4092/gring pixel_4092/VDD pixel_4092/GND pixel_4092/VREF pixel_4092/ROW_SEL
+ pixel_4092/NB1 pixel_4092/VBIAS pixel_4092/NB2 pixel_4092/AMP_IN pixel_4092/SF_IB
+ pixel_4092/PIX_OUT pixel_4092/CSA_VREF pixel
Xpixel_3391 pixel_3391/gring pixel_3391/VDD pixel_3391/GND pixel_3391/VREF pixel_3391/ROW_SEL
+ pixel_3391/NB1 pixel_3391/VBIAS pixel_3391/NB2 pixel_3391/AMP_IN pixel_3391/SF_IB
+ pixel_3391/PIX_OUT pixel_3391/CSA_VREF pixel
Xpixel_3380 pixel_3380/gring pixel_3380/VDD pixel_3380/GND pixel_3380/VREF pixel_3380/ROW_SEL
+ pixel_3380/NB1 pixel_3380/VBIAS pixel_3380/NB2 pixel_3380/AMP_IN pixel_3380/SF_IB
+ pixel_3380/PIX_OUT pixel_3380/CSA_VREF pixel
Xpixel_2690 pixel_2690/gring pixel_2690/VDD pixel_2690/GND pixel_2690/VREF pixel_2690/ROW_SEL
+ pixel_2690/NB1 pixel_2690/VBIAS pixel_2690/NB2 pixel_2690/AMP_IN pixel_2690/SF_IB
+ pixel_2690/PIX_OUT pixel_2690/CSA_VREF pixel
Xpixel_9004 pixel_9004/gring pixel_9004/VDD pixel_9004/GND pixel_9004/VREF pixel_9004/ROW_SEL
+ pixel_9004/NB1 pixel_9004/VBIAS pixel_9004/NB2 pixel_9004/AMP_IN pixel_9004/SF_IB
+ pixel_9004/PIX_OUT pixel_9004/CSA_VREF pixel
Xpixel_9037 pixel_9037/gring pixel_9037/VDD pixel_9037/GND pixel_9037/VREF pixel_9037/ROW_SEL
+ pixel_9037/NB1 pixel_9037/VBIAS pixel_9037/NB2 pixel_9037/AMP_IN pixel_9037/SF_IB
+ pixel_9037/PIX_OUT pixel_9037/CSA_VREF pixel
Xpixel_9026 pixel_9026/gring pixel_9026/VDD pixel_9026/GND pixel_9026/VREF pixel_9026/ROW_SEL
+ pixel_9026/NB1 pixel_9026/VBIAS pixel_9026/NB2 pixel_9026/AMP_IN pixel_9026/SF_IB
+ pixel_9026/PIX_OUT pixel_9026/CSA_VREF pixel
Xpixel_9015 pixel_9015/gring pixel_9015/VDD pixel_9015/GND pixel_9015/VREF pixel_9015/ROW_SEL
+ pixel_9015/NB1 pixel_9015/VBIAS pixel_9015/NB2 pixel_9015/AMP_IN pixel_9015/SF_IB
+ pixel_9015/PIX_OUT pixel_9015/CSA_VREF pixel
Xpixel_9059 pixel_9059/gring pixel_9059/VDD pixel_9059/GND pixel_9059/VREF pixel_9059/ROW_SEL
+ pixel_9059/NB1 pixel_9059/VBIAS pixel_9059/NB2 pixel_9059/AMP_IN pixel_9059/SF_IB
+ pixel_9059/PIX_OUT pixel_9059/CSA_VREF pixel
Xpixel_9048 pixel_9048/gring pixel_9048/VDD pixel_9048/GND pixel_9048/VREF pixel_9048/ROW_SEL
+ pixel_9048/NB1 pixel_9048/VBIAS pixel_9048/NB2 pixel_9048/AMP_IN pixel_9048/SF_IB
+ pixel_9048/PIX_OUT pixel_9048/CSA_VREF pixel
Xpixel_8303 pixel_8303/gring pixel_8303/VDD pixel_8303/GND pixel_8303/VREF pixel_8303/ROW_SEL
+ pixel_8303/NB1 pixel_8303/VBIAS pixel_8303/NB2 pixel_8303/AMP_IN pixel_8303/SF_IB
+ pixel_8303/PIX_OUT pixel_8303/CSA_VREF pixel
Xpixel_8314 pixel_8314/gring pixel_8314/VDD pixel_8314/GND pixel_8314/VREF pixel_8314/ROW_SEL
+ pixel_8314/NB1 pixel_8314/VBIAS pixel_8314/NB2 pixel_8314/AMP_IN pixel_8314/SF_IB
+ pixel_8314/PIX_OUT pixel_8314/CSA_VREF pixel
Xpixel_8325 pixel_8325/gring pixel_8325/VDD pixel_8325/GND pixel_8325/VREF pixel_8325/ROW_SEL
+ pixel_8325/NB1 pixel_8325/VBIAS pixel_8325/NB2 pixel_8325/AMP_IN pixel_8325/SF_IB
+ pixel_8325/PIX_OUT pixel_8325/CSA_VREF pixel
Xpixel_8336 pixel_8336/gring pixel_8336/VDD pixel_8336/GND pixel_8336/VREF pixel_8336/ROW_SEL
+ pixel_8336/NB1 pixel_8336/VBIAS pixel_8336/NB2 pixel_8336/AMP_IN pixel_8336/SF_IB
+ pixel_8336/PIX_OUT pixel_8336/CSA_VREF pixel
Xpixel_8347 pixel_8347/gring pixel_8347/VDD pixel_8347/GND pixel_8347/VREF pixel_8347/ROW_SEL
+ pixel_8347/NB1 pixel_8347/VBIAS pixel_8347/NB2 pixel_8347/AMP_IN pixel_8347/SF_IB
+ pixel_8347/PIX_OUT pixel_8347/CSA_VREF pixel
Xpixel_8358 pixel_8358/gring pixel_8358/VDD pixel_8358/GND pixel_8358/VREF pixel_8358/ROW_SEL
+ pixel_8358/NB1 pixel_8358/VBIAS pixel_8358/NB2 pixel_8358/AMP_IN pixel_8358/SF_IB
+ pixel_8358/PIX_OUT pixel_8358/CSA_VREF pixel
Xpixel_8369 pixel_8369/gring pixel_8369/VDD pixel_8369/GND pixel_8369/VREF pixel_8369/ROW_SEL
+ pixel_8369/NB1 pixel_8369/VBIAS pixel_8369/NB2 pixel_8369/AMP_IN pixel_8369/SF_IB
+ pixel_8369/PIX_OUT pixel_8369/CSA_VREF pixel
Xpixel_7602 pixel_7602/gring pixel_7602/VDD pixel_7602/GND pixel_7602/VREF pixel_7602/ROW_SEL
+ pixel_7602/NB1 pixel_7602/VBIAS pixel_7602/NB2 pixel_7602/AMP_IN pixel_7602/SF_IB
+ pixel_7602/PIX_OUT pixel_7602/CSA_VREF pixel
Xpixel_7613 pixel_7613/gring pixel_7613/VDD pixel_7613/GND pixel_7613/VREF pixel_7613/ROW_SEL
+ pixel_7613/NB1 pixel_7613/VBIAS pixel_7613/NB2 pixel_7613/AMP_IN pixel_7613/SF_IB
+ pixel_7613/PIX_OUT pixel_7613/CSA_VREF pixel
Xpixel_7624 pixel_7624/gring pixel_7624/VDD pixel_7624/GND pixel_7624/VREF pixel_7624/ROW_SEL
+ pixel_7624/NB1 pixel_7624/VBIAS pixel_7624/NB2 pixel_7624/AMP_IN pixel_7624/SF_IB
+ pixel_7624/PIX_OUT pixel_7624/CSA_VREF pixel
Xpixel_7635 pixel_7635/gring pixel_7635/VDD pixel_7635/GND pixel_7635/VREF pixel_7635/ROW_SEL
+ pixel_7635/NB1 pixel_7635/VBIAS pixel_7635/NB2 pixel_7635/AMP_IN pixel_7635/SF_IB
+ pixel_7635/PIX_OUT pixel_7635/CSA_VREF pixel
Xpixel_7646 pixel_7646/gring pixel_7646/VDD pixel_7646/GND pixel_7646/VREF pixel_7646/ROW_SEL
+ pixel_7646/NB1 pixel_7646/VBIAS pixel_7646/NB2 pixel_7646/AMP_IN pixel_7646/SF_IB
+ pixel_7646/PIX_OUT pixel_7646/CSA_VREF pixel
Xpixel_7657 pixel_7657/gring pixel_7657/VDD pixel_7657/GND pixel_7657/VREF pixel_7657/ROW_SEL
+ pixel_7657/NB1 pixel_7657/VBIAS pixel_7657/NB2 pixel_7657/AMP_IN pixel_7657/SF_IB
+ pixel_7657/PIX_OUT pixel_7657/CSA_VREF pixel
Xpixel_6901 pixel_6901/gring pixel_6901/VDD pixel_6901/GND pixel_6901/VREF pixel_6901/ROW_SEL
+ pixel_6901/NB1 pixel_6901/VBIAS pixel_6901/NB2 pixel_6901/AMP_IN pixel_6901/SF_IB
+ pixel_6901/PIX_OUT pixel_6901/CSA_VREF pixel
Xpixel_6912 pixel_6912/gring pixel_6912/VDD pixel_6912/GND pixel_6912/VREF pixel_6912/ROW_SEL
+ pixel_6912/NB1 pixel_6912/VBIAS pixel_6912/NB2 pixel_6912/AMP_IN pixel_6912/SF_IB
+ pixel_6912/PIX_OUT pixel_6912/CSA_VREF pixel
Xpixel_7668 pixel_7668/gring pixel_7668/VDD pixel_7668/GND pixel_7668/VREF pixel_7668/ROW_SEL
+ pixel_7668/NB1 pixel_7668/VBIAS pixel_7668/NB2 pixel_7668/AMP_IN pixel_7668/SF_IB
+ pixel_7668/PIX_OUT pixel_7668/CSA_VREF pixel
Xpixel_7679 pixel_7679/gring pixel_7679/VDD pixel_7679/GND pixel_7679/VREF pixel_7679/ROW_SEL
+ pixel_7679/NB1 pixel_7679/VBIAS pixel_7679/NB2 pixel_7679/AMP_IN pixel_7679/SF_IB
+ pixel_7679/PIX_OUT pixel_7679/CSA_VREF pixel
Xpixel_6923 pixel_6923/gring pixel_6923/VDD pixel_6923/GND pixel_6923/VREF pixel_6923/ROW_SEL
+ pixel_6923/NB1 pixel_6923/VBIAS pixel_6923/NB2 pixel_6923/AMP_IN pixel_6923/SF_IB
+ pixel_6923/PIX_OUT pixel_6923/CSA_VREF pixel
Xpixel_6934 pixel_6934/gring pixel_6934/VDD pixel_6934/GND pixel_6934/VREF pixel_6934/ROW_SEL
+ pixel_6934/NB1 pixel_6934/VBIAS pixel_6934/NB2 pixel_6934/AMP_IN pixel_6934/SF_IB
+ pixel_6934/PIX_OUT pixel_6934/CSA_VREF pixel
Xpixel_6945 pixel_6945/gring pixel_6945/VDD pixel_6945/GND pixel_6945/VREF pixel_6945/ROW_SEL
+ pixel_6945/NB1 pixel_6945/VBIAS pixel_6945/NB2 pixel_6945/AMP_IN pixel_6945/SF_IB
+ pixel_6945/PIX_OUT pixel_6945/CSA_VREF pixel
Xpixel_37 pixel_37/gring pixel_37/VDD pixel_37/GND pixel_37/VREF pixel_37/ROW_SEL
+ pixel_37/NB1 pixel_37/VBIAS pixel_37/NB2 pixel_37/AMP_IN pixel_37/SF_IB pixel_37/PIX_OUT
+ pixel_37/CSA_VREF pixel
Xpixel_26 pixel_26/gring pixel_26/VDD pixel_26/GND pixel_26/VREF pixel_26/ROW_SEL
+ pixel_26/NB1 pixel_26/VBIAS pixel_26/NB2 pixel_26/AMP_IN pixel_26/SF_IB pixel_26/PIX_OUT
+ pixel_26/CSA_VREF pixel
Xpixel_15 pixel_15/gring pixel_15/VDD pixel_15/GND pixel_15/VREF pixel_15/ROW_SEL
+ pixel_15/NB1 pixel_15/VBIAS pixel_15/NB2 pixel_15/AMP_IN pixel_15/SF_IB pixel_15/PIX_OUT
+ pixel_15/CSA_VREF pixel
Xpixel_6956 pixel_6956/gring pixel_6956/VDD pixel_6956/GND pixel_6956/VREF pixel_6956/ROW_SEL
+ pixel_6956/NB1 pixel_6956/VBIAS pixel_6956/NB2 pixel_6956/AMP_IN pixel_6956/SF_IB
+ pixel_6956/PIX_OUT pixel_6956/CSA_VREF pixel
Xpixel_6967 pixel_6967/gring pixel_6967/VDD pixel_6967/GND pixel_6967/VREF pixel_6967/ROW_SEL
+ pixel_6967/NB1 pixel_6967/VBIAS pixel_6967/NB2 pixel_6967/AMP_IN pixel_6967/SF_IB
+ pixel_6967/PIX_OUT pixel_6967/CSA_VREF pixel
Xpixel_6978 pixel_6978/gring pixel_6978/VDD pixel_6978/GND pixel_6978/VREF pixel_6978/ROW_SEL
+ pixel_6978/NB1 pixel_6978/VBIAS pixel_6978/NB2 pixel_6978/AMP_IN pixel_6978/SF_IB
+ pixel_6978/PIX_OUT pixel_6978/CSA_VREF pixel
Xpixel_6989 pixel_6989/gring pixel_6989/VDD pixel_6989/GND pixel_6989/VREF pixel_6989/ROW_SEL
+ pixel_6989/NB1 pixel_6989/VBIAS pixel_6989/NB2 pixel_6989/AMP_IN pixel_6989/SF_IB
+ pixel_6989/PIX_OUT pixel_6989/CSA_VREF pixel
Xpixel_59 pixel_59/gring pixel_59/VDD pixel_59/GND pixel_59/VREF pixel_59/ROW_SEL
+ pixel_59/NB1 pixel_59/VBIAS pixel_59/NB2 pixel_59/AMP_IN pixel_59/SF_IB pixel_59/PIX_OUT
+ pixel_59/CSA_VREF pixel
Xpixel_48 pixel_48/gring pixel_48/VDD pixel_48/GND pixel_48/VREF pixel_48/ROW_SEL
+ pixel_48/NB1 pixel_48/VBIAS pixel_48/NB2 pixel_48/AMP_IN pixel_48/SF_IB pixel_48/PIX_OUT
+ pixel_48/CSA_VREF pixel
Xpixel_1241 pixel_1241/gring pixel_1241/VDD pixel_1241/GND pixel_1241/VREF pixel_1241/ROW_SEL
+ pixel_1241/NB1 pixel_1241/VBIAS pixel_1241/NB2 pixel_1241/AMP_IN pixel_1241/SF_IB
+ pixel_1241/PIX_OUT pixel_1241/CSA_VREF pixel
Xpixel_1230 pixel_1230/gring pixel_1230/VDD pixel_1230/GND pixel_1230/VREF pixel_1230/ROW_SEL
+ pixel_1230/NB1 pixel_1230/VBIAS pixel_1230/NB2 pixel_1230/AMP_IN pixel_1230/SF_IB
+ pixel_1230/PIX_OUT pixel_1230/CSA_VREF pixel
Xpixel_1285 pixel_1285/gring pixel_1285/VDD pixel_1285/GND pixel_1285/VREF pixel_1285/ROW_SEL
+ pixel_1285/NB1 pixel_1285/VBIAS pixel_1285/NB2 pixel_1285/AMP_IN pixel_1285/SF_IB
+ pixel_1285/PIX_OUT pixel_1285/CSA_VREF pixel
Xpixel_1274 pixel_1274/gring pixel_1274/VDD pixel_1274/GND pixel_1274/VREF pixel_1274/ROW_SEL
+ pixel_1274/NB1 pixel_1274/VBIAS pixel_1274/NB2 pixel_1274/AMP_IN pixel_1274/SF_IB
+ pixel_1274/PIX_OUT pixel_1274/CSA_VREF pixel
Xpixel_1263 pixel_1263/gring pixel_1263/VDD pixel_1263/GND pixel_1263/VREF pixel_1263/ROW_SEL
+ pixel_1263/NB1 pixel_1263/VBIAS pixel_1263/NB2 pixel_1263/AMP_IN pixel_1263/SF_IB
+ pixel_1263/PIX_OUT pixel_1263/CSA_VREF pixel
Xpixel_1252 pixel_1252/gring pixel_1252/VDD pixel_1252/GND pixel_1252/VREF pixel_1252/ROW_SEL
+ pixel_1252/NB1 pixel_1252/VBIAS pixel_1252/NB2 pixel_1252/AMP_IN pixel_1252/SF_IB
+ pixel_1252/PIX_OUT pixel_1252/CSA_VREF pixel
Xpixel_1296 pixel_1296/gring pixel_1296/VDD pixel_1296/GND pixel_1296/VREF pixel_1296/ROW_SEL
+ pixel_1296/NB1 pixel_1296/VBIAS pixel_1296/NB2 pixel_1296/AMP_IN pixel_1296/SF_IB
+ pixel_1296/PIX_OUT pixel_1296/CSA_VREF pixel
Xpixel_9593 pixel_9593/gring pixel_9593/VDD pixel_9593/GND pixel_9593/VREF pixel_9593/ROW_SEL
+ pixel_9593/NB1 pixel_9593/VBIAS pixel_9593/NB2 pixel_9593/AMP_IN pixel_9593/SF_IB
+ pixel_9593/PIX_OUT pixel_9593/CSA_VREF pixel
Xpixel_9582 pixel_9582/gring pixel_9582/VDD pixel_9582/GND pixel_9582/VREF pixel_9582/ROW_SEL
+ pixel_9582/NB1 pixel_9582/VBIAS pixel_9582/NB2 pixel_9582/AMP_IN pixel_9582/SF_IB
+ pixel_9582/PIX_OUT pixel_9582/CSA_VREF pixel
Xpixel_9571 pixel_9571/gring pixel_9571/VDD pixel_9571/GND pixel_9571/VREF pixel_9571/ROW_SEL
+ pixel_9571/NB1 pixel_9571/VBIAS pixel_9571/NB2 pixel_9571/AMP_IN pixel_9571/SF_IB
+ pixel_9571/PIX_OUT pixel_9571/CSA_VREF pixel
Xpixel_9560 pixel_9560/gring pixel_9560/VDD pixel_9560/GND pixel_9560/VREF pixel_9560/ROW_SEL
+ pixel_9560/NB1 pixel_9560/VBIAS pixel_9560/NB2 pixel_9560/AMP_IN pixel_9560/SF_IB
+ pixel_9560/PIX_OUT pixel_9560/CSA_VREF pixel
Xpixel_8881 pixel_8881/gring pixel_8881/VDD pixel_8881/GND pixel_8881/VREF pixel_8881/ROW_SEL
+ pixel_8881/NB1 pixel_8881/VBIAS pixel_8881/NB2 pixel_8881/AMP_IN pixel_8881/SF_IB
+ pixel_8881/PIX_OUT pixel_8881/CSA_VREF pixel
Xpixel_8870 pixel_8870/gring pixel_8870/VDD pixel_8870/GND pixel_8870/VREF pixel_8870/ROW_SEL
+ pixel_8870/NB1 pixel_8870/VBIAS pixel_8870/NB2 pixel_8870/AMP_IN pixel_8870/SF_IB
+ pixel_8870/PIX_OUT pixel_8870/CSA_VREF pixel
Xpixel_8892 pixel_8892/gring pixel_8892/VDD pixel_8892/GND pixel_8892/VREF pixel_8892/ROW_SEL
+ pixel_8892/NB1 pixel_8892/VBIAS pixel_8892/NB2 pixel_8892/AMP_IN pixel_8892/SF_IB
+ pixel_8892/PIX_OUT pixel_8892/CSA_VREF pixel
Xpixel_6208 pixel_6208/gring pixel_6208/VDD pixel_6208/GND pixel_6208/VREF pixel_6208/ROW_SEL
+ pixel_6208/NB1 pixel_6208/VBIAS pixel_6208/NB2 pixel_6208/AMP_IN pixel_6208/SF_IB
+ pixel_6208/PIX_OUT pixel_6208/CSA_VREF pixel
Xpixel_6219 pixel_6219/gring pixel_6219/VDD pixel_6219/GND pixel_6219/VREF pixel_6219/ROW_SEL
+ pixel_6219/NB1 pixel_6219/VBIAS pixel_6219/NB2 pixel_6219/AMP_IN pixel_6219/SF_IB
+ pixel_6219/PIX_OUT pixel_6219/CSA_VREF pixel
Xpixel_5507 pixel_5507/gring pixel_5507/VDD pixel_5507/GND pixel_5507/VREF pixel_5507/ROW_SEL
+ pixel_5507/NB1 pixel_5507/VBIAS pixel_5507/NB2 pixel_5507/AMP_IN pixel_5507/SF_IB
+ pixel_5507/PIX_OUT pixel_5507/CSA_VREF pixel
Xpixel_5518 pixel_5518/gring pixel_5518/VDD pixel_5518/GND pixel_5518/VREF pixel_5518/ROW_SEL
+ pixel_5518/NB1 pixel_5518/VBIAS pixel_5518/NB2 pixel_5518/AMP_IN pixel_5518/SF_IB
+ pixel_5518/PIX_OUT pixel_5518/CSA_VREF pixel
Xpixel_5529 pixel_5529/gring pixel_5529/VDD pixel_5529/GND pixel_5529/VREF pixel_5529/ROW_SEL
+ pixel_5529/NB1 pixel_5529/VBIAS pixel_5529/NB2 pixel_5529/AMP_IN pixel_5529/SF_IB
+ pixel_5529/PIX_OUT pixel_5529/CSA_VREF pixel
Xpixel_823 pixel_823/gring pixel_823/VDD pixel_823/GND pixel_823/VREF pixel_823/ROW_SEL
+ pixel_823/NB1 pixel_823/VBIAS pixel_823/NB2 pixel_823/AMP_IN pixel_823/SF_IB pixel_823/PIX_OUT
+ pixel_823/CSA_VREF pixel
Xpixel_812 pixel_812/gring pixel_812/VDD pixel_812/GND pixel_812/VREF pixel_812/ROW_SEL
+ pixel_812/NB1 pixel_812/VBIAS pixel_812/NB2 pixel_812/AMP_IN pixel_812/SF_IB pixel_812/PIX_OUT
+ pixel_812/CSA_VREF pixel
Xpixel_801 pixel_801/gring pixel_801/VDD pixel_801/GND pixel_801/VREF pixel_801/ROW_SEL
+ pixel_801/NB1 pixel_801/VBIAS pixel_801/NB2 pixel_801/AMP_IN pixel_801/SF_IB pixel_801/PIX_OUT
+ pixel_801/CSA_VREF pixel
Xpixel_4806 pixel_4806/gring pixel_4806/VDD pixel_4806/GND pixel_4806/VREF pixel_4806/ROW_SEL
+ pixel_4806/NB1 pixel_4806/VBIAS pixel_4806/NB2 pixel_4806/AMP_IN pixel_4806/SF_IB
+ pixel_4806/PIX_OUT pixel_4806/CSA_VREF pixel
Xpixel_4817 pixel_4817/gring pixel_4817/VDD pixel_4817/GND pixel_4817/VREF pixel_4817/ROW_SEL
+ pixel_4817/NB1 pixel_4817/VBIAS pixel_4817/NB2 pixel_4817/AMP_IN pixel_4817/SF_IB
+ pixel_4817/PIX_OUT pixel_4817/CSA_VREF pixel
Xpixel_4828 pixel_4828/gring pixel_4828/VDD pixel_4828/GND pixel_4828/VREF pixel_4828/ROW_SEL
+ pixel_4828/NB1 pixel_4828/VBIAS pixel_4828/NB2 pixel_4828/AMP_IN pixel_4828/SF_IB
+ pixel_4828/PIX_OUT pixel_4828/CSA_VREF pixel
Xpixel_856 pixel_856/gring pixel_856/VDD pixel_856/GND pixel_856/VREF pixel_856/ROW_SEL
+ pixel_856/NB1 pixel_856/VBIAS pixel_856/NB2 pixel_856/AMP_IN pixel_856/SF_IB pixel_856/PIX_OUT
+ pixel_856/CSA_VREF pixel
Xpixel_845 pixel_845/gring pixel_845/VDD pixel_845/GND pixel_845/VREF pixel_845/ROW_SEL
+ pixel_845/NB1 pixel_845/VBIAS pixel_845/NB2 pixel_845/AMP_IN pixel_845/SF_IB pixel_845/PIX_OUT
+ pixel_845/CSA_VREF pixel
Xpixel_834 pixel_834/gring pixel_834/VDD pixel_834/GND pixel_834/VREF pixel_834/ROW_SEL
+ pixel_834/NB1 pixel_834/VBIAS pixel_834/NB2 pixel_834/AMP_IN pixel_834/SF_IB pixel_834/PIX_OUT
+ pixel_834/CSA_VREF pixel
Xpixel_4839 pixel_4839/gring pixel_4839/VDD pixel_4839/GND pixel_4839/VREF pixel_4839/ROW_SEL
+ pixel_4839/NB1 pixel_4839/VBIAS pixel_4839/NB2 pixel_4839/AMP_IN pixel_4839/SF_IB
+ pixel_4839/PIX_OUT pixel_4839/CSA_VREF pixel
Xpixel_889 pixel_889/gring pixel_889/VDD pixel_889/GND pixel_889/VREF pixel_889/ROW_SEL
+ pixel_889/NB1 pixel_889/VBIAS pixel_889/NB2 pixel_889/AMP_IN pixel_889/SF_IB pixel_889/PIX_OUT
+ pixel_889/CSA_VREF pixel
Xpixel_878 pixel_878/gring pixel_878/VDD pixel_878/GND pixel_878/VREF pixel_878/ROW_SEL
+ pixel_878/NB1 pixel_878/VBIAS pixel_878/NB2 pixel_878/AMP_IN pixel_878/SF_IB pixel_878/PIX_OUT
+ pixel_878/CSA_VREF pixel
Xpixel_867 pixel_867/gring pixel_867/VDD pixel_867/GND pixel_867/VREF pixel_867/ROW_SEL
+ pixel_867/NB1 pixel_867/VBIAS pixel_867/NB2 pixel_867/AMP_IN pixel_867/SF_IB pixel_867/PIX_OUT
+ pixel_867/CSA_VREF pixel
Xpixel_8100 pixel_8100/gring pixel_8100/VDD pixel_8100/GND pixel_8100/VREF pixel_8100/ROW_SEL
+ pixel_8100/NB1 pixel_8100/VBIAS pixel_8100/NB2 pixel_8100/AMP_IN pixel_8100/SF_IB
+ pixel_8100/PIX_OUT pixel_8100/CSA_VREF pixel
Xpixel_8111 pixel_8111/gring pixel_8111/VDD pixel_8111/GND pixel_8111/VREF pixel_8111/ROW_SEL
+ pixel_8111/NB1 pixel_8111/VBIAS pixel_8111/NB2 pixel_8111/AMP_IN pixel_8111/SF_IB
+ pixel_8111/PIX_OUT pixel_8111/CSA_VREF pixel
Xpixel_8122 pixel_8122/gring pixel_8122/VDD pixel_8122/GND pixel_8122/VREF pixel_8122/ROW_SEL
+ pixel_8122/NB1 pixel_8122/VBIAS pixel_8122/NB2 pixel_8122/AMP_IN pixel_8122/SF_IB
+ pixel_8122/PIX_OUT pixel_8122/CSA_VREF pixel
Xpixel_8133 pixel_8133/gring pixel_8133/VDD pixel_8133/GND pixel_8133/VREF pixel_8133/ROW_SEL
+ pixel_8133/NB1 pixel_8133/VBIAS pixel_8133/NB2 pixel_8133/AMP_IN pixel_8133/SF_IB
+ pixel_8133/PIX_OUT pixel_8133/CSA_VREF pixel
Xpixel_8144 pixel_8144/gring pixel_8144/VDD pixel_8144/GND pixel_8144/VREF pixel_8144/ROW_SEL
+ pixel_8144/NB1 pixel_8144/VBIAS pixel_8144/NB2 pixel_8144/AMP_IN pixel_8144/SF_IB
+ pixel_8144/PIX_OUT pixel_8144/CSA_VREF pixel
Xpixel_8155 pixel_8155/gring pixel_8155/VDD pixel_8155/GND pixel_8155/VREF pixel_8155/ROW_SEL
+ pixel_8155/NB1 pixel_8155/VBIAS pixel_8155/NB2 pixel_8155/AMP_IN pixel_8155/SF_IB
+ pixel_8155/PIX_OUT pixel_8155/CSA_VREF pixel
Xpixel_8166 pixel_8166/gring pixel_8166/VDD pixel_8166/GND pixel_8166/VREF pixel_8166/ROW_SEL
+ pixel_8166/NB1 pixel_8166/VBIAS pixel_8166/NB2 pixel_8166/AMP_IN pixel_8166/SF_IB
+ pixel_8166/PIX_OUT pixel_8166/CSA_VREF pixel
Xpixel_8177 pixel_8177/gring pixel_8177/VDD pixel_8177/GND pixel_8177/VREF pixel_8177/ROW_SEL
+ pixel_8177/NB1 pixel_8177/VBIAS pixel_8177/NB2 pixel_8177/AMP_IN pixel_8177/SF_IB
+ pixel_8177/PIX_OUT pixel_8177/CSA_VREF pixel
Xpixel_7410 pixel_7410/gring pixel_7410/VDD pixel_7410/GND pixel_7410/VREF pixel_7410/ROW_SEL
+ pixel_7410/NB1 pixel_7410/VBIAS pixel_7410/NB2 pixel_7410/AMP_IN pixel_7410/SF_IB
+ pixel_7410/PIX_OUT pixel_7410/CSA_VREF pixel
Xpixel_7421 pixel_7421/gring pixel_7421/VDD pixel_7421/GND pixel_7421/VREF pixel_7421/ROW_SEL
+ pixel_7421/NB1 pixel_7421/VBIAS pixel_7421/NB2 pixel_7421/AMP_IN pixel_7421/SF_IB
+ pixel_7421/PIX_OUT pixel_7421/CSA_VREF pixel
Xpixel_7432 pixel_7432/gring pixel_7432/VDD pixel_7432/GND pixel_7432/VREF pixel_7432/ROW_SEL
+ pixel_7432/NB1 pixel_7432/VBIAS pixel_7432/NB2 pixel_7432/AMP_IN pixel_7432/SF_IB
+ pixel_7432/PIX_OUT pixel_7432/CSA_VREF pixel
Xpixel_8188 pixel_8188/gring pixel_8188/VDD pixel_8188/GND pixel_8188/VREF pixel_8188/ROW_SEL
+ pixel_8188/NB1 pixel_8188/VBIAS pixel_8188/NB2 pixel_8188/AMP_IN pixel_8188/SF_IB
+ pixel_8188/PIX_OUT pixel_8188/CSA_VREF pixel
Xpixel_8199 pixel_8199/gring pixel_8199/VDD pixel_8199/GND pixel_8199/VREF pixel_8199/ROW_SEL
+ pixel_8199/NB1 pixel_8199/VBIAS pixel_8199/NB2 pixel_8199/AMP_IN pixel_8199/SF_IB
+ pixel_8199/PIX_OUT pixel_8199/CSA_VREF pixel
Xpixel_7443 pixel_7443/gring pixel_7443/VDD pixel_7443/GND pixel_7443/VREF pixel_7443/ROW_SEL
+ pixel_7443/NB1 pixel_7443/VBIAS pixel_7443/NB2 pixel_7443/AMP_IN pixel_7443/SF_IB
+ pixel_7443/PIX_OUT pixel_7443/CSA_VREF pixel
Xpixel_7454 pixel_7454/gring pixel_7454/VDD pixel_7454/GND pixel_7454/VREF pixel_7454/ROW_SEL
+ pixel_7454/NB1 pixel_7454/VBIAS pixel_7454/NB2 pixel_7454/AMP_IN pixel_7454/SF_IB
+ pixel_7454/PIX_OUT pixel_7454/CSA_VREF pixel
Xpixel_7465 pixel_7465/gring pixel_7465/VDD pixel_7465/GND pixel_7465/VREF pixel_7465/ROW_SEL
+ pixel_7465/NB1 pixel_7465/VBIAS pixel_7465/NB2 pixel_7465/AMP_IN pixel_7465/SF_IB
+ pixel_7465/PIX_OUT pixel_7465/CSA_VREF pixel
Xpixel_6720 pixel_6720/gring pixel_6720/VDD pixel_6720/GND pixel_6720/VREF pixel_6720/ROW_SEL
+ pixel_6720/NB1 pixel_6720/VBIAS pixel_6720/NB2 pixel_6720/AMP_IN pixel_6720/SF_IB
+ pixel_6720/PIX_OUT pixel_6720/CSA_VREF pixel
Xpixel_7476 pixel_7476/gring pixel_7476/VDD pixel_7476/GND pixel_7476/VREF pixel_7476/ROW_SEL
+ pixel_7476/NB1 pixel_7476/VBIAS pixel_7476/NB2 pixel_7476/AMP_IN pixel_7476/SF_IB
+ pixel_7476/PIX_OUT pixel_7476/CSA_VREF pixel
Xpixel_7487 pixel_7487/gring pixel_7487/VDD pixel_7487/GND pixel_7487/VREF pixel_7487/ROW_SEL
+ pixel_7487/NB1 pixel_7487/VBIAS pixel_7487/NB2 pixel_7487/AMP_IN pixel_7487/SF_IB
+ pixel_7487/PIX_OUT pixel_7487/CSA_VREF pixel
Xpixel_7498 pixel_7498/gring pixel_7498/VDD pixel_7498/GND pixel_7498/VREF pixel_7498/ROW_SEL
+ pixel_7498/NB1 pixel_7498/VBIAS pixel_7498/NB2 pixel_7498/AMP_IN pixel_7498/SF_IB
+ pixel_7498/PIX_OUT pixel_7498/CSA_VREF pixel
Xpixel_6731 pixel_6731/gring pixel_6731/VDD pixel_6731/GND pixel_6731/VREF pixel_6731/ROW_SEL
+ pixel_6731/NB1 pixel_6731/VBIAS pixel_6731/NB2 pixel_6731/AMP_IN pixel_6731/SF_IB
+ pixel_6731/PIX_OUT pixel_6731/CSA_VREF pixel
Xpixel_6742 pixel_6742/gring pixel_6742/VDD pixel_6742/GND pixel_6742/VREF pixel_6742/ROW_SEL
+ pixel_6742/NB1 pixel_6742/VBIAS pixel_6742/NB2 pixel_6742/AMP_IN pixel_6742/SF_IB
+ pixel_6742/PIX_OUT pixel_6742/CSA_VREF pixel
Xpixel_6753 pixel_6753/gring pixel_6753/VDD pixel_6753/GND pixel_6753/VREF pixel_6753/ROW_SEL
+ pixel_6753/NB1 pixel_6753/VBIAS pixel_6753/NB2 pixel_6753/AMP_IN pixel_6753/SF_IB
+ pixel_6753/PIX_OUT pixel_6753/CSA_VREF pixel
Xpixel_6764 pixel_6764/gring pixel_6764/VDD pixel_6764/GND pixel_6764/VREF pixel_6764/ROW_SEL
+ pixel_6764/NB1 pixel_6764/VBIAS pixel_6764/NB2 pixel_6764/AMP_IN pixel_6764/SF_IB
+ pixel_6764/PIX_OUT pixel_6764/CSA_VREF pixel
Xpixel_6775 pixel_6775/gring pixel_6775/VDD pixel_6775/GND pixel_6775/VREF pixel_6775/ROW_SEL
+ pixel_6775/NB1 pixel_6775/VBIAS pixel_6775/NB2 pixel_6775/AMP_IN pixel_6775/SF_IB
+ pixel_6775/PIX_OUT pixel_6775/CSA_VREF pixel
Xpixel_6786 pixel_6786/gring pixel_6786/VDD pixel_6786/GND pixel_6786/VREF pixel_6786/ROW_SEL
+ pixel_6786/NB1 pixel_6786/VBIAS pixel_6786/NB2 pixel_6786/AMP_IN pixel_6786/SF_IB
+ pixel_6786/PIX_OUT pixel_6786/CSA_VREF pixel
Xpixel_6797 pixel_6797/gring pixel_6797/VDD pixel_6797/GND pixel_6797/VREF pixel_6797/ROW_SEL
+ pixel_6797/NB1 pixel_6797/VBIAS pixel_6797/NB2 pixel_6797/AMP_IN pixel_6797/SF_IB
+ pixel_6797/PIX_OUT pixel_6797/CSA_VREF pixel
Xpixel_1060 pixel_1060/gring pixel_1060/VDD pixel_1060/GND pixel_1060/VREF pixel_1060/ROW_SEL
+ pixel_1060/NB1 pixel_1060/VBIAS pixel_1060/NB2 pixel_1060/AMP_IN pixel_1060/SF_IB
+ pixel_1060/PIX_OUT pixel_1060/CSA_VREF pixel
Xpixel_1093 pixel_1093/gring pixel_1093/VDD pixel_1093/GND pixel_1093/VREF pixel_1093/ROW_SEL
+ pixel_1093/NB1 pixel_1093/VBIAS pixel_1093/NB2 pixel_1093/AMP_IN pixel_1093/SF_IB
+ pixel_1093/PIX_OUT pixel_1093/CSA_VREF pixel
Xpixel_1082 pixel_1082/gring pixel_1082/VDD pixel_1082/GND pixel_1082/VREF pixel_1082/ROW_SEL
+ pixel_1082/NB1 pixel_1082/VBIAS pixel_1082/NB2 pixel_1082/AMP_IN pixel_1082/SF_IB
+ pixel_1082/PIX_OUT pixel_1082/CSA_VREF pixel
Xpixel_1071 pixel_1071/gring pixel_1071/VDD pixel_1071/GND pixel_1071/VREF pixel_1071/ROW_SEL
+ pixel_1071/NB1 pixel_1071/VBIAS pixel_1071/NB2 pixel_1071/AMP_IN pixel_1071/SF_IB
+ pixel_1071/PIX_OUT pixel_1071/CSA_VREF pixel
Xpixel_9390 pixel_9390/gring pixel_9390/VDD pixel_9390/GND pixel_9390/VREF pixel_9390/ROW_SEL
+ pixel_9390/NB1 pixel_9390/VBIAS pixel_9390/NB2 pixel_9390/AMP_IN pixel_9390/SF_IB
+ pixel_9390/PIX_OUT pixel_9390/CSA_VREF pixel
Xpixel_119 pixel_119/gring pixel_119/VDD pixel_119/GND pixel_119/VREF pixel_119/ROW_SEL
+ pixel_119/NB1 pixel_119/VBIAS pixel_119/NB2 pixel_119/AMP_IN pixel_119/SF_IB pixel_119/PIX_OUT
+ pixel_119/CSA_VREF pixel
Xpixel_108 pixel_108/gring pixel_108/VDD pixel_108/GND pixel_108/VREF pixel_108/ROW_SEL
+ pixel_108/NB1 pixel_108/VBIAS pixel_108/NB2 pixel_108/AMP_IN pixel_108/SF_IB pixel_108/PIX_OUT
+ pixel_108/CSA_VREF pixel
Xpixel_6005 pixel_6005/gring pixel_6005/VDD pixel_6005/GND pixel_6005/VREF pixel_6005/ROW_SEL
+ pixel_6005/NB1 pixel_6005/VBIAS pixel_6005/NB2 pixel_6005/AMP_IN pixel_6005/SF_IB
+ pixel_6005/PIX_OUT pixel_6005/CSA_VREF pixel
Xpixel_6016 pixel_6016/gring pixel_6016/VDD pixel_6016/GND pixel_6016/VREF pixel_6016/ROW_SEL
+ pixel_6016/NB1 pixel_6016/VBIAS pixel_6016/NB2 pixel_6016/AMP_IN pixel_6016/SF_IB
+ pixel_6016/PIX_OUT pixel_6016/CSA_VREF pixel
Xpixel_6027 pixel_6027/gring pixel_6027/VDD pixel_6027/GND pixel_6027/VREF pixel_6027/ROW_SEL
+ pixel_6027/NB1 pixel_6027/VBIAS pixel_6027/NB2 pixel_6027/AMP_IN pixel_6027/SF_IB
+ pixel_6027/PIX_OUT pixel_6027/CSA_VREF pixel
Xpixel_6038 pixel_6038/gring pixel_6038/VDD pixel_6038/GND pixel_6038/VREF pixel_6038/ROW_SEL
+ pixel_6038/NB1 pixel_6038/VBIAS pixel_6038/NB2 pixel_6038/AMP_IN pixel_6038/SF_IB
+ pixel_6038/PIX_OUT pixel_6038/CSA_VREF pixel
Xpixel_6049 pixel_6049/gring pixel_6049/VDD pixel_6049/GND pixel_6049/VREF pixel_6049/ROW_SEL
+ pixel_6049/NB1 pixel_6049/VBIAS pixel_6049/NB2 pixel_6049/AMP_IN pixel_6049/SF_IB
+ pixel_6049/PIX_OUT pixel_6049/CSA_VREF pixel
Xpixel_5304 pixel_5304/gring pixel_5304/VDD pixel_5304/GND pixel_5304/VREF pixel_5304/ROW_SEL
+ pixel_5304/NB1 pixel_5304/VBIAS pixel_5304/NB2 pixel_5304/AMP_IN pixel_5304/SF_IB
+ pixel_5304/PIX_OUT pixel_5304/CSA_VREF pixel
Xpixel_5315 pixel_5315/gring pixel_5315/VDD pixel_5315/GND pixel_5315/VREF pixel_5315/ROW_SEL
+ pixel_5315/NB1 pixel_5315/VBIAS pixel_5315/NB2 pixel_5315/AMP_IN pixel_5315/SF_IB
+ pixel_5315/PIX_OUT pixel_5315/CSA_VREF pixel
Xpixel_5326 pixel_5326/gring pixel_5326/VDD pixel_5326/GND pixel_5326/VREF pixel_5326/ROW_SEL
+ pixel_5326/NB1 pixel_5326/VBIAS pixel_5326/NB2 pixel_5326/AMP_IN pixel_5326/SF_IB
+ pixel_5326/PIX_OUT pixel_5326/CSA_VREF pixel
Xpixel_5337 pixel_5337/gring pixel_5337/VDD pixel_5337/GND pixel_5337/VREF pixel_5337/ROW_SEL
+ pixel_5337/NB1 pixel_5337/VBIAS pixel_5337/NB2 pixel_5337/AMP_IN pixel_5337/SF_IB
+ pixel_5337/PIX_OUT pixel_5337/CSA_VREF pixel
Xpixel_5348 pixel_5348/gring pixel_5348/VDD pixel_5348/GND pixel_5348/VREF pixel_5348/ROW_SEL
+ pixel_5348/NB1 pixel_5348/VBIAS pixel_5348/NB2 pixel_5348/AMP_IN pixel_5348/SF_IB
+ pixel_5348/PIX_OUT pixel_5348/CSA_VREF pixel
Xpixel_4603 pixel_4603/gring pixel_4603/VDD pixel_4603/GND pixel_4603/VREF pixel_4603/ROW_SEL
+ pixel_4603/NB1 pixel_4603/VBIAS pixel_4603/NB2 pixel_4603/AMP_IN pixel_4603/SF_IB
+ pixel_4603/PIX_OUT pixel_4603/CSA_VREF pixel
Xpixel_631 pixel_631/gring pixel_631/VDD pixel_631/GND pixel_631/VREF pixel_631/ROW_SEL
+ pixel_631/NB1 pixel_631/VBIAS pixel_631/NB2 pixel_631/AMP_IN pixel_631/SF_IB pixel_631/PIX_OUT
+ pixel_631/CSA_VREF pixel
Xpixel_620 pixel_620/gring pixel_620/VDD pixel_620/GND pixel_620/VREF pixel_620/ROW_SEL
+ pixel_620/NB1 pixel_620/VBIAS pixel_620/NB2 pixel_620/AMP_IN pixel_620/SF_IB pixel_620/PIX_OUT
+ pixel_620/CSA_VREF pixel
Xpixel_5359 pixel_5359/gring pixel_5359/VDD pixel_5359/GND pixel_5359/VREF pixel_5359/ROW_SEL
+ pixel_5359/NB1 pixel_5359/VBIAS pixel_5359/NB2 pixel_5359/AMP_IN pixel_5359/SF_IB
+ pixel_5359/PIX_OUT pixel_5359/CSA_VREF pixel
Xpixel_4614 pixel_4614/gring pixel_4614/VDD pixel_4614/GND pixel_4614/VREF pixel_4614/ROW_SEL
+ pixel_4614/NB1 pixel_4614/VBIAS pixel_4614/NB2 pixel_4614/AMP_IN pixel_4614/SF_IB
+ pixel_4614/PIX_OUT pixel_4614/CSA_VREF pixel
Xpixel_4625 pixel_4625/gring pixel_4625/VDD pixel_4625/GND pixel_4625/VREF pixel_4625/ROW_SEL
+ pixel_4625/NB1 pixel_4625/VBIAS pixel_4625/NB2 pixel_4625/AMP_IN pixel_4625/SF_IB
+ pixel_4625/PIX_OUT pixel_4625/CSA_VREF pixel
Xpixel_4636 pixel_4636/gring pixel_4636/VDD pixel_4636/GND pixel_4636/VREF pixel_4636/ROW_SEL
+ pixel_4636/NB1 pixel_4636/VBIAS pixel_4636/NB2 pixel_4636/AMP_IN pixel_4636/SF_IB
+ pixel_4636/PIX_OUT pixel_4636/CSA_VREF pixel
Xpixel_675 pixel_675/gring pixel_675/VDD pixel_675/GND pixel_675/VREF pixel_675/ROW_SEL
+ pixel_675/NB1 pixel_675/VBIAS pixel_675/NB2 pixel_675/AMP_IN pixel_675/SF_IB pixel_675/PIX_OUT
+ pixel_675/CSA_VREF pixel
Xpixel_664 pixel_664/gring pixel_664/VDD pixel_664/GND pixel_664/VREF pixel_664/ROW_SEL
+ pixel_664/NB1 pixel_664/VBIAS pixel_664/NB2 pixel_664/AMP_IN pixel_664/SF_IB pixel_664/PIX_OUT
+ pixel_664/CSA_VREF pixel
Xpixel_653 pixel_653/gring pixel_653/VDD pixel_653/GND pixel_653/VREF pixel_653/ROW_SEL
+ pixel_653/NB1 pixel_653/VBIAS pixel_653/NB2 pixel_653/AMP_IN pixel_653/SF_IB pixel_653/PIX_OUT
+ pixel_653/CSA_VREF pixel
Xpixel_642 pixel_642/gring pixel_642/VDD pixel_642/GND pixel_642/VREF pixel_642/ROW_SEL
+ pixel_642/NB1 pixel_642/VBIAS pixel_642/NB2 pixel_642/AMP_IN pixel_642/SF_IB pixel_642/PIX_OUT
+ pixel_642/CSA_VREF pixel
Xpixel_4647 pixel_4647/gring pixel_4647/VDD pixel_4647/GND pixel_4647/VREF pixel_4647/ROW_SEL
+ pixel_4647/NB1 pixel_4647/VBIAS pixel_4647/NB2 pixel_4647/AMP_IN pixel_4647/SF_IB
+ pixel_4647/PIX_OUT pixel_4647/CSA_VREF pixel
Xpixel_4658 pixel_4658/gring pixel_4658/VDD pixel_4658/GND pixel_4658/VREF pixel_4658/ROW_SEL
+ pixel_4658/NB1 pixel_4658/VBIAS pixel_4658/NB2 pixel_4658/AMP_IN pixel_4658/SF_IB
+ pixel_4658/PIX_OUT pixel_4658/CSA_VREF pixel
Xpixel_4669 pixel_4669/gring pixel_4669/VDD pixel_4669/GND pixel_4669/VREF pixel_4669/ROW_SEL
+ pixel_4669/NB1 pixel_4669/VBIAS pixel_4669/NB2 pixel_4669/AMP_IN pixel_4669/SF_IB
+ pixel_4669/PIX_OUT pixel_4669/CSA_VREF pixel
Xpixel_3902 pixel_3902/gring pixel_3902/VDD pixel_3902/GND pixel_3902/VREF pixel_3902/ROW_SEL
+ pixel_3902/NB1 pixel_3902/VBIAS pixel_3902/NB2 pixel_3902/AMP_IN pixel_3902/SF_IB
+ pixel_3902/PIX_OUT pixel_3902/CSA_VREF pixel
Xpixel_3913 pixel_3913/gring pixel_3913/VDD pixel_3913/GND pixel_3913/VREF pixel_3913/ROW_SEL
+ pixel_3913/NB1 pixel_3913/VBIAS pixel_3913/NB2 pixel_3913/AMP_IN pixel_3913/SF_IB
+ pixel_3913/PIX_OUT pixel_3913/CSA_VREF pixel
Xpixel_3924 pixel_3924/gring pixel_3924/VDD pixel_3924/GND pixel_3924/VREF pixel_3924/ROW_SEL
+ pixel_3924/NB1 pixel_3924/VBIAS pixel_3924/NB2 pixel_3924/AMP_IN pixel_3924/SF_IB
+ pixel_3924/PIX_OUT pixel_3924/CSA_VREF pixel
Xpixel_3935 pixel_3935/gring pixel_3935/VDD pixel_3935/GND pixel_3935/VREF pixel_3935/ROW_SEL
+ pixel_3935/NB1 pixel_3935/VBIAS pixel_3935/NB2 pixel_3935/AMP_IN pixel_3935/SF_IB
+ pixel_3935/PIX_OUT pixel_3935/CSA_VREF pixel
Xpixel_697 pixel_697/gring pixel_697/VDD pixel_697/GND pixel_697/VREF pixel_697/ROW_SEL
+ pixel_697/NB1 pixel_697/VBIAS pixel_697/NB2 pixel_697/AMP_IN pixel_697/SF_IB pixel_697/PIX_OUT
+ pixel_697/CSA_VREF pixel
Xpixel_686 pixel_686/gring pixel_686/VDD pixel_686/GND pixel_686/VREF pixel_686/ROW_SEL
+ pixel_686/NB1 pixel_686/VBIAS pixel_686/NB2 pixel_686/AMP_IN pixel_686/SF_IB pixel_686/PIX_OUT
+ pixel_686/CSA_VREF pixel
Xpixel_3946 pixel_3946/gring pixel_3946/VDD pixel_3946/GND pixel_3946/VREF pixel_3946/ROW_SEL
+ pixel_3946/NB1 pixel_3946/VBIAS pixel_3946/NB2 pixel_3946/AMP_IN pixel_3946/SF_IB
+ pixel_3946/PIX_OUT pixel_3946/CSA_VREF pixel
Xpixel_3957 pixel_3957/gring pixel_3957/VDD pixel_3957/GND pixel_3957/VREF pixel_3957/ROW_SEL
+ pixel_3957/NB1 pixel_3957/VBIAS pixel_3957/NB2 pixel_3957/AMP_IN pixel_3957/SF_IB
+ pixel_3957/PIX_OUT pixel_3957/CSA_VREF pixel
Xpixel_3968 pixel_3968/gring pixel_3968/VDD pixel_3968/GND pixel_3968/VREF pixel_3968/ROW_SEL
+ pixel_3968/NB1 pixel_3968/VBIAS pixel_3968/NB2 pixel_3968/AMP_IN pixel_3968/SF_IB
+ pixel_3968/PIX_OUT pixel_3968/CSA_VREF pixel
Xpixel_3979 pixel_3979/gring pixel_3979/VDD pixel_3979/GND pixel_3979/VREF pixel_3979/ROW_SEL
+ pixel_3979/NB1 pixel_3979/VBIAS pixel_3979/NB2 pixel_3979/AMP_IN pixel_3979/SF_IB
+ pixel_3979/PIX_OUT pixel_3979/CSA_VREF pixel
Xpixel_7240 pixel_7240/gring pixel_7240/VDD pixel_7240/GND pixel_7240/VREF pixel_7240/ROW_SEL
+ pixel_7240/NB1 pixel_7240/VBIAS pixel_7240/NB2 pixel_7240/AMP_IN pixel_7240/SF_IB
+ pixel_7240/PIX_OUT pixel_7240/CSA_VREF pixel
Xpixel_7251 pixel_7251/gring pixel_7251/VDD pixel_7251/GND pixel_7251/VREF pixel_7251/ROW_SEL
+ pixel_7251/NB1 pixel_7251/VBIAS pixel_7251/NB2 pixel_7251/AMP_IN pixel_7251/SF_IB
+ pixel_7251/PIX_OUT pixel_7251/CSA_VREF pixel
Xpixel_7262 pixel_7262/gring pixel_7262/VDD pixel_7262/GND pixel_7262/VREF pixel_7262/ROW_SEL
+ pixel_7262/NB1 pixel_7262/VBIAS pixel_7262/NB2 pixel_7262/AMP_IN pixel_7262/SF_IB
+ pixel_7262/PIX_OUT pixel_7262/CSA_VREF pixel
Xpixel_7273 pixel_7273/gring pixel_7273/VDD pixel_7273/GND pixel_7273/VREF pixel_7273/ROW_SEL
+ pixel_7273/NB1 pixel_7273/VBIAS pixel_7273/NB2 pixel_7273/AMP_IN pixel_7273/SF_IB
+ pixel_7273/PIX_OUT pixel_7273/CSA_VREF pixel
Xpixel_7284 pixel_7284/gring pixel_7284/VDD pixel_7284/GND pixel_7284/VREF pixel_7284/ROW_SEL
+ pixel_7284/NB1 pixel_7284/VBIAS pixel_7284/NB2 pixel_7284/AMP_IN pixel_7284/SF_IB
+ pixel_7284/PIX_OUT pixel_7284/CSA_VREF pixel
Xpixel_7295 pixel_7295/gring pixel_7295/VDD pixel_7295/GND pixel_7295/VREF pixel_7295/ROW_SEL
+ pixel_7295/NB1 pixel_7295/VBIAS pixel_7295/NB2 pixel_7295/AMP_IN pixel_7295/SF_IB
+ pixel_7295/PIX_OUT pixel_7295/CSA_VREF pixel
Xpixel_6550 pixel_6550/gring pixel_6550/VDD pixel_6550/GND pixel_6550/VREF pixel_6550/ROW_SEL
+ pixel_6550/NB1 pixel_6550/VBIAS pixel_6550/NB2 pixel_6550/AMP_IN pixel_6550/SF_IB
+ pixel_6550/PIX_OUT pixel_6550/CSA_VREF pixel
Xpixel_6561 pixel_6561/gring pixel_6561/VDD pixel_6561/GND pixel_6561/VREF pixel_6561/ROW_SEL
+ pixel_6561/NB1 pixel_6561/VBIAS pixel_6561/NB2 pixel_6561/AMP_IN pixel_6561/SF_IB
+ pixel_6561/PIX_OUT pixel_6561/CSA_VREF pixel
Xpixel_6572 pixel_6572/gring pixel_6572/VDD pixel_6572/GND pixel_6572/VREF pixel_6572/ROW_SEL
+ pixel_6572/NB1 pixel_6572/VBIAS pixel_6572/NB2 pixel_6572/AMP_IN pixel_6572/SF_IB
+ pixel_6572/PIX_OUT pixel_6572/CSA_VREF pixel
Xpixel_6583 pixel_6583/gring pixel_6583/VDD pixel_6583/GND pixel_6583/VREF pixel_6583/ROW_SEL
+ pixel_6583/NB1 pixel_6583/VBIAS pixel_6583/NB2 pixel_6583/AMP_IN pixel_6583/SF_IB
+ pixel_6583/PIX_OUT pixel_6583/CSA_VREF pixel
Xpixel_6594 pixel_6594/gring pixel_6594/VDD pixel_6594/GND pixel_6594/VREF pixel_6594/ROW_SEL
+ pixel_6594/NB1 pixel_6594/VBIAS pixel_6594/NB2 pixel_6594/AMP_IN pixel_6594/SF_IB
+ pixel_6594/PIX_OUT pixel_6594/CSA_VREF pixel
Xpixel_5860 pixel_5860/gring pixel_5860/VDD pixel_5860/GND pixel_5860/VREF pixel_5860/ROW_SEL
+ pixel_5860/NB1 pixel_5860/VBIAS pixel_5860/NB2 pixel_5860/AMP_IN pixel_5860/SF_IB
+ pixel_5860/PIX_OUT pixel_5860/CSA_VREF pixel
Xpixel_5871 pixel_5871/gring pixel_5871/VDD pixel_5871/GND pixel_5871/VREF pixel_5871/ROW_SEL
+ pixel_5871/NB1 pixel_5871/VBIAS pixel_5871/NB2 pixel_5871/AMP_IN pixel_5871/SF_IB
+ pixel_5871/PIX_OUT pixel_5871/CSA_VREF pixel
Xpixel_5882 pixel_5882/gring pixel_5882/VDD pixel_5882/GND pixel_5882/VREF pixel_5882/ROW_SEL
+ pixel_5882/NB1 pixel_5882/VBIAS pixel_5882/NB2 pixel_5882/AMP_IN pixel_5882/SF_IB
+ pixel_5882/PIX_OUT pixel_5882/CSA_VREF pixel
Xpixel_5893 pixel_5893/gring pixel_5893/VDD pixel_5893/GND pixel_5893/VREF pixel_5893/ROW_SEL
+ pixel_5893/NB1 pixel_5893/VBIAS pixel_5893/NB2 pixel_5893/AMP_IN pixel_5893/SF_IB
+ pixel_5893/PIX_OUT pixel_5893/CSA_VREF pixel
Xpixel_3209 pixel_3209/gring pixel_3209/VDD pixel_3209/GND pixel_3209/VREF pixel_3209/ROW_SEL
+ pixel_3209/NB1 pixel_3209/VBIAS pixel_3209/NB2 pixel_3209/AMP_IN pixel_3209/SF_IB
+ pixel_3209/PIX_OUT pixel_3209/CSA_VREF pixel
Xpixel_2519 pixel_2519/gring pixel_2519/VDD pixel_2519/GND pixel_2519/VREF pixel_2519/ROW_SEL
+ pixel_2519/NB1 pixel_2519/VBIAS pixel_2519/NB2 pixel_2519/AMP_IN pixel_2519/SF_IB
+ pixel_2519/PIX_OUT pixel_2519/CSA_VREF pixel
Xpixel_2508 pixel_2508/gring pixel_2508/VDD pixel_2508/GND pixel_2508/VREF pixel_2508/ROW_SEL
+ pixel_2508/NB1 pixel_2508/VBIAS pixel_2508/NB2 pixel_2508/AMP_IN pixel_2508/SF_IB
+ pixel_2508/PIX_OUT pixel_2508/CSA_VREF pixel
Xpixel_1807 pixel_1807/gring pixel_1807/VDD pixel_1807/GND pixel_1807/VREF pixel_1807/ROW_SEL
+ pixel_1807/NB1 pixel_1807/VBIAS pixel_1807/NB2 pixel_1807/AMP_IN pixel_1807/SF_IB
+ pixel_1807/PIX_OUT pixel_1807/CSA_VREF pixel
Xpixel_1829 pixel_1829/gring pixel_1829/VDD pixel_1829/GND pixel_1829/VREF pixel_1829/ROW_SEL
+ pixel_1829/NB1 pixel_1829/VBIAS pixel_1829/NB2 pixel_1829/AMP_IN pixel_1829/SF_IB
+ pixel_1829/PIX_OUT pixel_1829/CSA_VREF pixel
Xpixel_1818 pixel_1818/gring pixel_1818/VDD pixel_1818/GND pixel_1818/VREF pixel_1818/ROW_SEL
+ pixel_1818/NB1 pixel_1818/VBIAS pixel_1818/NB2 pixel_1818/AMP_IN pixel_1818/SF_IB
+ pixel_1818/PIX_OUT pixel_1818/CSA_VREF pixel
Xpixel_5101 pixel_5101/gring pixel_5101/VDD pixel_5101/GND pixel_5101/VREF pixel_5101/ROW_SEL
+ pixel_5101/NB1 pixel_5101/VBIAS pixel_5101/NB2 pixel_5101/AMP_IN pixel_5101/SF_IB
+ pixel_5101/PIX_OUT pixel_5101/CSA_VREF pixel
Xpixel_5112 pixel_5112/gring pixel_5112/VDD pixel_5112/GND pixel_5112/VREF pixel_5112/ROW_SEL
+ pixel_5112/NB1 pixel_5112/VBIAS pixel_5112/NB2 pixel_5112/AMP_IN pixel_5112/SF_IB
+ pixel_5112/PIX_OUT pixel_5112/CSA_VREF pixel
Xpixel_5123 pixel_5123/gring pixel_5123/VDD pixel_5123/GND pixel_5123/VREF pixel_5123/ROW_SEL
+ pixel_5123/NB1 pixel_5123/VBIAS pixel_5123/NB2 pixel_5123/AMP_IN pixel_5123/SF_IB
+ pixel_5123/PIX_OUT pixel_5123/CSA_VREF pixel
Xpixel_5134 pixel_5134/gring pixel_5134/VDD pixel_5134/GND pixel_5134/VREF pixel_5134/ROW_SEL
+ pixel_5134/NB1 pixel_5134/VBIAS pixel_5134/NB2 pixel_5134/AMP_IN pixel_5134/SF_IB
+ pixel_5134/PIX_OUT pixel_5134/CSA_VREF pixel
Xpixel_5145 pixel_5145/gring pixel_5145/VDD pixel_5145/GND pixel_5145/VREF pixel_5145/ROW_SEL
+ pixel_5145/NB1 pixel_5145/VBIAS pixel_5145/NB2 pixel_5145/AMP_IN pixel_5145/SF_IB
+ pixel_5145/PIX_OUT pixel_5145/CSA_VREF pixel
Xpixel_5156 pixel_5156/gring pixel_5156/VDD pixel_5156/GND pixel_5156/VREF pixel_5156/ROW_SEL
+ pixel_5156/NB1 pixel_5156/VBIAS pixel_5156/NB2 pixel_5156/AMP_IN pixel_5156/SF_IB
+ pixel_5156/PIX_OUT pixel_5156/CSA_VREF pixel
Xpixel_4400 pixel_4400/gring pixel_4400/VDD pixel_4400/GND pixel_4400/VREF pixel_4400/ROW_SEL
+ pixel_4400/NB1 pixel_4400/VBIAS pixel_4400/NB2 pixel_4400/AMP_IN pixel_4400/SF_IB
+ pixel_4400/PIX_OUT pixel_4400/CSA_VREF pixel
Xpixel_4411 pixel_4411/gring pixel_4411/VDD pixel_4411/GND pixel_4411/VREF pixel_4411/ROW_SEL
+ pixel_4411/NB1 pixel_4411/VBIAS pixel_4411/NB2 pixel_4411/AMP_IN pixel_4411/SF_IB
+ pixel_4411/PIX_OUT pixel_4411/CSA_VREF pixel
Xpixel_450 pixel_450/gring pixel_450/VDD pixel_450/GND pixel_450/VREF pixel_450/ROW_SEL
+ pixel_450/NB1 pixel_450/VBIAS pixel_450/NB2 pixel_450/AMP_IN pixel_450/SF_IB pixel_450/PIX_OUT
+ pixel_450/CSA_VREF pixel
Xpixel_3710 pixel_3710/gring pixel_3710/VDD pixel_3710/GND pixel_3710/VREF pixel_3710/ROW_SEL
+ pixel_3710/NB1 pixel_3710/VBIAS pixel_3710/NB2 pixel_3710/AMP_IN pixel_3710/SF_IB
+ pixel_3710/PIX_OUT pixel_3710/CSA_VREF pixel
Xpixel_5167 pixel_5167/gring pixel_5167/VDD pixel_5167/GND pixel_5167/VREF pixel_5167/ROW_SEL
+ pixel_5167/NB1 pixel_5167/VBIAS pixel_5167/NB2 pixel_5167/AMP_IN pixel_5167/SF_IB
+ pixel_5167/PIX_OUT pixel_5167/CSA_VREF pixel
Xpixel_5178 pixel_5178/gring pixel_5178/VDD pixel_5178/GND pixel_5178/VREF pixel_5178/ROW_SEL
+ pixel_5178/NB1 pixel_5178/VBIAS pixel_5178/NB2 pixel_5178/AMP_IN pixel_5178/SF_IB
+ pixel_5178/PIX_OUT pixel_5178/CSA_VREF pixel
Xpixel_5189 pixel_5189/gring pixel_5189/VDD pixel_5189/GND pixel_5189/VREF pixel_5189/ROW_SEL
+ pixel_5189/NB1 pixel_5189/VBIAS pixel_5189/NB2 pixel_5189/AMP_IN pixel_5189/SF_IB
+ pixel_5189/PIX_OUT pixel_5189/CSA_VREF pixel
Xpixel_4422 pixel_4422/gring pixel_4422/VDD pixel_4422/GND pixel_4422/VREF pixel_4422/ROW_SEL
+ pixel_4422/NB1 pixel_4422/VBIAS pixel_4422/NB2 pixel_4422/AMP_IN pixel_4422/SF_IB
+ pixel_4422/PIX_OUT pixel_4422/CSA_VREF pixel
Xpixel_4433 pixel_4433/gring pixel_4433/VDD pixel_4433/GND pixel_4433/VREF pixel_4433/ROW_SEL
+ pixel_4433/NB1 pixel_4433/VBIAS pixel_4433/NB2 pixel_4433/AMP_IN pixel_4433/SF_IB
+ pixel_4433/PIX_OUT pixel_4433/CSA_VREF pixel
Xpixel_4444 pixel_4444/gring pixel_4444/VDD pixel_4444/GND pixel_4444/VREF pixel_4444/ROW_SEL
+ pixel_4444/NB1 pixel_4444/VBIAS pixel_4444/NB2 pixel_4444/AMP_IN pixel_4444/SF_IB
+ pixel_4444/PIX_OUT pixel_4444/CSA_VREF pixel
Xpixel_483 pixel_483/gring pixel_483/VDD pixel_483/GND pixel_483/VREF pixel_483/ROW_SEL
+ pixel_483/NB1 pixel_483/VBIAS pixel_483/NB2 pixel_483/AMP_IN pixel_483/SF_IB pixel_483/PIX_OUT
+ pixel_483/CSA_VREF pixel
Xpixel_472 pixel_472/gring pixel_472/VDD pixel_472/GND pixel_472/VREF pixel_472/ROW_SEL
+ pixel_472/NB1 pixel_472/VBIAS pixel_472/NB2 pixel_472/AMP_IN pixel_472/SF_IB pixel_472/PIX_OUT
+ pixel_472/CSA_VREF pixel
Xpixel_461 pixel_461/gring pixel_461/VDD pixel_461/GND pixel_461/VREF pixel_461/ROW_SEL
+ pixel_461/NB1 pixel_461/VBIAS pixel_461/NB2 pixel_461/AMP_IN pixel_461/SF_IB pixel_461/PIX_OUT
+ pixel_461/CSA_VREF pixel
Xpixel_3743 pixel_3743/gring pixel_3743/VDD pixel_3743/GND pixel_3743/VREF pixel_3743/ROW_SEL
+ pixel_3743/NB1 pixel_3743/VBIAS pixel_3743/NB2 pixel_3743/AMP_IN pixel_3743/SF_IB
+ pixel_3743/PIX_OUT pixel_3743/CSA_VREF pixel
Xpixel_3732 pixel_3732/gring pixel_3732/VDD pixel_3732/GND pixel_3732/VREF pixel_3732/ROW_SEL
+ pixel_3732/NB1 pixel_3732/VBIAS pixel_3732/NB2 pixel_3732/AMP_IN pixel_3732/SF_IB
+ pixel_3732/PIX_OUT pixel_3732/CSA_VREF pixel
Xpixel_3721 pixel_3721/gring pixel_3721/VDD pixel_3721/GND pixel_3721/VREF pixel_3721/ROW_SEL
+ pixel_3721/NB1 pixel_3721/VBIAS pixel_3721/NB2 pixel_3721/AMP_IN pixel_3721/SF_IB
+ pixel_3721/PIX_OUT pixel_3721/CSA_VREF pixel
Xpixel_4455 pixel_4455/gring pixel_4455/VDD pixel_4455/GND pixel_4455/VREF pixel_4455/ROW_SEL
+ pixel_4455/NB1 pixel_4455/VBIAS pixel_4455/NB2 pixel_4455/AMP_IN pixel_4455/SF_IB
+ pixel_4455/PIX_OUT pixel_4455/CSA_VREF pixel
Xpixel_4466 pixel_4466/gring pixel_4466/VDD pixel_4466/GND pixel_4466/VREF pixel_4466/ROW_SEL
+ pixel_4466/NB1 pixel_4466/VBIAS pixel_4466/NB2 pixel_4466/AMP_IN pixel_4466/SF_IB
+ pixel_4466/PIX_OUT pixel_4466/CSA_VREF pixel
Xpixel_4477 pixel_4477/gring pixel_4477/VDD pixel_4477/GND pixel_4477/VREF pixel_4477/ROW_SEL
+ pixel_4477/NB1 pixel_4477/VBIAS pixel_4477/NB2 pixel_4477/AMP_IN pixel_4477/SF_IB
+ pixel_4477/PIX_OUT pixel_4477/CSA_VREF pixel
Xpixel_4488 pixel_4488/gring pixel_4488/VDD pixel_4488/GND pixel_4488/VREF pixel_4488/ROW_SEL
+ pixel_4488/NB1 pixel_4488/VBIAS pixel_4488/NB2 pixel_4488/AMP_IN pixel_4488/SF_IB
+ pixel_4488/PIX_OUT pixel_4488/CSA_VREF pixel
Xpixel_494 pixel_494/gring pixel_494/VDD pixel_494/GND pixel_494/VREF pixel_494/ROW_SEL
+ pixel_494/NB1 pixel_494/VBIAS pixel_494/NB2 pixel_494/AMP_IN pixel_494/SF_IB pixel_494/PIX_OUT
+ pixel_494/CSA_VREF pixel
Xpixel_3776 pixel_3776/gring pixel_3776/VDD pixel_3776/GND pixel_3776/VREF pixel_3776/ROW_SEL
+ pixel_3776/NB1 pixel_3776/VBIAS pixel_3776/NB2 pixel_3776/AMP_IN pixel_3776/SF_IB
+ pixel_3776/PIX_OUT pixel_3776/CSA_VREF pixel
Xpixel_3765 pixel_3765/gring pixel_3765/VDD pixel_3765/GND pixel_3765/VREF pixel_3765/ROW_SEL
+ pixel_3765/NB1 pixel_3765/VBIAS pixel_3765/NB2 pixel_3765/AMP_IN pixel_3765/SF_IB
+ pixel_3765/PIX_OUT pixel_3765/CSA_VREF pixel
Xpixel_3754 pixel_3754/gring pixel_3754/VDD pixel_3754/GND pixel_3754/VREF pixel_3754/ROW_SEL
+ pixel_3754/NB1 pixel_3754/VBIAS pixel_3754/NB2 pixel_3754/AMP_IN pixel_3754/SF_IB
+ pixel_3754/PIX_OUT pixel_3754/CSA_VREF pixel
Xpixel_4499 pixel_4499/gring pixel_4499/VDD pixel_4499/GND pixel_4499/VREF pixel_4499/ROW_SEL
+ pixel_4499/NB1 pixel_4499/VBIAS pixel_4499/NB2 pixel_4499/AMP_IN pixel_4499/SF_IB
+ pixel_4499/PIX_OUT pixel_4499/CSA_VREF pixel
Xpixel_3798 pixel_3798/gring pixel_3798/VDD pixel_3798/GND pixel_3798/VREF pixel_3798/ROW_SEL
+ pixel_3798/NB1 pixel_3798/VBIAS pixel_3798/NB2 pixel_3798/AMP_IN pixel_3798/SF_IB
+ pixel_3798/PIX_OUT pixel_3798/CSA_VREF pixel
Xpixel_3787 pixel_3787/gring pixel_3787/VDD pixel_3787/GND pixel_3787/VREF pixel_3787/ROW_SEL
+ pixel_3787/NB1 pixel_3787/VBIAS pixel_3787/NB2 pixel_3787/AMP_IN pixel_3787/SF_IB
+ pixel_3787/PIX_OUT pixel_3787/CSA_VREF pixel
Xpixel_7070 pixel_7070/gring pixel_7070/VDD pixel_7070/GND pixel_7070/VREF pixel_7070/ROW_SEL
+ pixel_7070/NB1 pixel_7070/VBIAS pixel_7070/NB2 pixel_7070/AMP_IN pixel_7070/SF_IB
+ pixel_7070/PIX_OUT pixel_7070/CSA_VREF pixel
Xpixel_7081 pixel_7081/gring pixel_7081/VDD pixel_7081/GND pixel_7081/VREF pixel_7081/ROW_SEL
+ pixel_7081/NB1 pixel_7081/VBIAS pixel_7081/NB2 pixel_7081/AMP_IN pixel_7081/SF_IB
+ pixel_7081/PIX_OUT pixel_7081/CSA_VREF pixel
Xpixel_7092 pixel_7092/gring pixel_7092/VDD pixel_7092/GND pixel_7092/VREF pixel_7092/ROW_SEL
+ pixel_7092/NB1 pixel_7092/VBIAS pixel_7092/NB2 pixel_7092/AMP_IN pixel_7092/SF_IB
+ pixel_7092/PIX_OUT pixel_7092/CSA_VREF pixel
Xpixel_6380 pixel_6380/gring pixel_6380/VDD pixel_6380/GND pixel_6380/VREF pixel_6380/ROW_SEL
+ pixel_6380/NB1 pixel_6380/VBIAS pixel_6380/NB2 pixel_6380/AMP_IN pixel_6380/SF_IB
+ pixel_6380/PIX_OUT pixel_6380/CSA_VREF pixel
Xpixel_6391 pixel_6391/gring pixel_6391/VDD pixel_6391/GND pixel_6391/VREF pixel_6391/ROW_SEL
+ pixel_6391/NB1 pixel_6391/VBIAS pixel_6391/NB2 pixel_6391/AMP_IN pixel_6391/SF_IB
+ pixel_6391/PIX_OUT pixel_6391/CSA_VREF pixel
Xpixel_5690 pixel_5690/gring pixel_5690/VDD pixel_5690/GND pixel_5690/VREF pixel_5690/ROW_SEL
+ pixel_5690/NB1 pixel_5690/VBIAS pixel_5690/NB2 pixel_5690/AMP_IN pixel_5690/SF_IB
+ pixel_5690/PIX_OUT pixel_5690/CSA_VREF pixel
Xpixel_3039 pixel_3039/gring pixel_3039/VDD pixel_3039/GND pixel_3039/VREF pixel_3039/ROW_SEL
+ pixel_3039/NB1 pixel_3039/VBIAS pixel_3039/NB2 pixel_3039/AMP_IN pixel_3039/SF_IB
+ pixel_3039/PIX_OUT pixel_3039/CSA_VREF pixel
Xpixel_3028 pixel_3028/gring pixel_3028/VDD pixel_3028/GND pixel_3028/VREF pixel_3028/ROW_SEL
+ pixel_3028/NB1 pixel_3028/VBIAS pixel_3028/NB2 pixel_3028/AMP_IN pixel_3028/SF_IB
+ pixel_3028/PIX_OUT pixel_3028/CSA_VREF pixel
Xpixel_3017 pixel_3017/gring pixel_3017/VDD pixel_3017/GND pixel_3017/VREF pixel_3017/ROW_SEL
+ pixel_3017/NB1 pixel_3017/VBIAS pixel_3017/NB2 pixel_3017/AMP_IN pixel_3017/SF_IB
+ pixel_3017/PIX_OUT pixel_3017/CSA_VREF pixel
Xpixel_3006 pixel_3006/gring pixel_3006/VDD pixel_3006/GND pixel_3006/VREF pixel_3006/ROW_SEL
+ pixel_3006/NB1 pixel_3006/VBIAS pixel_3006/NB2 pixel_3006/AMP_IN pixel_3006/SF_IB
+ pixel_3006/PIX_OUT pixel_3006/CSA_VREF pixel
Xpixel_2327 pixel_2327/gring pixel_2327/VDD pixel_2327/GND pixel_2327/VREF pixel_2327/ROW_SEL
+ pixel_2327/NB1 pixel_2327/VBIAS pixel_2327/NB2 pixel_2327/AMP_IN pixel_2327/SF_IB
+ pixel_2327/PIX_OUT pixel_2327/CSA_VREF pixel
Xpixel_2316 pixel_2316/gring pixel_2316/VDD pixel_2316/GND pixel_2316/VREF pixel_2316/ROW_SEL
+ pixel_2316/NB1 pixel_2316/VBIAS pixel_2316/NB2 pixel_2316/AMP_IN pixel_2316/SF_IB
+ pixel_2316/PIX_OUT pixel_2316/CSA_VREF pixel
Xpixel_2305 pixel_2305/gring pixel_2305/VDD pixel_2305/GND pixel_2305/VREF pixel_2305/ROW_SEL
+ pixel_2305/NB1 pixel_2305/VBIAS pixel_2305/NB2 pixel_2305/AMP_IN pixel_2305/SF_IB
+ pixel_2305/PIX_OUT pixel_2305/CSA_VREF pixel
Xpixel_1615 pixel_1615/gring pixel_1615/VDD pixel_1615/GND pixel_1615/VREF pixel_1615/ROW_SEL
+ pixel_1615/NB1 pixel_1615/VBIAS pixel_1615/NB2 pixel_1615/AMP_IN pixel_1615/SF_IB
+ pixel_1615/PIX_OUT pixel_1615/CSA_VREF pixel
Xpixel_1604 pixel_1604/gring pixel_1604/VDD pixel_1604/GND pixel_1604/VREF pixel_1604/ROW_SEL
+ pixel_1604/NB1 pixel_1604/VBIAS pixel_1604/NB2 pixel_1604/AMP_IN pixel_1604/SF_IB
+ pixel_1604/PIX_OUT pixel_1604/CSA_VREF pixel
Xpixel_2349 pixel_2349/gring pixel_2349/VDD pixel_2349/GND pixel_2349/VREF pixel_2349/ROW_SEL
+ pixel_2349/NB1 pixel_2349/VBIAS pixel_2349/NB2 pixel_2349/AMP_IN pixel_2349/SF_IB
+ pixel_2349/PIX_OUT pixel_2349/CSA_VREF pixel
Xpixel_2338 pixel_2338/gring pixel_2338/VDD pixel_2338/GND pixel_2338/VREF pixel_2338/ROW_SEL
+ pixel_2338/NB1 pixel_2338/VBIAS pixel_2338/NB2 pixel_2338/AMP_IN pixel_2338/SF_IB
+ pixel_2338/PIX_OUT pixel_2338/CSA_VREF pixel
Xpixel_1659 pixel_1659/gring pixel_1659/VDD pixel_1659/GND pixel_1659/VREF pixel_1659/ROW_SEL
+ pixel_1659/NB1 pixel_1659/VBIAS pixel_1659/NB2 pixel_1659/AMP_IN pixel_1659/SF_IB
+ pixel_1659/PIX_OUT pixel_1659/CSA_VREF pixel
Xpixel_1648 pixel_1648/gring pixel_1648/VDD pixel_1648/GND pixel_1648/VREF pixel_1648/ROW_SEL
+ pixel_1648/NB1 pixel_1648/VBIAS pixel_1648/NB2 pixel_1648/AMP_IN pixel_1648/SF_IB
+ pixel_1648/PIX_OUT pixel_1648/CSA_VREF pixel
Xpixel_1637 pixel_1637/gring pixel_1637/VDD pixel_1637/GND pixel_1637/VREF pixel_1637/ROW_SEL
+ pixel_1637/NB1 pixel_1637/VBIAS pixel_1637/NB2 pixel_1637/AMP_IN pixel_1637/SF_IB
+ pixel_1637/PIX_OUT pixel_1637/CSA_VREF pixel
Xpixel_1626 pixel_1626/gring pixel_1626/VDD pixel_1626/GND pixel_1626/VREF pixel_1626/ROW_SEL
+ pixel_1626/NB1 pixel_1626/VBIAS pixel_1626/NB2 pixel_1626/AMP_IN pixel_1626/SF_IB
+ pixel_1626/PIX_OUT pixel_1626/CSA_VREF pixel
Xpixel_9923 pixel_9923/gring pixel_9923/VDD pixel_9923/GND pixel_9923/VREF pixel_9923/ROW_SEL
+ pixel_9923/NB1 pixel_9923/VBIAS pixel_9923/NB2 pixel_9923/AMP_IN pixel_9923/SF_IB
+ pixel_9923/PIX_OUT pixel_9923/CSA_VREF pixel
Xpixel_9912 pixel_9912/gring pixel_9912/VDD pixel_9912/GND pixel_9912/VREF pixel_9912/ROW_SEL
+ pixel_9912/NB1 pixel_9912/VBIAS pixel_9912/NB2 pixel_9912/AMP_IN pixel_9912/SF_IB
+ pixel_9912/PIX_OUT pixel_9912/CSA_VREF pixel
Xpixel_9901 pixel_9901/gring pixel_9901/VDD pixel_9901/GND pixel_9901/VREF pixel_9901/ROW_SEL
+ pixel_9901/NB1 pixel_9901/VBIAS pixel_9901/NB2 pixel_9901/AMP_IN pixel_9901/SF_IB
+ pixel_9901/PIX_OUT pixel_9901/CSA_VREF pixel
Xpixel_9945 pixel_9945/gring pixel_9945/VDD pixel_9945/GND pixel_9945/VREF pixel_9945/ROW_SEL
+ pixel_9945/NB1 pixel_9945/VBIAS pixel_9945/NB2 pixel_9945/AMP_IN pixel_9945/SF_IB
+ pixel_9945/PIX_OUT pixel_9945/CSA_VREF pixel
Xpixel_9934 pixel_9934/gring pixel_9934/VDD pixel_9934/GND pixel_9934/VREF pixel_9934/ROW_SEL
+ pixel_9934/NB1 pixel_9934/VBIAS pixel_9934/NB2 pixel_9934/AMP_IN pixel_9934/SF_IB
+ pixel_9934/PIX_OUT pixel_9934/CSA_VREF pixel
Xpixel_9956 pixel_9956/gring pixel_9956/VDD pixel_9956/GND pixel_9956/VREF pixel_9956/ROW_SEL
+ pixel_9956/NB1 pixel_9956/VBIAS pixel_9956/NB2 pixel_9956/AMP_IN pixel_9956/SF_IB
+ pixel_9956/PIX_OUT pixel_9956/CSA_VREF pixel
Xpixel_9967 pixel_9967/gring pixel_9967/VDD pixel_9967/GND pixel_9967/VREF pixel_9967/ROW_SEL
+ pixel_9967/NB1 pixel_9967/VBIAS pixel_9967/NB2 pixel_9967/AMP_IN pixel_9967/SF_IB
+ pixel_9967/PIX_OUT pixel_9967/CSA_VREF pixel
Xpixel_9978 pixel_9978/gring pixel_9978/VDD pixel_9978/GND pixel_9978/VREF pixel_9978/ROW_SEL
+ pixel_9978/NB1 pixel_9978/VBIAS pixel_9978/NB2 pixel_9978/AMP_IN pixel_9978/SF_IB
+ pixel_9978/PIX_OUT pixel_9978/CSA_VREF pixel
Xpixel_9989 pixel_9989/gring pixel_9989/VDD pixel_9989/GND pixel_9989/VREF pixel_9989/ROW_SEL
+ pixel_9989/NB1 pixel_9989/VBIAS pixel_9989/NB2 pixel_9989/AMP_IN pixel_9989/SF_IB
+ pixel_9989/PIX_OUT pixel_9989/CSA_VREF pixel
Xpixel_4230 pixel_4230/gring pixel_4230/VDD pixel_4230/GND pixel_4230/VREF pixel_4230/ROW_SEL
+ pixel_4230/NB1 pixel_4230/VBIAS pixel_4230/NB2 pixel_4230/AMP_IN pixel_4230/SF_IB
+ pixel_4230/PIX_OUT pixel_4230/CSA_VREF pixel
Xpixel_4241 pixel_4241/gring pixel_4241/VDD pixel_4241/GND pixel_4241/VREF pixel_4241/ROW_SEL
+ pixel_4241/NB1 pixel_4241/VBIAS pixel_4241/NB2 pixel_4241/AMP_IN pixel_4241/SF_IB
+ pixel_4241/PIX_OUT pixel_4241/CSA_VREF pixel
Xpixel_4252 pixel_4252/gring pixel_4252/VDD pixel_4252/GND pixel_4252/VREF pixel_4252/ROW_SEL
+ pixel_4252/NB1 pixel_4252/VBIAS pixel_4252/NB2 pixel_4252/AMP_IN pixel_4252/SF_IB
+ pixel_4252/PIX_OUT pixel_4252/CSA_VREF pixel
Xpixel_4263 pixel_4263/gring pixel_4263/VDD pixel_4263/GND pixel_4263/VREF pixel_4263/ROW_SEL
+ pixel_4263/NB1 pixel_4263/VBIAS pixel_4263/NB2 pixel_4263/AMP_IN pixel_4263/SF_IB
+ pixel_4263/PIX_OUT pixel_4263/CSA_VREF pixel
Xpixel_291 pixel_291/gring pixel_291/VDD pixel_291/GND pixel_291/VREF pixel_291/ROW_SEL
+ pixel_291/NB1 pixel_291/VBIAS pixel_291/NB2 pixel_291/AMP_IN pixel_291/SF_IB pixel_291/PIX_OUT
+ pixel_291/CSA_VREF pixel
Xpixel_280 pixel_280/gring pixel_280/VDD pixel_280/GND pixel_280/VREF pixel_280/ROW_SEL
+ pixel_280/NB1 pixel_280/VBIAS pixel_280/NB2 pixel_280/AMP_IN pixel_280/SF_IB pixel_280/PIX_OUT
+ pixel_280/CSA_VREF pixel
Xpixel_3551 pixel_3551/gring pixel_3551/VDD pixel_3551/GND pixel_3551/VREF pixel_3551/ROW_SEL
+ pixel_3551/NB1 pixel_3551/VBIAS pixel_3551/NB2 pixel_3551/AMP_IN pixel_3551/SF_IB
+ pixel_3551/PIX_OUT pixel_3551/CSA_VREF pixel
Xpixel_3540 pixel_3540/gring pixel_3540/VDD pixel_3540/GND pixel_3540/VREF pixel_3540/ROW_SEL
+ pixel_3540/NB1 pixel_3540/VBIAS pixel_3540/NB2 pixel_3540/AMP_IN pixel_3540/SF_IB
+ pixel_3540/PIX_OUT pixel_3540/CSA_VREF pixel
Xpixel_4274 pixel_4274/gring pixel_4274/VDD pixel_4274/GND pixel_4274/VREF pixel_4274/ROW_SEL
+ pixel_4274/NB1 pixel_4274/VBIAS pixel_4274/NB2 pixel_4274/AMP_IN pixel_4274/SF_IB
+ pixel_4274/PIX_OUT pixel_4274/CSA_VREF pixel
Xpixel_4285 pixel_4285/gring pixel_4285/VDD pixel_4285/GND pixel_4285/VREF pixel_4285/ROW_SEL
+ pixel_4285/NB1 pixel_4285/VBIAS pixel_4285/NB2 pixel_4285/AMP_IN pixel_4285/SF_IB
+ pixel_4285/PIX_OUT pixel_4285/CSA_VREF pixel
Xpixel_4296 pixel_4296/gring pixel_4296/VDD pixel_4296/GND pixel_4296/VREF pixel_4296/ROW_SEL
+ pixel_4296/NB1 pixel_4296/VBIAS pixel_4296/NB2 pixel_4296/AMP_IN pixel_4296/SF_IB
+ pixel_4296/PIX_OUT pixel_4296/CSA_VREF pixel
Xpixel_2850 pixel_2850/gring pixel_2850/VDD pixel_2850/GND pixel_2850/VREF pixel_2850/ROW_SEL
+ pixel_2850/NB1 pixel_2850/VBIAS pixel_2850/NB2 pixel_2850/AMP_IN pixel_2850/SF_IB
+ pixel_2850/PIX_OUT pixel_2850/CSA_VREF pixel
Xpixel_3584 pixel_3584/gring pixel_3584/VDD pixel_3584/GND pixel_3584/VREF pixel_3584/ROW_SEL
+ pixel_3584/NB1 pixel_3584/VBIAS pixel_3584/NB2 pixel_3584/AMP_IN pixel_3584/SF_IB
+ pixel_3584/PIX_OUT pixel_3584/CSA_VREF pixel
Xpixel_3573 pixel_3573/gring pixel_3573/VDD pixel_3573/GND pixel_3573/VREF pixel_3573/ROW_SEL
+ pixel_3573/NB1 pixel_3573/VBIAS pixel_3573/NB2 pixel_3573/AMP_IN pixel_3573/SF_IB
+ pixel_3573/PIX_OUT pixel_3573/CSA_VREF pixel
Xpixel_3562 pixel_3562/gring pixel_3562/VDD pixel_3562/GND pixel_3562/VREF pixel_3562/ROW_SEL
+ pixel_3562/NB1 pixel_3562/VBIAS pixel_3562/NB2 pixel_3562/AMP_IN pixel_3562/SF_IB
+ pixel_3562/PIX_OUT pixel_3562/CSA_VREF pixel
Xpixel_2883 pixel_2883/gring pixel_2883/VDD pixel_2883/GND pixel_2883/VREF pixel_2883/ROW_SEL
+ pixel_2883/NB1 pixel_2883/VBIAS pixel_2883/NB2 pixel_2883/AMP_IN pixel_2883/SF_IB
+ pixel_2883/PIX_OUT pixel_2883/CSA_VREF pixel
Xpixel_2872 pixel_2872/gring pixel_2872/VDD pixel_2872/GND pixel_2872/VREF pixel_2872/ROW_SEL
+ pixel_2872/NB1 pixel_2872/VBIAS pixel_2872/NB2 pixel_2872/AMP_IN pixel_2872/SF_IB
+ pixel_2872/PIX_OUT pixel_2872/CSA_VREF pixel
Xpixel_2861 pixel_2861/gring pixel_2861/VDD pixel_2861/GND pixel_2861/VREF pixel_2861/ROW_SEL
+ pixel_2861/NB1 pixel_2861/VBIAS pixel_2861/NB2 pixel_2861/AMP_IN pixel_2861/SF_IB
+ pixel_2861/PIX_OUT pixel_2861/CSA_VREF pixel
Xpixel_3595 pixel_3595/gring pixel_3595/VDD pixel_3595/GND pixel_3595/VREF pixel_3595/ROW_SEL
+ pixel_3595/NB1 pixel_3595/VBIAS pixel_3595/NB2 pixel_3595/AMP_IN pixel_3595/SF_IB
+ pixel_3595/PIX_OUT pixel_3595/CSA_VREF pixel
Xpixel_2894 pixel_2894/gring pixel_2894/VDD pixel_2894/GND pixel_2894/VREF pixel_2894/ROW_SEL
+ pixel_2894/NB1 pixel_2894/VBIAS pixel_2894/NB2 pixel_2894/AMP_IN pixel_2894/SF_IB
+ pixel_2894/PIX_OUT pixel_2894/CSA_VREF pixel
Xpixel_9219 pixel_9219/gring pixel_9219/VDD pixel_9219/GND pixel_9219/VREF pixel_9219/ROW_SEL
+ pixel_9219/NB1 pixel_9219/VBIAS pixel_9219/NB2 pixel_9219/AMP_IN pixel_9219/SF_IB
+ pixel_9219/PIX_OUT pixel_9219/CSA_VREF pixel
Xpixel_9208 pixel_9208/gring pixel_9208/VDD pixel_9208/GND pixel_9208/VREF pixel_9208/ROW_SEL
+ pixel_9208/NB1 pixel_9208/VBIAS pixel_9208/NB2 pixel_9208/AMP_IN pixel_9208/SF_IB
+ pixel_9208/PIX_OUT pixel_9208/CSA_VREF pixel
Xpixel_8518 pixel_8518/gring pixel_8518/VDD pixel_8518/GND pixel_8518/VREF pixel_8518/ROW_SEL
+ pixel_8518/NB1 pixel_8518/VBIAS pixel_8518/NB2 pixel_8518/AMP_IN pixel_8518/SF_IB
+ pixel_8518/PIX_OUT pixel_8518/CSA_VREF pixel
Xpixel_8507 pixel_8507/gring pixel_8507/VDD pixel_8507/GND pixel_8507/VREF pixel_8507/ROW_SEL
+ pixel_8507/NB1 pixel_8507/VBIAS pixel_8507/NB2 pixel_8507/AMP_IN pixel_8507/SF_IB
+ pixel_8507/PIX_OUT pixel_8507/CSA_VREF pixel
Xpixel_8529 pixel_8529/gring pixel_8529/VDD pixel_8529/GND pixel_8529/VREF pixel_8529/ROW_SEL
+ pixel_8529/NB1 pixel_8529/VBIAS pixel_8529/NB2 pixel_8529/AMP_IN pixel_8529/SF_IB
+ pixel_8529/PIX_OUT pixel_8529/CSA_VREF pixel
Xpixel_7806 pixel_7806/gring pixel_7806/VDD pixel_7806/GND pixel_7806/VREF pixel_7806/ROW_SEL
+ pixel_7806/NB1 pixel_7806/VBIAS pixel_7806/NB2 pixel_7806/AMP_IN pixel_7806/SF_IB
+ pixel_7806/PIX_OUT pixel_7806/CSA_VREF pixel
Xpixel_7817 pixel_7817/gring pixel_7817/VDD pixel_7817/GND pixel_7817/VREF pixel_7817/ROW_SEL
+ pixel_7817/NB1 pixel_7817/VBIAS pixel_7817/NB2 pixel_7817/AMP_IN pixel_7817/SF_IB
+ pixel_7817/PIX_OUT pixel_7817/CSA_VREF pixel
Xpixel_7828 pixel_7828/gring pixel_7828/VDD pixel_7828/GND pixel_7828/VREF pixel_7828/ROW_SEL
+ pixel_7828/NB1 pixel_7828/VBIAS pixel_7828/NB2 pixel_7828/AMP_IN pixel_7828/SF_IB
+ pixel_7828/PIX_OUT pixel_7828/CSA_VREF pixel
Xpixel_7839 pixel_7839/gring pixel_7839/VDD pixel_7839/GND pixel_7839/VREF pixel_7839/ROW_SEL
+ pixel_7839/NB1 pixel_7839/VBIAS pixel_7839/NB2 pixel_7839/AMP_IN pixel_7839/SF_IB
+ pixel_7839/PIX_OUT pixel_7839/CSA_VREF pixel
Xpixel_2102 pixel_2102/gring pixel_2102/VDD pixel_2102/GND pixel_2102/VREF pixel_2102/ROW_SEL
+ pixel_2102/NB1 pixel_2102/VBIAS pixel_2102/NB2 pixel_2102/AMP_IN pixel_2102/SF_IB
+ pixel_2102/PIX_OUT pixel_2102/CSA_VREF pixel
Xpixel_2135 pixel_2135/gring pixel_2135/VDD pixel_2135/GND pixel_2135/VREF pixel_2135/ROW_SEL
+ pixel_2135/NB1 pixel_2135/VBIAS pixel_2135/NB2 pixel_2135/AMP_IN pixel_2135/SF_IB
+ pixel_2135/PIX_OUT pixel_2135/CSA_VREF pixel
Xpixel_2124 pixel_2124/gring pixel_2124/VDD pixel_2124/GND pixel_2124/VREF pixel_2124/ROW_SEL
+ pixel_2124/NB1 pixel_2124/VBIAS pixel_2124/NB2 pixel_2124/AMP_IN pixel_2124/SF_IB
+ pixel_2124/PIX_OUT pixel_2124/CSA_VREF pixel
Xpixel_2113 pixel_2113/gring pixel_2113/VDD pixel_2113/GND pixel_2113/VREF pixel_2113/ROW_SEL
+ pixel_2113/NB1 pixel_2113/VBIAS pixel_2113/NB2 pixel_2113/AMP_IN pixel_2113/SF_IB
+ pixel_2113/PIX_OUT pixel_2113/CSA_VREF pixel
Xpixel_1434 pixel_1434/gring pixel_1434/VDD pixel_1434/GND pixel_1434/VREF pixel_1434/ROW_SEL
+ pixel_1434/NB1 pixel_1434/VBIAS pixel_1434/NB2 pixel_1434/AMP_IN pixel_1434/SF_IB
+ pixel_1434/PIX_OUT pixel_1434/CSA_VREF pixel
Xpixel_1423 pixel_1423/gring pixel_1423/VDD pixel_1423/GND pixel_1423/VREF pixel_1423/ROW_SEL
+ pixel_1423/NB1 pixel_1423/VBIAS pixel_1423/NB2 pixel_1423/AMP_IN pixel_1423/SF_IB
+ pixel_1423/PIX_OUT pixel_1423/CSA_VREF pixel
Xpixel_1412 pixel_1412/gring pixel_1412/VDD pixel_1412/GND pixel_1412/VREF pixel_1412/ROW_SEL
+ pixel_1412/NB1 pixel_1412/VBIAS pixel_1412/NB2 pixel_1412/AMP_IN pixel_1412/SF_IB
+ pixel_1412/PIX_OUT pixel_1412/CSA_VREF pixel
Xpixel_1401 pixel_1401/gring pixel_1401/VDD pixel_1401/GND pixel_1401/VREF pixel_1401/ROW_SEL
+ pixel_1401/NB1 pixel_1401/VBIAS pixel_1401/NB2 pixel_1401/AMP_IN pixel_1401/SF_IB
+ pixel_1401/PIX_OUT pixel_1401/CSA_VREF pixel
Xpixel_2168 pixel_2168/gring pixel_2168/VDD pixel_2168/GND pixel_2168/VREF pixel_2168/ROW_SEL
+ pixel_2168/NB1 pixel_2168/VBIAS pixel_2168/NB2 pixel_2168/AMP_IN pixel_2168/SF_IB
+ pixel_2168/PIX_OUT pixel_2168/CSA_VREF pixel
Xpixel_2157 pixel_2157/gring pixel_2157/VDD pixel_2157/GND pixel_2157/VREF pixel_2157/ROW_SEL
+ pixel_2157/NB1 pixel_2157/VBIAS pixel_2157/NB2 pixel_2157/AMP_IN pixel_2157/SF_IB
+ pixel_2157/PIX_OUT pixel_2157/CSA_VREF pixel
Xpixel_2146 pixel_2146/gring pixel_2146/VDD pixel_2146/GND pixel_2146/VREF pixel_2146/ROW_SEL
+ pixel_2146/NB1 pixel_2146/VBIAS pixel_2146/NB2 pixel_2146/AMP_IN pixel_2146/SF_IB
+ pixel_2146/PIX_OUT pixel_2146/CSA_VREF pixel
Xpixel_1467 pixel_1467/gring pixel_1467/VDD pixel_1467/GND pixel_1467/VREF pixel_1467/ROW_SEL
+ pixel_1467/NB1 pixel_1467/VBIAS pixel_1467/NB2 pixel_1467/AMP_IN pixel_1467/SF_IB
+ pixel_1467/PIX_OUT pixel_1467/CSA_VREF pixel
Xpixel_1456 pixel_1456/gring pixel_1456/VDD pixel_1456/GND pixel_1456/VREF pixel_1456/ROW_SEL
+ pixel_1456/NB1 pixel_1456/VBIAS pixel_1456/NB2 pixel_1456/AMP_IN pixel_1456/SF_IB
+ pixel_1456/PIX_OUT pixel_1456/CSA_VREF pixel
Xpixel_1445 pixel_1445/gring pixel_1445/VDD pixel_1445/GND pixel_1445/VREF pixel_1445/ROW_SEL
+ pixel_1445/NB1 pixel_1445/VBIAS pixel_1445/NB2 pixel_1445/AMP_IN pixel_1445/SF_IB
+ pixel_1445/PIX_OUT pixel_1445/CSA_VREF pixel
Xpixel_2179 pixel_2179/gring pixel_2179/VDD pixel_2179/GND pixel_2179/VREF pixel_2179/ROW_SEL
+ pixel_2179/NB1 pixel_2179/VBIAS pixel_2179/NB2 pixel_2179/AMP_IN pixel_2179/SF_IB
+ pixel_2179/PIX_OUT pixel_2179/CSA_VREF pixel
Xpixel_1489 pixel_1489/gring pixel_1489/VDD pixel_1489/GND pixel_1489/VREF pixel_1489/ROW_SEL
+ pixel_1489/NB1 pixel_1489/VBIAS pixel_1489/NB2 pixel_1489/AMP_IN pixel_1489/SF_IB
+ pixel_1489/PIX_OUT pixel_1489/CSA_VREF pixel
Xpixel_1478 pixel_1478/gring pixel_1478/VDD pixel_1478/GND pixel_1478/VREF pixel_1478/ROW_SEL
+ pixel_1478/NB1 pixel_1478/VBIAS pixel_1478/NB2 pixel_1478/AMP_IN pixel_1478/SF_IB
+ pixel_1478/PIX_OUT pixel_1478/CSA_VREF pixel
Xpixel_9720 pixel_9720/gring pixel_9720/VDD pixel_9720/GND pixel_9720/VREF pixel_9720/ROW_SEL
+ pixel_9720/NB1 pixel_9720/VBIAS pixel_9720/NB2 pixel_9720/AMP_IN pixel_9720/SF_IB
+ pixel_9720/PIX_OUT pixel_9720/CSA_VREF pixel
Xpixel_9731 pixel_9731/gring pixel_9731/VDD pixel_9731/GND pixel_9731/VREF pixel_9731/ROW_SEL
+ pixel_9731/NB1 pixel_9731/VBIAS pixel_9731/NB2 pixel_9731/AMP_IN pixel_9731/SF_IB
+ pixel_9731/PIX_OUT pixel_9731/CSA_VREF pixel
Xpixel_9742 pixel_9742/gring pixel_9742/VDD pixel_9742/GND pixel_9742/VREF pixel_9742/ROW_SEL
+ pixel_9742/NB1 pixel_9742/VBIAS pixel_9742/NB2 pixel_9742/AMP_IN pixel_9742/SF_IB
+ pixel_9742/PIX_OUT pixel_9742/CSA_VREF pixel
Xpixel_9753 pixel_9753/gring pixel_9753/VDD pixel_9753/GND pixel_9753/VREF pixel_9753/ROW_SEL
+ pixel_9753/NB1 pixel_9753/VBIAS pixel_9753/NB2 pixel_9753/AMP_IN pixel_9753/SF_IB
+ pixel_9753/PIX_OUT pixel_9753/CSA_VREF pixel
Xpixel_9764 pixel_9764/gring pixel_9764/VDD pixel_9764/GND pixel_9764/VREF pixel_9764/ROW_SEL
+ pixel_9764/NB1 pixel_9764/VBIAS pixel_9764/NB2 pixel_9764/AMP_IN pixel_9764/SF_IB
+ pixel_9764/PIX_OUT pixel_9764/CSA_VREF pixel
Xpixel_9775 pixel_9775/gring pixel_9775/VDD pixel_9775/GND pixel_9775/VREF pixel_9775/ROW_SEL
+ pixel_9775/NB1 pixel_9775/VBIAS pixel_9775/NB2 pixel_9775/AMP_IN pixel_9775/SF_IB
+ pixel_9775/PIX_OUT pixel_9775/CSA_VREF pixel
Xpixel_9786 pixel_9786/gring pixel_9786/VDD pixel_9786/GND pixel_9786/VREF pixel_9786/ROW_SEL
+ pixel_9786/NB1 pixel_9786/VBIAS pixel_9786/NB2 pixel_9786/AMP_IN pixel_9786/SF_IB
+ pixel_9786/PIX_OUT pixel_9786/CSA_VREF pixel
Xpixel_9797 pixel_9797/gring pixel_9797/VDD pixel_9797/GND pixel_9797/VREF pixel_9797/ROW_SEL
+ pixel_9797/NB1 pixel_9797/VBIAS pixel_9797/NB2 pixel_9797/AMP_IN pixel_9797/SF_IB
+ pixel_9797/PIX_OUT pixel_9797/CSA_VREF pixel
Xpixel_4060 pixel_4060/gring pixel_4060/VDD pixel_4060/GND pixel_4060/VREF pixel_4060/ROW_SEL
+ pixel_4060/NB1 pixel_4060/VBIAS pixel_4060/NB2 pixel_4060/AMP_IN pixel_4060/SF_IB
+ pixel_4060/PIX_OUT pixel_4060/CSA_VREF pixel
Xpixel_4071 pixel_4071/gring pixel_4071/VDD pixel_4071/GND pixel_4071/VREF pixel_4071/ROW_SEL
+ pixel_4071/NB1 pixel_4071/VBIAS pixel_4071/NB2 pixel_4071/AMP_IN pixel_4071/SF_IB
+ pixel_4071/PIX_OUT pixel_4071/CSA_VREF pixel
Xpixel_4082 pixel_4082/gring pixel_4082/VDD pixel_4082/GND pixel_4082/VREF pixel_4082/ROW_SEL
+ pixel_4082/NB1 pixel_4082/VBIAS pixel_4082/NB2 pixel_4082/AMP_IN pixel_4082/SF_IB
+ pixel_4082/PIX_OUT pixel_4082/CSA_VREF pixel
Xpixel_4093 pixel_4093/gring pixel_4093/VDD pixel_4093/GND pixel_4093/VREF pixel_4093/ROW_SEL
+ pixel_4093/NB1 pixel_4093/VBIAS pixel_4093/NB2 pixel_4093/AMP_IN pixel_4093/SF_IB
+ pixel_4093/PIX_OUT pixel_4093/CSA_VREF pixel
Xpixel_3392 pixel_3392/gring pixel_3392/VDD pixel_3392/GND pixel_3392/VREF pixel_3392/ROW_SEL
+ pixel_3392/NB1 pixel_3392/VBIAS pixel_3392/NB2 pixel_3392/AMP_IN pixel_3392/SF_IB
+ pixel_3392/PIX_OUT pixel_3392/CSA_VREF pixel
Xpixel_3381 pixel_3381/gring pixel_3381/VDD pixel_3381/GND pixel_3381/VREF pixel_3381/ROW_SEL
+ pixel_3381/NB1 pixel_3381/VBIAS pixel_3381/NB2 pixel_3381/AMP_IN pixel_3381/SF_IB
+ pixel_3381/PIX_OUT pixel_3381/CSA_VREF pixel
Xpixel_3370 pixel_3370/gring pixel_3370/VDD pixel_3370/GND pixel_3370/VREF pixel_3370/ROW_SEL
+ pixel_3370/NB1 pixel_3370/VBIAS pixel_3370/NB2 pixel_3370/AMP_IN pixel_3370/SF_IB
+ pixel_3370/PIX_OUT pixel_3370/CSA_VREF pixel
Xpixel_2691 pixel_2691/gring pixel_2691/VDD pixel_2691/GND pixel_2691/VREF pixel_2691/ROW_SEL
+ pixel_2691/NB1 pixel_2691/VBIAS pixel_2691/NB2 pixel_2691/AMP_IN pixel_2691/SF_IB
+ pixel_2691/PIX_OUT pixel_2691/CSA_VREF pixel
Xpixel_2680 pixel_2680/gring pixel_2680/VDD pixel_2680/GND pixel_2680/VREF pixel_2680/ROW_SEL
+ pixel_2680/NB1 pixel_2680/VBIAS pixel_2680/NB2 pixel_2680/AMP_IN pixel_2680/SF_IB
+ pixel_2680/PIX_OUT pixel_2680/CSA_VREF pixel
Xpixel_1990 pixel_1990/gring pixel_1990/VDD pixel_1990/GND pixel_1990/VREF pixel_1990/ROW_SEL
+ pixel_1990/NB1 pixel_1990/VBIAS pixel_1990/NB2 pixel_1990/AMP_IN pixel_1990/SF_IB
+ pixel_1990/PIX_OUT pixel_1990/CSA_VREF pixel
Xpixel_9027 pixel_9027/gring pixel_9027/VDD pixel_9027/GND pixel_9027/VREF pixel_9027/ROW_SEL
+ pixel_9027/NB1 pixel_9027/VBIAS pixel_9027/NB2 pixel_9027/AMP_IN pixel_9027/SF_IB
+ pixel_9027/PIX_OUT pixel_9027/CSA_VREF pixel
Xpixel_9016 pixel_9016/gring pixel_9016/VDD pixel_9016/GND pixel_9016/VREF pixel_9016/ROW_SEL
+ pixel_9016/NB1 pixel_9016/VBIAS pixel_9016/NB2 pixel_9016/AMP_IN pixel_9016/SF_IB
+ pixel_9016/PIX_OUT pixel_9016/CSA_VREF pixel
Xpixel_9005 pixel_9005/gring pixel_9005/VDD pixel_9005/GND pixel_9005/VREF pixel_9005/ROW_SEL
+ pixel_9005/NB1 pixel_9005/VBIAS pixel_9005/NB2 pixel_9005/AMP_IN pixel_9005/SF_IB
+ pixel_9005/PIX_OUT pixel_9005/CSA_VREF pixel
Xpixel_9049 pixel_9049/gring pixel_9049/VDD pixel_9049/GND pixel_9049/VREF pixel_9049/ROW_SEL
+ pixel_9049/NB1 pixel_9049/VBIAS pixel_9049/NB2 pixel_9049/AMP_IN pixel_9049/SF_IB
+ pixel_9049/PIX_OUT pixel_9049/CSA_VREF pixel
Xpixel_9038 pixel_9038/gring pixel_9038/VDD pixel_9038/GND pixel_9038/VREF pixel_9038/ROW_SEL
+ pixel_9038/NB1 pixel_9038/VBIAS pixel_9038/NB2 pixel_9038/AMP_IN pixel_9038/SF_IB
+ pixel_9038/PIX_OUT pixel_9038/CSA_VREF pixel
Xpixel_8304 pixel_8304/gring pixel_8304/VDD pixel_8304/GND pixel_8304/VREF pixel_8304/ROW_SEL
+ pixel_8304/NB1 pixel_8304/VBIAS pixel_8304/NB2 pixel_8304/AMP_IN pixel_8304/SF_IB
+ pixel_8304/PIX_OUT pixel_8304/CSA_VREF pixel
Xpixel_8315 pixel_8315/gring pixel_8315/VDD pixel_8315/GND pixel_8315/VREF pixel_8315/ROW_SEL
+ pixel_8315/NB1 pixel_8315/VBIAS pixel_8315/NB2 pixel_8315/AMP_IN pixel_8315/SF_IB
+ pixel_8315/PIX_OUT pixel_8315/CSA_VREF pixel
Xpixel_8326 pixel_8326/gring pixel_8326/VDD pixel_8326/GND pixel_8326/VREF pixel_8326/ROW_SEL
+ pixel_8326/NB1 pixel_8326/VBIAS pixel_8326/NB2 pixel_8326/AMP_IN pixel_8326/SF_IB
+ pixel_8326/PIX_OUT pixel_8326/CSA_VREF pixel
Xpixel_8337 pixel_8337/gring pixel_8337/VDD pixel_8337/GND pixel_8337/VREF pixel_8337/ROW_SEL
+ pixel_8337/NB1 pixel_8337/VBIAS pixel_8337/NB2 pixel_8337/AMP_IN pixel_8337/SF_IB
+ pixel_8337/PIX_OUT pixel_8337/CSA_VREF pixel
Xpixel_8348 pixel_8348/gring pixel_8348/VDD pixel_8348/GND pixel_8348/VREF pixel_8348/ROW_SEL
+ pixel_8348/NB1 pixel_8348/VBIAS pixel_8348/NB2 pixel_8348/AMP_IN pixel_8348/SF_IB
+ pixel_8348/PIX_OUT pixel_8348/CSA_VREF pixel
Xpixel_8359 pixel_8359/gring pixel_8359/VDD pixel_8359/GND pixel_8359/VREF pixel_8359/ROW_SEL
+ pixel_8359/NB1 pixel_8359/VBIAS pixel_8359/NB2 pixel_8359/AMP_IN pixel_8359/SF_IB
+ pixel_8359/PIX_OUT pixel_8359/CSA_VREF pixel
Xpixel_7603 pixel_7603/gring pixel_7603/VDD pixel_7603/GND pixel_7603/VREF pixel_7603/ROW_SEL
+ pixel_7603/NB1 pixel_7603/VBIAS pixel_7603/NB2 pixel_7603/AMP_IN pixel_7603/SF_IB
+ pixel_7603/PIX_OUT pixel_7603/CSA_VREF pixel
Xpixel_7614 pixel_7614/gring pixel_7614/VDD pixel_7614/GND pixel_7614/VREF pixel_7614/ROW_SEL
+ pixel_7614/NB1 pixel_7614/VBIAS pixel_7614/NB2 pixel_7614/AMP_IN pixel_7614/SF_IB
+ pixel_7614/PIX_OUT pixel_7614/CSA_VREF pixel
Xpixel_7625 pixel_7625/gring pixel_7625/VDD pixel_7625/GND pixel_7625/VREF pixel_7625/ROW_SEL
+ pixel_7625/NB1 pixel_7625/VBIAS pixel_7625/NB2 pixel_7625/AMP_IN pixel_7625/SF_IB
+ pixel_7625/PIX_OUT pixel_7625/CSA_VREF pixel
Xpixel_7636 pixel_7636/gring pixel_7636/VDD pixel_7636/GND pixel_7636/VREF pixel_7636/ROW_SEL
+ pixel_7636/NB1 pixel_7636/VBIAS pixel_7636/NB2 pixel_7636/AMP_IN pixel_7636/SF_IB
+ pixel_7636/PIX_OUT pixel_7636/CSA_VREF pixel
Xpixel_7647 pixel_7647/gring pixel_7647/VDD pixel_7647/GND pixel_7647/VREF pixel_7647/ROW_SEL
+ pixel_7647/NB1 pixel_7647/VBIAS pixel_7647/NB2 pixel_7647/AMP_IN pixel_7647/SF_IB
+ pixel_7647/PIX_OUT pixel_7647/CSA_VREF pixel
Xpixel_6902 pixel_6902/gring pixel_6902/VDD pixel_6902/GND pixel_6902/VREF pixel_6902/ROW_SEL
+ pixel_6902/NB1 pixel_6902/VBIAS pixel_6902/NB2 pixel_6902/AMP_IN pixel_6902/SF_IB
+ pixel_6902/PIX_OUT pixel_6902/CSA_VREF pixel
Xpixel_6913 pixel_6913/gring pixel_6913/VDD pixel_6913/GND pixel_6913/VREF pixel_6913/ROW_SEL
+ pixel_6913/NB1 pixel_6913/VBIAS pixel_6913/NB2 pixel_6913/AMP_IN pixel_6913/SF_IB
+ pixel_6913/PIX_OUT pixel_6913/CSA_VREF pixel
Xpixel_7658 pixel_7658/gring pixel_7658/VDD pixel_7658/GND pixel_7658/VREF pixel_7658/ROW_SEL
+ pixel_7658/NB1 pixel_7658/VBIAS pixel_7658/NB2 pixel_7658/AMP_IN pixel_7658/SF_IB
+ pixel_7658/PIX_OUT pixel_7658/CSA_VREF pixel
Xpixel_7669 pixel_7669/gring pixel_7669/VDD pixel_7669/GND pixel_7669/VREF pixel_7669/ROW_SEL
+ pixel_7669/NB1 pixel_7669/VBIAS pixel_7669/NB2 pixel_7669/AMP_IN pixel_7669/SF_IB
+ pixel_7669/PIX_OUT pixel_7669/CSA_VREF pixel
Xpixel_6924 pixel_6924/gring pixel_6924/VDD pixel_6924/GND pixel_6924/VREF pixel_6924/ROW_SEL
+ pixel_6924/NB1 pixel_6924/VBIAS pixel_6924/NB2 pixel_6924/AMP_IN pixel_6924/SF_IB
+ pixel_6924/PIX_OUT pixel_6924/CSA_VREF pixel
Xpixel_6935 pixel_6935/gring pixel_6935/VDD pixel_6935/GND pixel_6935/VREF pixel_6935/ROW_SEL
+ pixel_6935/NB1 pixel_6935/VBIAS pixel_6935/NB2 pixel_6935/AMP_IN pixel_6935/SF_IB
+ pixel_6935/PIX_OUT pixel_6935/CSA_VREF pixel
Xpixel_6946 pixel_6946/gring pixel_6946/VDD pixel_6946/GND pixel_6946/VREF pixel_6946/ROW_SEL
+ pixel_6946/NB1 pixel_6946/VBIAS pixel_6946/NB2 pixel_6946/AMP_IN pixel_6946/SF_IB
+ pixel_6946/PIX_OUT pixel_6946/CSA_VREF pixel
Xpixel_27 pixel_27/gring pixel_27/VDD pixel_27/GND pixel_27/VREF pixel_27/ROW_SEL
+ pixel_27/NB1 pixel_27/VBIAS pixel_27/NB2 pixel_27/AMP_IN pixel_27/SF_IB pixel_27/PIX_OUT
+ pixel_27/CSA_VREF pixel
Xpixel_16 pixel_16/gring pixel_16/VDD pixel_16/GND pixel_16/VREF pixel_16/ROW_SEL
+ pixel_16/NB1 pixel_16/VBIAS pixel_16/NB2 pixel_16/AMP_IN pixel_16/SF_IB pixel_16/PIX_OUT
+ pixel_16/CSA_VREF pixel
Xpixel_6957 pixel_6957/gring pixel_6957/VDD pixel_6957/GND pixel_6957/VREF pixel_6957/ROW_SEL
+ pixel_6957/NB1 pixel_6957/VBIAS pixel_6957/NB2 pixel_6957/AMP_IN pixel_6957/SF_IB
+ pixel_6957/PIX_OUT pixel_6957/CSA_VREF pixel
Xpixel_6968 pixel_6968/gring pixel_6968/VDD pixel_6968/GND pixel_6968/VREF pixel_6968/ROW_SEL
+ pixel_6968/NB1 pixel_6968/VBIAS pixel_6968/NB2 pixel_6968/AMP_IN pixel_6968/SF_IB
+ pixel_6968/PIX_OUT pixel_6968/CSA_VREF pixel
Xpixel_6979 pixel_6979/gring pixel_6979/VDD pixel_6979/GND pixel_6979/VREF pixel_6979/ROW_SEL
+ pixel_6979/NB1 pixel_6979/VBIAS pixel_6979/NB2 pixel_6979/AMP_IN pixel_6979/SF_IB
+ pixel_6979/PIX_OUT pixel_6979/CSA_VREF pixel
Xpixel_49 pixel_49/gring pixel_49/VDD pixel_49/GND pixel_49/VREF pixel_49/ROW_SEL
+ pixel_49/NB1 pixel_49/VBIAS pixel_49/NB2 pixel_49/AMP_IN pixel_49/SF_IB pixel_49/PIX_OUT
+ pixel_49/CSA_VREF pixel
Xpixel_38 pixel_38/gring pixel_38/VDD pixel_38/GND pixel_38/VREF pixel_38/ROW_SEL
+ pixel_38/NB1 pixel_38/VBIAS pixel_38/NB2 pixel_38/AMP_IN pixel_38/SF_IB pixel_38/PIX_OUT
+ pixel_38/CSA_VREF pixel
Xpixel_1242 pixel_1242/gring pixel_1242/VDD pixel_1242/GND pixel_1242/VREF pixel_1242/ROW_SEL
+ pixel_1242/NB1 pixel_1242/VBIAS pixel_1242/NB2 pixel_1242/AMP_IN pixel_1242/SF_IB
+ pixel_1242/PIX_OUT pixel_1242/CSA_VREF pixel
Xpixel_1231 pixel_1231/gring pixel_1231/VDD pixel_1231/GND pixel_1231/VREF pixel_1231/ROW_SEL
+ pixel_1231/NB1 pixel_1231/VBIAS pixel_1231/NB2 pixel_1231/AMP_IN pixel_1231/SF_IB
+ pixel_1231/PIX_OUT pixel_1231/CSA_VREF pixel
Xpixel_1220 pixel_1220/gring pixel_1220/VDD pixel_1220/GND pixel_1220/VREF pixel_1220/ROW_SEL
+ pixel_1220/NB1 pixel_1220/VBIAS pixel_1220/NB2 pixel_1220/AMP_IN pixel_1220/SF_IB
+ pixel_1220/PIX_OUT pixel_1220/CSA_VREF pixel
Xpixel_1275 pixel_1275/gring pixel_1275/VDD pixel_1275/GND pixel_1275/VREF pixel_1275/ROW_SEL
+ pixel_1275/NB1 pixel_1275/VBIAS pixel_1275/NB2 pixel_1275/AMP_IN pixel_1275/SF_IB
+ pixel_1275/PIX_OUT pixel_1275/CSA_VREF pixel
Xpixel_1264 pixel_1264/gring pixel_1264/VDD pixel_1264/GND pixel_1264/VREF pixel_1264/ROW_SEL
+ pixel_1264/NB1 pixel_1264/VBIAS pixel_1264/NB2 pixel_1264/AMP_IN pixel_1264/SF_IB
+ pixel_1264/PIX_OUT pixel_1264/CSA_VREF pixel
Xpixel_1253 pixel_1253/gring pixel_1253/VDD pixel_1253/GND pixel_1253/VREF pixel_1253/ROW_SEL
+ pixel_1253/NB1 pixel_1253/VBIAS pixel_1253/NB2 pixel_1253/AMP_IN pixel_1253/SF_IB
+ pixel_1253/PIX_OUT pixel_1253/CSA_VREF pixel
Xpixel_1297 pixel_1297/gring pixel_1297/VDD pixel_1297/GND pixel_1297/VREF pixel_1297/ROW_SEL
+ pixel_1297/NB1 pixel_1297/VBIAS pixel_1297/NB2 pixel_1297/AMP_IN pixel_1297/SF_IB
+ pixel_1297/PIX_OUT pixel_1297/CSA_VREF pixel
Xpixel_1286 pixel_1286/gring pixel_1286/VDD pixel_1286/GND pixel_1286/VREF pixel_1286/ROW_SEL
+ pixel_1286/NB1 pixel_1286/VBIAS pixel_1286/NB2 pixel_1286/AMP_IN pixel_1286/SF_IB
+ pixel_1286/PIX_OUT pixel_1286/CSA_VREF pixel
Xpixel_9550 pixel_9550/gring pixel_9550/VDD pixel_9550/GND pixel_9550/VREF pixel_9550/ROW_SEL
+ pixel_9550/NB1 pixel_9550/VBIAS pixel_9550/NB2 pixel_9550/AMP_IN pixel_9550/SF_IB
+ pixel_9550/PIX_OUT pixel_9550/CSA_VREF pixel
Xpixel_9583 pixel_9583/gring pixel_9583/VDD pixel_9583/GND pixel_9583/VREF pixel_9583/ROW_SEL
+ pixel_9583/NB1 pixel_9583/VBIAS pixel_9583/NB2 pixel_9583/AMP_IN pixel_9583/SF_IB
+ pixel_9583/PIX_OUT pixel_9583/CSA_VREF pixel
Xpixel_9572 pixel_9572/gring pixel_9572/VDD pixel_9572/GND pixel_9572/VREF pixel_9572/ROW_SEL
+ pixel_9572/NB1 pixel_9572/VBIAS pixel_9572/NB2 pixel_9572/AMP_IN pixel_9572/SF_IB
+ pixel_9572/PIX_OUT pixel_9572/CSA_VREF pixel
Xpixel_9561 pixel_9561/gring pixel_9561/VDD pixel_9561/GND pixel_9561/VREF pixel_9561/ROW_SEL
+ pixel_9561/NB1 pixel_9561/VBIAS pixel_9561/NB2 pixel_9561/AMP_IN pixel_9561/SF_IB
+ pixel_9561/PIX_OUT pixel_9561/CSA_VREF pixel
Xpixel_8882 pixel_8882/gring pixel_8882/VDD pixel_8882/GND pixel_8882/VREF pixel_8882/ROW_SEL
+ pixel_8882/NB1 pixel_8882/VBIAS pixel_8882/NB2 pixel_8882/AMP_IN pixel_8882/SF_IB
+ pixel_8882/PIX_OUT pixel_8882/CSA_VREF pixel
Xpixel_8871 pixel_8871/gring pixel_8871/VDD pixel_8871/GND pixel_8871/VREF pixel_8871/ROW_SEL
+ pixel_8871/NB1 pixel_8871/VBIAS pixel_8871/NB2 pixel_8871/AMP_IN pixel_8871/SF_IB
+ pixel_8871/PIX_OUT pixel_8871/CSA_VREF pixel
Xpixel_8860 pixel_8860/gring pixel_8860/VDD pixel_8860/GND pixel_8860/VREF pixel_8860/ROW_SEL
+ pixel_8860/NB1 pixel_8860/VBIAS pixel_8860/NB2 pixel_8860/AMP_IN pixel_8860/SF_IB
+ pixel_8860/PIX_OUT pixel_8860/CSA_VREF pixel
Xpixel_9594 pixel_9594/gring pixel_9594/VDD pixel_9594/GND pixel_9594/VREF pixel_9594/ROW_SEL
+ pixel_9594/NB1 pixel_9594/VBIAS pixel_9594/NB2 pixel_9594/AMP_IN pixel_9594/SF_IB
+ pixel_9594/PIX_OUT pixel_9594/CSA_VREF pixel
Xpixel_8893 pixel_8893/gring pixel_8893/VDD pixel_8893/GND pixel_8893/VREF pixel_8893/ROW_SEL
+ pixel_8893/NB1 pixel_8893/VBIAS pixel_8893/NB2 pixel_8893/AMP_IN pixel_8893/SF_IB
+ pixel_8893/PIX_OUT pixel_8893/CSA_VREF pixel
Xpixel_6209 pixel_6209/gring pixel_6209/VDD pixel_6209/GND pixel_6209/VREF pixel_6209/ROW_SEL
+ pixel_6209/NB1 pixel_6209/VBIAS pixel_6209/NB2 pixel_6209/AMP_IN pixel_6209/SF_IB
+ pixel_6209/PIX_OUT pixel_6209/CSA_VREF pixel
Xpixel_5508 pixel_5508/gring pixel_5508/VDD pixel_5508/GND pixel_5508/VREF pixel_5508/ROW_SEL
+ pixel_5508/NB1 pixel_5508/VBIAS pixel_5508/NB2 pixel_5508/AMP_IN pixel_5508/SF_IB
+ pixel_5508/PIX_OUT pixel_5508/CSA_VREF pixel
Xpixel_5519 pixel_5519/gring pixel_5519/VDD pixel_5519/GND pixel_5519/VREF pixel_5519/ROW_SEL
+ pixel_5519/NB1 pixel_5519/VBIAS pixel_5519/NB2 pixel_5519/AMP_IN pixel_5519/SF_IB
+ pixel_5519/PIX_OUT pixel_5519/CSA_VREF pixel
Xpixel_824 pixel_824/gring pixel_824/VDD pixel_824/GND pixel_824/VREF pixel_824/ROW_SEL
+ pixel_824/NB1 pixel_824/VBIAS pixel_824/NB2 pixel_824/AMP_IN pixel_824/SF_IB pixel_824/PIX_OUT
+ pixel_824/CSA_VREF pixel
Xpixel_813 pixel_813/gring pixel_813/VDD pixel_813/GND pixel_813/VREF pixel_813/ROW_SEL
+ pixel_813/NB1 pixel_813/VBIAS pixel_813/NB2 pixel_813/AMP_IN pixel_813/SF_IB pixel_813/PIX_OUT
+ pixel_813/CSA_VREF pixel
Xpixel_802 pixel_802/gring pixel_802/VDD pixel_802/GND pixel_802/VREF pixel_802/ROW_SEL
+ pixel_802/NB1 pixel_802/VBIAS pixel_802/NB2 pixel_802/AMP_IN pixel_802/SF_IB pixel_802/PIX_OUT
+ pixel_802/CSA_VREF pixel
Xpixel_4807 pixel_4807/gring pixel_4807/VDD pixel_4807/GND pixel_4807/VREF pixel_4807/ROW_SEL
+ pixel_4807/NB1 pixel_4807/VBIAS pixel_4807/NB2 pixel_4807/AMP_IN pixel_4807/SF_IB
+ pixel_4807/PIX_OUT pixel_4807/CSA_VREF pixel
Xpixel_4818 pixel_4818/gring pixel_4818/VDD pixel_4818/GND pixel_4818/VREF pixel_4818/ROW_SEL
+ pixel_4818/NB1 pixel_4818/VBIAS pixel_4818/NB2 pixel_4818/AMP_IN pixel_4818/SF_IB
+ pixel_4818/PIX_OUT pixel_4818/CSA_VREF pixel
Xpixel_857 pixel_857/gring pixel_857/VDD pixel_857/GND pixel_857/VREF pixel_857/ROW_SEL
+ pixel_857/NB1 pixel_857/VBIAS pixel_857/NB2 pixel_857/AMP_IN pixel_857/SF_IB pixel_857/PIX_OUT
+ pixel_857/CSA_VREF pixel
Xpixel_846 pixel_846/gring pixel_846/VDD pixel_846/GND pixel_846/VREF pixel_846/ROW_SEL
+ pixel_846/NB1 pixel_846/VBIAS pixel_846/NB2 pixel_846/AMP_IN pixel_846/SF_IB pixel_846/PIX_OUT
+ pixel_846/CSA_VREF pixel
Xpixel_835 pixel_835/gring pixel_835/VDD pixel_835/GND pixel_835/VREF pixel_835/ROW_SEL
+ pixel_835/NB1 pixel_835/VBIAS pixel_835/NB2 pixel_835/AMP_IN pixel_835/SF_IB pixel_835/PIX_OUT
+ pixel_835/CSA_VREF pixel
Xpixel_4829 pixel_4829/gring pixel_4829/VDD pixel_4829/GND pixel_4829/VREF pixel_4829/ROW_SEL
+ pixel_4829/NB1 pixel_4829/VBIAS pixel_4829/NB2 pixel_4829/AMP_IN pixel_4829/SF_IB
+ pixel_4829/PIX_OUT pixel_4829/CSA_VREF pixel
Xpixel_879 pixel_879/gring pixel_879/VDD pixel_879/GND pixel_879/VREF pixel_879/ROW_SEL
+ pixel_879/NB1 pixel_879/VBIAS pixel_879/NB2 pixel_879/AMP_IN pixel_879/SF_IB pixel_879/PIX_OUT
+ pixel_879/CSA_VREF pixel
Xpixel_868 pixel_868/gring pixel_868/VDD pixel_868/GND pixel_868/VREF pixel_868/ROW_SEL
+ pixel_868/NB1 pixel_868/VBIAS pixel_868/NB2 pixel_868/AMP_IN pixel_868/SF_IB pixel_868/PIX_OUT
+ pixel_868/CSA_VREF pixel
Xpixel_8101 pixel_8101/gring pixel_8101/VDD pixel_8101/GND pixel_8101/VREF pixel_8101/ROW_SEL
+ pixel_8101/NB1 pixel_8101/VBIAS pixel_8101/NB2 pixel_8101/AMP_IN pixel_8101/SF_IB
+ pixel_8101/PIX_OUT pixel_8101/CSA_VREF pixel
Xpixel_8112 pixel_8112/gring pixel_8112/VDD pixel_8112/GND pixel_8112/VREF pixel_8112/ROW_SEL
+ pixel_8112/NB1 pixel_8112/VBIAS pixel_8112/NB2 pixel_8112/AMP_IN pixel_8112/SF_IB
+ pixel_8112/PIX_OUT pixel_8112/CSA_VREF pixel
Xpixel_8123 pixel_8123/gring pixel_8123/VDD pixel_8123/GND pixel_8123/VREF pixel_8123/ROW_SEL
+ pixel_8123/NB1 pixel_8123/VBIAS pixel_8123/NB2 pixel_8123/AMP_IN pixel_8123/SF_IB
+ pixel_8123/PIX_OUT pixel_8123/CSA_VREF pixel
Xpixel_8134 pixel_8134/gring pixel_8134/VDD pixel_8134/GND pixel_8134/VREF pixel_8134/ROW_SEL
+ pixel_8134/NB1 pixel_8134/VBIAS pixel_8134/NB2 pixel_8134/AMP_IN pixel_8134/SF_IB
+ pixel_8134/PIX_OUT pixel_8134/CSA_VREF pixel
Xpixel_8145 pixel_8145/gring pixel_8145/VDD pixel_8145/GND pixel_8145/VREF pixel_8145/ROW_SEL
+ pixel_8145/NB1 pixel_8145/VBIAS pixel_8145/NB2 pixel_8145/AMP_IN pixel_8145/SF_IB
+ pixel_8145/PIX_OUT pixel_8145/CSA_VREF pixel
Xpixel_8156 pixel_8156/gring pixel_8156/VDD pixel_8156/GND pixel_8156/VREF pixel_8156/ROW_SEL
+ pixel_8156/NB1 pixel_8156/VBIAS pixel_8156/NB2 pixel_8156/AMP_IN pixel_8156/SF_IB
+ pixel_8156/PIX_OUT pixel_8156/CSA_VREF pixel
Xpixel_8167 pixel_8167/gring pixel_8167/VDD pixel_8167/GND pixel_8167/VREF pixel_8167/ROW_SEL
+ pixel_8167/NB1 pixel_8167/VBIAS pixel_8167/NB2 pixel_8167/AMP_IN pixel_8167/SF_IB
+ pixel_8167/PIX_OUT pixel_8167/CSA_VREF pixel
Xpixel_7400 pixel_7400/gring pixel_7400/VDD pixel_7400/GND pixel_7400/VREF pixel_7400/ROW_SEL
+ pixel_7400/NB1 pixel_7400/VBIAS pixel_7400/NB2 pixel_7400/AMP_IN pixel_7400/SF_IB
+ pixel_7400/PIX_OUT pixel_7400/CSA_VREF pixel
Xpixel_7411 pixel_7411/gring pixel_7411/VDD pixel_7411/GND pixel_7411/VREF pixel_7411/ROW_SEL
+ pixel_7411/NB1 pixel_7411/VBIAS pixel_7411/NB2 pixel_7411/AMP_IN pixel_7411/SF_IB
+ pixel_7411/PIX_OUT pixel_7411/CSA_VREF pixel
Xpixel_7422 pixel_7422/gring pixel_7422/VDD pixel_7422/GND pixel_7422/VREF pixel_7422/ROW_SEL
+ pixel_7422/NB1 pixel_7422/VBIAS pixel_7422/NB2 pixel_7422/AMP_IN pixel_7422/SF_IB
+ pixel_7422/PIX_OUT pixel_7422/CSA_VREF pixel
Xpixel_8178 pixel_8178/gring pixel_8178/VDD pixel_8178/GND pixel_8178/VREF pixel_8178/ROW_SEL
+ pixel_8178/NB1 pixel_8178/VBIAS pixel_8178/NB2 pixel_8178/AMP_IN pixel_8178/SF_IB
+ pixel_8178/PIX_OUT pixel_8178/CSA_VREF pixel
Xpixel_8189 pixel_8189/gring pixel_8189/VDD pixel_8189/GND pixel_8189/VREF pixel_8189/ROW_SEL
+ pixel_8189/NB1 pixel_8189/VBIAS pixel_8189/NB2 pixel_8189/AMP_IN pixel_8189/SF_IB
+ pixel_8189/PIX_OUT pixel_8189/CSA_VREF pixel
Xpixel_7433 pixel_7433/gring pixel_7433/VDD pixel_7433/GND pixel_7433/VREF pixel_7433/ROW_SEL
+ pixel_7433/NB1 pixel_7433/VBIAS pixel_7433/NB2 pixel_7433/AMP_IN pixel_7433/SF_IB
+ pixel_7433/PIX_OUT pixel_7433/CSA_VREF pixel
Xpixel_7444 pixel_7444/gring pixel_7444/VDD pixel_7444/GND pixel_7444/VREF pixel_7444/ROW_SEL
+ pixel_7444/NB1 pixel_7444/VBIAS pixel_7444/NB2 pixel_7444/AMP_IN pixel_7444/SF_IB
+ pixel_7444/PIX_OUT pixel_7444/CSA_VREF pixel
Xpixel_7455 pixel_7455/gring pixel_7455/VDD pixel_7455/GND pixel_7455/VREF pixel_7455/ROW_SEL
+ pixel_7455/NB1 pixel_7455/VBIAS pixel_7455/NB2 pixel_7455/AMP_IN pixel_7455/SF_IB
+ pixel_7455/PIX_OUT pixel_7455/CSA_VREF pixel
Xpixel_7466 pixel_7466/gring pixel_7466/VDD pixel_7466/GND pixel_7466/VREF pixel_7466/ROW_SEL
+ pixel_7466/NB1 pixel_7466/VBIAS pixel_7466/NB2 pixel_7466/AMP_IN pixel_7466/SF_IB
+ pixel_7466/PIX_OUT pixel_7466/CSA_VREF pixel
Xpixel_6710 pixel_6710/gring pixel_6710/VDD pixel_6710/GND pixel_6710/VREF pixel_6710/ROW_SEL
+ pixel_6710/NB1 pixel_6710/VBIAS pixel_6710/NB2 pixel_6710/AMP_IN pixel_6710/SF_IB
+ pixel_6710/PIX_OUT pixel_6710/CSA_VREF pixel
Xpixel_6721 pixel_6721/gring pixel_6721/VDD pixel_6721/GND pixel_6721/VREF pixel_6721/ROW_SEL
+ pixel_6721/NB1 pixel_6721/VBIAS pixel_6721/NB2 pixel_6721/AMP_IN pixel_6721/SF_IB
+ pixel_6721/PIX_OUT pixel_6721/CSA_VREF pixel
Xpixel_7477 pixel_7477/gring pixel_7477/VDD pixel_7477/GND pixel_7477/VREF pixel_7477/ROW_SEL
+ pixel_7477/NB1 pixel_7477/VBIAS pixel_7477/NB2 pixel_7477/AMP_IN pixel_7477/SF_IB
+ pixel_7477/PIX_OUT pixel_7477/CSA_VREF pixel
Xpixel_7488 pixel_7488/gring pixel_7488/VDD pixel_7488/GND pixel_7488/VREF pixel_7488/ROW_SEL
+ pixel_7488/NB1 pixel_7488/VBIAS pixel_7488/NB2 pixel_7488/AMP_IN pixel_7488/SF_IB
+ pixel_7488/PIX_OUT pixel_7488/CSA_VREF pixel
Xpixel_7499 pixel_7499/gring pixel_7499/VDD pixel_7499/GND pixel_7499/VREF pixel_7499/ROW_SEL
+ pixel_7499/NB1 pixel_7499/VBIAS pixel_7499/NB2 pixel_7499/AMP_IN pixel_7499/SF_IB
+ pixel_7499/PIX_OUT pixel_7499/CSA_VREF pixel
Xpixel_6732 pixel_6732/gring pixel_6732/VDD pixel_6732/GND pixel_6732/VREF pixel_6732/ROW_SEL
+ pixel_6732/NB1 pixel_6732/VBIAS pixel_6732/NB2 pixel_6732/AMP_IN pixel_6732/SF_IB
+ pixel_6732/PIX_OUT pixel_6732/CSA_VREF pixel
Xpixel_6743 pixel_6743/gring pixel_6743/VDD pixel_6743/GND pixel_6743/VREF pixel_6743/ROW_SEL
+ pixel_6743/NB1 pixel_6743/VBIAS pixel_6743/NB2 pixel_6743/AMP_IN pixel_6743/SF_IB
+ pixel_6743/PIX_OUT pixel_6743/CSA_VREF pixel
Xpixel_6754 pixel_6754/gring pixel_6754/VDD pixel_6754/GND pixel_6754/VREF pixel_6754/ROW_SEL
+ pixel_6754/NB1 pixel_6754/VBIAS pixel_6754/NB2 pixel_6754/AMP_IN pixel_6754/SF_IB
+ pixel_6754/PIX_OUT pixel_6754/CSA_VREF pixel
Xpixel_6765 pixel_6765/gring pixel_6765/VDD pixel_6765/GND pixel_6765/VREF pixel_6765/ROW_SEL
+ pixel_6765/NB1 pixel_6765/VBIAS pixel_6765/NB2 pixel_6765/AMP_IN pixel_6765/SF_IB
+ pixel_6765/PIX_OUT pixel_6765/CSA_VREF pixel
Xpixel_6776 pixel_6776/gring pixel_6776/VDD pixel_6776/GND pixel_6776/VREF pixel_6776/ROW_SEL
+ pixel_6776/NB1 pixel_6776/VBIAS pixel_6776/NB2 pixel_6776/AMP_IN pixel_6776/SF_IB
+ pixel_6776/PIX_OUT pixel_6776/CSA_VREF pixel
Xpixel_6787 pixel_6787/gring pixel_6787/VDD pixel_6787/GND pixel_6787/VREF pixel_6787/ROW_SEL
+ pixel_6787/NB1 pixel_6787/VBIAS pixel_6787/NB2 pixel_6787/AMP_IN pixel_6787/SF_IB
+ pixel_6787/PIX_OUT pixel_6787/CSA_VREF pixel
Xpixel_6798 pixel_6798/gring pixel_6798/VDD pixel_6798/GND pixel_6798/VREF pixel_6798/ROW_SEL
+ pixel_6798/NB1 pixel_6798/VBIAS pixel_6798/NB2 pixel_6798/AMP_IN pixel_6798/SF_IB
+ pixel_6798/PIX_OUT pixel_6798/CSA_VREF pixel
Xpixel_1050 pixel_1050/gring pixel_1050/VDD pixel_1050/GND pixel_1050/VREF pixel_1050/ROW_SEL
+ pixel_1050/NB1 pixel_1050/VBIAS pixel_1050/NB2 pixel_1050/AMP_IN pixel_1050/SF_IB
+ pixel_1050/PIX_OUT pixel_1050/CSA_VREF pixel
Xpixel_1083 pixel_1083/gring pixel_1083/VDD pixel_1083/GND pixel_1083/VREF pixel_1083/ROW_SEL
+ pixel_1083/NB1 pixel_1083/VBIAS pixel_1083/NB2 pixel_1083/AMP_IN pixel_1083/SF_IB
+ pixel_1083/PIX_OUT pixel_1083/CSA_VREF pixel
Xpixel_1072 pixel_1072/gring pixel_1072/VDD pixel_1072/GND pixel_1072/VREF pixel_1072/ROW_SEL
+ pixel_1072/NB1 pixel_1072/VBIAS pixel_1072/NB2 pixel_1072/AMP_IN pixel_1072/SF_IB
+ pixel_1072/PIX_OUT pixel_1072/CSA_VREF pixel
Xpixel_1061 pixel_1061/gring pixel_1061/VDD pixel_1061/GND pixel_1061/VREF pixel_1061/ROW_SEL
+ pixel_1061/NB1 pixel_1061/VBIAS pixel_1061/NB2 pixel_1061/AMP_IN pixel_1061/SF_IB
+ pixel_1061/PIX_OUT pixel_1061/CSA_VREF pixel
Xpixel_1094 pixel_1094/gring pixel_1094/VDD pixel_1094/GND pixel_1094/VREF pixel_1094/ROW_SEL
+ pixel_1094/NB1 pixel_1094/VBIAS pixel_1094/NB2 pixel_1094/AMP_IN pixel_1094/SF_IB
+ pixel_1094/PIX_OUT pixel_1094/CSA_VREF pixel
Xpixel_9391 pixel_9391/gring pixel_9391/VDD pixel_9391/GND pixel_9391/VREF pixel_9391/ROW_SEL
+ pixel_9391/NB1 pixel_9391/VBIAS pixel_9391/NB2 pixel_9391/AMP_IN pixel_9391/SF_IB
+ pixel_9391/PIX_OUT pixel_9391/CSA_VREF pixel
Xpixel_9380 pixel_9380/gring pixel_9380/VDD pixel_9380/GND pixel_9380/VREF pixel_9380/ROW_SEL
+ pixel_9380/NB1 pixel_9380/VBIAS pixel_9380/NB2 pixel_9380/AMP_IN pixel_9380/SF_IB
+ pixel_9380/PIX_OUT pixel_9380/CSA_VREF pixel
Xpixel_8690 pixel_8690/gring pixel_8690/VDD pixel_8690/GND pixel_8690/VREF pixel_8690/ROW_SEL
+ pixel_8690/NB1 pixel_8690/VBIAS pixel_8690/NB2 pixel_8690/AMP_IN pixel_8690/SF_IB
+ pixel_8690/PIX_OUT pixel_8690/CSA_VREF pixel
Xpixel_109 pixel_109/gring pixel_109/VDD pixel_109/GND pixel_109/VREF pixel_109/ROW_SEL
+ pixel_109/NB1 pixel_109/VBIAS pixel_109/NB2 pixel_109/AMP_IN pixel_109/SF_IB pixel_109/PIX_OUT
+ pixel_109/CSA_VREF pixel
Xpixel_6006 pixel_6006/gring pixel_6006/VDD pixel_6006/GND pixel_6006/VREF pixel_6006/ROW_SEL
+ pixel_6006/NB1 pixel_6006/VBIAS pixel_6006/NB2 pixel_6006/AMP_IN pixel_6006/SF_IB
+ pixel_6006/PIX_OUT pixel_6006/CSA_VREF pixel
Xpixel_6017 pixel_6017/gring pixel_6017/VDD pixel_6017/GND pixel_6017/VREF pixel_6017/ROW_SEL
+ pixel_6017/NB1 pixel_6017/VBIAS pixel_6017/NB2 pixel_6017/AMP_IN pixel_6017/SF_IB
+ pixel_6017/PIX_OUT pixel_6017/CSA_VREF pixel
Xpixel_6028 pixel_6028/gring pixel_6028/VDD pixel_6028/GND pixel_6028/VREF pixel_6028/ROW_SEL
+ pixel_6028/NB1 pixel_6028/VBIAS pixel_6028/NB2 pixel_6028/AMP_IN pixel_6028/SF_IB
+ pixel_6028/PIX_OUT pixel_6028/CSA_VREF pixel
Xpixel_6039 pixel_6039/gring pixel_6039/VDD pixel_6039/GND pixel_6039/VREF pixel_6039/ROW_SEL
+ pixel_6039/NB1 pixel_6039/VBIAS pixel_6039/NB2 pixel_6039/AMP_IN pixel_6039/SF_IB
+ pixel_6039/PIX_OUT pixel_6039/CSA_VREF pixel
Xpixel_5305 pixel_5305/gring pixel_5305/VDD pixel_5305/GND pixel_5305/VREF pixel_5305/ROW_SEL
+ pixel_5305/NB1 pixel_5305/VBIAS pixel_5305/NB2 pixel_5305/AMP_IN pixel_5305/SF_IB
+ pixel_5305/PIX_OUT pixel_5305/CSA_VREF pixel
Xpixel_5316 pixel_5316/gring pixel_5316/VDD pixel_5316/GND pixel_5316/VREF pixel_5316/ROW_SEL
+ pixel_5316/NB1 pixel_5316/VBIAS pixel_5316/NB2 pixel_5316/AMP_IN pixel_5316/SF_IB
+ pixel_5316/PIX_OUT pixel_5316/CSA_VREF pixel
Xpixel_5327 pixel_5327/gring pixel_5327/VDD pixel_5327/GND pixel_5327/VREF pixel_5327/ROW_SEL
+ pixel_5327/NB1 pixel_5327/VBIAS pixel_5327/NB2 pixel_5327/AMP_IN pixel_5327/SF_IB
+ pixel_5327/PIX_OUT pixel_5327/CSA_VREF pixel
Xpixel_5338 pixel_5338/gring pixel_5338/VDD pixel_5338/GND pixel_5338/VREF pixel_5338/ROW_SEL
+ pixel_5338/NB1 pixel_5338/VBIAS pixel_5338/NB2 pixel_5338/AMP_IN pixel_5338/SF_IB
+ pixel_5338/PIX_OUT pixel_5338/CSA_VREF pixel
Xpixel_632 pixel_632/gring pixel_632/VDD pixel_632/GND pixel_632/VREF pixel_632/ROW_SEL
+ pixel_632/NB1 pixel_632/VBIAS pixel_632/NB2 pixel_632/AMP_IN pixel_632/SF_IB pixel_632/PIX_OUT
+ pixel_632/CSA_VREF pixel
Xpixel_621 pixel_621/gring pixel_621/VDD pixel_621/GND pixel_621/VREF pixel_621/ROW_SEL
+ pixel_621/NB1 pixel_621/VBIAS pixel_621/NB2 pixel_621/AMP_IN pixel_621/SF_IB pixel_621/PIX_OUT
+ pixel_621/CSA_VREF pixel
Xpixel_610 pixel_610/gring pixel_610/VDD pixel_610/GND pixel_610/VREF pixel_610/ROW_SEL
+ pixel_610/NB1 pixel_610/VBIAS pixel_610/NB2 pixel_610/AMP_IN pixel_610/SF_IB pixel_610/PIX_OUT
+ pixel_610/CSA_VREF pixel
Xpixel_5349 pixel_5349/gring pixel_5349/VDD pixel_5349/GND pixel_5349/VREF pixel_5349/ROW_SEL
+ pixel_5349/NB1 pixel_5349/VBIAS pixel_5349/NB2 pixel_5349/AMP_IN pixel_5349/SF_IB
+ pixel_5349/PIX_OUT pixel_5349/CSA_VREF pixel
Xpixel_4604 pixel_4604/gring pixel_4604/VDD pixel_4604/GND pixel_4604/VREF pixel_4604/ROW_SEL
+ pixel_4604/NB1 pixel_4604/VBIAS pixel_4604/NB2 pixel_4604/AMP_IN pixel_4604/SF_IB
+ pixel_4604/PIX_OUT pixel_4604/CSA_VREF pixel
Xpixel_4615 pixel_4615/gring pixel_4615/VDD pixel_4615/GND pixel_4615/VREF pixel_4615/ROW_SEL
+ pixel_4615/NB1 pixel_4615/VBIAS pixel_4615/NB2 pixel_4615/AMP_IN pixel_4615/SF_IB
+ pixel_4615/PIX_OUT pixel_4615/CSA_VREF pixel
Xpixel_4626 pixel_4626/gring pixel_4626/VDD pixel_4626/GND pixel_4626/VREF pixel_4626/ROW_SEL
+ pixel_4626/NB1 pixel_4626/VBIAS pixel_4626/NB2 pixel_4626/AMP_IN pixel_4626/SF_IB
+ pixel_4626/PIX_OUT pixel_4626/CSA_VREF pixel
Xpixel_4637 pixel_4637/gring pixel_4637/VDD pixel_4637/GND pixel_4637/VREF pixel_4637/ROW_SEL
+ pixel_4637/NB1 pixel_4637/VBIAS pixel_4637/NB2 pixel_4637/AMP_IN pixel_4637/SF_IB
+ pixel_4637/PIX_OUT pixel_4637/CSA_VREF pixel
Xpixel_665 pixel_665/gring pixel_665/VDD pixel_665/GND pixel_665/VREF pixel_665/ROW_SEL
+ pixel_665/NB1 pixel_665/VBIAS pixel_665/NB2 pixel_665/AMP_IN pixel_665/SF_IB pixel_665/PIX_OUT
+ pixel_665/CSA_VREF pixel
Xpixel_654 pixel_654/gring pixel_654/VDD pixel_654/GND pixel_654/VREF pixel_654/ROW_SEL
+ pixel_654/NB1 pixel_654/VBIAS pixel_654/NB2 pixel_654/AMP_IN pixel_654/SF_IB pixel_654/PIX_OUT
+ pixel_654/CSA_VREF pixel
Xpixel_643 pixel_643/gring pixel_643/VDD pixel_643/GND pixel_643/VREF pixel_643/ROW_SEL
+ pixel_643/NB1 pixel_643/VBIAS pixel_643/NB2 pixel_643/AMP_IN pixel_643/SF_IB pixel_643/PIX_OUT
+ pixel_643/CSA_VREF pixel
Xpixel_4648 pixel_4648/gring pixel_4648/VDD pixel_4648/GND pixel_4648/VREF pixel_4648/ROW_SEL
+ pixel_4648/NB1 pixel_4648/VBIAS pixel_4648/NB2 pixel_4648/AMP_IN pixel_4648/SF_IB
+ pixel_4648/PIX_OUT pixel_4648/CSA_VREF pixel
Xpixel_4659 pixel_4659/gring pixel_4659/VDD pixel_4659/GND pixel_4659/VREF pixel_4659/ROW_SEL
+ pixel_4659/NB1 pixel_4659/VBIAS pixel_4659/NB2 pixel_4659/AMP_IN pixel_4659/SF_IB
+ pixel_4659/PIX_OUT pixel_4659/CSA_VREF pixel
Xpixel_3903 pixel_3903/gring pixel_3903/VDD pixel_3903/GND pixel_3903/VREF pixel_3903/ROW_SEL
+ pixel_3903/NB1 pixel_3903/VBIAS pixel_3903/NB2 pixel_3903/AMP_IN pixel_3903/SF_IB
+ pixel_3903/PIX_OUT pixel_3903/CSA_VREF pixel
Xpixel_3914 pixel_3914/gring pixel_3914/VDD pixel_3914/GND pixel_3914/VREF pixel_3914/ROW_SEL
+ pixel_3914/NB1 pixel_3914/VBIAS pixel_3914/NB2 pixel_3914/AMP_IN pixel_3914/SF_IB
+ pixel_3914/PIX_OUT pixel_3914/CSA_VREF pixel
Xpixel_3925 pixel_3925/gring pixel_3925/VDD pixel_3925/GND pixel_3925/VREF pixel_3925/ROW_SEL
+ pixel_3925/NB1 pixel_3925/VBIAS pixel_3925/NB2 pixel_3925/AMP_IN pixel_3925/SF_IB
+ pixel_3925/PIX_OUT pixel_3925/CSA_VREF pixel
Xpixel_698 pixel_698/gring pixel_698/VDD pixel_698/GND pixel_698/VREF pixel_698/ROW_SEL
+ pixel_698/NB1 pixel_698/VBIAS pixel_698/NB2 pixel_698/AMP_IN pixel_698/SF_IB pixel_698/PIX_OUT
+ pixel_698/CSA_VREF pixel
Xpixel_687 pixel_687/gring pixel_687/VDD pixel_687/GND pixel_687/VREF pixel_687/ROW_SEL
+ pixel_687/NB1 pixel_687/VBIAS pixel_687/NB2 pixel_687/AMP_IN pixel_687/SF_IB pixel_687/PIX_OUT
+ pixel_687/CSA_VREF pixel
Xpixel_676 pixel_676/gring pixel_676/VDD pixel_676/GND pixel_676/VREF pixel_676/ROW_SEL
+ pixel_676/NB1 pixel_676/VBIAS pixel_676/NB2 pixel_676/AMP_IN pixel_676/SF_IB pixel_676/PIX_OUT
+ pixel_676/CSA_VREF pixel
Xpixel_3936 pixel_3936/gring pixel_3936/VDD pixel_3936/GND pixel_3936/VREF pixel_3936/ROW_SEL
+ pixel_3936/NB1 pixel_3936/VBIAS pixel_3936/NB2 pixel_3936/AMP_IN pixel_3936/SF_IB
+ pixel_3936/PIX_OUT pixel_3936/CSA_VREF pixel
Xpixel_3947 pixel_3947/gring pixel_3947/VDD pixel_3947/GND pixel_3947/VREF pixel_3947/ROW_SEL
+ pixel_3947/NB1 pixel_3947/VBIAS pixel_3947/NB2 pixel_3947/AMP_IN pixel_3947/SF_IB
+ pixel_3947/PIX_OUT pixel_3947/CSA_VREF pixel
Xpixel_3958 pixel_3958/gring pixel_3958/VDD pixel_3958/GND pixel_3958/VREF pixel_3958/ROW_SEL
+ pixel_3958/NB1 pixel_3958/VBIAS pixel_3958/NB2 pixel_3958/AMP_IN pixel_3958/SF_IB
+ pixel_3958/PIX_OUT pixel_3958/CSA_VREF pixel
Xpixel_3969 pixel_3969/gring pixel_3969/VDD pixel_3969/GND pixel_3969/VREF pixel_3969/ROW_SEL
+ pixel_3969/NB1 pixel_3969/VBIAS pixel_3969/NB2 pixel_3969/AMP_IN pixel_3969/SF_IB
+ pixel_3969/PIX_OUT pixel_3969/CSA_VREF pixel
Xpixel_7230 pixel_7230/gring pixel_7230/VDD pixel_7230/GND pixel_7230/VREF pixel_7230/ROW_SEL
+ pixel_7230/NB1 pixel_7230/VBIAS pixel_7230/NB2 pixel_7230/AMP_IN pixel_7230/SF_IB
+ pixel_7230/PIX_OUT pixel_7230/CSA_VREF pixel
Xpixel_7241 pixel_7241/gring pixel_7241/VDD pixel_7241/GND pixel_7241/VREF pixel_7241/ROW_SEL
+ pixel_7241/NB1 pixel_7241/VBIAS pixel_7241/NB2 pixel_7241/AMP_IN pixel_7241/SF_IB
+ pixel_7241/PIX_OUT pixel_7241/CSA_VREF pixel
Xpixel_7252 pixel_7252/gring pixel_7252/VDD pixel_7252/GND pixel_7252/VREF pixel_7252/ROW_SEL
+ pixel_7252/NB1 pixel_7252/VBIAS pixel_7252/NB2 pixel_7252/AMP_IN pixel_7252/SF_IB
+ pixel_7252/PIX_OUT pixel_7252/CSA_VREF pixel
Xpixel_7263 pixel_7263/gring pixel_7263/VDD pixel_7263/GND pixel_7263/VREF pixel_7263/ROW_SEL
+ pixel_7263/NB1 pixel_7263/VBIAS pixel_7263/NB2 pixel_7263/AMP_IN pixel_7263/SF_IB
+ pixel_7263/PIX_OUT pixel_7263/CSA_VREF pixel
Xpixel_7274 pixel_7274/gring pixel_7274/VDD pixel_7274/GND pixel_7274/VREF pixel_7274/ROW_SEL
+ pixel_7274/NB1 pixel_7274/VBIAS pixel_7274/NB2 pixel_7274/AMP_IN pixel_7274/SF_IB
+ pixel_7274/PIX_OUT pixel_7274/CSA_VREF pixel
Xpixel_7285 pixel_7285/gring pixel_7285/VDD pixel_7285/GND pixel_7285/VREF pixel_7285/ROW_SEL
+ pixel_7285/NB1 pixel_7285/VBIAS pixel_7285/NB2 pixel_7285/AMP_IN pixel_7285/SF_IB
+ pixel_7285/PIX_OUT pixel_7285/CSA_VREF pixel
Xpixel_7296 pixel_7296/gring pixel_7296/VDD pixel_7296/GND pixel_7296/VREF pixel_7296/ROW_SEL
+ pixel_7296/NB1 pixel_7296/VBIAS pixel_7296/NB2 pixel_7296/AMP_IN pixel_7296/SF_IB
+ pixel_7296/PIX_OUT pixel_7296/CSA_VREF pixel
Xpixel_6540 pixel_6540/gring pixel_6540/VDD pixel_6540/GND pixel_6540/VREF pixel_6540/ROW_SEL
+ pixel_6540/NB1 pixel_6540/VBIAS pixel_6540/NB2 pixel_6540/AMP_IN pixel_6540/SF_IB
+ pixel_6540/PIX_OUT pixel_6540/CSA_VREF pixel
Xpixel_6551 pixel_6551/gring pixel_6551/VDD pixel_6551/GND pixel_6551/VREF pixel_6551/ROW_SEL
+ pixel_6551/NB1 pixel_6551/VBIAS pixel_6551/NB2 pixel_6551/AMP_IN pixel_6551/SF_IB
+ pixel_6551/PIX_OUT pixel_6551/CSA_VREF pixel
Xpixel_6562 pixel_6562/gring pixel_6562/VDD pixel_6562/GND pixel_6562/VREF pixel_6562/ROW_SEL
+ pixel_6562/NB1 pixel_6562/VBIAS pixel_6562/NB2 pixel_6562/AMP_IN pixel_6562/SF_IB
+ pixel_6562/PIX_OUT pixel_6562/CSA_VREF pixel
Xpixel_6573 pixel_6573/gring pixel_6573/VDD pixel_6573/GND pixel_6573/VREF pixel_6573/ROW_SEL
+ pixel_6573/NB1 pixel_6573/VBIAS pixel_6573/NB2 pixel_6573/AMP_IN pixel_6573/SF_IB
+ pixel_6573/PIX_OUT pixel_6573/CSA_VREF pixel
Xpixel_6584 pixel_6584/gring pixel_6584/VDD pixel_6584/GND pixel_6584/VREF pixel_6584/ROW_SEL
+ pixel_6584/NB1 pixel_6584/VBIAS pixel_6584/NB2 pixel_6584/AMP_IN pixel_6584/SF_IB
+ pixel_6584/PIX_OUT pixel_6584/CSA_VREF pixel
Xpixel_6595 pixel_6595/gring pixel_6595/VDD pixel_6595/GND pixel_6595/VREF pixel_6595/ROW_SEL
+ pixel_6595/NB1 pixel_6595/VBIAS pixel_6595/NB2 pixel_6595/AMP_IN pixel_6595/SF_IB
+ pixel_6595/PIX_OUT pixel_6595/CSA_VREF pixel
Xpixel_5850 pixel_5850/gring pixel_5850/VDD pixel_5850/GND pixel_5850/VREF pixel_5850/ROW_SEL
+ pixel_5850/NB1 pixel_5850/VBIAS pixel_5850/NB2 pixel_5850/AMP_IN pixel_5850/SF_IB
+ pixel_5850/PIX_OUT pixel_5850/CSA_VREF pixel
Xpixel_5861 pixel_5861/gring pixel_5861/VDD pixel_5861/GND pixel_5861/VREF pixel_5861/ROW_SEL
+ pixel_5861/NB1 pixel_5861/VBIAS pixel_5861/NB2 pixel_5861/AMP_IN pixel_5861/SF_IB
+ pixel_5861/PIX_OUT pixel_5861/CSA_VREF pixel
Xpixel_5872 pixel_5872/gring pixel_5872/VDD pixel_5872/GND pixel_5872/VREF pixel_5872/ROW_SEL
+ pixel_5872/NB1 pixel_5872/VBIAS pixel_5872/NB2 pixel_5872/AMP_IN pixel_5872/SF_IB
+ pixel_5872/PIX_OUT pixel_5872/CSA_VREF pixel
Xpixel_5883 pixel_5883/gring pixel_5883/VDD pixel_5883/GND pixel_5883/VREF pixel_5883/ROW_SEL
+ pixel_5883/NB1 pixel_5883/VBIAS pixel_5883/NB2 pixel_5883/AMP_IN pixel_5883/SF_IB
+ pixel_5883/PIX_OUT pixel_5883/CSA_VREF pixel
Xpixel_5894 pixel_5894/gring pixel_5894/VDD pixel_5894/GND pixel_5894/VREF pixel_5894/ROW_SEL
+ pixel_5894/NB1 pixel_5894/VBIAS pixel_5894/NB2 pixel_5894/AMP_IN pixel_5894/SF_IB
+ pixel_5894/PIX_OUT pixel_5894/CSA_VREF pixel
Xpixel_2509 pixel_2509/gring pixel_2509/VDD pixel_2509/GND pixel_2509/VREF pixel_2509/ROW_SEL
+ pixel_2509/NB1 pixel_2509/VBIAS pixel_2509/NB2 pixel_2509/AMP_IN pixel_2509/SF_IB
+ pixel_2509/PIX_OUT pixel_2509/CSA_VREF pixel
Xpixel_1808 pixel_1808/gring pixel_1808/VDD pixel_1808/GND pixel_1808/VREF pixel_1808/ROW_SEL
+ pixel_1808/NB1 pixel_1808/VBIAS pixel_1808/NB2 pixel_1808/AMP_IN pixel_1808/SF_IB
+ pixel_1808/PIX_OUT pixel_1808/CSA_VREF pixel
Xpixel_1819 pixel_1819/gring pixel_1819/VDD pixel_1819/GND pixel_1819/VREF pixel_1819/ROW_SEL
+ pixel_1819/NB1 pixel_1819/VBIAS pixel_1819/NB2 pixel_1819/AMP_IN pixel_1819/SF_IB
+ pixel_1819/PIX_OUT pixel_1819/CSA_VREF pixel
Xpixel_5102 pixel_5102/gring pixel_5102/VDD pixel_5102/GND pixel_5102/VREF pixel_5102/ROW_SEL
+ pixel_5102/NB1 pixel_5102/VBIAS pixel_5102/NB2 pixel_5102/AMP_IN pixel_5102/SF_IB
+ pixel_5102/PIX_OUT pixel_5102/CSA_VREF pixel
Xpixel_5113 pixel_5113/gring pixel_5113/VDD pixel_5113/GND pixel_5113/VREF pixel_5113/ROW_SEL
+ pixel_5113/NB1 pixel_5113/VBIAS pixel_5113/NB2 pixel_5113/AMP_IN pixel_5113/SF_IB
+ pixel_5113/PIX_OUT pixel_5113/CSA_VREF pixel
Xpixel_5124 pixel_5124/gring pixel_5124/VDD pixel_5124/GND pixel_5124/VREF pixel_5124/ROW_SEL
+ pixel_5124/NB1 pixel_5124/VBIAS pixel_5124/NB2 pixel_5124/AMP_IN pixel_5124/SF_IB
+ pixel_5124/PIX_OUT pixel_5124/CSA_VREF pixel
Xpixel_5135 pixel_5135/gring pixel_5135/VDD pixel_5135/GND pixel_5135/VREF pixel_5135/ROW_SEL
+ pixel_5135/NB1 pixel_5135/VBIAS pixel_5135/NB2 pixel_5135/AMP_IN pixel_5135/SF_IB
+ pixel_5135/PIX_OUT pixel_5135/CSA_VREF pixel
Xpixel_5146 pixel_5146/gring pixel_5146/VDD pixel_5146/GND pixel_5146/VREF pixel_5146/ROW_SEL
+ pixel_5146/NB1 pixel_5146/VBIAS pixel_5146/NB2 pixel_5146/AMP_IN pixel_5146/SF_IB
+ pixel_5146/PIX_OUT pixel_5146/CSA_VREF pixel
Xpixel_4401 pixel_4401/gring pixel_4401/VDD pixel_4401/GND pixel_4401/VREF pixel_4401/ROW_SEL
+ pixel_4401/NB1 pixel_4401/VBIAS pixel_4401/NB2 pixel_4401/AMP_IN pixel_4401/SF_IB
+ pixel_4401/PIX_OUT pixel_4401/CSA_VREF pixel
Xpixel_4412 pixel_4412/gring pixel_4412/VDD pixel_4412/GND pixel_4412/VREF pixel_4412/ROW_SEL
+ pixel_4412/NB1 pixel_4412/VBIAS pixel_4412/NB2 pixel_4412/AMP_IN pixel_4412/SF_IB
+ pixel_4412/PIX_OUT pixel_4412/CSA_VREF pixel
Xpixel_440 pixel_440/gring pixel_440/VDD pixel_440/GND pixel_440/VREF pixel_440/ROW_SEL
+ pixel_440/NB1 pixel_440/VBIAS pixel_440/NB2 pixel_440/AMP_IN pixel_440/SF_IB pixel_440/PIX_OUT
+ pixel_440/CSA_VREF pixel
Xpixel_3700 pixel_3700/gring pixel_3700/VDD pixel_3700/GND pixel_3700/VREF pixel_3700/ROW_SEL
+ pixel_3700/NB1 pixel_3700/VBIAS pixel_3700/NB2 pixel_3700/AMP_IN pixel_3700/SF_IB
+ pixel_3700/PIX_OUT pixel_3700/CSA_VREF pixel
Xpixel_5157 pixel_5157/gring pixel_5157/VDD pixel_5157/GND pixel_5157/VREF pixel_5157/ROW_SEL
+ pixel_5157/NB1 pixel_5157/VBIAS pixel_5157/NB2 pixel_5157/AMP_IN pixel_5157/SF_IB
+ pixel_5157/PIX_OUT pixel_5157/CSA_VREF pixel
Xpixel_5168 pixel_5168/gring pixel_5168/VDD pixel_5168/GND pixel_5168/VREF pixel_5168/ROW_SEL
+ pixel_5168/NB1 pixel_5168/VBIAS pixel_5168/NB2 pixel_5168/AMP_IN pixel_5168/SF_IB
+ pixel_5168/PIX_OUT pixel_5168/CSA_VREF pixel
Xpixel_5179 pixel_5179/gring pixel_5179/VDD pixel_5179/GND pixel_5179/VREF pixel_5179/ROW_SEL
+ pixel_5179/NB1 pixel_5179/VBIAS pixel_5179/NB2 pixel_5179/AMP_IN pixel_5179/SF_IB
+ pixel_5179/PIX_OUT pixel_5179/CSA_VREF pixel
Xpixel_4423 pixel_4423/gring pixel_4423/VDD pixel_4423/GND pixel_4423/VREF pixel_4423/ROW_SEL
+ pixel_4423/NB1 pixel_4423/VBIAS pixel_4423/NB2 pixel_4423/AMP_IN pixel_4423/SF_IB
+ pixel_4423/PIX_OUT pixel_4423/CSA_VREF pixel
Xpixel_4434 pixel_4434/gring pixel_4434/VDD pixel_4434/GND pixel_4434/VREF pixel_4434/ROW_SEL
+ pixel_4434/NB1 pixel_4434/VBIAS pixel_4434/NB2 pixel_4434/AMP_IN pixel_4434/SF_IB
+ pixel_4434/PIX_OUT pixel_4434/CSA_VREF pixel
Xpixel_4445 pixel_4445/gring pixel_4445/VDD pixel_4445/GND pixel_4445/VREF pixel_4445/ROW_SEL
+ pixel_4445/NB1 pixel_4445/VBIAS pixel_4445/NB2 pixel_4445/AMP_IN pixel_4445/SF_IB
+ pixel_4445/PIX_OUT pixel_4445/CSA_VREF pixel
Xpixel_473 pixel_473/gring pixel_473/VDD pixel_473/GND pixel_473/VREF pixel_473/ROW_SEL
+ pixel_473/NB1 pixel_473/VBIAS pixel_473/NB2 pixel_473/AMP_IN pixel_473/SF_IB pixel_473/PIX_OUT
+ pixel_473/CSA_VREF pixel
Xpixel_462 pixel_462/gring pixel_462/VDD pixel_462/GND pixel_462/VREF pixel_462/ROW_SEL
+ pixel_462/NB1 pixel_462/VBIAS pixel_462/NB2 pixel_462/AMP_IN pixel_462/SF_IB pixel_462/PIX_OUT
+ pixel_462/CSA_VREF pixel
Xpixel_451 pixel_451/gring pixel_451/VDD pixel_451/GND pixel_451/VREF pixel_451/ROW_SEL
+ pixel_451/NB1 pixel_451/VBIAS pixel_451/NB2 pixel_451/AMP_IN pixel_451/SF_IB pixel_451/PIX_OUT
+ pixel_451/CSA_VREF pixel
Xpixel_3733 pixel_3733/gring pixel_3733/VDD pixel_3733/GND pixel_3733/VREF pixel_3733/ROW_SEL
+ pixel_3733/NB1 pixel_3733/VBIAS pixel_3733/NB2 pixel_3733/AMP_IN pixel_3733/SF_IB
+ pixel_3733/PIX_OUT pixel_3733/CSA_VREF pixel
Xpixel_3722 pixel_3722/gring pixel_3722/VDD pixel_3722/GND pixel_3722/VREF pixel_3722/ROW_SEL
+ pixel_3722/NB1 pixel_3722/VBIAS pixel_3722/NB2 pixel_3722/AMP_IN pixel_3722/SF_IB
+ pixel_3722/PIX_OUT pixel_3722/CSA_VREF pixel
Xpixel_3711 pixel_3711/gring pixel_3711/VDD pixel_3711/GND pixel_3711/VREF pixel_3711/ROW_SEL
+ pixel_3711/NB1 pixel_3711/VBIAS pixel_3711/NB2 pixel_3711/AMP_IN pixel_3711/SF_IB
+ pixel_3711/PIX_OUT pixel_3711/CSA_VREF pixel
Xpixel_4456 pixel_4456/gring pixel_4456/VDD pixel_4456/GND pixel_4456/VREF pixel_4456/ROW_SEL
+ pixel_4456/NB1 pixel_4456/VBIAS pixel_4456/NB2 pixel_4456/AMP_IN pixel_4456/SF_IB
+ pixel_4456/PIX_OUT pixel_4456/CSA_VREF pixel
Xpixel_4467 pixel_4467/gring pixel_4467/VDD pixel_4467/GND pixel_4467/VREF pixel_4467/ROW_SEL
+ pixel_4467/NB1 pixel_4467/VBIAS pixel_4467/NB2 pixel_4467/AMP_IN pixel_4467/SF_IB
+ pixel_4467/PIX_OUT pixel_4467/CSA_VREF pixel
Xpixel_4478 pixel_4478/gring pixel_4478/VDD pixel_4478/GND pixel_4478/VREF pixel_4478/ROW_SEL
+ pixel_4478/NB1 pixel_4478/VBIAS pixel_4478/NB2 pixel_4478/AMP_IN pixel_4478/SF_IB
+ pixel_4478/PIX_OUT pixel_4478/CSA_VREF pixel
Xpixel_495 pixel_495/gring pixel_495/VDD pixel_495/GND pixel_495/VREF pixel_495/ROW_SEL
+ pixel_495/NB1 pixel_495/VBIAS pixel_495/NB2 pixel_495/AMP_IN pixel_495/SF_IB pixel_495/PIX_OUT
+ pixel_495/CSA_VREF pixel
Xpixel_484 pixel_484/gring pixel_484/VDD pixel_484/GND pixel_484/VREF pixel_484/ROW_SEL
+ pixel_484/NB1 pixel_484/VBIAS pixel_484/NB2 pixel_484/AMP_IN pixel_484/SF_IB pixel_484/PIX_OUT
+ pixel_484/CSA_VREF pixel
Xpixel_3777 pixel_3777/gring pixel_3777/VDD pixel_3777/GND pixel_3777/VREF pixel_3777/ROW_SEL
+ pixel_3777/NB1 pixel_3777/VBIAS pixel_3777/NB2 pixel_3777/AMP_IN pixel_3777/SF_IB
+ pixel_3777/PIX_OUT pixel_3777/CSA_VREF pixel
Xpixel_3766 pixel_3766/gring pixel_3766/VDD pixel_3766/GND pixel_3766/VREF pixel_3766/ROW_SEL
+ pixel_3766/NB1 pixel_3766/VBIAS pixel_3766/NB2 pixel_3766/AMP_IN pixel_3766/SF_IB
+ pixel_3766/PIX_OUT pixel_3766/CSA_VREF pixel
Xpixel_3755 pixel_3755/gring pixel_3755/VDD pixel_3755/GND pixel_3755/VREF pixel_3755/ROW_SEL
+ pixel_3755/NB1 pixel_3755/VBIAS pixel_3755/NB2 pixel_3755/AMP_IN pixel_3755/SF_IB
+ pixel_3755/PIX_OUT pixel_3755/CSA_VREF pixel
Xpixel_3744 pixel_3744/gring pixel_3744/VDD pixel_3744/GND pixel_3744/VREF pixel_3744/ROW_SEL
+ pixel_3744/NB1 pixel_3744/VBIAS pixel_3744/NB2 pixel_3744/AMP_IN pixel_3744/SF_IB
+ pixel_3744/PIX_OUT pixel_3744/CSA_VREF pixel
Xpixel_4489 pixel_4489/gring pixel_4489/VDD pixel_4489/GND pixel_4489/VREF pixel_4489/ROW_SEL
+ pixel_4489/NB1 pixel_4489/VBIAS pixel_4489/NB2 pixel_4489/AMP_IN pixel_4489/SF_IB
+ pixel_4489/PIX_OUT pixel_4489/CSA_VREF pixel
Xpixel_3799 pixel_3799/gring pixel_3799/VDD pixel_3799/GND pixel_3799/VREF pixel_3799/ROW_SEL
+ pixel_3799/NB1 pixel_3799/VBIAS pixel_3799/NB2 pixel_3799/AMP_IN pixel_3799/SF_IB
+ pixel_3799/PIX_OUT pixel_3799/CSA_VREF pixel
Xpixel_3788 pixel_3788/gring pixel_3788/VDD pixel_3788/GND pixel_3788/VREF pixel_3788/ROW_SEL
+ pixel_3788/NB1 pixel_3788/VBIAS pixel_3788/NB2 pixel_3788/AMP_IN pixel_3788/SF_IB
+ pixel_3788/PIX_OUT pixel_3788/CSA_VREF pixel
Xpixel_7060 pixel_7060/gring pixel_7060/VDD pixel_7060/GND pixel_7060/VREF pixel_7060/ROW_SEL
+ pixel_7060/NB1 pixel_7060/VBIAS pixel_7060/NB2 pixel_7060/AMP_IN pixel_7060/SF_IB
+ pixel_7060/PIX_OUT pixel_7060/CSA_VREF pixel
Xpixel_7071 pixel_7071/gring pixel_7071/VDD pixel_7071/GND pixel_7071/VREF pixel_7071/ROW_SEL
+ pixel_7071/NB1 pixel_7071/VBIAS pixel_7071/NB2 pixel_7071/AMP_IN pixel_7071/SF_IB
+ pixel_7071/PIX_OUT pixel_7071/CSA_VREF pixel
Xpixel_7082 pixel_7082/gring pixel_7082/VDD pixel_7082/GND pixel_7082/VREF pixel_7082/ROW_SEL
+ pixel_7082/NB1 pixel_7082/VBIAS pixel_7082/NB2 pixel_7082/AMP_IN pixel_7082/SF_IB
+ pixel_7082/PIX_OUT pixel_7082/CSA_VREF pixel
Xpixel_7093 pixel_7093/gring pixel_7093/VDD pixel_7093/GND pixel_7093/VREF pixel_7093/ROW_SEL
+ pixel_7093/NB1 pixel_7093/VBIAS pixel_7093/NB2 pixel_7093/AMP_IN pixel_7093/SF_IB
+ pixel_7093/PIX_OUT pixel_7093/CSA_VREF pixel
Xpixel_6370 pixel_6370/gring pixel_6370/VDD pixel_6370/GND pixel_6370/VREF pixel_6370/ROW_SEL
+ pixel_6370/NB1 pixel_6370/VBIAS pixel_6370/NB2 pixel_6370/AMP_IN pixel_6370/SF_IB
+ pixel_6370/PIX_OUT pixel_6370/CSA_VREF pixel
Xpixel_6381 pixel_6381/gring pixel_6381/VDD pixel_6381/GND pixel_6381/VREF pixel_6381/ROW_SEL
+ pixel_6381/NB1 pixel_6381/VBIAS pixel_6381/NB2 pixel_6381/AMP_IN pixel_6381/SF_IB
+ pixel_6381/PIX_OUT pixel_6381/CSA_VREF pixel
Xpixel_6392 pixel_6392/gring pixel_6392/VDD pixel_6392/GND pixel_6392/VREF pixel_6392/ROW_SEL
+ pixel_6392/NB1 pixel_6392/VBIAS pixel_6392/NB2 pixel_6392/AMP_IN pixel_6392/SF_IB
+ pixel_6392/PIX_OUT pixel_6392/CSA_VREF pixel
Xpixel_5680 pixel_5680/gring pixel_5680/VDD pixel_5680/GND pixel_5680/VREF pixel_5680/ROW_SEL
+ pixel_5680/NB1 pixel_5680/VBIAS pixel_5680/NB2 pixel_5680/AMP_IN pixel_5680/SF_IB
+ pixel_5680/PIX_OUT pixel_5680/CSA_VREF pixel
Xpixel_5691 pixel_5691/gring pixel_5691/VDD pixel_5691/GND pixel_5691/VREF pixel_5691/ROW_SEL
+ pixel_5691/NB1 pixel_5691/VBIAS pixel_5691/NB2 pixel_5691/AMP_IN pixel_5691/SF_IB
+ pixel_5691/PIX_OUT pixel_5691/CSA_VREF pixel
Xpixel_4990 pixel_4990/gring pixel_4990/VDD pixel_4990/GND pixel_4990/VREF pixel_4990/ROW_SEL
+ pixel_4990/NB1 pixel_4990/VBIAS pixel_4990/NB2 pixel_4990/AMP_IN pixel_4990/SF_IB
+ pixel_4990/PIX_OUT pixel_4990/CSA_VREF pixel
Xpixel_3029 pixel_3029/gring pixel_3029/VDD pixel_3029/GND pixel_3029/VREF pixel_3029/ROW_SEL
+ pixel_3029/NB1 pixel_3029/VBIAS pixel_3029/NB2 pixel_3029/AMP_IN pixel_3029/SF_IB
+ pixel_3029/PIX_OUT pixel_3029/CSA_VREF pixel
Xpixel_3018 pixel_3018/gring pixel_3018/VDD pixel_3018/GND pixel_3018/VREF pixel_3018/ROW_SEL
+ pixel_3018/NB1 pixel_3018/VBIAS pixel_3018/NB2 pixel_3018/AMP_IN pixel_3018/SF_IB
+ pixel_3018/PIX_OUT pixel_3018/CSA_VREF pixel
Xpixel_3007 pixel_3007/gring pixel_3007/VDD pixel_3007/GND pixel_3007/VREF pixel_3007/ROW_SEL
+ pixel_3007/NB1 pixel_3007/VBIAS pixel_3007/NB2 pixel_3007/AMP_IN pixel_3007/SF_IB
+ pixel_3007/PIX_OUT pixel_3007/CSA_VREF pixel
Xpixel_2317 pixel_2317/gring pixel_2317/VDD pixel_2317/GND pixel_2317/VREF pixel_2317/ROW_SEL
+ pixel_2317/NB1 pixel_2317/VBIAS pixel_2317/NB2 pixel_2317/AMP_IN pixel_2317/SF_IB
+ pixel_2317/PIX_OUT pixel_2317/CSA_VREF pixel
Xpixel_2306 pixel_2306/gring pixel_2306/VDD pixel_2306/GND pixel_2306/VREF pixel_2306/ROW_SEL
+ pixel_2306/NB1 pixel_2306/VBIAS pixel_2306/NB2 pixel_2306/AMP_IN pixel_2306/SF_IB
+ pixel_2306/PIX_OUT pixel_2306/CSA_VREF pixel
Xpixel_1616 pixel_1616/gring pixel_1616/VDD pixel_1616/GND pixel_1616/VREF pixel_1616/ROW_SEL
+ pixel_1616/NB1 pixel_1616/VBIAS pixel_1616/NB2 pixel_1616/AMP_IN pixel_1616/SF_IB
+ pixel_1616/PIX_OUT pixel_1616/CSA_VREF pixel
Xpixel_1605 pixel_1605/gring pixel_1605/VDD pixel_1605/GND pixel_1605/VREF pixel_1605/ROW_SEL
+ pixel_1605/NB1 pixel_1605/VBIAS pixel_1605/NB2 pixel_1605/AMP_IN pixel_1605/SF_IB
+ pixel_1605/PIX_OUT pixel_1605/CSA_VREF pixel
Xpixel_2339 pixel_2339/gring pixel_2339/VDD pixel_2339/GND pixel_2339/VREF pixel_2339/ROW_SEL
+ pixel_2339/NB1 pixel_2339/VBIAS pixel_2339/NB2 pixel_2339/AMP_IN pixel_2339/SF_IB
+ pixel_2339/PIX_OUT pixel_2339/CSA_VREF pixel
Xpixel_2328 pixel_2328/gring pixel_2328/VDD pixel_2328/GND pixel_2328/VREF pixel_2328/ROW_SEL
+ pixel_2328/NB1 pixel_2328/VBIAS pixel_2328/NB2 pixel_2328/AMP_IN pixel_2328/SF_IB
+ pixel_2328/PIX_OUT pixel_2328/CSA_VREF pixel
Xpixel_1649 pixel_1649/gring pixel_1649/VDD pixel_1649/GND pixel_1649/VREF pixel_1649/ROW_SEL
+ pixel_1649/NB1 pixel_1649/VBIAS pixel_1649/NB2 pixel_1649/AMP_IN pixel_1649/SF_IB
+ pixel_1649/PIX_OUT pixel_1649/CSA_VREF pixel
Xpixel_1638 pixel_1638/gring pixel_1638/VDD pixel_1638/GND pixel_1638/VREF pixel_1638/ROW_SEL
+ pixel_1638/NB1 pixel_1638/VBIAS pixel_1638/NB2 pixel_1638/AMP_IN pixel_1638/SF_IB
+ pixel_1638/PIX_OUT pixel_1638/CSA_VREF pixel
Xpixel_1627 pixel_1627/gring pixel_1627/VDD pixel_1627/GND pixel_1627/VREF pixel_1627/ROW_SEL
+ pixel_1627/NB1 pixel_1627/VBIAS pixel_1627/NB2 pixel_1627/AMP_IN pixel_1627/SF_IB
+ pixel_1627/PIX_OUT pixel_1627/CSA_VREF pixel
Xpixel_9924 pixel_9924/gring pixel_9924/VDD pixel_9924/GND pixel_9924/VREF pixel_9924/ROW_SEL
+ pixel_9924/NB1 pixel_9924/VBIAS pixel_9924/NB2 pixel_9924/AMP_IN pixel_9924/SF_IB
+ pixel_9924/PIX_OUT pixel_9924/CSA_VREF pixel
Xpixel_9913 pixel_9913/gring pixel_9913/VDD pixel_9913/GND pixel_9913/VREF pixel_9913/ROW_SEL
+ pixel_9913/NB1 pixel_9913/VBIAS pixel_9913/NB2 pixel_9913/AMP_IN pixel_9913/SF_IB
+ pixel_9913/PIX_OUT pixel_9913/CSA_VREF pixel
Xpixel_9902 pixel_9902/gring pixel_9902/VDD pixel_9902/GND pixel_9902/VREF pixel_9902/ROW_SEL
+ pixel_9902/NB1 pixel_9902/VBIAS pixel_9902/NB2 pixel_9902/AMP_IN pixel_9902/SF_IB
+ pixel_9902/PIX_OUT pixel_9902/CSA_VREF pixel
Xpixel_9946 pixel_9946/gring pixel_9946/VDD pixel_9946/GND pixel_9946/VREF pixel_9946/ROW_SEL
+ pixel_9946/NB1 pixel_9946/VBIAS pixel_9946/NB2 pixel_9946/AMP_IN pixel_9946/SF_IB
+ pixel_9946/PIX_OUT pixel_9946/CSA_VREF pixel
Xpixel_9935 pixel_9935/gring pixel_9935/VDD pixel_9935/GND pixel_9935/VREF pixel_9935/ROW_SEL
+ pixel_9935/NB1 pixel_9935/VBIAS pixel_9935/NB2 pixel_9935/AMP_IN pixel_9935/SF_IB
+ pixel_9935/PIX_OUT pixel_9935/CSA_VREF pixel
Xpixel_9957 pixel_9957/gring pixel_9957/VDD pixel_9957/GND pixel_9957/VREF pixel_9957/ROW_SEL
+ pixel_9957/NB1 pixel_9957/VBIAS pixel_9957/NB2 pixel_9957/AMP_IN pixel_9957/SF_IB
+ pixel_9957/PIX_OUT pixel_9957/CSA_VREF pixel
Xpixel_9968 pixel_9968/gring pixel_9968/VDD pixel_9968/GND pixel_9968/VREF pixel_9968/ROW_SEL
+ pixel_9968/NB1 pixel_9968/VBIAS pixel_9968/NB2 pixel_9968/AMP_IN pixel_9968/SF_IB
+ pixel_9968/PIX_OUT pixel_9968/CSA_VREF pixel
Xpixel_9979 pixel_9979/gring pixel_9979/VDD pixel_9979/GND pixel_9979/VREF pixel_9979/ROW_SEL
+ pixel_9979/NB1 pixel_9979/VBIAS pixel_9979/NB2 pixel_9979/AMP_IN pixel_9979/SF_IB
+ pixel_9979/PIX_OUT pixel_9979/CSA_VREF pixel
Xpixel_4220 pixel_4220/gring pixel_4220/VDD pixel_4220/GND pixel_4220/VREF pixel_4220/ROW_SEL
+ pixel_4220/NB1 pixel_4220/VBIAS pixel_4220/NB2 pixel_4220/AMP_IN pixel_4220/SF_IB
+ pixel_4220/PIX_OUT pixel_4220/CSA_VREF pixel
Xpixel_4231 pixel_4231/gring pixel_4231/VDD pixel_4231/GND pixel_4231/VREF pixel_4231/ROW_SEL
+ pixel_4231/NB1 pixel_4231/VBIAS pixel_4231/NB2 pixel_4231/AMP_IN pixel_4231/SF_IB
+ pixel_4231/PIX_OUT pixel_4231/CSA_VREF pixel
Xpixel_4242 pixel_4242/gring pixel_4242/VDD pixel_4242/GND pixel_4242/VREF pixel_4242/ROW_SEL
+ pixel_4242/NB1 pixel_4242/VBIAS pixel_4242/NB2 pixel_4242/AMP_IN pixel_4242/SF_IB
+ pixel_4242/PIX_OUT pixel_4242/CSA_VREF pixel
Xpixel_4253 pixel_4253/gring pixel_4253/VDD pixel_4253/GND pixel_4253/VREF pixel_4253/ROW_SEL
+ pixel_4253/NB1 pixel_4253/VBIAS pixel_4253/NB2 pixel_4253/AMP_IN pixel_4253/SF_IB
+ pixel_4253/PIX_OUT pixel_4253/CSA_VREF pixel
Xpixel_292 pixel_292/gring pixel_292/VDD pixel_292/GND pixel_292/VREF pixel_292/ROW_SEL
+ pixel_292/NB1 pixel_292/VBIAS pixel_292/NB2 pixel_292/AMP_IN pixel_292/SF_IB pixel_292/PIX_OUT
+ pixel_292/CSA_VREF pixel
Xpixel_281 pixel_281/gring pixel_281/VDD pixel_281/GND pixel_281/VREF pixel_281/ROW_SEL
+ pixel_281/NB1 pixel_281/VBIAS pixel_281/NB2 pixel_281/AMP_IN pixel_281/SF_IB pixel_281/PIX_OUT
+ pixel_281/CSA_VREF pixel
Xpixel_270 pixel_270/gring pixel_270/VDD pixel_270/GND pixel_270/VREF pixel_270/ROW_SEL
+ pixel_270/NB1 pixel_270/VBIAS pixel_270/NB2 pixel_270/AMP_IN pixel_270/SF_IB pixel_270/PIX_OUT
+ pixel_270/CSA_VREF pixel
Xpixel_3552 pixel_3552/gring pixel_3552/VDD pixel_3552/GND pixel_3552/VREF pixel_3552/ROW_SEL
+ pixel_3552/NB1 pixel_3552/VBIAS pixel_3552/NB2 pixel_3552/AMP_IN pixel_3552/SF_IB
+ pixel_3552/PIX_OUT pixel_3552/CSA_VREF pixel
Xpixel_3541 pixel_3541/gring pixel_3541/VDD pixel_3541/GND pixel_3541/VREF pixel_3541/ROW_SEL
+ pixel_3541/NB1 pixel_3541/VBIAS pixel_3541/NB2 pixel_3541/AMP_IN pixel_3541/SF_IB
+ pixel_3541/PIX_OUT pixel_3541/CSA_VREF pixel
Xpixel_3530 pixel_3530/gring pixel_3530/VDD pixel_3530/GND pixel_3530/VREF pixel_3530/ROW_SEL
+ pixel_3530/NB1 pixel_3530/VBIAS pixel_3530/NB2 pixel_3530/AMP_IN pixel_3530/SF_IB
+ pixel_3530/PIX_OUT pixel_3530/CSA_VREF pixel
Xpixel_4264 pixel_4264/gring pixel_4264/VDD pixel_4264/GND pixel_4264/VREF pixel_4264/ROW_SEL
+ pixel_4264/NB1 pixel_4264/VBIAS pixel_4264/NB2 pixel_4264/AMP_IN pixel_4264/SF_IB
+ pixel_4264/PIX_OUT pixel_4264/CSA_VREF pixel
Xpixel_4275 pixel_4275/gring pixel_4275/VDD pixel_4275/GND pixel_4275/VREF pixel_4275/ROW_SEL
+ pixel_4275/NB1 pixel_4275/VBIAS pixel_4275/NB2 pixel_4275/AMP_IN pixel_4275/SF_IB
+ pixel_4275/PIX_OUT pixel_4275/CSA_VREF pixel
Xpixel_4286 pixel_4286/gring pixel_4286/VDD pixel_4286/GND pixel_4286/VREF pixel_4286/ROW_SEL
+ pixel_4286/NB1 pixel_4286/VBIAS pixel_4286/NB2 pixel_4286/AMP_IN pixel_4286/SF_IB
+ pixel_4286/PIX_OUT pixel_4286/CSA_VREF pixel
Xpixel_2840 pixel_2840/gring pixel_2840/VDD pixel_2840/GND pixel_2840/VREF pixel_2840/ROW_SEL
+ pixel_2840/NB1 pixel_2840/VBIAS pixel_2840/NB2 pixel_2840/AMP_IN pixel_2840/SF_IB
+ pixel_2840/PIX_OUT pixel_2840/CSA_VREF pixel
Xpixel_3585 pixel_3585/gring pixel_3585/VDD pixel_3585/GND pixel_3585/VREF pixel_3585/ROW_SEL
+ pixel_3585/NB1 pixel_3585/VBIAS pixel_3585/NB2 pixel_3585/AMP_IN pixel_3585/SF_IB
+ pixel_3585/PIX_OUT pixel_3585/CSA_VREF pixel
Xpixel_3574 pixel_3574/gring pixel_3574/VDD pixel_3574/GND pixel_3574/VREF pixel_3574/ROW_SEL
+ pixel_3574/NB1 pixel_3574/VBIAS pixel_3574/NB2 pixel_3574/AMP_IN pixel_3574/SF_IB
+ pixel_3574/PIX_OUT pixel_3574/CSA_VREF pixel
Xpixel_3563 pixel_3563/gring pixel_3563/VDD pixel_3563/GND pixel_3563/VREF pixel_3563/ROW_SEL
+ pixel_3563/NB1 pixel_3563/VBIAS pixel_3563/NB2 pixel_3563/AMP_IN pixel_3563/SF_IB
+ pixel_3563/PIX_OUT pixel_3563/CSA_VREF pixel
Xpixel_4297 pixel_4297/gring pixel_4297/VDD pixel_4297/GND pixel_4297/VREF pixel_4297/ROW_SEL
+ pixel_4297/NB1 pixel_4297/VBIAS pixel_4297/NB2 pixel_4297/AMP_IN pixel_4297/SF_IB
+ pixel_4297/PIX_OUT pixel_4297/CSA_VREF pixel
Xpixel_2873 pixel_2873/gring pixel_2873/VDD pixel_2873/GND pixel_2873/VREF pixel_2873/ROW_SEL
+ pixel_2873/NB1 pixel_2873/VBIAS pixel_2873/NB2 pixel_2873/AMP_IN pixel_2873/SF_IB
+ pixel_2873/PIX_OUT pixel_2873/CSA_VREF pixel
Xpixel_2862 pixel_2862/gring pixel_2862/VDD pixel_2862/GND pixel_2862/VREF pixel_2862/ROW_SEL
+ pixel_2862/NB1 pixel_2862/VBIAS pixel_2862/NB2 pixel_2862/AMP_IN pixel_2862/SF_IB
+ pixel_2862/PIX_OUT pixel_2862/CSA_VREF pixel
Xpixel_2851 pixel_2851/gring pixel_2851/VDD pixel_2851/GND pixel_2851/VREF pixel_2851/ROW_SEL
+ pixel_2851/NB1 pixel_2851/VBIAS pixel_2851/NB2 pixel_2851/AMP_IN pixel_2851/SF_IB
+ pixel_2851/PIX_OUT pixel_2851/CSA_VREF pixel
Xpixel_3596 pixel_3596/gring pixel_3596/VDD pixel_3596/GND pixel_3596/VREF pixel_3596/ROW_SEL
+ pixel_3596/NB1 pixel_3596/VBIAS pixel_3596/NB2 pixel_3596/AMP_IN pixel_3596/SF_IB
+ pixel_3596/PIX_OUT pixel_3596/CSA_VREF pixel
Xpixel_2895 pixel_2895/gring pixel_2895/VDD pixel_2895/GND pixel_2895/VREF pixel_2895/ROW_SEL
+ pixel_2895/NB1 pixel_2895/VBIAS pixel_2895/NB2 pixel_2895/AMP_IN pixel_2895/SF_IB
+ pixel_2895/PIX_OUT pixel_2895/CSA_VREF pixel
Xpixel_2884 pixel_2884/gring pixel_2884/VDD pixel_2884/GND pixel_2884/VREF pixel_2884/ROW_SEL
+ pixel_2884/NB1 pixel_2884/VBIAS pixel_2884/NB2 pixel_2884/AMP_IN pixel_2884/SF_IB
+ pixel_2884/PIX_OUT pixel_2884/CSA_VREF pixel
Xpixel_9209 pixel_9209/gring pixel_9209/VDD pixel_9209/GND pixel_9209/VREF pixel_9209/ROW_SEL
+ pixel_9209/NB1 pixel_9209/VBIAS pixel_9209/NB2 pixel_9209/AMP_IN pixel_9209/SF_IB
+ pixel_9209/PIX_OUT pixel_9209/CSA_VREF pixel
Xpixel_8508 pixel_8508/gring pixel_8508/VDD pixel_8508/GND pixel_8508/VREF pixel_8508/ROW_SEL
+ pixel_8508/NB1 pixel_8508/VBIAS pixel_8508/NB2 pixel_8508/AMP_IN pixel_8508/SF_IB
+ pixel_8508/PIX_OUT pixel_8508/CSA_VREF pixel
Xpixel_8519 pixel_8519/gring pixel_8519/VDD pixel_8519/GND pixel_8519/VREF pixel_8519/ROW_SEL
+ pixel_8519/NB1 pixel_8519/VBIAS pixel_8519/NB2 pixel_8519/AMP_IN pixel_8519/SF_IB
+ pixel_8519/PIX_OUT pixel_8519/CSA_VREF pixel
Xpixel_7807 pixel_7807/gring pixel_7807/VDD pixel_7807/GND pixel_7807/VREF pixel_7807/ROW_SEL
+ pixel_7807/NB1 pixel_7807/VBIAS pixel_7807/NB2 pixel_7807/AMP_IN pixel_7807/SF_IB
+ pixel_7807/PIX_OUT pixel_7807/CSA_VREF pixel
Xpixel_7818 pixel_7818/gring pixel_7818/VDD pixel_7818/GND pixel_7818/VREF pixel_7818/ROW_SEL
+ pixel_7818/NB1 pixel_7818/VBIAS pixel_7818/NB2 pixel_7818/AMP_IN pixel_7818/SF_IB
+ pixel_7818/PIX_OUT pixel_7818/CSA_VREF pixel
Xpixel_7829 pixel_7829/gring pixel_7829/VDD pixel_7829/GND pixel_7829/VREF pixel_7829/ROW_SEL
+ pixel_7829/NB1 pixel_7829/VBIAS pixel_7829/NB2 pixel_7829/AMP_IN pixel_7829/SF_IB
+ pixel_7829/PIX_OUT pixel_7829/CSA_VREF pixel
Xpixel_2136 pixel_2136/gring pixel_2136/VDD pixel_2136/GND pixel_2136/VREF pixel_2136/ROW_SEL
+ pixel_2136/NB1 pixel_2136/VBIAS pixel_2136/NB2 pixel_2136/AMP_IN pixel_2136/SF_IB
+ pixel_2136/PIX_OUT pixel_2136/CSA_VREF pixel
Xpixel_2125 pixel_2125/gring pixel_2125/VDD pixel_2125/GND pixel_2125/VREF pixel_2125/ROW_SEL
+ pixel_2125/NB1 pixel_2125/VBIAS pixel_2125/NB2 pixel_2125/AMP_IN pixel_2125/SF_IB
+ pixel_2125/PIX_OUT pixel_2125/CSA_VREF pixel
Xpixel_2114 pixel_2114/gring pixel_2114/VDD pixel_2114/GND pixel_2114/VREF pixel_2114/ROW_SEL
+ pixel_2114/NB1 pixel_2114/VBIAS pixel_2114/NB2 pixel_2114/AMP_IN pixel_2114/SF_IB
+ pixel_2114/PIX_OUT pixel_2114/CSA_VREF pixel
Xpixel_2103 pixel_2103/gring pixel_2103/VDD pixel_2103/GND pixel_2103/VREF pixel_2103/ROW_SEL
+ pixel_2103/NB1 pixel_2103/VBIAS pixel_2103/NB2 pixel_2103/AMP_IN pixel_2103/SF_IB
+ pixel_2103/PIX_OUT pixel_2103/CSA_VREF pixel
Xpixel_1424 pixel_1424/gring pixel_1424/VDD pixel_1424/GND pixel_1424/VREF pixel_1424/ROW_SEL
+ pixel_1424/NB1 pixel_1424/VBIAS pixel_1424/NB2 pixel_1424/AMP_IN pixel_1424/SF_IB
+ pixel_1424/PIX_OUT pixel_1424/CSA_VREF pixel
Xpixel_1413 pixel_1413/gring pixel_1413/VDD pixel_1413/GND pixel_1413/VREF pixel_1413/ROW_SEL
+ pixel_1413/NB1 pixel_1413/VBIAS pixel_1413/NB2 pixel_1413/AMP_IN pixel_1413/SF_IB
+ pixel_1413/PIX_OUT pixel_1413/CSA_VREF pixel
Xpixel_1402 pixel_1402/gring pixel_1402/VDD pixel_1402/GND pixel_1402/VREF pixel_1402/ROW_SEL
+ pixel_1402/NB1 pixel_1402/VBIAS pixel_1402/NB2 pixel_1402/AMP_IN pixel_1402/SF_IB
+ pixel_1402/PIX_OUT pixel_1402/CSA_VREF pixel
Xpixel_2169 pixel_2169/gring pixel_2169/VDD pixel_2169/GND pixel_2169/VREF pixel_2169/ROW_SEL
+ pixel_2169/NB1 pixel_2169/VBIAS pixel_2169/NB2 pixel_2169/AMP_IN pixel_2169/SF_IB
+ pixel_2169/PIX_OUT pixel_2169/CSA_VREF pixel
Xpixel_2158 pixel_2158/gring pixel_2158/VDD pixel_2158/GND pixel_2158/VREF pixel_2158/ROW_SEL
+ pixel_2158/NB1 pixel_2158/VBIAS pixel_2158/NB2 pixel_2158/AMP_IN pixel_2158/SF_IB
+ pixel_2158/PIX_OUT pixel_2158/CSA_VREF pixel
Xpixel_2147 pixel_2147/gring pixel_2147/VDD pixel_2147/GND pixel_2147/VREF pixel_2147/ROW_SEL
+ pixel_2147/NB1 pixel_2147/VBIAS pixel_2147/NB2 pixel_2147/AMP_IN pixel_2147/SF_IB
+ pixel_2147/PIX_OUT pixel_2147/CSA_VREF pixel
Xpixel_1457 pixel_1457/gring pixel_1457/VDD pixel_1457/GND pixel_1457/VREF pixel_1457/ROW_SEL
+ pixel_1457/NB1 pixel_1457/VBIAS pixel_1457/NB2 pixel_1457/AMP_IN pixel_1457/SF_IB
+ pixel_1457/PIX_OUT pixel_1457/CSA_VREF pixel
Xpixel_1446 pixel_1446/gring pixel_1446/VDD pixel_1446/GND pixel_1446/VREF pixel_1446/ROW_SEL
+ pixel_1446/NB1 pixel_1446/VBIAS pixel_1446/NB2 pixel_1446/AMP_IN pixel_1446/SF_IB
+ pixel_1446/PIX_OUT pixel_1446/CSA_VREF pixel
Xpixel_1435 pixel_1435/gring pixel_1435/VDD pixel_1435/GND pixel_1435/VREF pixel_1435/ROW_SEL
+ pixel_1435/NB1 pixel_1435/VBIAS pixel_1435/NB2 pixel_1435/AMP_IN pixel_1435/SF_IB
+ pixel_1435/PIX_OUT pixel_1435/CSA_VREF pixel
Xpixel_1479 pixel_1479/gring pixel_1479/VDD pixel_1479/GND pixel_1479/VREF pixel_1479/ROW_SEL
+ pixel_1479/NB1 pixel_1479/VBIAS pixel_1479/NB2 pixel_1479/AMP_IN pixel_1479/SF_IB
+ pixel_1479/PIX_OUT pixel_1479/CSA_VREF pixel
Xpixel_1468 pixel_1468/gring pixel_1468/VDD pixel_1468/GND pixel_1468/VREF pixel_1468/ROW_SEL
+ pixel_1468/NB1 pixel_1468/VBIAS pixel_1468/NB2 pixel_1468/AMP_IN pixel_1468/SF_IB
+ pixel_1468/PIX_OUT pixel_1468/CSA_VREF pixel
Xpixel_9710 pixel_9710/gring pixel_9710/VDD pixel_9710/GND pixel_9710/VREF pixel_9710/ROW_SEL
+ pixel_9710/NB1 pixel_9710/VBIAS pixel_9710/NB2 pixel_9710/AMP_IN pixel_9710/SF_IB
+ pixel_9710/PIX_OUT pixel_9710/CSA_VREF pixel
Xpixel_9721 pixel_9721/gring pixel_9721/VDD pixel_9721/GND pixel_9721/VREF pixel_9721/ROW_SEL
+ pixel_9721/NB1 pixel_9721/VBIAS pixel_9721/NB2 pixel_9721/AMP_IN pixel_9721/SF_IB
+ pixel_9721/PIX_OUT pixel_9721/CSA_VREF pixel
Xpixel_9732 pixel_9732/gring pixel_9732/VDD pixel_9732/GND pixel_9732/VREF pixel_9732/ROW_SEL
+ pixel_9732/NB1 pixel_9732/VBIAS pixel_9732/NB2 pixel_9732/AMP_IN pixel_9732/SF_IB
+ pixel_9732/PIX_OUT pixel_9732/CSA_VREF pixel
Xpixel_9743 pixel_9743/gring pixel_9743/VDD pixel_9743/GND pixel_9743/VREF pixel_9743/ROW_SEL
+ pixel_9743/NB1 pixel_9743/VBIAS pixel_9743/NB2 pixel_9743/AMP_IN pixel_9743/SF_IB
+ pixel_9743/PIX_OUT pixel_9743/CSA_VREF pixel
Xpixel_9754 pixel_9754/gring pixel_9754/VDD pixel_9754/GND pixel_9754/VREF pixel_9754/ROW_SEL
+ pixel_9754/NB1 pixel_9754/VBIAS pixel_9754/NB2 pixel_9754/AMP_IN pixel_9754/SF_IB
+ pixel_9754/PIX_OUT pixel_9754/CSA_VREF pixel
Xpixel_9765 pixel_9765/gring pixel_9765/VDD pixel_9765/GND pixel_9765/VREF pixel_9765/ROW_SEL
+ pixel_9765/NB1 pixel_9765/VBIAS pixel_9765/NB2 pixel_9765/AMP_IN pixel_9765/SF_IB
+ pixel_9765/PIX_OUT pixel_9765/CSA_VREF pixel
Xpixel_9776 pixel_9776/gring pixel_9776/VDD pixel_9776/GND pixel_9776/VREF pixel_9776/ROW_SEL
+ pixel_9776/NB1 pixel_9776/VBIAS pixel_9776/NB2 pixel_9776/AMP_IN pixel_9776/SF_IB
+ pixel_9776/PIX_OUT pixel_9776/CSA_VREF pixel
Xpixel_9787 pixel_9787/gring pixel_9787/VDD pixel_9787/GND pixel_9787/VREF pixel_9787/ROW_SEL
+ pixel_9787/NB1 pixel_9787/VBIAS pixel_9787/NB2 pixel_9787/AMP_IN pixel_9787/SF_IB
+ pixel_9787/PIX_OUT pixel_9787/CSA_VREF pixel
Xpixel_9798 pixel_9798/gring pixel_9798/VDD pixel_9798/GND pixel_9798/VREF pixel_9798/ROW_SEL
+ pixel_9798/NB1 pixel_9798/VBIAS pixel_9798/NB2 pixel_9798/AMP_IN pixel_9798/SF_IB
+ pixel_9798/PIX_OUT pixel_9798/CSA_VREF pixel
Xpixel_4050 pixel_4050/gring pixel_4050/VDD pixel_4050/GND pixel_4050/VREF pixel_4050/ROW_SEL
+ pixel_4050/NB1 pixel_4050/VBIAS pixel_4050/NB2 pixel_4050/AMP_IN pixel_4050/SF_IB
+ pixel_4050/PIX_OUT pixel_4050/CSA_VREF pixel
Xpixel_4061 pixel_4061/gring pixel_4061/VDD pixel_4061/GND pixel_4061/VREF pixel_4061/ROW_SEL
+ pixel_4061/NB1 pixel_4061/VBIAS pixel_4061/NB2 pixel_4061/AMP_IN pixel_4061/SF_IB
+ pixel_4061/PIX_OUT pixel_4061/CSA_VREF pixel
Xpixel_3360 pixel_3360/gring pixel_3360/VDD pixel_3360/GND pixel_3360/VREF pixel_3360/ROW_SEL
+ pixel_3360/NB1 pixel_3360/VBIAS pixel_3360/NB2 pixel_3360/AMP_IN pixel_3360/SF_IB
+ pixel_3360/PIX_OUT pixel_3360/CSA_VREF pixel
Xpixel_4072 pixel_4072/gring pixel_4072/VDD pixel_4072/GND pixel_4072/VREF pixel_4072/ROW_SEL
+ pixel_4072/NB1 pixel_4072/VBIAS pixel_4072/NB2 pixel_4072/AMP_IN pixel_4072/SF_IB
+ pixel_4072/PIX_OUT pixel_4072/CSA_VREF pixel
Xpixel_4083 pixel_4083/gring pixel_4083/VDD pixel_4083/GND pixel_4083/VREF pixel_4083/ROW_SEL
+ pixel_4083/NB1 pixel_4083/VBIAS pixel_4083/NB2 pixel_4083/AMP_IN pixel_4083/SF_IB
+ pixel_4083/PIX_OUT pixel_4083/CSA_VREF pixel
Xpixel_4094 pixel_4094/gring pixel_4094/VDD pixel_4094/GND pixel_4094/VREF pixel_4094/ROW_SEL
+ pixel_4094/NB1 pixel_4094/VBIAS pixel_4094/NB2 pixel_4094/AMP_IN pixel_4094/SF_IB
+ pixel_4094/PIX_OUT pixel_4094/CSA_VREF pixel
Xpixel_3393 pixel_3393/gring pixel_3393/VDD pixel_3393/GND pixel_3393/VREF pixel_3393/ROW_SEL
+ pixel_3393/NB1 pixel_3393/VBIAS pixel_3393/NB2 pixel_3393/AMP_IN pixel_3393/SF_IB
+ pixel_3393/PIX_OUT pixel_3393/CSA_VREF pixel
Xpixel_3382 pixel_3382/gring pixel_3382/VDD pixel_3382/GND pixel_3382/VREF pixel_3382/ROW_SEL
+ pixel_3382/NB1 pixel_3382/VBIAS pixel_3382/NB2 pixel_3382/AMP_IN pixel_3382/SF_IB
+ pixel_3382/PIX_OUT pixel_3382/CSA_VREF pixel
Xpixel_3371 pixel_3371/gring pixel_3371/VDD pixel_3371/GND pixel_3371/VREF pixel_3371/ROW_SEL
+ pixel_3371/NB1 pixel_3371/VBIAS pixel_3371/NB2 pixel_3371/AMP_IN pixel_3371/SF_IB
+ pixel_3371/PIX_OUT pixel_3371/CSA_VREF pixel
Xpixel_2692 pixel_2692/gring pixel_2692/VDD pixel_2692/GND pixel_2692/VREF pixel_2692/ROW_SEL
+ pixel_2692/NB1 pixel_2692/VBIAS pixel_2692/NB2 pixel_2692/AMP_IN pixel_2692/SF_IB
+ pixel_2692/PIX_OUT pixel_2692/CSA_VREF pixel
Xpixel_2681 pixel_2681/gring pixel_2681/VDD pixel_2681/GND pixel_2681/VREF pixel_2681/ROW_SEL
+ pixel_2681/NB1 pixel_2681/VBIAS pixel_2681/NB2 pixel_2681/AMP_IN pixel_2681/SF_IB
+ pixel_2681/PIX_OUT pixel_2681/CSA_VREF pixel
Xpixel_2670 pixel_2670/gring pixel_2670/VDD pixel_2670/GND pixel_2670/VREF pixel_2670/ROW_SEL
+ pixel_2670/NB1 pixel_2670/VBIAS pixel_2670/NB2 pixel_2670/AMP_IN pixel_2670/SF_IB
+ pixel_2670/PIX_OUT pixel_2670/CSA_VREF pixel
Xpixel_1980 pixel_1980/gring pixel_1980/VDD pixel_1980/GND pixel_1980/VREF pixel_1980/ROW_SEL
+ pixel_1980/NB1 pixel_1980/VBIAS pixel_1980/NB2 pixel_1980/AMP_IN pixel_1980/SF_IB
+ pixel_1980/PIX_OUT pixel_1980/CSA_VREF pixel
Xpixel_1991 pixel_1991/gring pixel_1991/VDD pixel_1991/GND pixel_1991/VREF pixel_1991/ROW_SEL
+ pixel_1991/NB1 pixel_1991/VBIAS pixel_1991/NB2 pixel_1991/AMP_IN pixel_1991/SF_IB
+ pixel_1991/PIX_OUT pixel_1991/CSA_VREF pixel
Xpixel_9028 pixel_9028/gring pixel_9028/VDD pixel_9028/GND pixel_9028/VREF pixel_9028/ROW_SEL
+ pixel_9028/NB1 pixel_9028/VBIAS pixel_9028/NB2 pixel_9028/AMP_IN pixel_9028/SF_IB
+ pixel_9028/PIX_OUT pixel_9028/CSA_VREF pixel
Xpixel_9017 pixel_9017/gring pixel_9017/VDD pixel_9017/GND pixel_9017/VREF pixel_9017/ROW_SEL
+ pixel_9017/NB1 pixel_9017/VBIAS pixel_9017/NB2 pixel_9017/AMP_IN pixel_9017/SF_IB
+ pixel_9017/PIX_OUT pixel_9017/CSA_VREF pixel
Xpixel_9006 pixel_9006/gring pixel_9006/VDD pixel_9006/GND pixel_9006/VREF pixel_9006/ROW_SEL
+ pixel_9006/NB1 pixel_9006/VBIAS pixel_9006/NB2 pixel_9006/AMP_IN pixel_9006/SF_IB
+ pixel_9006/PIX_OUT pixel_9006/CSA_VREF pixel
Xpixel_9039 pixel_9039/gring pixel_9039/VDD pixel_9039/GND pixel_9039/VREF pixel_9039/ROW_SEL
+ pixel_9039/NB1 pixel_9039/VBIAS pixel_9039/NB2 pixel_9039/AMP_IN pixel_9039/SF_IB
+ pixel_9039/PIX_OUT pixel_9039/CSA_VREF pixel
Xpixel_8305 pixel_8305/gring pixel_8305/VDD pixel_8305/GND pixel_8305/VREF pixel_8305/ROW_SEL
+ pixel_8305/NB1 pixel_8305/VBIAS pixel_8305/NB2 pixel_8305/AMP_IN pixel_8305/SF_IB
+ pixel_8305/PIX_OUT pixel_8305/CSA_VREF pixel
Xpixel_8316 pixel_8316/gring pixel_8316/VDD pixel_8316/GND pixel_8316/VREF pixel_8316/ROW_SEL
+ pixel_8316/NB1 pixel_8316/VBIAS pixel_8316/NB2 pixel_8316/AMP_IN pixel_8316/SF_IB
+ pixel_8316/PIX_OUT pixel_8316/CSA_VREF pixel
Xpixel_8327 pixel_8327/gring pixel_8327/VDD pixel_8327/GND pixel_8327/VREF pixel_8327/ROW_SEL
+ pixel_8327/NB1 pixel_8327/VBIAS pixel_8327/NB2 pixel_8327/AMP_IN pixel_8327/SF_IB
+ pixel_8327/PIX_OUT pixel_8327/CSA_VREF pixel
Xpixel_8338 pixel_8338/gring pixel_8338/VDD pixel_8338/GND pixel_8338/VREF pixel_8338/ROW_SEL
+ pixel_8338/NB1 pixel_8338/VBIAS pixel_8338/NB2 pixel_8338/AMP_IN pixel_8338/SF_IB
+ pixel_8338/PIX_OUT pixel_8338/CSA_VREF pixel
Xpixel_8349 pixel_8349/gring pixel_8349/VDD pixel_8349/GND pixel_8349/VREF pixel_8349/ROW_SEL
+ pixel_8349/NB1 pixel_8349/VBIAS pixel_8349/NB2 pixel_8349/AMP_IN pixel_8349/SF_IB
+ pixel_8349/PIX_OUT pixel_8349/CSA_VREF pixel
Xpixel_7604 pixel_7604/gring pixel_7604/VDD pixel_7604/GND pixel_7604/VREF pixel_7604/ROW_SEL
+ pixel_7604/NB1 pixel_7604/VBIAS pixel_7604/NB2 pixel_7604/AMP_IN pixel_7604/SF_IB
+ pixel_7604/PIX_OUT pixel_7604/CSA_VREF pixel
Xpixel_7615 pixel_7615/gring pixel_7615/VDD pixel_7615/GND pixel_7615/VREF pixel_7615/ROW_SEL
+ pixel_7615/NB1 pixel_7615/VBIAS pixel_7615/NB2 pixel_7615/AMP_IN pixel_7615/SF_IB
+ pixel_7615/PIX_OUT pixel_7615/CSA_VREF pixel
Xpixel_7626 pixel_7626/gring pixel_7626/VDD pixel_7626/GND pixel_7626/VREF pixel_7626/ROW_SEL
+ pixel_7626/NB1 pixel_7626/VBIAS pixel_7626/NB2 pixel_7626/AMP_IN pixel_7626/SF_IB
+ pixel_7626/PIX_OUT pixel_7626/CSA_VREF pixel
Xpixel_7637 pixel_7637/gring pixel_7637/VDD pixel_7637/GND pixel_7637/VREF pixel_7637/ROW_SEL
+ pixel_7637/NB1 pixel_7637/VBIAS pixel_7637/NB2 pixel_7637/AMP_IN pixel_7637/SF_IB
+ pixel_7637/PIX_OUT pixel_7637/CSA_VREF pixel
Xpixel_7648 pixel_7648/gring pixel_7648/VDD pixel_7648/GND pixel_7648/VREF pixel_7648/ROW_SEL
+ pixel_7648/NB1 pixel_7648/VBIAS pixel_7648/NB2 pixel_7648/AMP_IN pixel_7648/SF_IB
+ pixel_7648/PIX_OUT pixel_7648/CSA_VREF pixel
Xpixel_6903 pixel_6903/gring pixel_6903/VDD pixel_6903/GND pixel_6903/VREF pixel_6903/ROW_SEL
+ pixel_6903/NB1 pixel_6903/VBIAS pixel_6903/NB2 pixel_6903/AMP_IN pixel_6903/SF_IB
+ pixel_6903/PIX_OUT pixel_6903/CSA_VREF pixel
Xpixel_7659 pixel_7659/gring pixel_7659/VDD pixel_7659/GND pixel_7659/VREF pixel_7659/ROW_SEL
+ pixel_7659/NB1 pixel_7659/VBIAS pixel_7659/NB2 pixel_7659/AMP_IN pixel_7659/SF_IB
+ pixel_7659/PIX_OUT pixel_7659/CSA_VREF pixel
Xpixel_6914 pixel_6914/gring pixel_6914/VDD pixel_6914/GND pixel_6914/VREF pixel_6914/ROW_SEL
+ pixel_6914/NB1 pixel_6914/VBIAS pixel_6914/NB2 pixel_6914/AMP_IN pixel_6914/SF_IB
+ pixel_6914/PIX_OUT pixel_6914/CSA_VREF pixel
Xpixel_6925 pixel_6925/gring pixel_6925/VDD pixel_6925/GND pixel_6925/VREF pixel_6925/ROW_SEL
+ pixel_6925/NB1 pixel_6925/VBIAS pixel_6925/NB2 pixel_6925/AMP_IN pixel_6925/SF_IB
+ pixel_6925/PIX_OUT pixel_6925/CSA_VREF pixel
Xpixel_6936 pixel_6936/gring pixel_6936/VDD pixel_6936/GND pixel_6936/VREF pixel_6936/ROW_SEL
+ pixel_6936/NB1 pixel_6936/VBIAS pixel_6936/NB2 pixel_6936/AMP_IN pixel_6936/SF_IB
+ pixel_6936/PIX_OUT pixel_6936/CSA_VREF pixel
Xpixel_28 pixel_28/gring pixel_28/VDD pixel_28/GND pixel_28/VREF pixel_28/ROW_SEL
+ pixel_28/NB1 pixel_28/VBIAS pixel_28/NB2 pixel_28/AMP_IN pixel_28/SF_IB pixel_28/PIX_OUT
+ pixel_28/CSA_VREF pixel
Xpixel_17 pixel_17/gring pixel_17/VDD pixel_17/GND pixel_17/VREF pixel_17/ROW_SEL
+ pixel_17/NB1 pixel_17/VBIAS pixel_17/NB2 pixel_17/AMP_IN pixel_17/SF_IB pixel_17/PIX_OUT
+ pixel_17/CSA_VREF pixel
Xpixel_6947 pixel_6947/gring pixel_6947/VDD pixel_6947/GND pixel_6947/VREF pixel_6947/ROW_SEL
+ pixel_6947/NB1 pixel_6947/VBIAS pixel_6947/NB2 pixel_6947/AMP_IN pixel_6947/SF_IB
+ pixel_6947/PIX_OUT pixel_6947/CSA_VREF pixel
Xpixel_6958 pixel_6958/gring pixel_6958/VDD pixel_6958/GND pixel_6958/VREF pixel_6958/ROW_SEL
+ pixel_6958/NB1 pixel_6958/VBIAS pixel_6958/NB2 pixel_6958/AMP_IN pixel_6958/SF_IB
+ pixel_6958/PIX_OUT pixel_6958/CSA_VREF pixel
Xpixel_6969 pixel_6969/gring pixel_6969/VDD pixel_6969/GND pixel_6969/VREF pixel_6969/ROW_SEL
+ pixel_6969/NB1 pixel_6969/VBIAS pixel_6969/NB2 pixel_6969/AMP_IN pixel_6969/SF_IB
+ pixel_6969/PIX_OUT pixel_6969/CSA_VREF pixel
Xpixel_39 pixel_39/gring pixel_39/VDD pixel_39/GND pixel_39/VREF pixel_39/ROW_SEL
+ pixel_39/NB1 pixel_39/VBIAS pixel_39/NB2 pixel_39/AMP_IN pixel_39/SF_IB pixel_39/PIX_OUT
+ pixel_39/CSA_VREF pixel
Xpixel_1232 pixel_1232/gring pixel_1232/VDD pixel_1232/GND pixel_1232/VREF pixel_1232/ROW_SEL
+ pixel_1232/NB1 pixel_1232/VBIAS pixel_1232/NB2 pixel_1232/AMP_IN pixel_1232/SF_IB
+ pixel_1232/PIX_OUT pixel_1232/CSA_VREF pixel
Xpixel_1221 pixel_1221/gring pixel_1221/VDD pixel_1221/GND pixel_1221/VREF pixel_1221/ROW_SEL
+ pixel_1221/NB1 pixel_1221/VBIAS pixel_1221/NB2 pixel_1221/AMP_IN pixel_1221/SF_IB
+ pixel_1221/PIX_OUT pixel_1221/CSA_VREF pixel
Xpixel_1210 pixel_1210/gring pixel_1210/VDD pixel_1210/GND pixel_1210/VREF pixel_1210/ROW_SEL
+ pixel_1210/NB1 pixel_1210/VBIAS pixel_1210/NB2 pixel_1210/AMP_IN pixel_1210/SF_IB
+ pixel_1210/PIX_OUT pixel_1210/CSA_VREF pixel
Xpixel_1276 pixel_1276/gring pixel_1276/VDD pixel_1276/GND pixel_1276/VREF pixel_1276/ROW_SEL
+ pixel_1276/NB1 pixel_1276/VBIAS pixel_1276/NB2 pixel_1276/AMP_IN pixel_1276/SF_IB
+ pixel_1276/PIX_OUT pixel_1276/CSA_VREF pixel
Xpixel_1265 pixel_1265/gring pixel_1265/VDD pixel_1265/GND pixel_1265/VREF pixel_1265/ROW_SEL
+ pixel_1265/NB1 pixel_1265/VBIAS pixel_1265/NB2 pixel_1265/AMP_IN pixel_1265/SF_IB
+ pixel_1265/PIX_OUT pixel_1265/CSA_VREF pixel
Xpixel_1254 pixel_1254/gring pixel_1254/VDD pixel_1254/GND pixel_1254/VREF pixel_1254/ROW_SEL
+ pixel_1254/NB1 pixel_1254/VBIAS pixel_1254/NB2 pixel_1254/AMP_IN pixel_1254/SF_IB
+ pixel_1254/PIX_OUT pixel_1254/CSA_VREF pixel
Xpixel_1243 pixel_1243/gring pixel_1243/VDD pixel_1243/GND pixel_1243/VREF pixel_1243/ROW_SEL
+ pixel_1243/NB1 pixel_1243/VBIAS pixel_1243/NB2 pixel_1243/AMP_IN pixel_1243/SF_IB
+ pixel_1243/PIX_OUT pixel_1243/CSA_VREF pixel
Xpixel_1298 pixel_1298/gring pixel_1298/VDD pixel_1298/GND pixel_1298/VREF pixel_1298/ROW_SEL
+ pixel_1298/NB1 pixel_1298/VBIAS pixel_1298/NB2 pixel_1298/AMP_IN pixel_1298/SF_IB
+ pixel_1298/PIX_OUT pixel_1298/CSA_VREF pixel
Xpixel_1287 pixel_1287/gring pixel_1287/VDD pixel_1287/GND pixel_1287/VREF pixel_1287/ROW_SEL
+ pixel_1287/NB1 pixel_1287/VBIAS pixel_1287/NB2 pixel_1287/AMP_IN pixel_1287/SF_IB
+ pixel_1287/PIX_OUT pixel_1287/CSA_VREF pixel
Xpixel_9540 pixel_9540/gring pixel_9540/VDD pixel_9540/GND pixel_9540/VREF pixel_9540/ROW_SEL
+ pixel_9540/NB1 pixel_9540/VBIAS pixel_9540/NB2 pixel_9540/AMP_IN pixel_9540/SF_IB
+ pixel_9540/PIX_OUT pixel_9540/CSA_VREF pixel
Xpixel_9584 pixel_9584/gring pixel_9584/VDD pixel_9584/GND pixel_9584/VREF pixel_9584/ROW_SEL
+ pixel_9584/NB1 pixel_9584/VBIAS pixel_9584/NB2 pixel_9584/AMP_IN pixel_9584/SF_IB
+ pixel_9584/PIX_OUT pixel_9584/CSA_VREF pixel
Xpixel_9573 pixel_9573/gring pixel_9573/VDD pixel_9573/GND pixel_9573/VREF pixel_9573/ROW_SEL
+ pixel_9573/NB1 pixel_9573/VBIAS pixel_9573/NB2 pixel_9573/AMP_IN pixel_9573/SF_IB
+ pixel_9573/PIX_OUT pixel_9573/CSA_VREF pixel
Xpixel_9562 pixel_9562/gring pixel_9562/VDD pixel_9562/GND pixel_9562/VREF pixel_9562/ROW_SEL
+ pixel_9562/NB1 pixel_9562/VBIAS pixel_9562/NB2 pixel_9562/AMP_IN pixel_9562/SF_IB
+ pixel_9562/PIX_OUT pixel_9562/CSA_VREF pixel
Xpixel_9551 pixel_9551/gring pixel_9551/VDD pixel_9551/GND pixel_9551/VREF pixel_9551/ROW_SEL
+ pixel_9551/NB1 pixel_9551/VBIAS pixel_9551/NB2 pixel_9551/AMP_IN pixel_9551/SF_IB
+ pixel_9551/PIX_OUT pixel_9551/CSA_VREF pixel
Xpixel_8872 pixel_8872/gring pixel_8872/VDD pixel_8872/GND pixel_8872/VREF pixel_8872/ROW_SEL
+ pixel_8872/NB1 pixel_8872/VBIAS pixel_8872/NB2 pixel_8872/AMP_IN pixel_8872/SF_IB
+ pixel_8872/PIX_OUT pixel_8872/CSA_VREF pixel
Xpixel_8861 pixel_8861/gring pixel_8861/VDD pixel_8861/GND pixel_8861/VREF pixel_8861/ROW_SEL
+ pixel_8861/NB1 pixel_8861/VBIAS pixel_8861/NB2 pixel_8861/AMP_IN pixel_8861/SF_IB
+ pixel_8861/PIX_OUT pixel_8861/CSA_VREF pixel
Xpixel_8850 pixel_8850/gring pixel_8850/VDD pixel_8850/GND pixel_8850/VREF pixel_8850/ROW_SEL
+ pixel_8850/NB1 pixel_8850/VBIAS pixel_8850/NB2 pixel_8850/AMP_IN pixel_8850/SF_IB
+ pixel_8850/PIX_OUT pixel_8850/CSA_VREF pixel
Xpixel_9595 pixel_9595/gring pixel_9595/VDD pixel_9595/GND pixel_9595/VREF pixel_9595/ROW_SEL
+ pixel_9595/NB1 pixel_9595/VBIAS pixel_9595/NB2 pixel_9595/AMP_IN pixel_9595/SF_IB
+ pixel_9595/PIX_OUT pixel_9595/CSA_VREF pixel
Xpixel_8894 pixel_8894/gring pixel_8894/VDD pixel_8894/GND pixel_8894/VREF pixel_8894/ROW_SEL
+ pixel_8894/NB1 pixel_8894/VBIAS pixel_8894/NB2 pixel_8894/AMP_IN pixel_8894/SF_IB
+ pixel_8894/PIX_OUT pixel_8894/CSA_VREF pixel
Xpixel_8883 pixel_8883/gring pixel_8883/VDD pixel_8883/GND pixel_8883/VREF pixel_8883/ROW_SEL
+ pixel_8883/NB1 pixel_8883/VBIAS pixel_8883/NB2 pixel_8883/AMP_IN pixel_8883/SF_IB
+ pixel_8883/PIX_OUT pixel_8883/CSA_VREF pixel
Xpixel_3190 pixel_3190/gring pixel_3190/VDD pixel_3190/GND pixel_3190/VREF pixel_3190/ROW_SEL
+ pixel_3190/NB1 pixel_3190/VBIAS pixel_3190/NB2 pixel_3190/AMP_IN pixel_3190/SF_IB
+ pixel_3190/PIX_OUT pixel_3190/CSA_VREF pixel
Xpixel_5509 pixel_5509/gring pixel_5509/VDD pixel_5509/GND pixel_5509/VREF pixel_5509/ROW_SEL
+ pixel_5509/NB1 pixel_5509/VBIAS pixel_5509/NB2 pixel_5509/AMP_IN pixel_5509/SF_IB
+ pixel_5509/PIX_OUT pixel_5509/CSA_VREF pixel
Xpixel_814 pixel_814/gring pixel_814/VDD pixel_814/GND pixel_814/VREF pixel_814/ROW_SEL
+ pixel_814/NB1 pixel_814/VBIAS pixel_814/NB2 pixel_814/AMP_IN pixel_814/SF_IB pixel_814/PIX_OUT
+ pixel_814/CSA_VREF pixel
Xpixel_803 pixel_803/gring pixel_803/VDD pixel_803/GND pixel_803/VREF pixel_803/ROW_SEL
+ pixel_803/NB1 pixel_803/VBIAS pixel_803/NB2 pixel_803/AMP_IN pixel_803/SF_IB pixel_803/PIX_OUT
+ pixel_803/CSA_VREF pixel
Xpixel_4808 pixel_4808/gring pixel_4808/VDD pixel_4808/GND pixel_4808/VREF pixel_4808/ROW_SEL
+ pixel_4808/NB1 pixel_4808/VBIAS pixel_4808/NB2 pixel_4808/AMP_IN pixel_4808/SF_IB
+ pixel_4808/PIX_OUT pixel_4808/CSA_VREF pixel
Xpixel_4819 pixel_4819/gring pixel_4819/VDD pixel_4819/GND pixel_4819/VREF pixel_4819/ROW_SEL
+ pixel_4819/NB1 pixel_4819/VBIAS pixel_4819/NB2 pixel_4819/AMP_IN pixel_4819/SF_IB
+ pixel_4819/PIX_OUT pixel_4819/CSA_VREF pixel
Xpixel_847 pixel_847/gring pixel_847/VDD pixel_847/GND pixel_847/VREF pixel_847/ROW_SEL
+ pixel_847/NB1 pixel_847/VBIAS pixel_847/NB2 pixel_847/AMP_IN pixel_847/SF_IB pixel_847/PIX_OUT
+ pixel_847/CSA_VREF pixel
Xpixel_836 pixel_836/gring pixel_836/VDD pixel_836/GND pixel_836/VREF pixel_836/ROW_SEL
+ pixel_836/NB1 pixel_836/VBIAS pixel_836/NB2 pixel_836/AMP_IN pixel_836/SF_IB pixel_836/PIX_OUT
+ pixel_836/CSA_VREF pixel
Xpixel_825 pixel_825/gring pixel_825/VDD pixel_825/GND pixel_825/VREF pixel_825/ROW_SEL
+ pixel_825/NB1 pixel_825/VBIAS pixel_825/NB2 pixel_825/AMP_IN pixel_825/SF_IB pixel_825/PIX_OUT
+ pixel_825/CSA_VREF pixel
Xpixel_869 pixel_869/gring pixel_869/VDD pixel_869/GND pixel_869/VREF pixel_869/ROW_SEL
+ pixel_869/NB1 pixel_869/VBIAS pixel_869/NB2 pixel_869/AMP_IN pixel_869/SF_IB pixel_869/PIX_OUT
+ pixel_869/CSA_VREF pixel
Xpixel_858 pixel_858/gring pixel_858/VDD pixel_858/GND pixel_858/VREF pixel_858/ROW_SEL
+ pixel_858/NB1 pixel_858/VBIAS pixel_858/NB2 pixel_858/AMP_IN pixel_858/SF_IB pixel_858/PIX_OUT
+ pixel_858/CSA_VREF pixel
Xpixel_8102 pixel_8102/gring pixel_8102/VDD pixel_8102/GND pixel_8102/VREF pixel_8102/ROW_SEL
+ pixel_8102/NB1 pixel_8102/VBIAS pixel_8102/NB2 pixel_8102/AMP_IN pixel_8102/SF_IB
+ pixel_8102/PIX_OUT pixel_8102/CSA_VREF pixel
Xpixel_8113 pixel_8113/gring pixel_8113/VDD pixel_8113/GND pixel_8113/VREF pixel_8113/ROW_SEL
+ pixel_8113/NB1 pixel_8113/VBIAS pixel_8113/NB2 pixel_8113/AMP_IN pixel_8113/SF_IB
+ pixel_8113/PIX_OUT pixel_8113/CSA_VREF pixel
Xpixel_8124 pixel_8124/gring pixel_8124/VDD pixel_8124/GND pixel_8124/VREF pixel_8124/ROW_SEL
+ pixel_8124/NB1 pixel_8124/VBIAS pixel_8124/NB2 pixel_8124/AMP_IN pixel_8124/SF_IB
+ pixel_8124/PIX_OUT pixel_8124/CSA_VREF pixel
Xpixel_8135 pixel_8135/gring pixel_8135/VDD pixel_8135/GND pixel_8135/VREF pixel_8135/ROW_SEL
+ pixel_8135/NB1 pixel_8135/VBIAS pixel_8135/NB2 pixel_8135/AMP_IN pixel_8135/SF_IB
+ pixel_8135/PIX_OUT pixel_8135/CSA_VREF pixel
Xpixel_8146 pixel_8146/gring pixel_8146/VDD pixel_8146/GND pixel_8146/VREF pixel_8146/ROW_SEL
+ pixel_8146/NB1 pixel_8146/VBIAS pixel_8146/NB2 pixel_8146/AMP_IN pixel_8146/SF_IB
+ pixel_8146/PIX_OUT pixel_8146/CSA_VREF pixel
Xpixel_8157 pixel_8157/gring pixel_8157/VDD pixel_8157/GND pixel_8157/VREF pixel_8157/ROW_SEL
+ pixel_8157/NB1 pixel_8157/VBIAS pixel_8157/NB2 pixel_8157/AMP_IN pixel_8157/SF_IB
+ pixel_8157/PIX_OUT pixel_8157/CSA_VREF pixel
Xpixel_8168 pixel_8168/gring pixel_8168/VDD pixel_8168/GND pixel_8168/VREF pixel_8168/ROW_SEL
+ pixel_8168/NB1 pixel_8168/VBIAS pixel_8168/NB2 pixel_8168/AMP_IN pixel_8168/SF_IB
+ pixel_8168/PIX_OUT pixel_8168/CSA_VREF pixel
Xpixel_7401 pixel_7401/gring pixel_7401/VDD pixel_7401/GND pixel_7401/VREF pixel_7401/ROW_SEL
+ pixel_7401/NB1 pixel_7401/VBIAS pixel_7401/NB2 pixel_7401/AMP_IN pixel_7401/SF_IB
+ pixel_7401/PIX_OUT pixel_7401/CSA_VREF pixel
Xpixel_7412 pixel_7412/gring pixel_7412/VDD pixel_7412/GND pixel_7412/VREF pixel_7412/ROW_SEL
+ pixel_7412/NB1 pixel_7412/VBIAS pixel_7412/NB2 pixel_7412/AMP_IN pixel_7412/SF_IB
+ pixel_7412/PIX_OUT pixel_7412/CSA_VREF pixel
Xpixel_7423 pixel_7423/gring pixel_7423/VDD pixel_7423/GND pixel_7423/VREF pixel_7423/ROW_SEL
+ pixel_7423/NB1 pixel_7423/VBIAS pixel_7423/NB2 pixel_7423/AMP_IN pixel_7423/SF_IB
+ pixel_7423/PIX_OUT pixel_7423/CSA_VREF pixel
Xpixel_8179 pixel_8179/gring pixel_8179/VDD pixel_8179/GND pixel_8179/VREF pixel_8179/ROW_SEL
+ pixel_8179/NB1 pixel_8179/VBIAS pixel_8179/NB2 pixel_8179/AMP_IN pixel_8179/SF_IB
+ pixel_8179/PIX_OUT pixel_8179/CSA_VREF pixel
Xpixel_7434 pixel_7434/gring pixel_7434/VDD pixel_7434/GND pixel_7434/VREF pixel_7434/ROW_SEL
+ pixel_7434/NB1 pixel_7434/VBIAS pixel_7434/NB2 pixel_7434/AMP_IN pixel_7434/SF_IB
+ pixel_7434/PIX_OUT pixel_7434/CSA_VREF pixel
Xpixel_7445 pixel_7445/gring pixel_7445/VDD pixel_7445/GND pixel_7445/VREF pixel_7445/ROW_SEL
+ pixel_7445/NB1 pixel_7445/VBIAS pixel_7445/NB2 pixel_7445/AMP_IN pixel_7445/SF_IB
+ pixel_7445/PIX_OUT pixel_7445/CSA_VREF pixel
Xpixel_7456 pixel_7456/gring pixel_7456/VDD pixel_7456/GND pixel_7456/VREF pixel_7456/ROW_SEL
+ pixel_7456/NB1 pixel_7456/VBIAS pixel_7456/NB2 pixel_7456/AMP_IN pixel_7456/SF_IB
+ pixel_7456/PIX_OUT pixel_7456/CSA_VREF pixel
Xpixel_6700 pixel_6700/gring pixel_6700/VDD pixel_6700/GND pixel_6700/VREF pixel_6700/ROW_SEL
+ pixel_6700/NB1 pixel_6700/VBIAS pixel_6700/NB2 pixel_6700/AMP_IN pixel_6700/SF_IB
+ pixel_6700/PIX_OUT pixel_6700/CSA_VREF pixel
Xpixel_6711 pixel_6711/gring pixel_6711/VDD pixel_6711/GND pixel_6711/VREF pixel_6711/ROW_SEL
+ pixel_6711/NB1 pixel_6711/VBIAS pixel_6711/NB2 pixel_6711/AMP_IN pixel_6711/SF_IB
+ pixel_6711/PIX_OUT pixel_6711/CSA_VREF pixel
Xpixel_7467 pixel_7467/gring pixel_7467/VDD pixel_7467/GND pixel_7467/VREF pixel_7467/ROW_SEL
+ pixel_7467/NB1 pixel_7467/VBIAS pixel_7467/NB2 pixel_7467/AMP_IN pixel_7467/SF_IB
+ pixel_7467/PIX_OUT pixel_7467/CSA_VREF pixel
Xpixel_7478 pixel_7478/gring pixel_7478/VDD pixel_7478/GND pixel_7478/VREF pixel_7478/ROW_SEL
+ pixel_7478/NB1 pixel_7478/VBIAS pixel_7478/NB2 pixel_7478/AMP_IN pixel_7478/SF_IB
+ pixel_7478/PIX_OUT pixel_7478/CSA_VREF pixel
Xpixel_7489 pixel_7489/gring pixel_7489/VDD pixel_7489/GND pixel_7489/VREF pixel_7489/ROW_SEL
+ pixel_7489/NB1 pixel_7489/VBIAS pixel_7489/NB2 pixel_7489/AMP_IN pixel_7489/SF_IB
+ pixel_7489/PIX_OUT pixel_7489/CSA_VREF pixel
Xpixel_6722 pixel_6722/gring pixel_6722/VDD pixel_6722/GND pixel_6722/VREF pixel_6722/ROW_SEL
+ pixel_6722/NB1 pixel_6722/VBIAS pixel_6722/NB2 pixel_6722/AMP_IN pixel_6722/SF_IB
+ pixel_6722/PIX_OUT pixel_6722/CSA_VREF pixel
Xpixel_6733 pixel_6733/gring pixel_6733/VDD pixel_6733/GND pixel_6733/VREF pixel_6733/ROW_SEL
+ pixel_6733/NB1 pixel_6733/VBIAS pixel_6733/NB2 pixel_6733/AMP_IN pixel_6733/SF_IB
+ pixel_6733/PIX_OUT pixel_6733/CSA_VREF pixel
Xpixel_6744 pixel_6744/gring pixel_6744/VDD pixel_6744/GND pixel_6744/VREF pixel_6744/ROW_SEL
+ pixel_6744/NB1 pixel_6744/VBIAS pixel_6744/NB2 pixel_6744/AMP_IN pixel_6744/SF_IB
+ pixel_6744/PIX_OUT pixel_6744/CSA_VREF pixel
Xpixel_6755 pixel_6755/gring pixel_6755/VDD pixel_6755/GND pixel_6755/VREF pixel_6755/ROW_SEL
+ pixel_6755/NB1 pixel_6755/VBIAS pixel_6755/NB2 pixel_6755/AMP_IN pixel_6755/SF_IB
+ pixel_6755/PIX_OUT pixel_6755/CSA_VREF pixel
Xpixel_6766 pixel_6766/gring pixel_6766/VDD pixel_6766/GND pixel_6766/VREF pixel_6766/ROW_SEL
+ pixel_6766/NB1 pixel_6766/VBIAS pixel_6766/NB2 pixel_6766/AMP_IN pixel_6766/SF_IB
+ pixel_6766/PIX_OUT pixel_6766/CSA_VREF pixel
Xpixel_6777 pixel_6777/gring pixel_6777/VDD pixel_6777/GND pixel_6777/VREF pixel_6777/ROW_SEL
+ pixel_6777/NB1 pixel_6777/VBIAS pixel_6777/NB2 pixel_6777/AMP_IN pixel_6777/SF_IB
+ pixel_6777/PIX_OUT pixel_6777/CSA_VREF pixel
Xpixel_6788 pixel_6788/gring pixel_6788/VDD pixel_6788/GND pixel_6788/VREF pixel_6788/ROW_SEL
+ pixel_6788/NB1 pixel_6788/VBIAS pixel_6788/NB2 pixel_6788/AMP_IN pixel_6788/SF_IB
+ pixel_6788/PIX_OUT pixel_6788/CSA_VREF pixel
Xpixel_6799 pixel_6799/gring pixel_6799/VDD pixel_6799/GND pixel_6799/VREF pixel_6799/ROW_SEL
+ pixel_6799/NB1 pixel_6799/VBIAS pixel_6799/NB2 pixel_6799/AMP_IN pixel_6799/SF_IB
+ pixel_6799/PIX_OUT pixel_6799/CSA_VREF pixel
Xpixel_1051 pixel_1051/gring pixel_1051/VDD pixel_1051/GND pixel_1051/VREF pixel_1051/ROW_SEL
+ pixel_1051/NB1 pixel_1051/VBIAS pixel_1051/NB2 pixel_1051/AMP_IN pixel_1051/SF_IB
+ pixel_1051/PIX_OUT pixel_1051/CSA_VREF pixel
Xpixel_1040 pixel_1040/gring pixel_1040/VDD pixel_1040/GND pixel_1040/VREF pixel_1040/ROW_SEL
+ pixel_1040/NB1 pixel_1040/VBIAS pixel_1040/NB2 pixel_1040/AMP_IN pixel_1040/SF_IB
+ pixel_1040/PIX_OUT pixel_1040/CSA_VREF pixel
Xpixel_1084 pixel_1084/gring pixel_1084/VDD pixel_1084/GND pixel_1084/VREF pixel_1084/ROW_SEL
+ pixel_1084/NB1 pixel_1084/VBIAS pixel_1084/NB2 pixel_1084/AMP_IN pixel_1084/SF_IB
+ pixel_1084/PIX_OUT pixel_1084/CSA_VREF pixel
Xpixel_1073 pixel_1073/gring pixel_1073/VDD pixel_1073/GND pixel_1073/VREF pixel_1073/ROW_SEL
+ pixel_1073/NB1 pixel_1073/VBIAS pixel_1073/NB2 pixel_1073/AMP_IN pixel_1073/SF_IB
+ pixel_1073/PIX_OUT pixel_1073/CSA_VREF pixel
Xpixel_1062 pixel_1062/gring pixel_1062/VDD pixel_1062/GND pixel_1062/VREF pixel_1062/ROW_SEL
+ pixel_1062/NB1 pixel_1062/VBIAS pixel_1062/NB2 pixel_1062/AMP_IN pixel_1062/SF_IB
+ pixel_1062/PIX_OUT pixel_1062/CSA_VREF pixel
Xpixel_1095 pixel_1095/gring pixel_1095/VDD pixel_1095/GND pixel_1095/VREF pixel_1095/ROW_SEL
+ pixel_1095/NB1 pixel_1095/VBIAS pixel_1095/NB2 pixel_1095/AMP_IN pixel_1095/SF_IB
+ pixel_1095/PIX_OUT pixel_1095/CSA_VREF pixel
Xpixel_9392 pixel_9392/gring pixel_9392/VDD pixel_9392/GND pixel_9392/VREF pixel_9392/ROW_SEL
+ pixel_9392/NB1 pixel_9392/VBIAS pixel_9392/NB2 pixel_9392/AMP_IN pixel_9392/SF_IB
+ pixel_9392/PIX_OUT pixel_9392/CSA_VREF pixel
Xpixel_9381 pixel_9381/gring pixel_9381/VDD pixel_9381/GND pixel_9381/VREF pixel_9381/ROW_SEL
+ pixel_9381/NB1 pixel_9381/VBIAS pixel_9381/NB2 pixel_9381/AMP_IN pixel_9381/SF_IB
+ pixel_9381/PIX_OUT pixel_9381/CSA_VREF pixel
Xpixel_9370 pixel_9370/gring pixel_9370/VDD pixel_9370/GND pixel_9370/VREF pixel_9370/ROW_SEL
+ pixel_9370/NB1 pixel_9370/VBIAS pixel_9370/NB2 pixel_9370/AMP_IN pixel_9370/SF_IB
+ pixel_9370/PIX_OUT pixel_9370/CSA_VREF pixel
Xpixel_8680 pixel_8680/gring pixel_8680/VDD pixel_8680/GND pixel_8680/VREF pixel_8680/ROW_SEL
+ pixel_8680/NB1 pixel_8680/VBIAS pixel_8680/NB2 pixel_8680/AMP_IN pixel_8680/SF_IB
+ pixel_8680/PIX_OUT pixel_8680/CSA_VREF pixel
Xpixel_8691 pixel_8691/gring pixel_8691/VDD pixel_8691/GND pixel_8691/VREF pixel_8691/ROW_SEL
+ pixel_8691/NB1 pixel_8691/VBIAS pixel_8691/NB2 pixel_8691/AMP_IN pixel_8691/SF_IB
+ pixel_8691/PIX_OUT pixel_8691/CSA_VREF pixel
Xpixel_7990 pixel_7990/gring pixel_7990/VDD pixel_7990/GND pixel_7990/VREF pixel_7990/ROW_SEL
+ pixel_7990/NB1 pixel_7990/VBIAS pixel_7990/NB2 pixel_7990/AMP_IN pixel_7990/SF_IB
+ pixel_7990/PIX_OUT pixel_7990/CSA_VREF pixel
Xpixel_6007 pixel_6007/gring pixel_6007/VDD pixel_6007/GND pixel_6007/VREF pixel_6007/ROW_SEL
+ pixel_6007/NB1 pixel_6007/VBIAS pixel_6007/NB2 pixel_6007/AMP_IN pixel_6007/SF_IB
+ pixel_6007/PIX_OUT pixel_6007/CSA_VREF pixel
Xpixel_6018 pixel_6018/gring pixel_6018/VDD pixel_6018/GND pixel_6018/VREF pixel_6018/ROW_SEL
+ pixel_6018/NB1 pixel_6018/VBIAS pixel_6018/NB2 pixel_6018/AMP_IN pixel_6018/SF_IB
+ pixel_6018/PIX_OUT pixel_6018/CSA_VREF pixel
Xpixel_6029 pixel_6029/gring pixel_6029/VDD pixel_6029/GND pixel_6029/VREF pixel_6029/ROW_SEL
+ pixel_6029/NB1 pixel_6029/VBIAS pixel_6029/NB2 pixel_6029/AMP_IN pixel_6029/SF_IB
+ pixel_6029/PIX_OUT pixel_6029/CSA_VREF pixel
Xpixel_5306 pixel_5306/gring pixel_5306/VDD pixel_5306/GND pixel_5306/VREF pixel_5306/ROW_SEL
+ pixel_5306/NB1 pixel_5306/VBIAS pixel_5306/NB2 pixel_5306/AMP_IN pixel_5306/SF_IB
+ pixel_5306/PIX_OUT pixel_5306/CSA_VREF pixel
Xpixel_5317 pixel_5317/gring pixel_5317/VDD pixel_5317/GND pixel_5317/VREF pixel_5317/ROW_SEL
+ pixel_5317/NB1 pixel_5317/VBIAS pixel_5317/NB2 pixel_5317/AMP_IN pixel_5317/SF_IB
+ pixel_5317/PIX_OUT pixel_5317/CSA_VREF pixel
Xpixel_5328 pixel_5328/gring pixel_5328/VDD pixel_5328/GND pixel_5328/VREF pixel_5328/ROW_SEL
+ pixel_5328/NB1 pixel_5328/VBIAS pixel_5328/NB2 pixel_5328/AMP_IN pixel_5328/SF_IB
+ pixel_5328/PIX_OUT pixel_5328/CSA_VREF pixel
Xpixel_5339 pixel_5339/gring pixel_5339/VDD pixel_5339/GND pixel_5339/VREF pixel_5339/ROW_SEL
+ pixel_5339/NB1 pixel_5339/VBIAS pixel_5339/NB2 pixel_5339/AMP_IN pixel_5339/SF_IB
+ pixel_5339/PIX_OUT pixel_5339/CSA_VREF pixel
Xpixel_622 pixel_622/gring pixel_622/VDD pixel_622/GND pixel_622/VREF pixel_622/ROW_SEL
+ pixel_622/NB1 pixel_622/VBIAS pixel_622/NB2 pixel_622/AMP_IN pixel_622/SF_IB pixel_622/PIX_OUT
+ pixel_622/CSA_VREF pixel
Xpixel_611 pixel_611/gring pixel_611/VDD pixel_611/GND pixel_611/VREF pixel_611/ROW_SEL
+ pixel_611/NB1 pixel_611/VBIAS pixel_611/NB2 pixel_611/AMP_IN pixel_611/SF_IB pixel_611/PIX_OUT
+ pixel_611/CSA_VREF pixel
Xpixel_600 pixel_600/gring pixel_600/VDD pixel_600/GND pixel_600/VREF pixel_600/ROW_SEL
+ pixel_600/NB1 pixel_600/VBIAS pixel_600/NB2 pixel_600/AMP_IN pixel_600/SF_IB pixel_600/PIX_OUT
+ pixel_600/CSA_VREF pixel
Xpixel_4605 pixel_4605/gring pixel_4605/VDD pixel_4605/GND pixel_4605/VREF pixel_4605/ROW_SEL
+ pixel_4605/NB1 pixel_4605/VBIAS pixel_4605/NB2 pixel_4605/AMP_IN pixel_4605/SF_IB
+ pixel_4605/PIX_OUT pixel_4605/CSA_VREF pixel
Xpixel_4616 pixel_4616/gring pixel_4616/VDD pixel_4616/GND pixel_4616/VREF pixel_4616/ROW_SEL
+ pixel_4616/NB1 pixel_4616/VBIAS pixel_4616/NB2 pixel_4616/AMP_IN pixel_4616/SF_IB
+ pixel_4616/PIX_OUT pixel_4616/CSA_VREF pixel
Xpixel_4627 pixel_4627/gring pixel_4627/VDD pixel_4627/GND pixel_4627/VREF pixel_4627/ROW_SEL
+ pixel_4627/NB1 pixel_4627/VBIAS pixel_4627/NB2 pixel_4627/AMP_IN pixel_4627/SF_IB
+ pixel_4627/PIX_OUT pixel_4627/CSA_VREF pixel
Xpixel_666 pixel_666/gring pixel_666/VDD pixel_666/GND pixel_666/VREF pixel_666/ROW_SEL
+ pixel_666/NB1 pixel_666/VBIAS pixel_666/NB2 pixel_666/AMP_IN pixel_666/SF_IB pixel_666/PIX_OUT
+ pixel_666/CSA_VREF pixel
Xpixel_655 pixel_655/gring pixel_655/VDD pixel_655/GND pixel_655/VREF pixel_655/ROW_SEL
+ pixel_655/NB1 pixel_655/VBIAS pixel_655/NB2 pixel_655/AMP_IN pixel_655/SF_IB pixel_655/PIX_OUT
+ pixel_655/CSA_VREF pixel
Xpixel_644 pixel_644/gring pixel_644/VDD pixel_644/GND pixel_644/VREF pixel_644/ROW_SEL
+ pixel_644/NB1 pixel_644/VBIAS pixel_644/NB2 pixel_644/AMP_IN pixel_644/SF_IB pixel_644/PIX_OUT
+ pixel_644/CSA_VREF pixel
Xpixel_633 pixel_633/gring pixel_633/VDD pixel_633/GND pixel_633/VREF pixel_633/ROW_SEL
+ pixel_633/NB1 pixel_633/VBIAS pixel_633/NB2 pixel_633/AMP_IN pixel_633/SF_IB pixel_633/PIX_OUT
+ pixel_633/CSA_VREF pixel
Xpixel_4638 pixel_4638/gring pixel_4638/VDD pixel_4638/GND pixel_4638/VREF pixel_4638/ROW_SEL
+ pixel_4638/NB1 pixel_4638/VBIAS pixel_4638/NB2 pixel_4638/AMP_IN pixel_4638/SF_IB
+ pixel_4638/PIX_OUT pixel_4638/CSA_VREF pixel
Xpixel_4649 pixel_4649/gring pixel_4649/VDD pixel_4649/GND pixel_4649/VREF pixel_4649/ROW_SEL
+ pixel_4649/NB1 pixel_4649/VBIAS pixel_4649/NB2 pixel_4649/AMP_IN pixel_4649/SF_IB
+ pixel_4649/PIX_OUT pixel_4649/CSA_VREF pixel
Xpixel_3904 pixel_3904/gring pixel_3904/VDD pixel_3904/GND pixel_3904/VREF pixel_3904/ROW_SEL
+ pixel_3904/NB1 pixel_3904/VBIAS pixel_3904/NB2 pixel_3904/AMP_IN pixel_3904/SF_IB
+ pixel_3904/PIX_OUT pixel_3904/CSA_VREF pixel
Xpixel_3915 pixel_3915/gring pixel_3915/VDD pixel_3915/GND pixel_3915/VREF pixel_3915/ROW_SEL
+ pixel_3915/NB1 pixel_3915/VBIAS pixel_3915/NB2 pixel_3915/AMP_IN pixel_3915/SF_IB
+ pixel_3915/PIX_OUT pixel_3915/CSA_VREF pixel
Xpixel_3926 pixel_3926/gring pixel_3926/VDD pixel_3926/GND pixel_3926/VREF pixel_3926/ROW_SEL
+ pixel_3926/NB1 pixel_3926/VBIAS pixel_3926/NB2 pixel_3926/AMP_IN pixel_3926/SF_IB
+ pixel_3926/PIX_OUT pixel_3926/CSA_VREF pixel
Xpixel_699 pixel_699/gring pixel_699/VDD pixel_699/GND pixel_699/VREF pixel_699/ROW_SEL
+ pixel_699/NB1 pixel_699/VBIAS pixel_699/NB2 pixel_699/AMP_IN pixel_699/SF_IB pixel_699/PIX_OUT
+ pixel_699/CSA_VREF pixel
Xpixel_688 pixel_688/gring pixel_688/VDD pixel_688/GND pixel_688/VREF pixel_688/ROW_SEL
+ pixel_688/NB1 pixel_688/VBIAS pixel_688/NB2 pixel_688/AMP_IN pixel_688/SF_IB pixel_688/PIX_OUT
+ pixel_688/CSA_VREF pixel
Xpixel_677 pixel_677/gring pixel_677/VDD pixel_677/GND pixel_677/VREF pixel_677/ROW_SEL
+ pixel_677/NB1 pixel_677/VBIAS pixel_677/NB2 pixel_677/AMP_IN pixel_677/SF_IB pixel_677/PIX_OUT
+ pixel_677/CSA_VREF pixel
Xpixel_3937 pixel_3937/gring pixel_3937/VDD pixel_3937/GND pixel_3937/VREF pixel_3937/ROW_SEL
+ pixel_3937/NB1 pixel_3937/VBIAS pixel_3937/NB2 pixel_3937/AMP_IN pixel_3937/SF_IB
+ pixel_3937/PIX_OUT pixel_3937/CSA_VREF pixel
Xpixel_3948 pixel_3948/gring pixel_3948/VDD pixel_3948/GND pixel_3948/VREF pixel_3948/ROW_SEL
+ pixel_3948/NB1 pixel_3948/VBIAS pixel_3948/NB2 pixel_3948/AMP_IN pixel_3948/SF_IB
+ pixel_3948/PIX_OUT pixel_3948/CSA_VREF pixel
Xpixel_3959 pixel_3959/gring pixel_3959/VDD pixel_3959/GND pixel_3959/VREF pixel_3959/ROW_SEL
+ pixel_3959/NB1 pixel_3959/VBIAS pixel_3959/NB2 pixel_3959/AMP_IN pixel_3959/SF_IB
+ pixel_3959/PIX_OUT pixel_3959/CSA_VREF pixel
Xpixel_7220 pixel_7220/gring pixel_7220/VDD pixel_7220/GND pixel_7220/VREF pixel_7220/ROW_SEL
+ pixel_7220/NB1 pixel_7220/VBIAS pixel_7220/NB2 pixel_7220/AMP_IN pixel_7220/SF_IB
+ pixel_7220/PIX_OUT pixel_7220/CSA_VREF pixel
Xpixel_7231 pixel_7231/gring pixel_7231/VDD pixel_7231/GND pixel_7231/VREF pixel_7231/ROW_SEL
+ pixel_7231/NB1 pixel_7231/VBIAS pixel_7231/NB2 pixel_7231/AMP_IN pixel_7231/SF_IB
+ pixel_7231/PIX_OUT pixel_7231/CSA_VREF pixel
Xpixel_7242 pixel_7242/gring pixel_7242/VDD pixel_7242/GND pixel_7242/VREF pixel_7242/ROW_SEL
+ pixel_7242/NB1 pixel_7242/VBIAS pixel_7242/NB2 pixel_7242/AMP_IN pixel_7242/SF_IB
+ pixel_7242/PIX_OUT pixel_7242/CSA_VREF pixel
Xpixel_7253 pixel_7253/gring pixel_7253/VDD pixel_7253/GND pixel_7253/VREF pixel_7253/ROW_SEL
+ pixel_7253/NB1 pixel_7253/VBIAS pixel_7253/NB2 pixel_7253/AMP_IN pixel_7253/SF_IB
+ pixel_7253/PIX_OUT pixel_7253/CSA_VREF pixel
Xpixel_7264 pixel_7264/gring pixel_7264/VDD pixel_7264/GND pixel_7264/VREF pixel_7264/ROW_SEL
+ pixel_7264/NB1 pixel_7264/VBIAS pixel_7264/NB2 pixel_7264/AMP_IN pixel_7264/SF_IB
+ pixel_7264/PIX_OUT pixel_7264/CSA_VREF pixel
Xpixel_6530 pixel_6530/gring pixel_6530/VDD pixel_6530/GND pixel_6530/VREF pixel_6530/ROW_SEL
+ pixel_6530/NB1 pixel_6530/VBIAS pixel_6530/NB2 pixel_6530/AMP_IN pixel_6530/SF_IB
+ pixel_6530/PIX_OUT pixel_6530/CSA_VREF pixel
Xpixel_7275 pixel_7275/gring pixel_7275/VDD pixel_7275/GND pixel_7275/VREF pixel_7275/ROW_SEL
+ pixel_7275/NB1 pixel_7275/VBIAS pixel_7275/NB2 pixel_7275/AMP_IN pixel_7275/SF_IB
+ pixel_7275/PIX_OUT pixel_7275/CSA_VREF pixel
Xpixel_7286 pixel_7286/gring pixel_7286/VDD pixel_7286/GND pixel_7286/VREF pixel_7286/ROW_SEL
+ pixel_7286/NB1 pixel_7286/VBIAS pixel_7286/NB2 pixel_7286/AMP_IN pixel_7286/SF_IB
+ pixel_7286/PIX_OUT pixel_7286/CSA_VREF pixel
Xpixel_7297 pixel_7297/gring pixel_7297/VDD pixel_7297/GND pixel_7297/VREF pixel_7297/ROW_SEL
+ pixel_7297/NB1 pixel_7297/VBIAS pixel_7297/NB2 pixel_7297/AMP_IN pixel_7297/SF_IB
+ pixel_7297/PIX_OUT pixel_7297/CSA_VREF pixel
Xpixel_6541 pixel_6541/gring pixel_6541/VDD pixel_6541/GND pixel_6541/VREF pixel_6541/ROW_SEL
+ pixel_6541/NB1 pixel_6541/VBIAS pixel_6541/NB2 pixel_6541/AMP_IN pixel_6541/SF_IB
+ pixel_6541/PIX_OUT pixel_6541/CSA_VREF pixel
Xpixel_6552 pixel_6552/gring pixel_6552/VDD pixel_6552/GND pixel_6552/VREF pixel_6552/ROW_SEL
+ pixel_6552/NB1 pixel_6552/VBIAS pixel_6552/NB2 pixel_6552/AMP_IN pixel_6552/SF_IB
+ pixel_6552/PIX_OUT pixel_6552/CSA_VREF pixel
Xpixel_6563 pixel_6563/gring pixel_6563/VDD pixel_6563/GND pixel_6563/VREF pixel_6563/ROW_SEL
+ pixel_6563/NB1 pixel_6563/VBIAS pixel_6563/NB2 pixel_6563/AMP_IN pixel_6563/SF_IB
+ pixel_6563/PIX_OUT pixel_6563/CSA_VREF pixel
Xpixel_6574 pixel_6574/gring pixel_6574/VDD pixel_6574/GND pixel_6574/VREF pixel_6574/ROW_SEL
+ pixel_6574/NB1 pixel_6574/VBIAS pixel_6574/NB2 pixel_6574/AMP_IN pixel_6574/SF_IB
+ pixel_6574/PIX_OUT pixel_6574/CSA_VREF pixel
Xpixel_6585 pixel_6585/gring pixel_6585/VDD pixel_6585/GND pixel_6585/VREF pixel_6585/ROW_SEL
+ pixel_6585/NB1 pixel_6585/VBIAS pixel_6585/NB2 pixel_6585/AMP_IN pixel_6585/SF_IB
+ pixel_6585/PIX_OUT pixel_6585/CSA_VREF pixel
Xpixel_6596 pixel_6596/gring pixel_6596/VDD pixel_6596/GND pixel_6596/VREF pixel_6596/ROW_SEL
+ pixel_6596/NB1 pixel_6596/VBIAS pixel_6596/NB2 pixel_6596/AMP_IN pixel_6596/SF_IB
+ pixel_6596/PIX_OUT pixel_6596/CSA_VREF pixel
Xpixel_5840 pixel_5840/gring pixel_5840/VDD pixel_5840/GND pixel_5840/VREF pixel_5840/ROW_SEL
+ pixel_5840/NB1 pixel_5840/VBIAS pixel_5840/NB2 pixel_5840/AMP_IN pixel_5840/SF_IB
+ pixel_5840/PIX_OUT pixel_5840/CSA_VREF pixel
Xpixel_5851 pixel_5851/gring pixel_5851/VDD pixel_5851/GND pixel_5851/VREF pixel_5851/ROW_SEL
+ pixel_5851/NB1 pixel_5851/VBIAS pixel_5851/NB2 pixel_5851/AMP_IN pixel_5851/SF_IB
+ pixel_5851/PIX_OUT pixel_5851/CSA_VREF pixel
Xpixel_5862 pixel_5862/gring pixel_5862/VDD pixel_5862/GND pixel_5862/VREF pixel_5862/ROW_SEL
+ pixel_5862/NB1 pixel_5862/VBIAS pixel_5862/NB2 pixel_5862/AMP_IN pixel_5862/SF_IB
+ pixel_5862/PIX_OUT pixel_5862/CSA_VREF pixel
Xpixel_5873 pixel_5873/gring pixel_5873/VDD pixel_5873/GND pixel_5873/VREF pixel_5873/ROW_SEL
+ pixel_5873/NB1 pixel_5873/VBIAS pixel_5873/NB2 pixel_5873/AMP_IN pixel_5873/SF_IB
+ pixel_5873/PIX_OUT pixel_5873/CSA_VREF pixel
Xpixel_5884 pixel_5884/gring pixel_5884/VDD pixel_5884/GND pixel_5884/VREF pixel_5884/ROW_SEL
+ pixel_5884/NB1 pixel_5884/VBIAS pixel_5884/NB2 pixel_5884/AMP_IN pixel_5884/SF_IB
+ pixel_5884/PIX_OUT pixel_5884/CSA_VREF pixel
Xpixel_5895 pixel_5895/gring pixel_5895/VDD pixel_5895/GND pixel_5895/VREF pixel_5895/ROW_SEL
+ pixel_5895/NB1 pixel_5895/VBIAS pixel_5895/NB2 pixel_5895/AMP_IN pixel_5895/SF_IB
+ pixel_5895/PIX_OUT pixel_5895/CSA_VREF pixel
Xpixel_1809 pixel_1809/gring pixel_1809/VDD pixel_1809/GND pixel_1809/VREF pixel_1809/ROW_SEL
+ pixel_1809/NB1 pixel_1809/VBIAS pixel_1809/NB2 pixel_1809/AMP_IN pixel_1809/SF_IB
+ pixel_1809/PIX_OUT pixel_1809/CSA_VREF pixel
Xpixel_5103 pixel_5103/gring pixel_5103/VDD pixel_5103/GND pixel_5103/VREF pixel_5103/ROW_SEL
+ pixel_5103/NB1 pixel_5103/VBIAS pixel_5103/NB2 pixel_5103/AMP_IN pixel_5103/SF_IB
+ pixel_5103/PIX_OUT pixel_5103/CSA_VREF pixel
Xpixel_5114 pixel_5114/gring pixel_5114/VDD pixel_5114/GND pixel_5114/VREF pixel_5114/ROW_SEL
+ pixel_5114/NB1 pixel_5114/VBIAS pixel_5114/NB2 pixel_5114/AMP_IN pixel_5114/SF_IB
+ pixel_5114/PIX_OUT pixel_5114/CSA_VREF pixel
Xpixel_5125 pixel_5125/gring pixel_5125/VDD pixel_5125/GND pixel_5125/VREF pixel_5125/ROW_SEL
+ pixel_5125/NB1 pixel_5125/VBIAS pixel_5125/NB2 pixel_5125/AMP_IN pixel_5125/SF_IB
+ pixel_5125/PIX_OUT pixel_5125/CSA_VREF pixel
Xpixel_5136 pixel_5136/gring pixel_5136/VDD pixel_5136/GND pixel_5136/VREF pixel_5136/ROW_SEL
+ pixel_5136/NB1 pixel_5136/VBIAS pixel_5136/NB2 pixel_5136/AMP_IN pixel_5136/SF_IB
+ pixel_5136/PIX_OUT pixel_5136/CSA_VREF pixel
Xpixel_5147 pixel_5147/gring pixel_5147/VDD pixel_5147/GND pixel_5147/VREF pixel_5147/ROW_SEL
+ pixel_5147/NB1 pixel_5147/VBIAS pixel_5147/NB2 pixel_5147/AMP_IN pixel_5147/SF_IB
+ pixel_5147/PIX_OUT pixel_5147/CSA_VREF pixel
Xpixel_4402 pixel_4402/gring pixel_4402/VDD pixel_4402/GND pixel_4402/VREF pixel_4402/ROW_SEL
+ pixel_4402/NB1 pixel_4402/VBIAS pixel_4402/NB2 pixel_4402/AMP_IN pixel_4402/SF_IB
+ pixel_4402/PIX_OUT pixel_4402/CSA_VREF pixel
Xpixel_441 pixel_441/gring pixel_441/VDD pixel_441/GND pixel_441/VREF pixel_441/ROW_SEL
+ pixel_441/NB1 pixel_441/VBIAS pixel_441/NB2 pixel_441/AMP_IN pixel_441/SF_IB pixel_441/PIX_OUT
+ pixel_441/CSA_VREF pixel
Xpixel_430 pixel_430/gring pixel_430/VDD pixel_430/GND pixel_430/VREF pixel_430/ROW_SEL
+ pixel_430/NB1 pixel_430/VBIAS pixel_430/NB2 pixel_430/AMP_IN pixel_430/SF_IB pixel_430/PIX_OUT
+ pixel_430/CSA_VREF pixel
Xpixel_3701 pixel_3701/gring pixel_3701/VDD pixel_3701/GND pixel_3701/VREF pixel_3701/ROW_SEL
+ pixel_3701/NB1 pixel_3701/VBIAS pixel_3701/NB2 pixel_3701/AMP_IN pixel_3701/SF_IB
+ pixel_3701/PIX_OUT pixel_3701/CSA_VREF pixel
Xpixel_5158 pixel_5158/gring pixel_5158/VDD pixel_5158/GND pixel_5158/VREF pixel_5158/ROW_SEL
+ pixel_5158/NB1 pixel_5158/VBIAS pixel_5158/NB2 pixel_5158/AMP_IN pixel_5158/SF_IB
+ pixel_5158/PIX_OUT pixel_5158/CSA_VREF pixel
Xpixel_5169 pixel_5169/gring pixel_5169/VDD pixel_5169/GND pixel_5169/VREF pixel_5169/ROW_SEL
+ pixel_5169/NB1 pixel_5169/VBIAS pixel_5169/NB2 pixel_5169/AMP_IN pixel_5169/SF_IB
+ pixel_5169/PIX_OUT pixel_5169/CSA_VREF pixel
Xpixel_4413 pixel_4413/gring pixel_4413/VDD pixel_4413/GND pixel_4413/VREF pixel_4413/ROW_SEL
+ pixel_4413/NB1 pixel_4413/VBIAS pixel_4413/NB2 pixel_4413/AMP_IN pixel_4413/SF_IB
+ pixel_4413/PIX_OUT pixel_4413/CSA_VREF pixel
Xpixel_4424 pixel_4424/gring pixel_4424/VDD pixel_4424/GND pixel_4424/VREF pixel_4424/ROW_SEL
+ pixel_4424/NB1 pixel_4424/VBIAS pixel_4424/NB2 pixel_4424/AMP_IN pixel_4424/SF_IB
+ pixel_4424/PIX_OUT pixel_4424/CSA_VREF pixel
Xpixel_4435 pixel_4435/gring pixel_4435/VDD pixel_4435/GND pixel_4435/VREF pixel_4435/ROW_SEL
+ pixel_4435/NB1 pixel_4435/VBIAS pixel_4435/NB2 pixel_4435/AMP_IN pixel_4435/SF_IB
+ pixel_4435/PIX_OUT pixel_4435/CSA_VREF pixel
Xpixel_474 pixel_474/gring pixel_474/VDD pixel_474/GND pixel_474/VREF pixel_474/ROW_SEL
+ pixel_474/NB1 pixel_474/VBIAS pixel_474/NB2 pixel_474/AMP_IN pixel_474/SF_IB pixel_474/PIX_OUT
+ pixel_474/CSA_VREF pixel
Xpixel_463 pixel_463/gring pixel_463/VDD pixel_463/GND pixel_463/VREF pixel_463/ROW_SEL
+ pixel_463/NB1 pixel_463/VBIAS pixel_463/NB2 pixel_463/AMP_IN pixel_463/SF_IB pixel_463/PIX_OUT
+ pixel_463/CSA_VREF pixel
Xpixel_452 pixel_452/gring pixel_452/VDD pixel_452/GND pixel_452/VREF pixel_452/ROW_SEL
+ pixel_452/NB1 pixel_452/VBIAS pixel_452/NB2 pixel_452/AMP_IN pixel_452/SF_IB pixel_452/PIX_OUT
+ pixel_452/CSA_VREF pixel
Xpixel_3734 pixel_3734/gring pixel_3734/VDD pixel_3734/GND pixel_3734/VREF pixel_3734/ROW_SEL
+ pixel_3734/NB1 pixel_3734/VBIAS pixel_3734/NB2 pixel_3734/AMP_IN pixel_3734/SF_IB
+ pixel_3734/PIX_OUT pixel_3734/CSA_VREF pixel
Xpixel_3723 pixel_3723/gring pixel_3723/VDD pixel_3723/GND pixel_3723/VREF pixel_3723/ROW_SEL
+ pixel_3723/NB1 pixel_3723/VBIAS pixel_3723/NB2 pixel_3723/AMP_IN pixel_3723/SF_IB
+ pixel_3723/PIX_OUT pixel_3723/CSA_VREF pixel
Xpixel_3712 pixel_3712/gring pixel_3712/VDD pixel_3712/GND pixel_3712/VREF pixel_3712/ROW_SEL
+ pixel_3712/NB1 pixel_3712/VBIAS pixel_3712/NB2 pixel_3712/AMP_IN pixel_3712/SF_IB
+ pixel_3712/PIX_OUT pixel_3712/CSA_VREF pixel
Xpixel_4446 pixel_4446/gring pixel_4446/VDD pixel_4446/GND pixel_4446/VREF pixel_4446/ROW_SEL
+ pixel_4446/NB1 pixel_4446/VBIAS pixel_4446/NB2 pixel_4446/AMP_IN pixel_4446/SF_IB
+ pixel_4446/PIX_OUT pixel_4446/CSA_VREF pixel
Xpixel_4457 pixel_4457/gring pixel_4457/VDD pixel_4457/GND pixel_4457/VREF pixel_4457/ROW_SEL
+ pixel_4457/NB1 pixel_4457/VBIAS pixel_4457/NB2 pixel_4457/AMP_IN pixel_4457/SF_IB
+ pixel_4457/PIX_OUT pixel_4457/CSA_VREF pixel
Xpixel_4468 pixel_4468/gring pixel_4468/VDD pixel_4468/GND pixel_4468/VREF pixel_4468/ROW_SEL
+ pixel_4468/NB1 pixel_4468/VBIAS pixel_4468/NB2 pixel_4468/AMP_IN pixel_4468/SF_IB
+ pixel_4468/PIX_OUT pixel_4468/CSA_VREF pixel
Xpixel_4479 pixel_4479/gring pixel_4479/VDD pixel_4479/GND pixel_4479/VREF pixel_4479/ROW_SEL
+ pixel_4479/NB1 pixel_4479/VBIAS pixel_4479/NB2 pixel_4479/AMP_IN pixel_4479/SF_IB
+ pixel_4479/PIX_OUT pixel_4479/CSA_VREF pixel
Xpixel_496 pixel_496/gring pixel_496/VDD pixel_496/GND pixel_496/VREF pixel_496/ROW_SEL
+ pixel_496/NB1 pixel_496/VBIAS pixel_496/NB2 pixel_496/AMP_IN pixel_496/SF_IB pixel_496/PIX_OUT
+ pixel_496/CSA_VREF pixel
Xpixel_485 pixel_485/gring pixel_485/VDD pixel_485/GND pixel_485/VREF pixel_485/ROW_SEL
+ pixel_485/NB1 pixel_485/VBIAS pixel_485/NB2 pixel_485/AMP_IN pixel_485/SF_IB pixel_485/PIX_OUT
+ pixel_485/CSA_VREF pixel
Xpixel_3767 pixel_3767/gring pixel_3767/VDD pixel_3767/GND pixel_3767/VREF pixel_3767/ROW_SEL
+ pixel_3767/NB1 pixel_3767/VBIAS pixel_3767/NB2 pixel_3767/AMP_IN pixel_3767/SF_IB
+ pixel_3767/PIX_OUT pixel_3767/CSA_VREF pixel
Xpixel_3756 pixel_3756/gring pixel_3756/VDD pixel_3756/GND pixel_3756/VREF pixel_3756/ROW_SEL
+ pixel_3756/NB1 pixel_3756/VBIAS pixel_3756/NB2 pixel_3756/AMP_IN pixel_3756/SF_IB
+ pixel_3756/PIX_OUT pixel_3756/CSA_VREF pixel
Xpixel_3745 pixel_3745/gring pixel_3745/VDD pixel_3745/GND pixel_3745/VREF pixel_3745/ROW_SEL
+ pixel_3745/NB1 pixel_3745/VBIAS pixel_3745/NB2 pixel_3745/AMP_IN pixel_3745/SF_IB
+ pixel_3745/PIX_OUT pixel_3745/CSA_VREF pixel
Xpixel_3789 pixel_3789/gring pixel_3789/VDD pixel_3789/GND pixel_3789/VREF pixel_3789/ROW_SEL
+ pixel_3789/NB1 pixel_3789/VBIAS pixel_3789/NB2 pixel_3789/AMP_IN pixel_3789/SF_IB
+ pixel_3789/PIX_OUT pixel_3789/CSA_VREF pixel
Xpixel_3778 pixel_3778/gring pixel_3778/VDD pixel_3778/GND pixel_3778/VREF pixel_3778/ROW_SEL
+ pixel_3778/NB1 pixel_3778/VBIAS pixel_3778/NB2 pixel_3778/AMP_IN pixel_3778/SF_IB
+ pixel_3778/PIX_OUT pixel_3778/CSA_VREF pixel
Xpixel_7050 pixel_7050/gring pixel_7050/VDD pixel_7050/GND pixel_7050/VREF pixel_7050/ROW_SEL
+ pixel_7050/NB1 pixel_7050/VBIAS pixel_7050/NB2 pixel_7050/AMP_IN pixel_7050/SF_IB
+ pixel_7050/PIX_OUT pixel_7050/CSA_VREF pixel
Xpixel_7061 pixel_7061/gring pixel_7061/VDD pixel_7061/GND pixel_7061/VREF pixel_7061/ROW_SEL
+ pixel_7061/NB1 pixel_7061/VBIAS pixel_7061/NB2 pixel_7061/AMP_IN pixel_7061/SF_IB
+ pixel_7061/PIX_OUT pixel_7061/CSA_VREF pixel
Xpixel_7072 pixel_7072/gring pixel_7072/VDD pixel_7072/GND pixel_7072/VREF pixel_7072/ROW_SEL
+ pixel_7072/NB1 pixel_7072/VBIAS pixel_7072/NB2 pixel_7072/AMP_IN pixel_7072/SF_IB
+ pixel_7072/PIX_OUT pixel_7072/CSA_VREF pixel
Xpixel_7083 pixel_7083/gring pixel_7083/VDD pixel_7083/GND pixel_7083/VREF pixel_7083/ROW_SEL
+ pixel_7083/NB1 pixel_7083/VBIAS pixel_7083/NB2 pixel_7083/AMP_IN pixel_7083/SF_IB
+ pixel_7083/PIX_OUT pixel_7083/CSA_VREF pixel
Xpixel_7094 pixel_7094/gring pixel_7094/VDD pixel_7094/GND pixel_7094/VREF pixel_7094/ROW_SEL
+ pixel_7094/NB1 pixel_7094/VBIAS pixel_7094/NB2 pixel_7094/AMP_IN pixel_7094/SF_IB
+ pixel_7094/PIX_OUT pixel_7094/CSA_VREF pixel
Xpixel_6360 pixel_6360/gring pixel_6360/VDD pixel_6360/GND pixel_6360/VREF pixel_6360/ROW_SEL
+ pixel_6360/NB1 pixel_6360/VBIAS pixel_6360/NB2 pixel_6360/AMP_IN pixel_6360/SF_IB
+ pixel_6360/PIX_OUT pixel_6360/CSA_VREF pixel
Xpixel_6371 pixel_6371/gring pixel_6371/VDD pixel_6371/GND pixel_6371/VREF pixel_6371/ROW_SEL
+ pixel_6371/NB1 pixel_6371/VBIAS pixel_6371/NB2 pixel_6371/AMP_IN pixel_6371/SF_IB
+ pixel_6371/PIX_OUT pixel_6371/CSA_VREF pixel
Xpixel_6382 pixel_6382/gring pixel_6382/VDD pixel_6382/GND pixel_6382/VREF pixel_6382/ROW_SEL
+ pixel_6382/NB1 pixel_6382/VBIAS pixel_6382/NB2 pixel_6382/AMP_IN pixel_6382/SF_IB
+ pixel_6382/PIX_OUT pixel_6382/CSA_VREF pixel
Xpixel_6393 pixel_6393/gring pixel_6393/VDD pixel_6393/GND pixel_6393/VREF pixel_6393/ROW_SEL
+ pixel_6393/NB1 pixel_6393/VBIAS pixel_6393/NB2 pixel_6393/AMP_IN pixel_6393/SF_IB
+ pixel_6393/PIX_OUT pixel_6393/CSA_VREF pixel
Xpixel_5670 pixel_5670/gring pixel_5670/VDD pixel_5670/GND pixel_5670/VREF pixel_5670/ROW_SEL
+ pixel_5670/NB1 pixel_5670/VBIAS pixel_5670/NB2 pixel_5670/AMP_IN pixel_5670/SF_IB
+ pixel_5670/PIX_OUT pixel_5670/CSA_VREF pixel
Xpixel_5681 pixel_5681/gring pixel_5681/VDD pixel_5681/GND pixel_5681/VREF pixel_5681/ROW_SEL
+ pixel_5681/NB1 pixel_5681/VBIAS pixel_5681/NB2 pixel_5681/AMP_IN pixel_5681/SF_IB
+ pixel_5681/PIX_OUT pixel_5681/CSA_VREF pixel
Xpixel_5692 pixel_5692/gring pixel_5692/VDD pixel_5692/GND pixel_5692/VREF pixel_5692/ROW_SEL
+ pixel_5692/NB1 pixel_5692/VBIAS pixel_5692/NB2 pixel_5692/AMP_IN pixel_5692/SF_IB
+ pixel_5692/PIX_OUT pixel_5692/CSA_VREF pixel
Xpixel_4980 pixel_4980/gring pixel_4980/VDD pixel_4980/GND pixel_4980/VREF pixel_4980/ROW_SEL
+ pixel_4980/NB1 pixel_4980/VBIAS pixel_4980/NB2 pixel_4980/AMP_IN pixel_4980/SF_IB
+ pixel_4980/PIX_OUT pixel_4980/CSA_VREF pixel
Xpixel_4991 pixel_4991/gring pixel_4991/VDD pixel_4991/GND pixel_4991/VREF pixel_4991/ROW_SEL
+ pixel_4991/NB1 pixel_4991/VBIAS pixel_4991/NB2 pixel_4991/AMP_IN pixel_4991/SF_IB
+ pixel_4991/PIX_OUT pixel_4991/CSA_VREF pixel
Xpixel_3019 pixel_3019/gring pixel_3019/VDD pixel_3019/GND pixel_3019/VREF pixel_3019/ROW_SEL
+ pixel_3019/NB1 pixel_3019/VBIAS pixel_3019/NB2 pixel_3019/AMP_IN pixel_3019/SF_IB
+ pixel_3019/PIX_OUT pixel_3019/CSA_VREF pixel
Xpixel_3008 pixel_3008/gring pixel_3008/VDD pixel_3008/GND pixel_3008/VREF pixel_3008/ROW_SEL
+ pixel_3008/NB1 pixel_3008/VBIAS pixel_3008/NB2 pixel_3008/AMP_IN pixel_3008/SF_IB
+ pixel_3008/PIX_OUT pixel_3008/CSA_VREF pixel
Xpixel_2318 pixel_2318/gring pixel_2318/VDD pixel_2318/GND pixel_2318/VREF pixel_2318/ROW_SEL
+ pixel_2318/NB1 pixel_2318/VBIAS pixel_2318/NB2 pixel_2318/AMP_IN pixel_2318/SF_IB
+ pixel_2318/PIX_OUT pixel_2318/CSA_VREF pixel
Xpixel_2307 pixel_2307/gring pixel_2307/VDD pixel_2307/GND pixel_2307/VREF pixel_2307/ROW_SEL
+ pixel_2307/NB1 pixel_2307/VBIAS pixel_2307/NB2 pixel_2307/AMP_IN pixel_2307/SF_IB
+ pixel_2307/PIX_OUT pixel_2307/CSA_VREF pixel
Xpixel_1606 pixel_1606/gring pixel_1606/VDD pixel_1606/GND pixel_1606/VREF pixel_1606/ROW_SEL
+ pixel_1606/NB1 pixel_1606/VBIAS pixel_1606/NB2 pixel_1606/AMP_IN pixel_1606/SF_IB
+ pixel_1606/PIX_OUT pixel_1606/CSA_VREF pixel
Xpixel_2329 pixel_2329/gring pixel_2329/VDD pixel_2329/GND pixel_2329/VREF pixel_2329/ROW_SEL
+ pixel_2329/NB1 pixel_2329/VBIAS pixel_2329/NB2 pixel_2329/AMP_IN pixel_2329/SF_IB
+ pixel_2329/PIX_OUT pixel_2329/CSA_VREF pixel
Xpixel_1639 pixel_1639/gring pixel_1639/VDD pixel_1639/GND pixel_1639/VREF pixel_1639/ROW_SEL
+ pixel_1639/NB1 pixel_1639/VBIAS pixel_1639/NB2 pixel_1639/AMP_IN pixel_1639/SF_IB
+ pixel_1639/PIX_OUT pixel_1639/CSA_VREF pixel
Xpixel_1628 pixel_1628/gring pixel_1628/VDD pixel_1628/GND pixel_1628/VREF pixel_1628/ROW_SEL
+ pixel_1628/NB1 pixel_1628/VBIAS pixel_1628/NB2 pixel_1628/AMP_IN pixel_1628/SF_IB
+ pixel_1628/PIX_OUT pixel_1628/CSA_VREF pixel
Xpixel_1617 pixel_1617/gring pixel_1617/VDD pixel_1617/GND pixel_1617/VREF pixel_1617/ROW_SEL
+ pixel_1617/NB1 pixel_1617/VBIAS pixel_1617/NB2 pixel_1617/AMP_IN pixel_1617/SF_IB
+ pixel_1617/PIX_OUT pixel_1617/CSA_VREF pixel
Xpixel_9914 pixel_9914/gring pixel_9914/VDD pixel_9914/GND pixel_9914/VREF pixel_9914/ROW_SEL
+ pixel_9914/NB1 pixel_9914/VBIAS pixel_9914/NB2 pixel_9914/AMP_IN pixel_9914/SF_IB
+ pixel_9914/PIX_OUT pixel_9914/CSA_VREF pixel
Xpixel_9903 pixel_9903/gring pixel_9903/VDD pixel_9903/GND pixel_9903/VREF pixel_9903/ROW_SEL
+ pixel_9903/NB1 pixel_9903/VBIAS pixel_9903/NB2 pixel_9903/AMP_IN pixel_9903/SF_IB
+ pixel_9903/PIX_OUT pixel_9903/CSA_VREF pixel
Xpixel_9947 pixel_9947/gring pixel_9947/VDD pixel_9947/GND pixel_9947/VREF pixel_9947/ROW_SEL
+ pixel_9947/NB1 pixel_9947/VBIAS pixel_9947/NB2 pixel_9947/AMP_IN pixel_9947/SF_IB
+ pixel_9947/PIX_OUT pixel_9947/CSA_VREF pixel
Xpixel_9936 pixel_9936/gring pixel_9936/VDD pixel_9936/GND pixel_9936/VREF pixel_9936/ROW_SEL
+ pixel_9936/NB1 pixel_9936/VBIAS pixel_9936/NB2 pixel_9936/AMP_IN pixel_9936/SF_IB
+ pixel_9936/PIX_OUT pixel_9936/CSA_VREF pixel
Xpixel_9925 pixel_9925/gring pixel_9925/VDD pixel_9925/GND pixel_9925/VREF pixel_9925/ROW_SEL
+ pixel_9925/NB1 pixel_9925/VBIAS pixel_9925/NB2 pixel_9925/AMP_IN pixel_9925/SF_IB
+ pixel_9925/PIX_OUT pixel_9925/CSA_VREF pixel
Xpixel_9958 pixel_9958/gring pixel_9958/VDD pixel_9958/GND pixel_9958/VREF pixel_9958/ROW_SEL
+ pixel_9958/NB1 pixel_9958/VBIAS pixel_9958/NB2 pixel_9958/AMP_IN pixel_9958/SF_IB
+ pixel_9958/PIX_OUT pixel_9958/CSA_VREF pixel
Xpixel_9969 pixel_9969/gring pixel_9969/VDD pixel_9969/GND pixel_9969/VREF pixel_9969/ROW_SEL
+ pixel_9969/NB1 pixel_9969/VBIAS pixel_9969/NB2 pixel_9969/AMP_IN pixel_9969/SF_IB
+ pixel_9969/PIX_OUT pixel_9969/CSA_VREF pixel
Xpixel_4210 pixel_4210/gring pixel_4210/VDD pixel_4210/GND pixel_4210/VREF pixel_4210/ROW_SEL
+ pixel_4210/NB1 pixel_4210/VBIAS pixel_4210/NB2 pixel_4210/AMP_IN pixel_4210/SF_IB
+ pixel_4210/PIX_OUT pixel_4210/CSA_VREF pixel
Xpixel_4221 pixel_4221/gring pixel_4221/VDD pixel_4221/GND pixel_4221/VREF pixel_4221/ROW_SEL
+ pixel_4221/NB1 pixel_4221/VBIAS pixel_4221/NB2 pixel_4221/AMP_IN pixel_4221/SF_IB
+ pixel_4221/PIX_OUT pixel_4221/CSA_VREF pixel
Xpixel_4232 pixel_4232/gring pixel_4232/VDD pixel_4232/GND pixel_4232/VREF pixel_4232/ROW_SEL
+ pixel_4232/NB1 pixel_4232/VBIAS pixel_4232/NB2 pixel_4232/AMP_IN pixel_4232/SF_IB
+ pixel_4232/PIX_OUT pixel_4232/CSA_VREF pixel
Xpixel_4243 pixel_4243/gring pixel_4243/VDD pixel_4243/GND pixel_4243/VREF pixel_4243/ROW_SEL
+ pixel_4243/NB1 pixel_4243/VBIAS pixel_4243/NB2 pixel_4243/AMP_IN pixel_4243/SF_IB
+ pixel_4243/PIX_OUT pixel_4243/CSA_VREF pixel
Xpixel_4254 pixel_4254/gring pixel_4254/VDD pixel_4254/GND pixel_4254/VREF pixel_4254/ROW_SEL
+ pixel_4254/NB1 pixel_4254/VBIAS pixel_4254/NB2 pixel_4254/AMP_IN pixel_4254/SF_IB
+ pixel_4254/PIX_OUT pixel_4254/CSA_VREF pixel
Xpixel_282 pixel_282/gring pixel_282/VDD pixel_282/GND pixel_282/VREF pixel_282/ROW_SEL
+ pixel_282/NB1 pixel_282/VBIAS pixel_282/NB2 pixel_282/AMP_IN pixel_282/SF_IB pixel_282/PIX_OUT
+ pixel_282/CSA_VREF pixel
Xpixel_271 pixel_271/gring pixel_271/VDD pixel_271/GND pixel_271/VREF pixel_271/ROW_SEL
+ pixel_271/NB1 pixel_271/VBIAS pixel_271/NB2 pixel_271/AMP_IN pixel_271/SF_IB pixel_271/PIX_OUT
+ pixel_271/CSA_VREF pixel
Xpixel_260 pixel_260/gring pixel_260/VDD pixel_260/GND pixel_260/VREF pixel_260/ROW_SEL
+ pixel_260/NB1 pixel_260/VBIAS pixel_260/NB2 pixel_260/AMP_IN pixel_260/SF_IB pixel_260/PIX_OUT
+ pixel_260/CSA_VREF pixel
Xpixel_3542 pixel_3542/gring pixel_3542/VDD pixel_3542/GND pixel_3542/VREF pixel_3542/ROW_SEL
+ pixel_3542/NB1 pixel_3542/VBIAS pixel_3542/NB2 pixel_3542/AMP_IN pixel_3542/SF_IB
+ pixel_3542/PIX_OUT pixel_3542/CSA_VREF pixel
Xpixel_3531 pixel_3531/gring pixel_3531/VDD pixel_3531/GND pixel_3531/VREF pixel_3531/ROW_SEL
+ pixel_3531/NB1 pixel_3531/VBIAS pixel_3531/NB2 pixel_3531/AMP_IN pixel_3531/SF_IB
+ pixel_3531/PIX_OUT pixel_3531/CSA_VREF pixel
Xpixel_3520 pixel_3520/gring pixel_3520/VDD pixel_3520/GND pixel_3520/VREF pixel_3520/ROW_SEL
+ pixel_3520/NB1 pixel_3520/VBIAS pixel_3520/NB2 pixel_3520/AMP_IN pixel_3520/SF_IB
+ pixel_3520/PIX_OUT pixel_3520/CSA_VREF pixel
Xpixel_4265 pixel_4265/gring pixel_4265/VDD pixel_4265/GND pixel_4265/VREF pixel_4265/ROW_SEL
+ pixel_4265/NB1 pixel_4265/VBIAS pixel_4265/NB2 pixel_4265/AMP_IN pixel_4265/SF_IB
+ pixel_4265/PIX_OUT pixel_4265/CSA_VREF pixel
Xpixel_4276 pixel_4276/gring pixel_4276/VDD pixel_4276/GND pixel_4276/VREF pixel_4276/ROW_SEL
+ pixel_4276/NB1 pixel_4276/VBIAS pixel_4276/NB2 pixel_4276/AMP_IN pixel_4276/SF_IB
+ pixel_4276/PIX_OUT pixel_4276/CSA_VREF pixel
Xpixel_4287 pixel_4287/gring pixel_4287/VDD pixel_4287/GND pixel_4287/VREF pixel_4287/ROW_SEL
+ pixel_4287/NB1 pixel_4287/VBIAS pixel_4287/NB2 pixel_4287/AMP_IN pixel_4287/SF_IB
+ pixel_4287/PIX_OUT pixel_4287/CSA_VREF pixel
Xpixel_293 pixel_293/gring pixel_293/VDD pixel_293/GND pixel_293/VREF pixel_293/ROW_SEL
+ pixel_293/NB1 pixel_293/VBIAS pixel_293/NB2 pixel_293/AMP_IN pixel_293/SF_IB pixel_293/PIX_OUT
+ pixel_293/CSA_VREF pixel
Xpixel_2841 pixel_2841/gring pixel_2841/VDD pixel_2841/GND pixel_2841/VREF pixel_2841/ROW_SEL
+ pixel_2841/NB1 pixel_2841/VBIAS pixel_2841/NB2 pixel_2841/AMP_IN pixel_2841/SF_IB
+ pixel_2841/PIX_OUT pixel_2841/CSA_VREF pixel
Xpixel_2830 pixel_2830/gring pixel_2830/VDD pixel_2830/GND pixel_2830/VREF pixel_2830/ROW_SEL
+ pixel_2830/NB1 pixel_2830/VBIAS pixel_2830/NB2 pixel_2830/AMP_IN pixel_2830/SF_IB
+ pixel_2830/PIX_OUT pixel_2830/CSA_VREF pixel
Xpixel_3575 pixel_3575/gring pixel_3575/VDD pixel_3575/GND pixel_3575/VREF pixel_3575/ROW_SEL
+ pixel_3575/NB1 pixel_3575/VBIAS pixel_3575/NB2 pixel_3575/AMP_IN pixel_3575/SF_IB
+ pixel_3575/PIX_OUT pixel_3575/CSA_VREF pixel
Xpixel_3564 pixel_3564/gring pixel_3564/VDD pixel_3564/GND pixel_3564/VREF pixel_3564/ROW_SEL
+ pixel_3564/NB1 pixel_3564/VBIAS pixel_3564/NB2 pixel_3564/AMP_IN pixel_3564/SF_IB
+ pixel_3564/PIX_OUT pixel_3564/CSA_VREF pixel
Xpixel_3553 pixel_3553/gring pixel_3553/VDD pixel_3553/GND pixel_3553/VREF pixel_3553/ROW_SEL
+ pixel_3553/NB1 pixel_3553/VBIAS pixel_3553/NB2 pixel_3553/AMP_IN pixel_3553/SF_IB
+ pixel_3553/PIX_OUT pixel_3553/CSA_VREF pixel
Xpixel_4298 pixel_4298/gring pixel_4298/VDD pixel_4298/GND pixel_4298/VREF pixel_4298/ROW_SEL
+ pixel_4298/NB1 pixel_4298/VBIAS pixel_4298/NB2 pixel_4298/AMP_IN pixel_4298/SF_IB
+ pixel_4298/PIX_OUT pixel_4298/CSA_VREF pixel
Xpixel_2874 pixel_2874/gring pixel_2874/VDD pixel_2874/GND pixel_2874/VREF pixel_2874/ROW_SEL
+ pixel_2874/NB1 pixel_2874/VBIAS pixel_2874/NB2 pixel_2874/AMP_IN pixel_2874/SF_IB
+ pixel_2874/PIX_OUT pixel_2874/CSA_VREF pixel
Xpixel_2863 pixel_2863/gring pixel_2863/VDD pixel_2863/GND pixel_2863/VREF pixel_2863/ROW_SEL
+ pixel_2863/NB1 pixel_2863/VBIAS pixel_2863/NB2 pixel_2863/AMP_IN pixel_2863/SF_IB
+ pixel_2863/PIX_OUT pixel_2863/CSA_VREF pixel
Xpixel_2852 pixel_2852/gring pixel_2852/VDD pixel_2852/GND pixel_2852/VREF pixel_2852/ROW_SEL
+ pixel_2852/NB1 pixel_2852/VBIAS pixel_2852/NB2 pixel_2852/AMP_IN pixel_2852/SF_IB
+ pixel_2852/PIX_OUT pixel_2852/CSA_VREF pixel
Xpixel_3597 pixel_3597/gring pixel_3597/VDD pixel_3597/GND pixel_3597/VREF pixel_3597/ROW_SEL
+ pixel_3597/NB1 pixel_3597/VBIAS pixel_3597/NB2 pixel_3597/AMP_IN pixel_3597/SF_IB
+ pixel_3597/PIX_OUT pixel_3597/CSA_VREF pixel
Xpixel_3586 pixel_3586/gring pixel_3586/VDD pixel_3586/GND pixel_3586/VREF pixel_3586/ROW_SEL
+ pixel_3586/NB1 pixel_3586/VBIAS pixel_3586/NB2 pixel_3586/AMP_IN pixel_3586/SF_IB
+ pixel_3586/PIX_OUT pixel_3586/CSA_VREF pixel
Xpixel_2896 pixel_2896/gring pixel_2896/VDD pixel_2896/GND pixel_2896/VREF pixel_2896/ROW_SEL
+ pixel_2896/NB1 pixel_2896/VBIAS pixel_2896/NB2 pixel_2896/AMP_IN pixel_2896/SF_IB
+ pixel_2896/PIX_OUT pixel_2896/CSA_VREF pixel
Xpixel_2885 pixel_2885/gring pixel_2885/VDD pixel_2885/GND pixel_2885/VREF pixel_2885/ROW_SEL
+ pixel_2885/NB1 pixel_2885/VBIAS pixel_2885/NB2 pixel_2885/AMP_IN pixel_2885/SF_IB
+ pixel_2885/PIX_OUT pixel_2885/CSA_VREF pixel
Xpixel_6190 pixel_6190/gring pixel_6190/VDD pixel_6190/GND pixel_6190/VREF pixel_6190/ROW_SEL
+ pixel_6190/NB1 pixel_6190/VBIAS pixel_6190/NB2 pixel_6190/AMP_IN pixel_6190/SF_IB
+ pixel_6190/PIX_OUT pixel_6190/CSA_VREF pixel
Xpixel_8509 pixel_8509/gring pixel_8509/VDD pixel_8509/GND pixel_8509/VREF pixel_8509/ROW_SEL
+ pixel_8509/NB1 pixel_8509/VBIAS pixel_8509/NB2 pixel_8509/AMP_IN pixel_8509/SF_IB
+ pixel_8509/PIX_OUT pixel_8509/CSA_VREF pixel
Xpixel_7808 pixel_7808/gring pixel_7808/VDD pixel_7808/GND pixel_7808/VREF pixel_7808/ROW_SEL
+ pixel_7808/NB1 pixel_7808/VBIAS pixel_7808/NB2 pixel_7808/AMP_IN pixel_7808/SF_IB
+ pixel_7808/PIX_OUT pixel_7808/CSA_VREF pixel
Xpixel_7819 pixel_7819/gring pixel_7819/VDD pixel_7819/GND pixel_7819/VREF pixel_7819/ROW_SEL
+ pixel_7819/NB1 pixel_7819/VBIAS pixel_7819/NB2 pixel_7819/AMP_IN pixel_7819/SF_IB
+ pixel_7819/PIX_OUT pixel_7819/CSA_VREF pixel
Xpixel_2126 pixel_2126/gring pixel_2126/VDD pixel_2126/GND pixel_2126/VREF pixel_2126/ROW_SEL
+ pixel_2126/NB1 pixel_2126/VBIAS pixel_2126/NB2 pixel_2126/AMP_IN pixel_2126/SF_IB
+ pixel_2126/PIX_OUT pixel_2126/CSA_VREF pixel
Xpixel_2115 pixel_2115/gring pixel_2115/VDD pixel_2115/GND pixel_2115/VREF pixel_2115/ROW_SEL
+ pixel_2115/NB1 pixel_2115/VBIAS pixel_2115/NB2 pixel_2115/AMP_IN pixel_2115/SF_IB
+ pixel_2115/PIX_OUT pixel_2115/CSA_VREF pixel
Xpixel_2104 pixel_2104/gring pixel_2104/VDD pixel_2104/GND pixel_2104/VREF pixel_2104/ROW_SEL
+ pixel_2104/NB1 pixel_2104/VBIAS pixel_2104/NB2 pixel_2104/AMP_IN pixel_2104/SF_IB
+ pixel_2104/PIX_OUT pixel_2104/CSA_VREF pixel
Xpixel_1425 pixel_1425/gring pixel_1425/VDD pixel_1425/GND pixel_1425/VREF pixel_1425/ROW_SEL
+ pixel_1425/NB1 pixel_1425/VBIAS pixel_1425/NB2 pixel_1425/AMP_IN pixel_1425/SF_IB
+ pixel_1425/PIX_OUT pixel_1425/CSA_VREF pixel
Xpixel_1414 pixel_1414/gring pixel_1414/VDD pixel_1414/GND pixel_1414/VREF pixel_1414/ROW_SEL
+ pixel_1414/NB1 pixel_1414/VBIAS pixel_1414/NB2 pixel_1414/AMP_IN pixel_1414/SF_IB
+ pixel_1414/PIX_OUT pixel_1414/CSA_VREF pixel
Xpixel_1403 pixel_1403/gring pixel_1403/VDD pixel_1403/GND pixel_1403/VREF pixel_1403/ROW_SEL
+ pixel_1403/NB1 pixel_1403/VBIAS pixel_1403/NB2 pixel_1403/AMP_IN pixel_1403/SF_IB
+ pixel_1403/PIX_OUT pixel_1403/CSA_VREF pixel
Xpixel_2159 pixel_2159/gring pixel_2159/VDD pixel_2159/GND pixel_2159/VREF pixel_2159/ROW_SEL
+ pixel_2159/NB1 pixel_2159/VBIAS pixel_2159/NB2 pixel_2159/AMP_IN pixel_2159/SF_IB
+ pixel_2159/PIX_OUT pixel_2159/CSA_VREF pixel
Xpixel_2148 pixel_2148/gring pixel_2148/VDD pixel_2148/GND pixel_2148/VREF pixel_2148/ROW_SEL
+ pixel_2148/NB1 pixel_2148/VBIAS pixel_2148/NB2 pixel_2148/AMP_IN pixel_2148/SF_IB
+ pixel_2148/PIX_OUT pixel_2148/CSA_VREF pixel
Xpixel_2137 pixel_2137/gring pixel_2137/VDD pixel_2137/GND pixel_2137/VREF pixel_2137/ROW_SEL
+ pixel_2137/NB1 pixel_2137/VBIAS pixel_2137/NB2 pixel_2137/AMP_IN pixel_2137/SF_IB
+ pixel_2137/PIX_OUT pixel_2137/CSA_VREF pixel
Xpixel_1458 pixel_1458/gring pixel_1458/VDD pixel_1458/GND pixel_1458/VREF pixel_1458/ROW_SEL
+ pixel_1458/NB1 pixel_1458/VBIAS pixel_1458/NB2 pixel_1458/AMP_IN pixel_1458/SF_IB
+ pixel_1458/PIX_OUT pixel_1458/CSA_VREF pixel
Xpixel_1447 pixel_1447/gring pixel_1447/VDD pixel_1447/GND pixel_1447/VREF pixel_1447/ROW_SEL
+ pixel_1447/NB1 pixel_1447/VBIAS pixel_1447/NB2 pixel_1447/AMP_IN pixel_1447/SF_IB
+ pixel_1447/PIX_OUT pixel_1447/CSA_VREF pixel
Xpixel_1436 pixel_1436/gring pixel_1436/VDD pixel_1436/GND pixel_1436/VREF pixel_1436/ROW_SEL
+ pixel_1436/NB1 pixel_1436/VBIAS pixel_1436/NB2 pixel_1436/AMP_IN pixel_1436/SF_IB
+ pixel_1436/PIX_OUT pixel_1436/CSA_VREF pixel
Xpixel_1469 pixel_1469/gring pixel_1469/VDD pixel_1469/GND pixel_1469/VREF pixel_1469/ROW_SEL
+ pixel_1469/NB1 pixel_1469/VBIAS pixel_1469/NB2 pixel_1469/AMP_IN pixel_1469/SF_IB
+ pixel_1469/PIX_OUT pixel_1469/CSA_VREF pixel
Xpixel_9700 pixel_9700/gring pixel_9700/VDD pixel_9700/GND pixel_9700/VREF pixel_9700/ROW_SEL
+ pixel_9700/NB1 pixel_9700/VBIAS pixel_9700/NB2 pixel_9700/AMP_IN pixel_9700/SF_IB
+ pixel_9700/PIX_OUT pixel_9700/CSA_VREF pixel
Xpixel_9711 pixel_9711/gring pixel_9711/VDD pixel_9711/GND pixel_9711/VREF pixel_9711/ROW_SEL
+ pixel_9711/NB1 pixel_9711/VBIAS pixel_9711/NB2 pixel_9711/AMP_IN pixel_9711/SF_IB
+ pixel_9711/PIX_OUT pixel_9711/CSA_VREF pixel
Xpixel_9722 pixel_9722/gring pixel_9722/VDD pixel_9722/GND pixel_9722/VREF pixel_9722/ROW_SEL
+ pixel_9722/NB1 pixel_9722/VBIAS pixel_9722/NB2 pixel_9722/AMP_IN pixel_9722/SF_IB
+ pixel_9722/PIX_OUT pixel_9722/CSA_VREF pixel
Xpixel_9733 pixel_9733/gring pixel_9733/VDD pixel_9733/GND pixel_9733/VREF pixel_9733/ROW_SEL
+ pixel_9733/NB1 pixel_9733/VBIAS pixel_9733/NB2 pixel_9733/AMP_IN pixel_9733/SF_IB
+ pixel_9733/PIX_OUT pixel_9733/CSA_VREF pixel
Xpixel_9744 pixel_9744/gring pixel_9744/VDD pixel_9744/GND pixel_9744/VREF pixel_9744/ROW_SEL
+ pixel_9744/NB1 pixel_9744/VBIAS pixel_9744/NB2 pixel_9744/AMP_IN pixel_9744/SF_IB
+ pixel_9744/PIX_OUT pixel_9744/CSA_VREF pixel
Xpixel_9755 pixel_9755/gring pixel_9755/VDD pixel_9755/GND pixel_9755/VREF pixel_9755/ROW_SEL
+ pixel_9755/NB1 pixel_9755/VBIAS pixel_9755/NB2 pixel_9755/AMP_IN pixel_9755/SF_IB
+ pixel_9755/PIX_OUT pixel_9755/CSA_VREF pixel
Xpixel_9766 pixel_9766/gring pixel_9766/VDD pixel_9766/GND pixel_9766/VREF pixel_9766/ROW_SEL
+ pixel_9766/NB1 pixel_9766/VBIAS pixel_9766/NB2 pixel_9766/AMP_IN pixel_9766/SF_IB
+ pixel_9766/PIX_OUT pixel_9766/CSA_VREF pixel
Xpixel_9777 pixel_9777/gring pixel_9777/VDD pixel_9777/GND pixel_9777/VREF pixel_9777/ROW_SEL
+ pixel_9777/NB1 pixel_9777/VBIAS pixel_9777/NB2 pixel_9777/AMP_IN pixel_9777/SF_IB
+ pixel_9777/PIX_OUT pixel_9777/CSA_VREF pixel
Xpixel_9788 pixel_9788/gring pixel_9788/VDD pixel_9788/GND pixel_9788/VREF pixel_9788/ROW_SEL
+ pixel_9788/NB1 pixel_9788/VBIAS pixel_9788/NB2 pixel_9788/AMP_IN pixel_9788/SF_IB
+ pixel_9788/PIX_OUT pixel_9788/CSA_VREF pixel
Xpixel_9799 pixel_9799/gring pixel_9799/VDD pixel_9799/GND pixel_9799/VREF pixel_9799/ROW_SEL
+ pixel_9799/NB1 pixel_9799/VBIAS pixel_9799/NB2 pixel_9799/AMP_IN pixel_9799/SF_IB
+ pixel_9799/PIX_OUT pixel_9799/CSA_VREF pixel
Xpixel_4040 pixel_4040/gring pixel_4040/VDD pixel_4040/GND pixel_4040/VREF pixel_4040/ROW_SEL
+ pixel_4040/NB1 pixel_4040/VBIAS pixel_4040/NB2 pixel_4040/AMP_IN pixel_4040/SF_IB
+ pixel_4040/PIX_OUT pixel_4040/CSA_VREF pixel
Xpixel_4051 pixel_4051/gring pixel_4051/VDD pixel_4051/GND pixel_4051/VREF pixel_4051/ROW_SEL
+ pixel_4051/NB1 pixel_4051/VBIAS pixel_4051/NB2 pixel_4051/AMP_IN pixel_4051/SF_IB
+ pixel_4051/PIX_OUT pixel_4051/CSA_VREF pixel
Xpixel_4062 pixel_4062/gring pixel_4062/VDD pixel_4062/GND pixel_4062/VREF pixel_4062/ROW_SEL
+ pixel_4062/NB1 pixel_4062/VBIAS pixel_4062/NB2 pixel_4062/AMP_IN pixel_4062/SF_IB
+ pixel_4062/PIX_OUT pixel_4062/CSA_VREF pixel
Xpixel_3350 pixel_3350/gring pixel_3350/VDD pixel_3350/GND pixel_3350/VREF pixel_3350/ROW_SEL
+ pixel_3350/NB1 pixel_3350/VBIAS pixel_3350/NB2 pixel_3350/AMP_IN pixel_3350/SF_IB
+ pixel_3350/PIX_OUT pixel_3350/CSA_VREF pixel
Xpixel_4073 pixel_4073/gring pixel_4073/VDD pixel_4073/GND pixel_4073/VREF pixel_4073/ROW_SEL
+ pixel_4073/NB1 pixel_4073/VBIAS pixel_4073/NB2 pixel_4073/AMP_IN pixel_4073/SF_IB
+ pixel_4073/PIX_OUT pixel_4073/CSA_VREF pixel
Xpixel_4084 pixel_4084/gring pixel_4084/VDD pixel_4084/GND pixel_4084/VREF pixel_4084/ROW_SEL
+ pixel_4084/NB1 pixel_4084/VBIAS pixel_4084/NB2 pixel_4084/AMP_IN pixel_4084/SF_IB
+ pixel_4084/PIX_OUT pixel_4084/CSA_VREF pixel
Xpixel_4095 pixel_4095/gring pixel_4095/VDD pixel_4095/GND pixel_4095/VREF pixel_4095/ROW_SEL
+ pixel_4095/NB1 pixel_4095/VBIAS pixel_4095/NB2 pixel_4095/AMP_IN pixel_4095/SF_IB
+ pixel_4095/PIX_OUT pixel_4095/CSA_VREF pixel
Xpixel_3394 pixel_3394/gring pixel_3394/VDD pixel_3394/GND pixel_3394/VREF pixel_3394/ROW_SEL
+ pixel_3394/NB1 pixel_3394/VBIAS pixel_3394/NB2 pixel_3394/AMP_IN pixel_3394/SF_IB
+ pixel_3394/PIX_OUT pixel_3394/CSA_VREF pixel
Xpixel_3383 pixel_3383/gring pixel_3383/VDD pixel_3383/GND pixel_3383/VREF pixel_3383/ROW_SEL
+ pixel_3383/NB1 pixel_3383/VBIAS pixel_3383/NB2 pixel_3383/AMP_IN pixel_3383/SF_IB
+ pixel_3383/PIX_OUT pixel_3383/CSA_VREF pixel
Xpixel_3372 pixel_3372/gring pixel_3372/VDD pixel_3372/GND pixel_3372/VREF pixel_3372/ROW_SEL
+ pixel_3372/NB1 pixel_3372/VBIAS pixel_3372/NB2 pixel_3372/AMP_IN pixel_3372/SF_IB
+ pixel_3372/PIX_OUT pixel_3372/CSA_VREF pixel
Xpixel_3361 pixel_3361/gring pixel_3361/VDD pixel_3361/GND pixel_3361/VREF pixel_3361/ROW_SEL
+ pixel_3361/NB1 pixel_3361/VBIAS pixel_3361/NB2 pixel_3361/AMP_IN pixel_3361/SF_IB
+ pixel_3361/PIX_OUT pixel_3361/CSA_VREF pixel
Xpixel_2682 pixel_2682/gring pixel_2682/VDD pixel_2682/GND pixel_2682/VREF pixel_2682/ROW_SEL
+ pixel_2682/NB1 pixel_2682/VBIAS pixel_2682/NB2 pixel_2682/AMP_IN pixel_2682/SF_IB
+ pixel_2682/PIX_OUT pixel_2682/CSA_VREF pixel
Xpixel_2671 pixel_2671/gring pixel_2671/VDD pixel_2671/GND pixel_2671/VREF pixel_2671/ROW_SEL
+ pixel_2671/NB1 pixel_2671/VBIAS pixel_2671/NB2 pixel_2671/AMP_IN pixel_2671/SF_IB
+ pixel_2671/PIX_OUT pixel_2671/CSA_VREF pixel
Xpixel_2660 pixel_2660/gring pixel_2660/VDD pixel_2660/GND pixel_2660/VREF pixel_2660/ROW_SEL
+ pixel_2660/NB1 pixel_2660/VBIAS pixel_2660/NB2 pixel_2660/AMP_IN pixel_2660/SF_IB
+ pixel_2660/PIX_OUT pixel_2660/CSA_VREF pixel
Xpixel_1970 pixel_1970/gring pixel_1970/VDD pixel_1970/GND pixel_1970/VREF pixel_1970/ROW_SEL
+ pixel_1970/NB1 pixel_1970/VBIAS pixel_1970/NB2 pixel_1970/AMP_IN pixel_1970/SF_IB
+ pixel_1970/PIX_OUT pixel_1970/CSA_VREF pixel
Xpixel_2693 pixel_2693/gring pixel_2693/VDD pixel_2693/GND pixel_2693/VREF pixel_2693/ROW_SEL
+ pixel_2693/NB1 pixel_2693/VBIAS pixel_2693/NB2 pixel_2693/AMP_IN pixel_2693/SF_IB
+ pixel_2693/PIX_OUT pixel_2693/CSA_VREF pixel
Xpixel_1992 pixel_1992/gring pixel_1992/VDD pixel_1992/GND pixel_1992/VREF pixel_1992/ROW_SEL
+ pixel_1992/NB1 pixel_1992/VBIAS pixel_1992/NB2 pixel_1992/AMP_IN pixel_1992/SF_IB
+ pixel_1992/PIX_OUT pixel_1992/CSA_VREF pixel
Xpixel_1981 pixel_1981/gring pixel_1981/VDD pixel_1981/GND pixel_1981/VREF pixel_1981/ROW_SEL
+ pixel_1981/NB1 pixel_1981/VBIAS pixel_1981/NB2 pixel_1981/AMP_IN pixel_1981/SF_IB
+ pixel_1981/PIX_OUT pixel_1981/CSA_VREF pixel
Xpixel_9018 pixel_9018/gring pixel_9018/VDD pixel_9018/GND pixel_9018/VREF pixel_9018/ROW_SEL
+ pixel_9018/NB1 pixel_9018/VBIAS pixel_9018/NB2 pixel_9018/AMP_IN pixel_9018/SF_IB
+ pixel_9018/PIX_OUT pixel_9018/CSA_VREF pixel
Xpixel_9007 pixel_9007/gring pixel_9007/VDD pixel_9007/GND pixel_9007/VREF pixel_9007/ROW_SEL
+ pixel_9007/NB1 pixel_9007/VBIAS pixel_9007/NB2 pixel_9007/AMP_IN pixel_9007/SF_IB
+ pixel_9007/PIX_OUT pixel_9007/CSA_VREF pixel
Xpixel_9029 pixel_9029/gring pixel_9029/VDD pixel_9029/GND pixel_9029/VREF pixel_9029/ROW_SEL
+ pixel_9029/NB1 pixel_9029/VBIAS pixel_9029/NB2 pixel_9029/AMP_IN pixel_9029/SF_IB
+ pixel_9029/PIX_OUT pixel_9029/CSA_VREF pixel
Xpixel_8306 pixel_8306/gring pixel_8306/VDD pixel_8306/GND pixel_8306/VREF pixel_8306/ROW_SEL
+ pixel_8306/NB1 pixel_8306/VBIAS pixel_8306/NB2 pixel_8306/AMP_IN pixel_8306/SF_IB
+ pixel_8306/PIX_OUT pixel_8306/CSA_VREF pixel
Xpixel_8317 pixel_8317/gring pixel_8317/VDD pixel_8317/GND pixel_8317/VREF pixel_8317/ROW_SEL
+ pixel_8317/NB1 pixel_8317/VBIAS pixel_8317/NB2 pixel_8317/AMP_IN pixel_8317/SF_IB
+ pixel_8317/PIX_OUT pixel_8317/CSA_VREF pixel
Xpixel_8328 pixel_8328/gring pixel_8328/VDD pixel_8328/GND pixel_8328/VREF pixel_8328/ROW_SEL
+ pixel_8328/NB1 pixel_8328/VBIAS pixel_8328/NB2 pixel_8328/AMP_IN pixel_8328/SF_IB
+ pixel_8328/PIX_OUT pixel_8328/CSA_VREF pixel
Xpixel_8339 pixel_8339/gring pixel_8339/VDD pixel_8339/GND pixel_8339/VREF pixel_8339/ROW_SEL
+ pixel_8339/NB1 pixel_8339/VBIAS pixel_8339/NB2 pixel_8339/AMP_IN pixel_8339/SF_IB
+ pixel_8339/PIX_OUT pixel_8339/CSA_VREF pixel
Xpixel_7605 pixel_7605/gring pixel_7605/VDD pixel_7605/GND pixel_7605/VREF pixel_7605/ROW_SEL
+ pixel_7605/NB1 pixel_7605/VBIAS pixel_7605/NB2 pixel_7605/AMP_IN pixel_7605/SF_IB
+ pixel_7605/PIX_OUT pixel_7605/CSA_VREF pixel
Xpixel_7616 pixel_7616/gring pixel_7616/VDD pixel_7616/GND pixel_7616/VREF pixel_7616/ROW_SEL
+ pixel_7616/NB1 pixel_7616/VBIAS pixel_7616/NB2 pixel_7616/AMP_IN pixel_7616/SF_IB
+ pixel_7616/PIX_OUT pixel_7616/CSA_VREF pixel
Xpixel_7627 pixel_7627/gring pixel_7627/VDD pixel_7627/GND pixel_7627/VREF pixel_7627/ROW_SEL
+ pixel_7627/NB1 pixel_7627/VBIAS pixel_7627/NB2 pixel_7627/AMP_IN pixel_7627/SF_IB
+ pixel_7627/PIX_OUT pixel_7627/CSA_VREF pixel
Xpixel_7638 pixel_7638/gring pixel_7638/VDD pixel_7638/GND pixel_7638/VREF pixel_7638/ROW_SEL
+ pixel_7638/NB1 pixel_7638/VBIAS pixel_7638/NB2 pixel_7638/AMP_IN pixel_7638/SF_IB
+ pixel_7638/PIX_OUT pixel_7638/CSA_VREF pixel
Xpixel_6904 pixel_6904/gring pixel_6904/VDD pixel_6904/GND pixel_6904/VREF pixel_6904/ROW_SEL
+ pixel_6904/NB1 pixel_6904/VBIAS pixel_6904/NB2 pixel_6904/AMP_IN pixel_6904/SF_IB
+ pixel_6904/PIX_OUT pixel_6904/CSA_VREF pixel
Xpixel_7649 pixel_7649/gring pixel_7649/VDD pixel_7649/GND pixel_7649/VREF pixel_7649/ROW_SEL
+ pixel_7649/NB1 pixel_7649/VBIAS pixel_7649/NB2 pixel_7649/AMP_IN pixel_7649/SF_IB
+ pixel_7649/PIX_OUT pixel_7649/CSA_VREF pixel
Xpixel_6915 pixel_6915/gring pixel_6915/VDD pixel_6915/GND pixel_6915/VREF pixel_6915/ROW_SEL
+ pixel_6915/NB1 pixel_6915/VBIAS pixel_6915/NB2 pixel_6915/AMP_IN pixel_6915/SF_IB
+ pixel_6915/PIX_OUT pixel_6915/CSA_VREF pixel
Xpixel_6926 pixel_6926/gring pixel_6926/VDD pixel_6926/GND pixel_6926/VREF pixel_6926/ROW_SEL
+ pixel_6926/NB1 pixel_6926/VBIAS pixel_6926/NB2 pixel_6926/AMP_IN pixel_6926/SF_IB
+ pixel_6926/PIX_OUT pixel_6926/CSA_VREF pixel
Xpixel_6937 pixel_6937/gring pixel_6937/VDD pixel_6937/GND pixel_6937/VREF pixel_6937/ROW_SEL
+ pixel_6937/NB1 pixel_6937/VBIAS pixel_6937/NB2 pixel_6937/AMP_IN pixel_6937/SF_IB
+ pixel_6937/PIX_OUT pixel_6937/CSA_VREF pixel
Xpixel_18 pixel_18/gring pixel_18/VDD pixel_18/GND pixel_18/VREF pixel_18/ROW_SEL
+ pixel_18/NB1 pixel_18/VBIAS pixel_18/NB2 pixel_18/AMP_IN pixel_18/SF_IB pixel_18/PIX_OUT
+ pixel_18/CSA_VREF pixel
Xpixel_6948 pixel_6948/gring pixel_6948/VDD pixel_6948/GND pixel_6948/VREF pixel_6948/ROW_SEL
+ pixel_6948/NB1 pixel_6948/VBIAS pixel_6948/NB2 pixel_6948/AMP_IN pixel_6948/SF_IB
+ pixel_6948/PIX_OUT pixel_6948/CSA_VREF pixel
Xpixel_6959 pixel_6959/gring pixel_6959/VDD pixel_6959/GND pixel_6959/VREF pixel_6959/ROW_SEL
+ pixel_6959/NB1 pixel_6959/VBIAS pixel_6959/NB2 pixel_6959/AMP_IN pixel_6959/SF_IB
+ pixel_6959/PIX_OUT pixel_6959/CSA_VREF pixel
Xpixel_29 pixel_29/gring pixel_29/VDD pixel_29/GND pixel_29/VREF pixel_29/ROW_SEL
+ pixel_29/NB1 pixel_29/VBIAS pixel_29/NB2 pixel_29/AMP_IN pixel_29/SF_IB pixel_29/PIX_OUT
+ pixel_29/CSA_VREF pixel
Xpixel_1200 pixel_1200/gring pixel_1200/VDD pixel_1200/GND pixel_1200/VREF pixel_1200/ROW_SEL
+ pixel_1200/NB1 pixel_1200/VBIAS pixel_1200/NB2 pixel_1200/AMP_IN pixel_1200/SF_IB
+ pixel_1200/PIX_OUT pixel_1200/CSA_VREF pixel
Xpixel_1233 pixel_1233/gring pixel_1233/VDD pixel_1233/GND pixel_1233/VREF pixel_1233/ROW_SEL
+ pixel_1233/NB1 pixel_1233/VBIAS pixel_1233/NB2 pixel_1233/AMP_IN pixel_1233/SF_IB
+ pixel_1233/PIX_OUT pixel_1233/CSA_VREF pixel
Xpixel_1222 pixel_1222/gring pixel_1222/VDD pixel_1222/GND pixel_1222/VREF pixel_1222/ROW_SEL
+ pixel_1222/NB1 pixel_1222/VBIAS pixel_1222/NB2 pixel_1222/AMP_IN pixel_1222/SF_IB
+ pixel_1222/PIX_OUT pixel_1222/CSA_VREF pixel
Xpixel_1211 pixel_1211/gring pixel_1211/VDD pixel_1211/GND pixel_1211/VREF pixel_1211/ROW_SEL
+ pixel_1211/NB1 pixel_1211/VBIAS pixel_1211/NB2 pixel_1211/AMP_IN pixel_1211/SF_IB
+ pixel_1211/PIX_OUT pixel_1211/CSA_VREF pixel
Xpixel_1266 pixel_1266/gring pixel_1266/VDD pixel_1266/GND pixel_1266/VREF pixel_1266/ROW_SEL
+ pixel_1266/NB1 pixel_1266/VBIAS pixel_1266/NB2 pixel_1266/AMP_IN pixel_1266/SF_IB
+ pixel_1266/PIX_OUT pixel_1266/CSA_VREF pixel
Xpixel_1255 pixel_1255/gring pixel_1255/VDD pixel_1255/GND pixel_1255/VREF pixel_1255/ROW_SEL
+ pixel_1255/NB1 pixel_1255/VBIAS pixel_1255/NB2 pixel_1255/AMP_IN pixel_1255/SF_IB
+ pixel_1255/PIX_OUT pixel_1255/CSA_VREF pixel
Xpixel_1244 pixel_1244/gring pixel_1244/VDD pixel_1244/GND pixel_1244/VREF pixel_1244/ROW_SEL
+ pixel_1244/NB1 pixel_1244/VBIAS pixel_1244/NB2 pixel_1244/AMP_IN pixel_1244/SF_IB
+ pixel_1244/PIX_OUT pixel_1244/CSA_VREF pixel
Xpixel_1299 pixel_1299/gring pixel_1299/VDD pixel_1299/GND pixel_1299/VREF pixel_1299/ROW_SEL
+ pixel_1299/NB1 pixel_1299/VBIAS pixel_1299/NB2 pixel_1299/AMP_IN pixel_1299/SF_IB
+ pixel_1299/PIX_OUT pixel_1299/CSA_VREF pixel
Xpixel_1288 pixel_1288/gring pixel_1288/VDD pixel_1288/GND pixel_1288/VREF pixel_1288/ROW_SEL
+ pixel_1288/NB1 pixel_1288/VBIAS pixel_1288/NB2 pixel_1288/AMP_IN pixel_1288/SF_IB
+ pixel_1288/PIX_OUT pixel_1288/CSA_VREF pixel
Xpixel_1277 pixel_1277/gring pixel_1277/VDD pixel_1277/GND pixel_1277/VREF pixel_1277/ROW_SEL
+ pixel_1277/NB1 pixel_1277/VBIAS pixel_1277/NB2 pixel_1277/AMP_IN pixel_1277/SF_IB
+ pixel_1277/PIX_OUT pixel_1277/CSA_VREF pixel
Xpixel_9541 pixel_9541/gring pixel_9541/VDD pixel_9541/GND pixel_9541/VREF pixel_9541/ROW_SEL
+ pixel_9541/NB1 pixel_9541/VBIAS pixel_9541/NB2 pixel_9541/AMP_IN pixel_9541/SF_IB
+ pixel_9541/PIX_OUT pixel_9541/CSA_VREF pixel
Xpixel_9530 pixel_9530/gring pixel_9530/VDD pixel_9530/GND pixel_9530/VREF pixel_9530/ROW_SEL
+ pixel_9530/NB1 pixel_9530/VBIAS pixel_9530/NB2 pixel_9530/AMP_IN pixel_9530/SF_IB
+ pixel_9530/PIX_OUT pixel_9530/CSA_VREF pixel
Xpixel_9574 pixel_9574/gring pixel_9574/VDD pixel_9574/GND pixel_9574/VREF pixel_9574/ROW_SEL
+ pixel_9574/NB1 pixel_9574/VBIAS pixel_9574/NB2 pixel_9574/AMP_IN pixel_9574/SF_IB
+ pixel_9574/PIX_OUT pixel_9574/CSA_VREF pixel
Xpixel_9563 pixel_9563/gring pixel_9563/VDD pixel_9563/GND pixel_9563/VREF pixel_9563/ROW_SEL
+ pixel_9563/NB1 pixel_9563/VBIAS pixel_9563/NB2 pixel_9563/AMP_IN pixel_9563/SF_IB
+ pixel_9563/PIX_OUT pixel_9563/CSA_VREF pixel
Xpixel_9552 pixel_9552/gring pixel_9552/VDD pixel_9552/GND pixel_9552/VREF pixel_9552/ROW_SEL
+ pixel_9552/NB1 pixel_9552/VBIAS pixel_9552/NB2 pixel_9552/AMP_IN pixel_9552/SF_IB
+ pixel_9552/PIX_OUT pixel_9552/CSA_VREF pixel
Xpixel_8873 pixel_8873/gring pixel_8873/VDD pixel_8873/GND pixel_8873/VREF pixel_8873/ROW_SEL
+ pixel_8873/NB1 pixel_8873/VBIAS pixel_8873/NB2 pixel_8873/AMP_IN pixel_8873/SF_IB
+ pixel_8873/PIX_OUT pixel_8873/CSA_VREF pixel
Xpixel_8862 pixel_8862/gring pixel_8862/VDD pixel_8862/GND pixel_8862/VREF pixel_8862/ROW_SEL
+ pixel_8862/NB1 pixel_8862/VBIAS pixel_8862/NB2 pixel_8862/AMP_IN pixel_8862/SF_IB
+ pixel_8862/PIX_OUT pixel_8862/CSA_VREF pixel
Xpixel_8851 pixel_8851/gring pixel_8851/VDD pixel_8851/GND pixel_8851/VREF pixel_8851/ROW_SEL
+ pixel_8851/NB1 pixel_8851/VBIAS pixel_8851/NB2 pixel_8851/AMP_IN pixel_8851/SF_IB
+ pixel_8851/PIX_OUT pixel_8851/CSA_VREF pixel
Xpixel_8840 pixel_8840/gring pixel_8840/VDD pixel_8840/GND pixel_8840/VREF pixel_8840/ROW_SEL
+ pixel_8840/NB1 pixel_8840/VBIAS pixel_8840/NB2 pixel_8840/AMP_IN pixel_8840/SF_IB
+ pixel_8840/PIX_OUT pixel_8840/CSA_VREF pixel
Xpixel_9596 pixel_9596/gring pixel_9596/VDD pixel_9596/GND pixel_9596/VREF pixel_9596/ROW_SEL
+ pixel_9596/NB1 pixel_9596/VBIAS pixel_9596/NB2 pixel_9596/AMP_IN pixel_9596/SF_IB
+ pixel_9596/PIX_OUT pixel_9596/CSA_VREF pixel
Xpixel_9585 pixel_9585/gring pixel_9585/VDD pixel_9585/GND pixel_9585/VREF pixel_9585/ROW_SEL
+ pixel_9585/NB1 pixel_9585/VBIAS pixel_9585/NB2 pixel_9585/AMP_IN pixel_9585/SF_IB
+ pixel_9585/PIX_OUT pixel_9585/CSA_VREF pixel
Xpixel_8895 pixel_8895/gring pixel_8895/VDD pixel_8895/GND pixel_8895/VREF pixel_8895/ROW_SEL
+ pixel_8895/NB1 pixel_8895/VBIAS pixel_8895/NB2 pixel_8895/AMP_IN pixel_8895/SF_IB
+ pixel_8895/PIX_OUT pixel_8895/CSA_VREF pixel
Xpixel_8884 pixel_8884/gring pixel_8884/VDD pixel_8884/GND pixel_8884/VREF pixel_8884/ROW_SEL
+ pixel_8884/NB1 pixel_8884/VBIAS pixel_8884/NB2 pixel_8884/AMP_IN pixel_8884/SF_IB
+ pixel_8884/PIX_OUT pixel_8884/CSA_VREF pixel
Xpixel_3191 pixel_3191/gring pixel_3191/VDD pixel_3191/GND pixel_3191/VREF pixel_3191/ROW_SEL
+ pixel_3191/NB1 pixel_3191/VBIAS pixel_3191/NB2 pixel_3191/AMP_IN pixel_3191/SF_IB
+ pixel_3191/PIX_OUT pixel_3191/CSA_VREF pixel
Xpixel_3180 pixel_3180/gring pixel_3180/VDD pixel_3180/GND pixel_3180/VREF pixel_3180/ROW_SEL
+ pixel_3180/NB1 pixel_3180/VBIAS pixel_3180/NB2 pixel_3180/AMP_IN pixel_3180/SF_IB
+ pixel_3180/PIX_OUT pixel_3180/CSA_VREF pixel
Xpixel_2490 pixel_2490/gring pixel_2490/VDD pixel_2490/GND pixel_2490/VREF pixel_2490/ROW_SEL
+ pixel_2490/NB1 pixel_2490/VBIAS pixel_2490/NB2 pixel_2490/AMP_IN pixel_2490/SF_IB
+ pixel_2490/PIX_OUT pixel_2490/CSA_VREF pixel
Xpixel_815 pixel_815/gring pixel_815/VDD pixel_815/GND pixel_815/VREF pixel_815/ROW_SEL
+ pixel_815/NB1 pixel_815/VBIAS pixel_815/NB2 pixel_815/AMP_IN pixel_815/SF_IB pixel_815/PIX_OUT
+ pixel_815/CSA_VREF pixel
Xpixel_804 pixel_804/gring pixel_804/VDD pixel_804/GND pixel_804/VREF pixel_804/ROW_SEL
+ pixel_804/NB1 pixel_804/VBIAS pixel_804/NB2 pixel_804/AMP_IN pixel_804/SF_IB pixel_804/PIX_OUT
+ pixel_804/CSA_VREF pixel
Xpixel_4809 pixel_4809/gring pixel_4809/VDD pixel_4809/GND pixel_4809/VREF pixel_4809/ROW_SEL
+ pixel_4809/NB1 pixel_4809/VBIAS pixel_4809/NB2 pixel_4809/AMP_IN pixel_4809/SF_IB
+ pixel_4809/PIX_OUT pixel_4809/CSA_VREF pixel
Xpixel_848 pixel_848/gring pixel_848/VDD pixel_848/GND pixel_848/VREF pixel_848/ROW_SEL
+ pixel_848/NB1 pixel_848/VBIAS pixel_848/NB2 pixel_848/AMP_IN pixel_848/SF_IB pixel_848/PIX_OUT
+ pixel_848/CSA_VREF pixel
Xpixel_837 pixel_837/gring pixel_837/VDD pixel_837/GND pixel_837/VREF pixel_837/ROW_SEL
+ pixel_837/NB1 pixel_837/VBIAS pixel_837/NB2 pixel_837/AMP_IN pixel_837/SF_IB pixel_837/PIX_OUT
+ pixel_837/CSA_VREF pixel
Xpixel_826 pixel_826/gring pixel_826/VDD pixel_826/GND pixel_826/VREF pixel_826/ROW_SEL
+ pixel_826/NB1 pixel_826/VBIAS pixel_826/NB2 pixel_826/AMP_IN pixel_826/SF_IB pixel_826/PIX_OUT
+ pixel_826/CSA_VREF pixel
Xpixel_859 pixel_859/gring pixel_859/VDD pixel_859/GND pixel_859/VREF pixel_859/ROW_SEL
+ pixel_859/NB1 pixel_859/VBIAS pixel_859/NB2 pixel_859/AMP_IN pixel_859/SF_IB pixel_859/PIX_OUT
+ pixel_859/CSA_VREF pixel
Xpixel_8103 pixel_8103/gring pixel_8103/VDD pixel_8103/GND pixel_8103/VREF pixel_8103/ROW_SEL
+ pixel_8103/NB1 pixel_8103/VBIAS pixel_8103/NB2 pixel_8103/AMP_IN pixel_8103/SF_IB
+ pixel_8103/PIX_OUT pixel_8103/CSA_VREF pixel
Xpixel_8114 pixel_8114/gring pixel_8114/VDD pixel_8114/GND pixel_8114/VREF pixel_8114/ROW_SEL
+ pixel_8114/NB1 pixel_8114/VBIAS pixel_8114/NB2 pixel_8114/AMP_IN pixel_8114/SF_IB
+ pixel_8114/PIX_OUT pixel_8114/CSA_VREF pixel
Xpixel_8125 pixel_8125/gring pixel_8125/VDD pixel_8125/GND pixel_8125/VREF pixel_8125/ROW_SEL
+ pixel_8125/NB1 pixel_8125/VBIAS pixel_8125/NB2 pixel_8125/AMP_IN pixel_8125/SF_IB
+ pixel_8125/PIX_OUT pixel_8125/CSA_VREF pixel
Xpixel_8136 pixel_8136/gring pixel_8136/VDD pixel_8136/GND pixel_8136/VREF pixel_8136/ROW_SEL
+ pixel_8136/NB1 pixel_8136/VBIAS pixel_8136/NB2 pixel_8136/AMP_IN pixel_8136/SF_IB
+ pixel_8136/PIX_OUT pixel_8136/CSA_VREF pixel
Xpixel_8147 pixel_8147/gring pixel_8147/VDD pixel_8147/GND pixel_8147/VREF pixel_8147/ROW_SEL
+ pixel_8147/NB1 pixel_8147/VBIAS pixel_8147/NB2 pixel_8147/AMP_IN pixel_8147/SF_IB
+ pixel_8147/PIX_OUT pixel_8147/CSA_VREF pixel
Xpixel_8158 pixel_8158/gring pixel_8158/VDD pixel_8158/GND pixel_8158/VREF pixel_8158/ROW_SEL
+ pixel_8158/NB1 pixel_8158/VBIAS pixel_8158/NB2 pixel_8158/AMP_IN pixel_8158/SF_IB
+ pixel_8158/PIX_OUT pixel_8158/CSA_VREF pixel
Xpixel_7402 pixel_7402/gring pixel_7402/VDD pixel_7402/GND pixel_7402/VREF pixel_7402/ROW_SEL
+ pixel_7402/NB1 pixel_7402/VBIAS pixel_7402/NB2 pixel_7402/AMP_IN pixel_7402/SF_IB
+ pixel_7402/PIX_OUT pixel_7402/CSA_VREF pixel
Xpixel_7413 pixel_7413/gring pixel_7413/VDD pixel_7413/GND pixel_7413/VREF pixel_7413/ROW_SEL
+ pixel_7413/NB1 pixel_7413/VBIAS pixel_7413/NB2 pixel_7413/AMP_IN pixel_7413/SF_IB
+ pixel_7413/PIX_OUT pixel_7413/CSA_VREF pixel
Xpixel_8169 pixel_8169/gring pixel_8169/VDD pixel_8169/GND pixel_8169/VREF pixel_8169/ROW_SEL
+ pixel_8169/NB1 pixel_8169/VBIAS pixel_8169/NB2 pixel_8169/AMP_IN pixel_8169/SF_IB
+ pixel_8169/PIX_OUT pixel_8169/CSA_VREF pixel
Xpixel_7424 pixel_7424/gring pixel_7424/VDD pixel_7424/GND pixel_7424/VREF pixel_7424/ROW_SEL
+ pixel_7424/NB1 pixel_7424/VBIAS pixel_7424/NB2 pixel_7424/AMP_IN pixel_7424/SF_IB
+ pixel_7424/PIX_OUT pixel_7424/CSA_VREF pixel
Xpixel_7435 pixel_7435/gring pixel_7435/VDD pixel_7435/GND pixel_7435/VREF pixel_7435/ROW_SEL
+ pixel_7435/NB1 pixel_7435/VBIAS pixel_7435/NB2 pixel_7435/AMP_IN pixel_7435/SF_IB
+ pixel_7435/PIX_OUT pixel_7435/CSA_VREF pixel
Xpixel_7446 pixel_7446/gring pixel_7446/VDD pixel_7446/GND pixel_7446/VREF pixel_7446/ROW_SEL
+ pixel_7446/NB1 pixel_7446/VBIAS pixel_7446/NB2 pixel_7446/AMP_IN pixel_7446/SF_IB
+ pixel_7446/PIX_OUT pixel_7446/CSA_VREF pixel
Xpixel_7457 pixel_7457/gring pixel_7457/VDD pixel_7457/GND pixel_7457/VREF pixel_7457/ROW_SEL
+ pixel_7457/NB1 pixel_7457/VBIAS pixel_7457/NB2 pixel_7457/AMP_IN pixel_7457/SF_IB
+ pixel_7457/PIX_OUT pixel_7457/CSA_VREF pixel
Xpixel_6701 pixel_6701/gring pixel_6701/VDD pixel_6701/GND pixel_6701/VREF pixel_6701/ROW_SEL
+ pixel_6701/NB1 pixel_6701/VBIAS pixel_6701/NB2 pixel_6701/AMP_IN pixel_6701/SF_IB
+ pixel_6701/PIX_OUT pixel_6701/CSA_VREF pixel
Xpixel_6712 pixel_6712/gring pixel_6712/VDD pixel_6712/GND pixel_6712/VREF pixel_6712/ROW_SEL
+ pixel_6712/NB1 pixel_6712/VBIAS pixel_6712/NB2 pixel_6712/AMP_IN pixel_6712/SF_IB
+ pixel_6712/PIX_OUT pixel_6712/CSA_VREF pixel
Xpixel_7468 pixel_7468/gring pixel_7468/VDD pixel_7468/GND pixel_7468/VREF pixel_7468/ROW_SEL
+ pixel_7468/NB1 pixel_7468/VBIAS pixel_7468/NB2 pixel_7468/AMP_IN pixel_7468/SF_IB
+ pixel_7468/PIX_OUT pixel_7468/CSA_VREF pixel
Xpixel_7479 pixel_7479/gring pixel_7479/VDD pixel_7479/GND pixel_7479/VREF pixel_7479/ROW_SEL
+ pixel_7479/NB1 pixel_7479/VBIAS pixel_7479/NB2 pixel_7479/AMP_IN pixel_7479/SF_IB
+ pixel_7479/PIX_OUT pixel_7479/CSA_VREF pixel
Xpixel_6723 pixel_6723/gring pixel_6723/VDD pixel_6723/GND pixel_6723/VREF pixel_6723/ROW_SEL
+ pixel_6723/NB1 pixel_6723/VBIAS pixel_6723/NB2 pixel_6723/AMP_IN pixel_6723/SF_IB
+ pixel_6723/PIX_OUT pixel_6723/CSA_VREF pixel
Xpixel_6734 pixel_6734/gring pixel_6734/VDD pixel_6734/GND pixel_6734/VREF pixel_6734/ROW_SEL
+ pixel_6734/NB1 pixel_6734/VBIAS pixel_6734/NB2 pixel_6734/AMP_IN pixel_6734/SF_IB
+ pixel_6734/PIX_OUT pixel_6734/CSA_VREF pixel
Xpixel_6745 pixel_6745/gring pixel_6745/VDD pixel_6745/GND pixel_6745/VREF pixel_6745/ROW_SEL
+ pixel_6745/NB1 pixel_6745/VBIAS pixel_6745/NB2 pixel_6745/AMP_IN pixel_6745/SF_IB
+ pixel_6745/PIX_OUT pixel_6745/CSA_VREF pixel
Xpixel_6756 pixel_6756/gring pixel_6756/VDD pixel_6756/GND pixel_6756/VREF pixel_6756/ROW_SEL
+ pixel_6756/NB1 pixel_6756/VBIAS pixel_6756/NB2 pixel_6756/AMP_IN pixel_6756/SF_IB
+ pixel_6756/PIX_OUT pixel_6756/CSA_VREF pixel
Xpixel_6767 pixel_6767/gring pixel_6767/VDD pixel_6767/GND pixel_6767/VREF pixel_6767/ROW_SEL
+ pixel_6767/NB1 pixel_6767/VBIAS pixel_6767/NB2 pixel_6767/AMP_IN pixel_6767/SF_IB
+ pixel_6767/PIX_OUT pixel_6767/CSA_VREF pixel
Xpixel_6778 pixel_6778/gring pixel_6778/VDD pixel_6778/GND pixel_6778/VREF pixel_6778/ROW_SEL
+ pixel_6778/NB1 pixel_6778/VBIAS pixel_6778/NB2 pixel_6778/AMP_IN pixel_6778/SF_IB
+ pixel_6778/PIX_OUT pixel_6778/CSA_VREF pixel
Xpixel_6789 pixel_6789/gring pixel_6789/VDD pixel_6789/GND pixel_6789/VREF pixel_6789/ROW_SEL
+ pixel_6789/NB1 pixel_6789/VBIAS pixel_6789/NB2 pixel_6789/AMP_IN pixel_6789/SF_IB
+ pixel_6789/PIX_OUT pixel_6789/CSA_VREF pixel
Xpixel_1041 pixel_1041/gring pixel_1041/VDD pixel_1041/GND pixel_1041/VREF pixel_1041/ROW_SEL
+ pixel_1041/NB1 pixel_1041/VBIAS pixel_1041/NB2 pixel_1041/AMP_IN pixel_1041/SF_IB
+ pixel_1041/PIX_OUT pixel_1041/CSA_VREF pixel
Xpixel_1030 pixel_1030/gring pixel_1030/VDD pixel_1030/GND pixel_1030/VREF pixel_1030/ROW_SEL
+ pixel_1030/NB1 pixel_1030/VBIAS pixel_1030/NB2 pixel_1030/AMP_IN pixel_1030/SF_IB
+ pixel_1030/PIX_OUT pixel_1030/CSA_VREF pixel
Xpixel_1074 pixel_1074/gring pixel_1074/VDD pixel_1074/GND pixel_1074/VREF pixel_1074/ROW_SEL
+ pixel_1074/NB1 pixel_1074/VBIAS pixel_1074/NB2 pixel_1074/AMP_IN pixel_1074/SF_IB
+ pixel_1074/PIX_OUT pixel_1074/CSA_VREF pixel
Xpixel_1063 pixel_1063/gring pixel_1063/VDD pixel_1063/GND pixel_1063/VREF pixel_1063/ROW_SEL
+ pixel_1063/NB1 pixel_1063/VBIAS pixel_1063/NB2 pixel_1063/AMP_IN pixel_1063/SF_IB
+ pixel_1063/PIX_OUT pixel_1063/CSA_VREF pixel
Xpixel_1052 pixel_1052/gring pixel_1052/VDD pixel_1052/GND pixel_1052/VREF pixel_1052/ROW_SEL
+ pixel_1052/NB1 pixel_1052/VBIAS pixel_1052/NB2 pixel_1052/AMP_IN pixel_1052/SF_IB
+ pixel_1052/PIX_OUT pixel_1052/CSA_VREF pixel
Xpixel_1096 pixel_1096/gring pixel_1096/VDD pixel_1096/GND pixel_1096/VREF pixel_1096/ROW_SEL
+ pixel_1096/NB1 pixel_1096/VBIAS pixel_1096/NB2 pixel_1096/AMP_IN pixel_1096/SF_IB
+ pixel_1096/PIX_OUT pixel_1096/CSA_VREF pixel
Xpixel_1085 pixel_1085/gring pixel_1085/VDD pixel_1085/GND pixel_1085/VREF pixel_1085/ROW_SEL
+ pixel_1085/NB1 pixel_1085/VBIAS pixel_1085/NB2 pixel_1085/AMP_IN pixel_1085/SF_IB
+ pixel_1085/PIX_OUT pixel_1085/CSA_VREF pixel
Xpixel_9382 pixel_9382/gring pixel_9382/VDD pixel_9382/GND pixel_9382/VREF pixel_9382/ROW_SEL
+ pixel_9382/NB1 pixel_9382/VBIAS pixel_9382/NB2 pixel_9382/AMP_IN pixel_9382/SF_IB
+ pixel_9382/PIX_OUT pixel_9382/CSA_VREF pixel
Xpixel_9371 pixel_9371/gring pixel_9371/VDD pixel_9371/GND pixel_9371/VREF pixel_9371/ROW_SEL
+ pixel_9371/NB1 pixel_9371/VBIAS pixel_9371/NB2 pixel_9371/AMP_IN pixel_9371/SF_IB
+ pixel_9371/PIX_OUT pixel_9371/CSA_VREF pixel
Xpixel_9360 pixel_9360/gring pixel_9360/VDD pixel_9360/GND pixel_9360/VREF pixel_9360/ROW_SEL
+ pixel_9360/NB1 pixel_9360/VBIAS pixel_9360/NB2 pixel_9360/AMP_IN pixel_9360/SF_IB
+ pixel_9360/PIX_OUT pixel_9360/CSA_VREF pixel
Xpixel_8681 pixel_8681/gring pixel_8681/VDD pixel_8681/GND pixel_8681/VREF pixel_8681/ROW_SEL
+ pixel_8681/NB1 pixel_8681/VBIAS pixel_8681/NB2 pixel_8681/AMP_IN pixel_8681/SF_IB
+ pixel_8681/PIX_OUT pixel_8681/CSA_VREF pixel
Xpixel_8670 pixel_8670/gring pixel_8670/VDD pixel_8670/GND pixel_8670/VREF pixel_8670/ROW_SEL
+ pixel_8670/NB1 pixel_8670/VBIAS pixel_8670/NB2 pixel_8670/AMP_IN pixel_8670/SF_IB
+ pixel_8670/PIX_OUT pixel_8670/CSA_VREF pixel
Xpixel_9393 pixel_9393/gring pixel_9393/VDD pixel_9393/GND pixel_9393/VREF pixel_9393/ROW_SEL
+ pixel_9393/NB1 pixel_9393/VBIAS pixel_9393/NB2 pixel_9393/AMP_IN pixel_9393/SF_IB
+ pixel_9393/PIX_OUT pixel_9393/CSA_VREF pixel
Xpixel_8692 pixel_8692/gring pixel_8692/VDD pixel_8692/GND pixel_8692/VREF pixel_8692/ROW_SEL
+ pixel_8692/NB1 pixel_8692/VBIAS pixel_8692/NB2 pixel_8692/AMP_IN pixel_8692/SF_IB
+ pixel_8692/PIX_OUT pixel_8692/CSA_VREF pixel
Xpixel_7980 pixel_7980/gring pixel_7980/VDD pixel_7980/GND pixel_7980/VREF pixel_7980/ROW_SEL
+ pixel_7980/NB1 pixel_7980/VBIAS pixel_7980/NB2 pixel_7980/AMP_IN pixel_7980/SF_IB
+ pixel_7980/PIX_OUT pixel_7980/CSA_VREF pixel
Xpixel_7991 pixel_7991/gring pixel_7991/VDD pixel_7991/GND pixel_7991/VREF pixel_7991/ROW_SEL
+ pixel_7991/NB1 pixel_7991/VBIAS pixel_7991/NB2 pixel_7991/AMP_IN pixel_7991/SF_IB
+ pixel_7991/PIX_OUT pixel_7991/CSA_VREF pixel
Xpixel_6008 pixel_6008/gring pixel_6008/VDD pixel_6008/GND pixel_6008/VREF pixel_6008/ROW_SEL
+ pixel_6008/NB1 pixel_6008/VBIAS pixel_6008/NB2 pixel_6008/AMP_IN pixel_6008/SF_IB
+ pixel_6008/PIX_OUT pixel_6008/CSA_VREF pixel
Xpixel_6019 pixel_6019/gring pixel_6019/VDD pixel_6019/GND pixel_6019/VREF pixel_6019/ROW_SEL
+ pixel_6019/NB1 pixel_6019/VBIAS pixel_6019/NB2 pixel_6019/AMP_IN pixel_6019/SF_IB
+ pixel_6019/PIX_OUT pixel_6019/CSA_VREF pixel
Xpixel_5307 pixel_5307/gring pixel_5307/VDD pixel_5307/GND pixel_5307/VREF pixel_5307/ROW_SEL
+ pixel_5307/NB1 pixel_5307/VBIAS pixel_5307/NB2 pixel_5307/AMP_IN pixel_5307/SF_IB
+ pixel_5307/PIX_OUT pixel_5307/CSA_VREF pixel
Xpixel_5318 pixel_5318/gring pixel_5318/VDD pixel_5318/GND pixel_5318/VREF pixel_5318/ROW_SEL
+ pixel_5318/NB1 pixel_5318/VBIAS pixel_5318/NB2 pixel_5318/AMP_IN pixel_5318/SF_IB
+ pixel_5318/PIX_OUT pixel_5318/CSA_VREF pixel
Xpixel_5329 pixel_5329/gring pixel_5329/VDD pixel_5329/GND pixel_5329/VREF pixel_5329/ROW_SEL
+ pixel_5329/NB1 pixel_5329/VBIAS pixel_5329/NB2 pixel_5329/AMP_IN pixel_5329/SF_IB
+ pixel_5329/PIX_OUT pixel_5329/CSA_VREF pixel
Xpixel_623 pixel_623/gring pixel_623/VDD pixel_623/GND pixel_623/VREF pixel_623/ROW_SEL
+ pixel_623/NB1 pixel_623/VBIAS pixel_623/NB2 pixel_623/AMP_IN pixel_623/SF_IB pixel_623/PIX_OUT
+ pixel_623/CSA_VREF pixel
Xpixel_612 pixel_612/gring pixel_612/VDD pixel_612/GND pixel_612/VREF pixel_612/ROW_SEL
+ pixel_612/NB1 pixel_612/VBIAS pixel_612/NB2 pixel_612/AMP_IN pixel_612/SF_IB pixel_612/PIX_OUT
+ pixel_612/CSA_VREF pixel
Xpixel_601 pixel_601/gring pixel_601/VDD pixel_601/GND pixel_601/VREF pixel_601/ROW_SEL
+ pixel_601/NB1 pixel_601/VBIAS pixel_601/NB2 pixel_601/AMP_IN pixel_601/SF_IB pixel_601/PIX_OUT
+ pixel_601/CSA_VREF pixel
Xpixel_4606 pixel_4606/gring pixel_4606/VDD pixel_4606/GND pixel_4606/VREF pixel_4606/ROW_SEL
+ pixel_4606/NB1 pixel_4606/VBIAS pixel_4606/NB2 pixel_4606/AMP_IN pixel_4606/SF_IB
+ pixel_4606/PIX_OUT pixel_4606/CSA_VREF pixel
Xpixel_4617 pixel_4617/gring pixel_4617/VDD pixel_4617/GND pixel_4617/VREF pixel_4617/ROW_SEL
+ pixel_4617/NB1 pixel_4617/VBIAS pixel_4617/NB2 pixel_4617/AMP_IN pixel_4617/SF_IB
+ pixel_4617/PIX_OUT pixel_4617/CSA_VREF pixel
Xpixel_4628 pixel_4628/gring pixel_4628/VDD pixel_4628/GND pixel_4628/VREF pixel_4628/ROW_SEL
+ pixel_4628/NB1 pixel_4628/VBIAS pixel_4628/NB2 pixel_4628/AMP_IN pixel_4628/SF_IB
+ pixel_4628/PIX_OUT pixel_4628/CSA_VREF pixel
Xpixel_656 pixel_656/gring pixel_656/VDD pixel_656/GND pixel_656/VREF pixel_656/ROW_SEL
+ pixel_656/NB1 pixel_656/VBIAS pixel_656/NB2 pixel_656/AMP_IN pixel_656/SF_IB pixel_656/PIX_OUT
+ pixel_656/CSA_VREF pixel
Xpixel_645 pixel_645/gring pixel_645/VDD pixel_645/GND pixel_645/VREF pixel_645/ROW_SEL
+ pixel_645/NB1 pixel_645/VBIAS pixel_645/NB2 pixel_645/AMP_IN pixel_645/SF_IB pixel_645/PIX_OUT
+ pixel_645/CSA_VREF pixel
Xpixel_634 pixel_634/gring pixel_634/VDD pixel_634/GND pixel_634/VREF pixel_634/ROW_SEL
+ pixel_634/NB1 pixel_634/VBIAS pixel_634/NB2 pixel_634/AMP_IN pixel_634/SF_IB pixel_634/PIX_OUT
+ pixel_634/CSA_VREF pixel
Xpixel_4639 pixel_4639/gring pixel_4639/VDD pixel_4639/GND pixel_4639/VREF pixel_4639/ROW_SEL
+ pixel_4639/NB1 pixel_4639/VBIAS pixel_4639/NB2 pixel_4639/AMP_IN pixel_4639/SF_IB
+ pixel_4639/PIX_OUT pixel_4639/CSA_VREF pixel
Xpixel_3905 pixel_3905/gring pixel_3905/VDD pixel_3905/GND pixel_3905/VREF pixel_3905/ROW_SEL
+ pixel_3905/NB1 pixel_3905/VBIAS pixel_3905/NB2 pixel_3905/AMP_IN pixel_3905/SF_IB
+ pixel_3905/PIX_OUT pixel_3905/CSA_VREF pixel
Xpixel_3916 pixel_3916/gring pixel_3916/VDD pixel_3916/GND pixel_3916/VREF pixel_3916/ROW_SEL
+ pixel_3916/NB1 pixel_3916/VBIAS pixel_3916/NB2 pixel_3916/AMP_IN pixel_3916/SF_IB
+ pixel_3916/PIX_OUT pixel_3916/CSA_VREF pixel
Xpixel_689 pixel_689/gring pixel_689/VDD pixel_689/GND pixel_689/VREF pixel_689/ROW_SEL
+ pixel_689/NB1 pixel_689/VBIAS pixel_689/NB2 pixel_689/AMP_IN pixel_689/SF_IB pixel_689/PIX_OUT
+ pixel_689/CSA_VREF pixel
Xpixel_678 pixel_678/gring pixel_678/VDD pixel_678/GND pixel_678/VREF pixel_678/ROW_SEL
+ pixel_678/NB1 pixel_678/VBIAS pixel_678/NB2 pixel_678/AMP_IN pixel_678/SF_IB pixel_678/PIX_OUT
+ pixel_678/CSA_VREF pixel
Xpixel_667 pixel_667/gring pixel_667/VDD pixel_667/GND pixel_667/VREF pixel_667/ROW_SEL
+ pixel_667/NB1 pixel_667/VBIAS pixel_667/NB2 pixel_667/AMP_IN pixel_667/SF_IB pixel_667/PIX_OUT
+ pixel_667/CSA_VREF pixel
Xpixel_3927 pixel_3927/gring pixel_3927/VDD pixel_3927/GND pixel_3927/VREF pixel_3927/ROW_SEL
+ pixel_3927/NB1 pixel_3927/VBIAS pixel_3927/NB2 pixel_3927/AMP_IN pixel_3927/SF_IB
+ pixel_3927/PIX_OUT pixel_3927/CSA_VREF pixel
Xpixel_3938 pixel_3938/gring pixel_3938/VDD pixel_3938/GND pixel_3938/VREF pixel_3938/ROW_SEL
+ pixel_3938/NB1 pixel_3938/VBIAS pixel_3938/NB2 pixel_3938/AMP_IN pixel_3938/SF_IB
+ pixel_3938/PIX_OUT pixel_3938/CSA_VREF pixel
Xpixel_3949 pixel_3949/gring pixel_3949/VDD pixel_3949/GND pixel_3949/VREF pixel_3949/ROW_SEL
+ pixel_3949/NB1 pixel_3949/VBIAS pixel_3949/NB2 pixel_3949/AMP_IN pixel_3949/SF_IB
+ pixel_3949/PIX_OUT pixel_3949/CSA_VREF pixel
Xpixel_7210 pixel_7210/gring pixel_7210/VDD pixel_7210/GND pixel_7210/VREF pixel_7210/ROW_SEL
+ pixel_7210/NB1 pixel_7210/VBIAS pixel_7210/NB2 pixel_7210/AMP_IN pixel_7210/SF_IB
+ pixel_7210/PIX_OUT pixel_7210/CSA_VREF pixel
Xpixel_7221 pixel_7221/gring pixel_7221/VDD pixel_7221/GND pixel_7221/VREF pixel_7221/ROW_SEL
+ pixel_7221/NB1 pixel_7221/VBIAS pixel_7221/NB2 pixel_7221/AMP_IN pixel_7221/SF_IB
+ pixel_7221/PIX_OUT pixel_7221/CSA_VREF pixel
Xpixel_7232 pixel_7232/gring pixel_7232/VDD pixel_7232/GND pixel_7232/VREF pixel_7232/ROW_SEL
+ pixel_7232/NB1 pixel_7232/VBIAS pixel_7232/NB2 pixel_7232/AMP_IN pixel_7232/SF_IB
+ pixel_7232/PIX_OUT pixel_7232/CSA_VREF pixel
Xpixel_7243 pixel_7243/gring pixel_7243/VDD pixel_7243/GND pixel_7243/VREF pixel_7243/ROW_SEL
+ pixel_7243/NB1 pixel_7243/VBIAS pixel_7243/NB2 pixel_7243/AMP_IN pixel_7243/SF_IB
+ pixel_7243/PIX_OUT pixel_7243/CSA_VREF pixel
Xpixel_7254 pixel_7254/gring pixel_7254/VDD pixel_7254/GND pixel_7254/VREF pixel_7254/ROW_SEL
+ pixel_7254/NB1 pixel_7254/VBIAS pixel_7254/NB2 pixel_7254/AMP_IN pixel_7254/SF_IB
+ pixel_7254/PIX_OUT pixel_7254/CSA_VREF pixel
Xpixel_7265 pixel_7265/gring pixel_7265/VDD pixel_7265/GND pixel_7265/VREF pixel_7265/ROW_SEL
+ pixel_7265/NB1 pixel_7265/VBIAS pixel_7265/NB2 pixel_7265/AMP_IN pixel_7265/SF_IB
+ pixel_7265/PIX_OUT pixel_7265/CSA_VREF pixel
Xpixel_6520 pixel_6520/gring pixel_6520/VDD pixel_6520/GND pixel_6520/VREF pixel_6520/ROW_SEL
+ pixel_6520/NB1 pixel_6520/VBIAS pixel_6520/NB2 pixel_6520/AMP_IN pixel_6520/SF_IB
+ pixel_6520/PIX_OUT pixel_6520/CSA_VREF pixel
Xpixel_7276 pixel_7276/gring pixel_7276/VDD pixel_7276/GND pixel_7276/VREF pixel_7276/ROW_SEL
+ pixel_7276/NB1 pixel_7276/VBIAS pixel_7276/NB2 pixel_7276/AMP_IN pixel_7276/SF_IB
+ pixel_7276/PIX_OUT pixel_7276/CSA_VREF pixel
Xpixel_7287 pixel_7287/gring pixel_7287/VDD pixel_7287/GND pixel_7287/VREF pixel_7287/ROW_SEL
+ pixel_7287/NB1 pixel_7287/VBIAS pixel_7287/NB2 pixel_7287/AMP_IN pixel_7287/SF_IB
+ pixel_7287/PIX_OUT pixel_7287/CSA_VREF pixel
Xpixel_7298 pixel_7298/gring pixel_7298/VDD pixel_7298/GND pixel_7298/VREF pixel_7298/ROW_SEL
+ pixel_7298/NB1 pixel_7298/VBIAS pixel_7298/NB2 pixel_7298/AMP_IN pixel_7298/SF_IB
+ pixel_7298/PIX_OUT pixel_7298/CSA_VREF pixel
Xpixel_6531 pixel_6531/gring pixel_6531/VDD pixel_6531/GND pixel_6531/VREF pixel_6531/ROW_SEL
+ pixel_6531/NB1 pixel_6531/VBIAS pixel_6531/NB2 pixel_6531/AMP_IN pixel_6531/SF_IB
+ pixel_6531/PIX_OUT pixel_6531/CSA_VREF pixel
Xpixel_6542 pixel_6542/gring pixel_6542/VDD pixel_6542/GND pixel_6542/VREF pixel_6542/ROW_SEL
+ pixel_6542/NB1 pixel_6542/VBIAS pixel_6542/NB2 pixel_6542/AMP_IN pixel_6542/SF_IB
+ pixel_6542/PIX_OUT pixel_6542/CSA_VREF pixel
Xpixel_6553 pixel_6553/gring pixel_6553/VDD pixel_6553/GND pixel_6553/VREF pixel_6553/ROW_SEL
+ pixel_6553/NB1 pixel_6553/VBIAS pixel_6553/NB2 pixel_6553/AMP_IN pixel_6553/SF_IB
+ pixel_6553/PIX_OUT pixel_6553/CSA_VREF pixel
Xpixel_6564 pixel_6564/gring pixel_6564/VDD pixel_6564/GND pixel_6564/VREF pixel_6564/ROW_SEL
+ pixel_6564/NB1 pixel_6564/VBIAS pixel_6564/NB2 pixel_6564/AMP_IN pixel_6564/SF_IB
+ pixel_6564/PIX_OUT pixel_6564/CSA_VREF pixel
Xpixel_6575 pixel_6575/gring pixel_6575/VDD pixel_6575/GND pixel_6575/VREF pixel_6575/ROW_SEL
+ pixel_6575/NB1 pixel_6575/VBIAS pixel_6575/NB2 pixel_6575/AMP_IN pixel_6575/SF_IB
+ pixel_6575/PIX_OUT pixel_6575/CSA_VREF pixel
Xpixel_6586 pixel_6586/gring pixel_6586/VDD pixel_6586/GND pixel_6586/VREF pixel_6586/ROW_SEL
+ pixel_6586/NB1 pixel_6586/VBIAS pixel_6586/NB2 pixel_6586/AMP_IN pixel_6586/SF_IB
+ pixel_6586/PIX_OUT pixel_6586/CSA_VREF pixel
Xpixel_6597 pixel_6597/gring pixel_6597/VDD pixel_6597/GND pixel_6597/VREF pixel_6597/ROW_SEL
+ pixel_6597/NB1 pixel_6597/VBIAS pixel_6597/NB2 pixel_6597/AMP_IN pixel_6597/SF_IB
+ pixel_6597/PIX_OUT pixel_6597/CSA_VREF pixel
Xpixel_5830 pixel_5830/gring pixel_5830/VDD pixel_5830/GND pixel_5830/VREF pixel_5830/ROW_SEL
+ pixel_5830/NB1 pixel_5830/VBIAS pixel_5830/NB2 pixel_5830/AMP_IN pixel_5830/SF_IB
+ pixel_5830/PIX_OUT pixel_5830/CSA_VREF pixel
Xpixel_5841 pixel_5841/gring pixel_5841/VDD pixel_5841/GND pixel_5841/VREF pixel_5841/ROW_SEL
+ pixel_5841/NB1 pixel_5841/VBIAS pixel_5841/NB2 pixel_5841/AMP_IN pixel_5841/SF_IB
+ pixel_5841/PIX_OUT pixel_5841/CSA_VREF pixel
Xpixel_5852 pixel_5852/gring pixel_5852/VDD pixel_5852/GND pixel_5852/VREF pixel_5852/ROW_SEL
+ pixel_5852/NB1 pixel_5852/VBIAS pixel_5852/NB2 pixel_5852/AMP_IN pixel_5852/SF_IB
+ pixel_5852/PIX_OUT pixel_5852/CSA_VREF pixel
Xpixel_5863 pixel_5863/gring pixel_5863/VDD pixel_5863/GND pixel_5863/VREF pixel_5863/ROW_SEL
+ pixel_5863/NB1 pixel_5863/VBIAS pixel_5863/NB2 pixel_5863/AMP_IN pixel_5863/SF_IB
+ pixel_5863/PIX_OUT pixel_5863/CSA_VREF pixel
Xpixel_5874 pixel_5874/gring pixel_5874/VDD pixel_5874/GND pixel_5874/VREF pixel_5874/ROW_SEL
+ pixel_5874/NB1 pixel_5874/VBIAS pixel_5874/NB2 pixel_5874/AMP_IN pixel_5874/SF_IB
+ pixel_5874/PIX_OUT pixel_5874/CSA_VREF pixel
Xpixel_5885 pixel_5885/gring pixel_5885/VDD pixel_5885/GND pixel_5885/VREF pixel_5885/ROW_SEL
+ pixel_5885/NB1 pixel_5885/VBIAS pixel_5885/NB2 pixel_5885/AMP_IN pixel_5885/SF_IB
+ pixel_5885/PIX_OUT pixel_5885/CSA_VREF pixel
Xpixel_5896 pixel_5896/gring pixel_5896/VDD pixel_5896/GND pixel_5896/VREF pixel_5896/ROW_SEL
+ pixel_5896/NB1 pixel_5896/VBIAS pixel_5896/NB2 pixel_5896/AMP_IN pixel_5896/SF_IB
+ pixel_5896/PIX_OUT pixel_5896/CSA_VREF pixel
Xpixel_9190 pixel_9190/gring pixel_9190/VDD pixel_9190/GND pixel_9190/VREF pixel_9190/ROW_SEL
+ pixel_9190/NB1 pixel_9190/VBIAS pixel_9190/NB2 pixel_9190/AMP_IN pixel_9190/SF_IB
+ pixel_9190/PIX_OUT pixel_9190/CSA_VREF pixel
Xpixel_5104 pixel_5104/gring pixel_5104/VDD pixel_5104/GND pixel_5104/VREF pixel_5104/ROW_SEL
+ pixel_5104/NB1 pixel_5104/VBIAS pixel_5104/NB2 pixel_5104/AMP_IN pixel_5104/SF_IB
+ pixel_5104/PIX_OUT pixel_5104/CSA_VREF pixel
Xpixel_5115 pixel_5115/gring pixel_5115/VDD pixel_5115/GND pixel_5115/VREF pixel_5115/ROW_SEL
+ pixel_5115/NB1 pixel_5115/VBIAS pixel_5115/NB2 pixel_5115/AMP_IN pixel_5115/SF_IB
+ pixel_5115/PIX_OUT pixel_5115/CSA_VREF pixel
Xpixel_5126 pixel_5126/gring pixel_5126/VDD pixel_5126/GND pixel_5126/VREF pixel_5126/ROW_SEL
+ pixel_5126/NB1 pixel_5126/VBIAS pixel_5126/NB2 pixel_5126/AMP_IN pixel_5126/SF_IB
+ pixel_5126/PIX_OUT pixel_5126/CSA_VREF pixel
Xpixel_5137 pixel_5137/gring pixel_5137/VDD pixel_5137/GND pixel_5137/VREF pixel_5137/ROW_SEL
+ pixel_5137/NB1 pixel_5137/VBIAS pixel_5137/NB2 pixel_5137/AMP_IN pixel_5137/SF_IB
+ pixel_5137/PIX_OUT pixel_5137/CSA_VREF pixel
Xpixel_4403 pixel_4403/gring pixel_4403/VDD pixel_4403/GND pixel_4403/VREF pixel_4403/ROW_SEL
+ pixel_4403/NB1 pixel_4403/VBIAS pixel_4403/NB2 pixel_4403/AMP_IN pixel_4403/SF_IB
+ pixel_4403/PIX_OUT pixel_4403/CSA_VREF pixel
Xpixel_431 pixel_431/gring pixel_431/VDD pixel_431/GND pixel_431/VREF pixel_431/ROW_SEL
+ pixel_431/NB1 pixel_431/VBIAS pixel_431/NB2 pixel_431/AMP_IN pixel_431/SF_IB pixel_431/PIX_OUT
+ pixel_431/CSA_VREF pixel
Xpixel_420 pixel_420/gring pixel_420/VDD pixel_420/GND pixel_420/VREF pixel_420/ROW_SEL
+ pixel_420/NB1 pixel_420/VBIAS pixel_420/NB2 pixel_420/AMP_IN pixel_420/SF_IB pixel_420/PIX_OUT
+ pixel_420/CSA_VREF pixel
Xpixel_5148 pixel_5148/gring pixel_5148/VDD pixel_5148/GND pixel_5148/VREF pixel_5148/ROW_SEL
+ pixel_5148/NB1 pixel_5148/VBIAS pixel_5148/NB2 pixel_5148/AMP_IN pixel_5148/SF_IB
+ pixel_5148/PIX_OUT pixel_5148/CSA_VREF pixel
Xpixel_5159 pixel_5159/gring pixel_5159/VDD pixel_5159/GND pixel_5159/VREF pixel_5159/ROW_SEL
+ pixel_5159/NB1 pixel_5159/VBIAS pixel_5159/NB2 pixel_5159/AMP_IN pixel_5159/SF_IB
+ pixel_5159/PIX_OUT pixel_5159/CSA_VREF pixel
Xpixel_4414 pixel_4414/gring pixel_4414/VDD pixel_4414/GND pixel_4414/VREF pixel_4414/ROW_SEL
+ pixel_4414/NB1 pixel_4414/VBIAS pixel_4414/NB2 pixel_4414/AMP_IN pixel_4414/SF_IB
+ pixel_4414/PIX_OUT pixel_4414/CSA_VREF pixel
Xpixel_4425 pixel_4425/gring pixel_4425/VDD pixel_4425/GND pixel_4425/VREF pixel_4425/ROW_SEL
+ pixel_4425/NB1 pixel_4425/VBIAS pixel_4425/NB2 pixel_4425/AMP_IN pixel_4425/SF_IB
+ pixel_4425/PIX_OUT pixel_4425/CSA_VREF pixel
Xpixel_4436 pixel_4436/gring pixel_4436/VDD pixel_4436/GND pixel_4436/VREF pixel_4436/ROW_SEL
+ pixel_4436/NB1 pixel_4436/VBIAS pixel_4436/NB2 pixel_4436/AMP_IN pixel_4436/SF_IB
+ pixel_4436/PIX_OUT pixel_4436/CSA_VREF pixel
Xpixel_464 pixel_464/gring pixel_464/VDD pixel_464/GND pixel_464/VREF pixel_464/ROW_SEL
+ pixel_464/NB1 pixel_464/VBIAS pixel_464/NB2 pixel_464/AMP_IN pixel_464/SF_IB pixel_464/PIX_OUT
+ pixel_464/CSA_VREF pixel
Xpixel_453 pixel_453/gring pixel_453/VDD pixel_453/GND pixel_453/VREF pixel_453/ROW_SEL
+ pixel_453/NB1 pixel_453/VBIAS pixel_453/NB2 pixel_453/AMP_IN pixel_453/SF_IB pixel_453/PIX_OUT
+ pixel_453/CSA_VREF pixel
Xpixel_442 pixel_442/gring pixel_442/VDD pixel_442/GND pixel_442/VREF pixel_442/ROW_SEL
+ pixel_442/NB1 pixel_442/VBIAS pixel_442/NB2 pixel_442/AMP_IN pixel_442/SF_IB pixel_442/PIX_OUT
+ pixel_442/CSA_VREF pixel
Xpixel_3724 pixel_3724/gring pixel_3724/VDD pixel_3724/GND pixel_3724/VREF pixel_3724/ROW_SEL
+ pixel_3724/NB1 pixel_3724/VBIAS pixel_3724/NB2 pixel_3724/AMP_IN pixel_3724/SF_IB
+ pixel_3724/PIX_OUT pixel_3724/CSA_VREF pixel
Xpixel_3713 pixel_3713/gring pixel_3713/VDD pixel_3713/GND pixel_3713/VREF pixel_3713/ROW_SEL
+ pixel_3713/NB1 pixel_3713/VBIAS pixel_3713/NB2 pixel_3713/AMP_IN pixel_3713/SF_IB
+ pixel_3713/PIX_OUT pixel_3713/CSA_VREF pixel
Xpixel_3702 pixel_3702/gring pixel_3702/VDD pixel_3702/GND pixel_3702/VREF pixel_3702/ROW_SEL
+ pixel_3702/NB1 pixel_3702/VBIAS pixel_3702/NB2 pixel_3702/AMP_IN pixel_3702/SF_IB
+ pixel_3702/PIX_OUT pixel_3702/CSA_VREF pixel
Xpixel_4447 pixel_4447/gring pixel_4447/VDD pixel_4447/GND pixel_4447/VREF pixel_4447/ROW_SEL
+ pixel_4447/NB1 pixel_4447/VBIAS pixel_4447/NB2 pixel_4447/AMP_IN pixel_4447/SF_IB
+ pixel_4447/PIX_OUT pixel_4447/CSA_VREF pixel
Xpixel_4458 pixel_4458/gring pixel_4458/VDD pixel_4458/GND pixel_4458/VREF pixel_4458/ROW_SEL
+ pixel_4458/NB1 pixel_4458/VBIAS pixel_4458/NB2 pixel_4458/AMP_IN pixel_4458/SF_IB
+ pixel_4458/PIX_OUT pixel_4458/CSA_VREF pixel
Xpixel_4469 pixel_4469/gring pixel_4469/VDD pixel_4469/GND pixel_4469/VREF pixel_4469/ROW_SEL
+ pixel_4469/NB1 pixel_4469/VBIAS pixel_4469/NB2 pixel_4469/AMP_IN pixel_4469/SF_IB
+ pixel_4469/PIX_OUT pixel_4469/CSA_VREF pixel
Xpixel_497 pixel_497/gring pixel_497/VDD pixel_497/GND pixel_497/VREF pixel_497/ROW_SEL
+ pixel_497/NB1 pixel_497/VBIAS pixel_497/NB2 pixel_497/AMP_IN pixel_497/SF_IB pixel_497/PIX_OUT
+ pixel_497/CSA_VREF pixel
Xpixel_486 pixel_486/gring pixel_486/VDD pixel_486/GND pixel_486/VREF pixel_486/ROW_SEL
+ pixel_486/NB1 pixel_486/VBIAS pixel_486/NB2 pixel_486/AMP_IN pixel_486/SF_IB pixel_486/PIX_OUT
+ pixel_486/CSA_VREF pixel
Xpixel_475 pixel_475/gring pixel_475/VDD pixel_475/GND pixel_475/VREF pixel_475/ROW_SEL
+ pixel_475/NB1 pixel_475/VBIAS pixel_475/NB2 pixel_475/AMP_IN pixel_475/SF_IB pixel_475/PIX_OUT
+ pixel_475/CSA_VREF pixel
Xpixel_3768 pixel_3768/gring pixel_3768/VDD pixel_3768/GND pixel_3768/VREF pixel_3768/ROW_SEL
+ pixel_3768/NB1 pixel_3768/VBIAS pixel_3768/NB2 pixel_3768/AMP_IN pixel_3768/SF_IB
+ pixel_3768/PIX_OUT pixel_3768/CSA_VREF pixel
Xpixel_3757 pixel_3757/gring pixel_3757/VDD pixel_3757/GND pixel_3757/VREF pixel_3757/ROW_SEL
+ pixel_3757/NB1 pixel_3757/VBIAS pixel_3757/NB2 pixel_3757/AMP_IN pixel_3757/SF_IB
+ pixel_3757/PIX_OUT pixel_3757/CSA_VREF pixel
Xpixel_3746 pixel_3746/gring pixel_3746/VDD pixel_3746/GND pixel_3746/VREF pixel_3746/ROW_SEL
+ pixel_3746/NB1 pixel_3746/VBIAS pixel_3746/NB2 pixel_3746/AMP_IN pixel_3746/SF_IB
+ pixel_3746/PIX_OUT pixel_3746/CSA_VREF pixel
Xpixel_3735 pixel_3735/gring pixel_3735/VDD pixel_3735/GND pixel_3735/VREF pixel_3735/ROW_SEL
+ pixel_3735/NB1 pixel_3735/VBIAS pixel_3735/NB2 pixel_3735/AMP_IN pixel_3735/SF_IB
+ pixel_3735/PIX_OUT pixel_3735/CSA_VREF pixel
Xpixel_3779 pixel_3779/gring pixel_3779/VDD pixel_3779/GND pixel_3779/VREF pixel_3779/ROW_SEL
+ pixel_3779/NB1 pixel_3779/VBIAS pixel_3779/NB2 pixel_3779/AMP_IN pixel_3779/SF_IB
+ pixel_3779/PIX_OUT pixel_3779/CSA_VREF pixel
Xpixel_7040 pixel_7040/gring pixel_7040/VDD pixel_7040/GND pixel_7040/VREF pixel_7040/ROW_SEL
+ pixel_7040/NB1 pixel_7040/VBIAS pixel_7040/NB2 pixel_7040/AMP_IN pixel_7040/SF_IB
+ pixel_7040/PIX_OUT pixel_7040/CSA_VREF pixel
Xpixel_7051 pixel_7051/gring pixel_7051/VDD pixel_7051/GND pixel_7051/VREF pixel_7051/ROW_SEL
+ pixel_7051/NB1 pixel_7051/VBIAS pixel_7051/NB2 pixel_7051/AMP_IN pixel_7051/SF_IB
+ pixel_7051/PIX_OUT pixel_7051/CSA_VREF pixel
Xpixel_7062 pixel_7062/gring pixel_7062/VDD pixel_7062/GND pixel_7062/VREF pixel_7062/ROW_SEL
+ pixel_7062/NB1 pixel_7062/VBIAS pixel_7062/NB2 pixel_7062/AMP_IN pixel_7062/SF_IB
+ pixel_7062/PIX_OUT pixel_7062/CSA_VREF pixel
Xpixel_7073 pixel_7073/gring pixel_7073/VDD pixel_7073/GND pixel_7073/VREF pixel_7073/ROW_SEL
+ pixel_7073/NB1 pixel_7073/VBIAS pixel_7073/NB2 pixel_7073/AMP_IN pixel_7073/SF_IB
+ pixel_7073/PIX_OUT pixel_7073/CSA_VREF pixel
Xpixel_7084 pixel_7084/gring pixel_7084/VDD pixel_7084/GND pixel_7084/VREF pixel_7084/ROW_SEL
+ pixel_7084/NB1 pixel_7084/VBIAS pixel_7084/NB2 pixel_7084/AMP_IN pixel_7084/SF_IB
+ pixel_7084/PIX_OUT pixel_7084/CSA_VREF pixel
Xpixel_7095 pixel_7095/gring pixel_7095/VDD pixel_7095/GND pixel_7095/VREF pixel_7095/ROW_SEL
+ pixel_7095/NB1 pixel_7095/VBIAS pixel_7095/NB2 pixel_7095/AMP_IN pixel_7095/SF_IB
+ pixel_7095/PIX_OUT pixel_7095/CSA_VREF pixel
Xpixel_6350 pixel_6350/gring pixel_6350/VDD pixel_6350/GND pixel_6350/VREF pixel_6350/ROW_SEL
+ pixel_6350/NB1 pixel_6350/VBIAS pixel_6350/NB2 pixel_6350/AMP_IN pixel_6350/SF_IB
+ pixel_6350/PIX_OUT pixel_6350/CSA_VREF pixel
Xpixel_6361 pixel_6361/gring pixel_6361/VDD pixel_6361/GND pixel_6361/VREF pixel_6361/ROW_SEL
+ pixel_6361/NB1 pixel_6361/VBIAS pixel_6361/NB2 pixel_6361/AMP_IN pixel_6361/SF_IB
+ pixel_6361/PIX_OUT pixel_6361/CSA_VREF pixel
Xpixel_6372 pixel_6372/gring pixel_6372/VDD pixel_6372/GND pixel_6372/VREF pixel_6372/ROW_SEL
+ pixel_6372/NB1 pixel_6372/VBIAS pixel_6372/NB2 pixel_6372/AMP_IN pixel_6372/SF_IB
+ pixel_6372/PIX_OUT pixel_6372/CSA_VREF pixel
Xpixel_6383 pixel_6383/gring pixel_6383/VDD pixel_6383/GND pixel_6383/VREF pixel_6383/ROW_SEL
+ pixel_6383/NB1 pixel_6383/VBIAS pixel_6383/NB2 pixel_6383/AMP_IN pixel_6383/SF_IB
+ pixel_6383/PIX_OUT pixel_6383/CSA_VREF pixel
Xpixel_6394 pixel_6394/gring pixel_6394/VDD pixel_6394/GND pixel_6394/VREF pixel_6394/ROW_SEL
+ pixel_6394/NB1 pixel_6394/VBIAS pixel_6394/NB2 pixel_6394/AMP_IN pixel_6394/SF_IB
+ pixel_6394/PIX_OUT pixel_6394/CSA_VREF pixel
Xpixel_5660 pixel_5660/gring pixel_5660/VDD pixel_5660/GND pixel_5660/VREF pixel_5660/ROW_SEL
+ pixel_5660/NB1 pixel_5660/VBIAS pixel_5660/NB2 pixel_5660/AMP_IN pixel_5660/SF_IB
+ pixel_5660/PIX_OUT pixel_5660/CSA_VREF pixel
Xpixel_5671 pixel_5671/gring pixel_5671/VDD pixel_5671/GND pixel_5671/VREF pixel_5671/ROW_SEL
+ pixel_5671/NB1 pixel_5671/VBIAS pixel_5671/NB2 pixel_5671/AMP_IN pixel_5671/SF_IB
+ pixel_5671/PIX_OUT pixel_5671/CSA_VREF pixel
Xpixel_5682 pixel_5682/gring pixel_5682/VDD pixel_5682/GND pixel_5682/VREF pixel_5682/ROW_SEL
+ pixel_5682/NB1 pixel_5682/VBIAS pixel_5682/NB2 pixel_5682/AMP_IN pixel_5682/SF_IB
+ pixel_5682/PIX_OUT pixel_5682/CSA_VREF pixel
Xpixel_5693 pixel_5693/gring pixel_5693/VDD pixel_5693/GND pixel_5693/VREF pixel_5693/ROW_SEL
+ pixel_5693/NB1 pixel_5693/VBIAS pixel_5693/NB2 pixel_5693/AMP_IN pixel_5693/SF_IB
+ pixel_5693/PIX_OUT pixel_5693/CSA_VREF pixel
Xpixel_4970 pixel_4970/gring pixel_4970/VDD pixel_4970/GND pixel_4970/VREF pixel_4970/ROW_SEL
+ pixel_4970/NB1 pixel_4970/VBIAS pixel_4970/NB2 pixel_4970/AMP_IN pixel_4970/SF_IB
+ pixel_4970/PIX_OUT pixel_4970/CSA_VREF pixel
Xpixel_4981 pixel_4981/gring pixel_4981/VDD pixel_4981/GND pixel_4981/VREF pixel_4981/ROW_SEL
+ pixel_4981/NB1 pixel_4981/VBIAS pixel_4981/NB2 pixel_4981/AMP_IN pixel_4981/SF_IB
+ pixel_4981/PIX_OUT pixel_4981/CSA_VREF pixel
Xpixel_4992 pixel_4992/gring pixel_4992/VDD pixel_4992/GND pixel_4992/VREF pixel_4992/ROW_SEL
+ pixel_4992/NB1 pixel_4992/VBIAS pixel_4992/NB2 pixel_4992/AMP_IN pixel_4992/SF_IB
+ pixel_4992/PIX_OUT pixel_4992/CSA_VREF pixel
Xpixel_3009 pixel_3009/gring pixel_3009/VDD pixel_3009/GND pixel_3009/VREF pixel_3009/ROW_SEL
+ pixel_3009/NB1 pixel_3009/VBIAS pixel_3009/NB2 pixel_3009/AMP_IN pixel_3009/SF_IB
+ pixel_3009/PIX_OUT pixel_3009/CSA_VREF pixel
Xpixel_2308 pixel_2308/gring pixel_2308/VDD pixel_2308/GND pixel_2308/VREF pixel_2308/ROW_SEL
+ pixel_2308/NB1 pixel_2308/VBIAS pixel_2308/NB2 pixel_2308/AMP_IN pixel_2308/SF_IB
+ pixel_2308/PIX_OUT pixel_2308/CSA_VREF pixel
Xpixel_1607 pixel_1607/gring pixel_1607/VDD pixel_1607/GND pixel_1607/VREF pixel_1607/ROW_SEL
+ pixel_1607/NB1 pixel_1607/VBIAS pixel_1607/NB2 pixel_1607/AMP_IN pixel_1607/SF_IB
+ pixel_1607/PIX_OUT pixel_1607/CSA_VREF pixel
Xpixel_2319 pixel_2319/gring pixel_2319/VDD pixel_2319/GND pixel_2319/VREF pixel_2319/ROW_SEL
+ pixel_2319/NB1 pixel_2319/VBIAS pixel_2319/NB2 pixel_2319/AMP_IN pixel_2319/SF_IB
+ pixel_2319/PIX_OUT pixel_2319/CSA_VREF pixel
Xpixel_1629 pixel_1629/gring pixel_1629/VDD pixel_1629/GND pixel_1629/VREF pixel_1629/ROW_SEL
+ pixel_1629/NB1 pixel_1629/VBIAS pixel_1629/NB2 pixel_1629/AMP_IN pixel_1629/SF_IB
+ pixel_1629/PIX_OUT pixel_1629/CSA_VREF pixel
Xpixel_1618 pixel_1618/gring pixel_1618/VDD pixel_1618/GND pixel_1618/VREF pixel_1618/ROW_SEL
+ pixel_1618/NB1 pixel_1618/VBIAS pixel_1618/NB2 pixel_1618/AMP_IN pixel_1618/SF_IB
+ pixel_1618/PIX_OUT pixel_1618/CSA_VREF pixel
Xpixel_9915 pixel_9915/gring pixel_9915/VDD pixel_9915/GND pixel_9915/VREF pixel_9915/ROW_SEL
+ pixel_9915/NB1 pixel_9915/VBIAS pixel_9915/NB2 pixel_9915/AMP_IN pixel_9915/SF_IB
+ pixel_9915/PIX_OUT pixel_9915/CSA_VREF pixel
Xpixel_9904 pixel_9904/gring pixel_9904/VDD pixel_9904/GND pixel_9904/VREF pixel_9904/ROW_SEL
+ pixel_9904/NB1 pixel_9904/VBIAS pixel_9904/NB2 pixel_9904/AMP_IN pixel_9904/SF_IB
+ pixel_9904/PIX_OUT pixel_9904/CSA_VREF pixel
Xpixel_9937 pixel_9937/gring pixel_9937/VDD pixel_9937/GND pixel_9937/VREF pixel_9937/ROW_SEL
+ pixel_9937/NB1 pixel_9937/VBIAS pixel_9937/NB2 pixel_9937/AMP_IN pixel_9937/SF_IB
+ pixel_9937/PIX_OUT pixel_9937/CSA_VREF pixel
Xpixel_9926 pixel_9926/gring pixel_9926/VDD pixel_9926/GND pixel_9926/VREF pixel_9926/ROW_SEL
+ pixel_9926/NB1 pixel_9926/VBIAS pixel_9926/NB2 pixel_9926/AMP_IN pixel_9926/SF_IB
+ pixel_9926/PIX_OUT pixel_9926/CSA_VREF pixel
Xpixel_9948 pixel_9948/gring pixel_9948/VDD pixel_9948/GND pixel_9948/VREF pixel_9948/ROW_SEL
+ pixel_9948/NB1 pixel_9948/VBIAS pixel_9948/NB2 pixel_9948/AMP_IN pixel_9948/SF_IB
+ pixel_9948/PIX_OUT pixel_9948/CSA_VREF pixel
Xpixel_9959 pixel_9959/gring pixel_9959/VDD pixel_9959/GND pixel_9959/VREF pixel_9959/ROW_SEL
+ pixel_9959/NB1 pixel_9959/VBIAS pixel_9959/NB2 pixel_9959/AMP_IN pixel_9959/SF_IB
+ pixel_9959/PIX_OUT pixel_9959/CSA_VREF pixel
Xpixel_4200 pixel_4200/gring pixel_4200/VDD pixel_4200/GND pixel_4200/VREF pixel_4200/ROW_SEL
+ pixel_4200/NB1 pixel_4200/VBIAS pixel_4200/NB2 pixel_4200/AMP_IN pixel_4200/SF_IB
+ pixel_4200/PIX_OUT pixel_4200/CSA_VREF pixel
Xpixel_4211 pixel_4211/gring pixel_4211/VDD pixel_4211/GND pixel_4211/VREF pixel_4211/ROW_SEL
+ pixel_4211/NB1 pixel_4211/VBIAS pixel_4211/NB2 pixel_4211/AMP_IN pixel_4211/SF_IB
+ pixel_4211/PIX_OUT pixel_4211/CSA_VREF pixel
Xpixel_4222 pixel_4222/gring pixel_4222/VDD pixel_4222/GND pixel_4222/VREF pixel_4222/ROW_SEL
+ pixel_4222/NB1 pixel_4222/VBIAS pixel_4222/NB2 pixel_4222/AMP_IN pixel_4222/SF_IB
+ pixel_4222/PIX_OUT pixel_4222/CSA_VREF pixel
Xpixel_4233 pixel_4233/gring pixel_4233/VDD pixel_4233/GND pixel_4233/VREF pixel_4233/ROW_SEL
+ pixel_4233/NB1 pixel_4233/VBIAS pixel_4233/NB2 pixel_4233/AMP_IN pixel_4233/SF_IB
+ pixel_4233/PIX_OUT pixel_4233/CSA_VREF pixel
Xpixel_4244 pixel_4244/gring pixel_4244/VDD pixel_4244/GND pixel_4244/VREF pixel_4244/ROW_SEL
+ pixel_4244/NB1 pixel_4244/VBIAS pixel_4244/NB2 pixel_4244/AMP_IN pixel_4244/SF_IB
+ pixel_4244/PIX_OUT pixel_4244/CSA_VREF pixel
Xpixel_283 pixel_283/gring pixel_283/VDD pixel_283/GND pixel_283/VREF pixel_283/ROW_SEL
+ pixel_283/NB1 pixel_283/VBIAS pixel_283/NB2 pixel_283/AMP_IN pixel_283/SF_IB pixel_283/PIX_OUT
+ pixel_283/CSA_VREF pixel
Xpixel_272 pixel_272/gring pixel_272/VDD pixel_272/GND pixel_272/VREF pixel_272/ROW_SEL
+ pixel_272/NB1 pixel_272/VBIAS pixel_272/NB2 pixel_272/AMP_IN pixel_272/SF_IB pixel_272/PIX_OUT
+ pixel_272/CSA_VREF pixel
Xpixel_261 pixel_261/gring pixel_261/VDD pixel_261/GND pixel_261/VREF pixel_261/ROW_SEL
+ pixel_261/NB1 pixel_261/VBIAS pixel_261/NB2 pixel_261/AMP_IN pixel_261/SF_IB pixel_261/PIX_OUT
+ pixel_261/CSA_VREF pixel
Xpixel_250 pixel_250/gring pixel_250/VDD pixel_250/GND pixel_250/VREF pixel_250/ROW_SEL
+ pixel_250/NB1 pixel_250/VBIAS pixel_250/NB2 pixel_250/AMP_IN pixel_250/SF_IB pixel_250/PIX_OUT
+ pixel_250/CSA_VREF pixel
Xpixel_3543 pixel_3543/gring pixel_3543/VDD pixel_3543/GND pixel_3543/VREF pixel_3543/ROW_SEL
+ pixel_3543/NB1 pixel_3543/VBIAS pixel_3543/NB2 pixel_3543/AMP_IN pixel_3543/SF_IB
+ pixel_3543/PIX_OUT pixel_3543/CSA_VREF pixel
Xpixel_3532 pixel_3532/gring pixel_3532/VDD pixel_3532/GND pixel_3532/VREF pixel_3532/ROW_SEL
+ pixel_3532/NB1 pixel_3532/VBIAS pixel_3532/NB2 pixel_3532/AMP_IN pixel_3532/SF_IB
+ pixel_3532/PIX_OUT pixel_3532/CSA_VREF pixel
Xpixel_3521 pixel_3521/gring pixel_3521/VDD pixel_3521/GND pixel_3521/VREF pixel_3521/ROW_SEL
+ pixel_3521/NB1 pixel_3521/VBIAS pixel_3521/NB2 pixel_3521/AMP_IN pixel_3521/SF_IB
+ pixel_3521/PIX_OUT pixel_3521/CSA_VREF pixel
Xpixel_3510 pixel_3510/gring pixel_3510/VDD pixel_3510/GND pixel_3510/VREF pixel_3510/ROW_SEL
+ pixel_3510/NB1 pixel_3510/VBIAS pixel_3510/NB2 pixel_3510/AMP_IN pixel_3510/SF_IB
+ pixel_3510/PIX_OUT pixel_3510/CSA_VREF pixel
Xpixel_4255 pixel_4255/gring pixel_4255/VDD pixel_4255/GND pixel_4255/VREF pixel_4255/ROW_SEL
+ pixel_4255/NB1 pixel_4255/VBIAS pixel_4255/NB2 pixel_4255/AMP_IN pixel_4255/SF_IB
+ pixel_4255/PIX_OUT pixel_4255/CSA_VREF pixel
Xpixel_4266 pixel_4266/gring pixel_4266/VDD pixel_4266/GND pixel_4266/VREF pixel_4266/ROW_SEL
+ pixel_4266/NB1 pixel_4266/VBIAS pixel_4266/NB2 pixel_4266/AMP_IN pixel_4266/SF_IB
+ pixel_4266/PIX_OUT pixel_4266/CSA_VREF pixel
Xpixel_4277 pixel_4277/gring pixel_4277/VDD pixel_4277/GND pixel_4277/VREF pixel_4277/ROW_SEL
+ pixel_4277/NB1 pixel_4277/VBIAS pixel_4277/NB2 pixel_4277/AMP_IN pixel_4277/SF_IB
+ pixel_4277/PIX_OUT pixel_4277/CSA_VREF pixel
Xpixel_294 pixel_294/gring pixel_294/VDD pixel_294/GND pixel_294/VREF pixel_294/ROW_SEL
+ pixel_294/NB1 pixel_294/VBIAS pixel_294/NB2 pixel_294/AMP_IN pixel_294/SF_IB pixel_294/PIX_OUT
+ pixel_294/CSA_VREF pixel
Xpixel_2831 pixel_2831/gring pixel_2831/VDD pixel_2831/GND pixel_2831/VREF pixel_2831/ROW_SEL
+ pixel_2831/NB1 pixel_2831/VBIAS pixel_2831/NB2 pixel_2831/AMP_IN pixel_2831/SF_IB
+ pixel_2831/PIX_OUT pixel_2831/CSA_VREF pixel
Xpixel_2820 pixel_2820/gring pixel_2820/VDD pixel_2820/GND pixel_2820/VREF pixel_2820/ROW_SEL
+ pixel_2820/NB1 pixel_2820/VBIAS pixel_2820/NB2 pixel_2820/AMP_IN pixel_2820/SF_IB
+ pixel_2820/PIX_OUT pixel_2820/CSA_VREF pixel
Xpixel_3576 pixel_3576/gring pixel_3576/VDD pixel_3576/GND pixel_3576/VREF pixel_3576/ROW_SEL
+ pixel_3576/NB1 pixel_3576/VBIAS pixel_3576/NB2 pixel_3576/AMP_IN pixel_3576/SF_IB
+ pixel_3576/PIX_OUT pixel_3576/CSA_VREF pixel
Xpixel_3565 pixel_3565/gring pixel_3565/VDD pixel_3565/GND pixel_3565/VREF pixel_3565/ROW_SEL
+ pixel_3565/NB1 pixel_3565/VBIAS pixel_3565/NB2 pixel_3565/AMP_IN pixel_3565/SF_IB
+ pixel_3565/PIX_OUT pixel_3565/CSA_VREF pixel
Xpixel_3554 pixel_3554/gring pixel_3554/VDD pixel_3554/GND pixel_3554/VREF pixel_3554/ROW_SEL
+ pixel_3554/NB1 pixel_3554/VBIAS pixel_3554/NB2 pixel_3554/AMP_IN pixel_3554/SF_IB
+ pixel_3554/PIX_OUT pixel_3554/CSA_VREF pixel
Xpixel_4288 pixel_4288/gring pixel_4288/VDD pixel_4288/GND pixel_4288/VREF pixel_4288/ROW_SEL
+ pixel_4288/NB1 pixel_4288/VBIAS pixel_4288/NB2 pixel_4288/AMP_IN pixel_4288/SF_IB
+ pixel_4288/PIX_OUT pixel_4288/CSA_VREF pixel
Xpixel_4299 pixel_4299/gring pixel_4299/VDD pixel_4299/GND pixel_4299/VREF pixel_4299/ROW_SEL
+ pixel_4299/NB1 pixel_4299/VBIAS pixel_4299/NB2 pixel_4299/AMP_IN pixel_4299/SF_IB
+ pixel_4299/PIX_OUT pixel_4299/CSA_VREF pixel
Xpixel_2864 pixel_2864/gring pixel_2864/VDD pixel_2864/GND pixel_2864/VREF pixel_2864/ROW_SEL
+ pixel_2864/NB1 pixel_2864/VBIAS pixel_2864/NB2 pixel_2864/AMP_IN pixel_2864/SF_IB
+ pixel_2864/PIX_OUT pixel_2864/CSA_VREF pixel
Xpixel_2853 pixel_2853/gring pixel_2853/VDD pixel_2853/GND pixel_2853/VREF pixel_2853/ROW_SEL
+ pixel_2853/NB1 pixel_2853/VBIAS pixel_2853/NB2 pixel_2853/AMP_IN pixel_2853/SF_IB
+ pixel_2853/PIX_OUT pixel_2853/CSA_VREF pixel
Xpixel_2842 pixel_2842/gring pixel_2842/VDD pixel_2842/GND pixel_2842/VREF pixel_2842/ROW_SEL
+ pixel_2842/NB1 pixel_2842/VBIAS pixel_2842/NB2 pixel_2842/AMP_IN pixel_2842/SF_IB
+ pixel_2842/PIX_OUT pixel_2842/CSA_VREF pixel
Xpixel_3598 pixel_3598/gring pixel_3598/VDD pixel_3598/GND pixel_3598/VREF pixel_3598/ROW_SEL
+ pixel_3598/NB1 pixel_3598/VBIAS pixel_3598/NB2 pixel_3598/AMP_IN pixel_3598/SF_IB
+ pixel_3598/PIX_OUT pixel_3598/CSA_VREF pixel
Xpixel_3587 pixel_3587/gring pixel_3587/VDD pixel_3587/GND pixel_3587/VREF pixel_3587/ROW_SEL
+ pixel_3587/NB1 pixel_3587/VBIAS pixel_3587/NB2 pixel_3587/AMP_IN pixel_3587/SF_IB
+ pixel_3587/PIX_OUT pixel_3587/CSA_VREF pixel
Xpixel_2897 pixel_2897/gring pixel_2897/VDD pixel_2897/GND pixel_2897/VREF pixel_2897/ROW_SEL
+ pixel_2897/NB1 pixel_2897/VBIAS pixel_2897/NB2 pixel_2897/AMP_IN pixel_2897/SF_IB
+ pixel_2897/PIX_OUT pixel_2897/CSA_VREF pixel
Xpixel_2886 pixel_2886/gring pixel_2886/VDD pixel_2886/GND pixel_2886/VREF pixel_2886/ROW_SEL
+ pixel_2886/NB1 pixel_2886/VBIAS pixel_2886/NB2 pixel_2886/AMP_IN pixel_2886/SF_IB
+ pixel_2886/PIX_OUT pixel_2886/CSA_VREF pixel
Xpixel_2875 pixel_2875/gring pixel_2875/VDD pixel_2875/GND pixel_2875/VREF pixel_2875/ROW_SEL
+ pixel_2875/NB1 pixel_2875/VBIAS pixel_2875/NB2 pixel_2875/AMP_IN pixel_2875/SF_IB
+ pixel_2875/PIX_OUT pixel_2875/CSA_VREF pixel
Xpixel_6180 pixel_6180/gring pixel_6180/VDD pixel_6180/GND pixel_6180/VREF pixel_6180/ROW_SEL
+ pixel_6180/NB1 pixel_6180/VBIAS pixel_6180/NB2 pixel_6180/AMP_IN pixel_6180/SF_IB
+ pixel_6180/PIX_OUT pixel_6180/CSA_VREF pixel
Xpixel_6191 pixel_6191/gring pixel_6191/VDD pixel_6191/GND pixel_6191/VREF pixel_6191/ROW_SEL
+ pixel_6191/NB1 pixel_6191/VBIAS pixel_6191/NB2 pixel_6191/AMP_IN pixel_6191/SF_IB
+ pixel_6191/PIX_OUT pixel_6191/CSA_VREF pixel
Xpixel_5490 pixel_5490/gring pixel_5490/VDD pixel_5490/GND pixel_5490/VREF pixel_5490/ROW_SEL
+ pixel_5490/NB1 pixel_5490/VBIAS pixel_5490/NB2 pixel_5490/AMP_IN pixel_5490/SF_IB
+ pixel_5490/PIX_OUT pixel_5490/CSA_VREF pixel
Xpixel_7809 pixel_7809/gring pixel_7809/VDD pixel_7809/GND pixel_7809/VREF pixel_7809/ROW_SEL
+ pixel_7809/NB1 pixel_7809/VBIAS pixel_7809/NB2 pixel_7809/AMP_IN pixel_7809/SF_IB
+ pixel_7809/PIX_OUT pixel_7809/CSA_VREF pixel
Xpixel_2127 pixel_2127/gring pixel_2127/VDD pixel_2127/GND pixel_2127/VREF pixel_2127/ROW_SEL
+ pixel_2127/NB1 pixel_2127/VBIAS pixel_2127/NB2 pixel_2127/AMP_IN pixel_2127/SF_IB
+ pixel_2127/PIX_OUT pixel_2127/CSA_VREF pixel
Xpixel_2116 pixel_2116/gring pixel_2116/VDD pixel_2116/GND pixel_2116/VREF pixel_2116/ROW_SEL
+ pixel_2116/NB1 pixel_2116/VBIAS pixel_2116/NB2 pixel_2116/AMP_IN pixel_2116/SF_IB
+ pixel_2116/PIX_OUT pixel_2116/CSA_VREF pixel
Xpixel_2105 pixel_2105/gring pixel_2105/VDD pixel_2105/GND pixel_2105/VREF pixel_2105/ROW_SEL
+ pixel_2105/NB1 pixel_2105/VBIAS pixel_2105/NB2 pixel_2105/AMP_IN pixel_2105/SF_IB
+ pixel_2105/PIX_OUT pixel_2105/CSA_VREF pixel
Xpixel_1415 pixel_1415/gring pixel_1415/VDD pixel_1415/GND pixel_1415/VREF pixel_1415/ROW_SEL
+ pixel_1415/NB1 pixel_1415/VBIAS pixel_1415/NB2 pixel_1415/AMP_IN pixel_1415/SF_IB
+ pixel_1415/PIX_OUT pixel_1415/CSA_VREF pixel
Xpixel_1404 pixel_1404/gring pixel_1404/VDD pixel_1404/GND pixel_1404/VREF pixel_1404/ROW_SEL
+ pixel_1404/NB1 pixel_1404/VBIAS pixel_1404/NB2 pixel_1404/AMP_IN pixel_1404/SF_IB
+ pixel_1404/PIX_OUT pixel_1404/CSA_VREF pixel
Xpixel_2149 pixel_2149/gring pixel_2149/VDD pixel_2149/GND pixel_2149/VREF pixel_2149/ROW_SEL
+ pixel_2149/NB1 pixel_2149/VBIAS pixel_2149/NB2 pixel_2149/AMP_IN pixel_2149/SF_IB
+ pixel_2149/PIX_OUT pixel_2149/CSA_VREF pixel
Xpixel_2138 pixel_2138/gring pixel_2138/VDD pixel_2138/GND pixel_2138/VREF pixel_2138/ROW_SEL
+ pixel_2138/NB1 pixel_2138/VBIAS pixel_2138/NB2 pixel_2138/AMP_IN pixel_2138/SF_IB
+ pixel_2138/PIX_OUT pixel_2138/CSA_VREF pixel
Xpixel_1448 pixel_1448/gring pixel_1448/VDD pixel_1448/GND pixel_1448/VREF pixel_1448/ROW_SEL
+ pixel_1448/NB1 pixel_1448/VBIAS pixel_1448/NB2 pixel_1448/AMP_IN pixel_1448/SF_IB
+ pixel_1448/PIX_OUT pixel_1448/CSA_VREF pixel
Xpixel_1437 pixel_1437/gring pixel_1437/VDD pixel_1437/GND pixel_1437/VREF pixel_1437/ROW_SEL
+ pixel_1437/NB1 pixel_1437/VBIAS pixel_1437/NB2 pixel_1437/AMP_IN pixel_1437/SF_IB
+ pixel_1437/PIX_OUT pixel_1437/CSA_VREF pixel
Xpixel_1426 pixel_1426/gring pixel_1426/VDD pixel_1426/GND pixel_1426/VREF pixel_1426/ROW_SEL
+ pixel_1426/NB1 pixel_1426/VBIAS pixel_1426/NB2 pixel_1426/AMP_IN pixel_1426/SF_IB
+ pixel_1426/PIX_OUT pixel_1426/CSA_VREF pixel
Xpixel_1459 pixel_1459/gring pixel_1459/VDD pixel_1459/GND pixel_1459/VREF pixel_1459/ROW_SEL
+ pixel_1459/NB1 pixel_1459/VBIAS pixel_1459/NB2 pixel_1459/AMP_IN pixel_1459/SF_IB
+ pixel_1459/PIX_OUT pixel_1459/CSA_VREF pixel
Xpixel_9701 pixel_9701/gring pixel_9701/VDD pixel_9701/GND pixel_9701/VREF pixel_9701/ROW_SEL
+ pixel_9701/NB1 pixel_9701/VBIAS pixel_9701/NB2 pixel_9701/AMP_IN pixel_9701/SF_IB
+ pixel_9701/PIX_OUT pixel_9701/CSA_VREF pixel
Xpixel_9712 pixel_9712/gring pixel_9712/VDD pixel_9712/GND pixel_9712/VREF pixel_9712/ROW_SEL
+ pixel_9712/NB1 pixel_9712/VBIAS pixel_9712/NB2 pixel_9712/AMP_IN pixel_9712/SF_IB
+ pixel_9712/PIX_OUT pixel_9712/CSA_VREF pixel
Xpixel_9723 pixel_9723/gring pixel_9723/VDD pixel_9723/GND pixel_9723/VREF pixel_9723/ROW_SEL
+ pixel_9723/NB1 pixel_9723/VBIAS pixel_9723/NB2 pixel_9723/AMP_IN pixel_9723/SF_IB
+ pixel_9723/PIX_OUT pixel_9723/CSA_VREF pixel
Xpixel_9734 pixel_9734/gring pixel_9734/VDD pixel_9734/GND pixel_9734/VREF pixel_9734/ROW_SEL
+ pixel_9734/NB1 pixel_9734/VBIAS pixel_9734/NB2 pixel_9734/AMP_IN pixel_9734/SF_IB
+ pixel_9734/PIX_OUT pixel_9734/CSA_VREF pixel
Xpixel_9745 pixel_9745/gring pixel_9745/VDD pixel_9745/GND pixel_9745/VREF pixel_9745/ROW_SEL
+ pixel_9745/NB1 pixel_9745/VBIAS pixel_9745/NB2 pixel_9745/AMP_IN pixel_9745/SF_IB
+ pixel_9745/PIX_OUT pixel_9745/CSA_VREF pixel
Xpixel_9756 pixel_9756/gring pixel_9756/VDD pixel_9756/GND pixel_9756/VREF pixel_9756/ROW_SEL
+ pixel_9756/NB1 pixel_9756/VBIAS pixel_9756/NB2 pixel_9756/AMP_IN pixel_9756/SF_IB
+ pixel_9756/PIX_OUT pixel_9756/CSA_VREF pixel
Xpixel_9767 pixel_9767/gring pixel_9767/VDD pixel_9767/GND pixel_9767/VREF pixel_9767/ROW_SEL
+ pixel_9767/NB1 pixel_9767/VBIAS pixel_9767/NB2 pixel_9767/AMP_IN pixel_9767/SF_IB
+ pixel_9767/PIX_OUT pixel_9767/CSA_VREF pixel
Xpixel_9778 pixel_9778/gring pixel_9778/VDD pixel_9778/GND pixel_9778/VREF pixel_9778/ROW_SEL
+ pixel_9778/NB1 pixel_9778/VBIAS pixel_9778/NB2 pixel_9778/AMP_IN pixel_9778/SF_IB
+ pixel_9778/PIX_OUT pixel_9778/CSA_VREF pixel
Xpixel_9789 pixel_9789/gring pixel_9789/VDD pixel_9789/GND pixel_9789/VREF pixel_9789/ROW_SEL
+ pixel_9789/NB1 pixel_9789/VBIAS pixel_9789/NB2 pixel_9789/AMP_IN pixel_9789/SF_IB
+ pixel_9789/PIX_OUT pixel_9789/CSA_VREF pixel
Xpixel_4030 pixel_4030/gring pixel_4030/VDD pixel_4030/GND pixel_4030/VREF pixel_4030/ROW_SEL
+ pixel_4030/NB1 pixel_4030/VBIAS pixel_4030/NB2 pixel_4030/AMP_IN pixel_4030/SF_IB
+ pixel_4030/PIX_OUT pixel_4030/CSA_VREF pixel
Xpixel_4041 pixel_4041/gring pixel_4041/VDD pixel_4041/GND pixel_4041/VREF pixel_4041/ROW_SEL
+ pixel_4041/NB1 pixel_4041/VBIAS pixel_4041/NB2 pixel_4041/AMP_IN pixel_4041/SF_IB
+ pixel_4041/PIX_OUT pixel_4041/CSA_VREF pixel
Xpixel_4052 pixel_4052/gring pixel_4052/VDD pixel_4052/GND pixel_4052/VREF pixel_4052/ROW_SEL
+ pixel_4052/NB1 pixel_4052/VBIAS pixel_4052/NB2 pixel_4052/AMP_IN pixel_4052/SF_IB
+ pixel_4052/PIX_OUT pixel_4052/CSA_VREF pixel
Xpixel_3351 pixel_3351/gring pixel_3351/VDD pixel_3351/GND pixel_3351/VREF pixel_3351/ROW_SEL
+ pixel_3351/NB1 pixel_3351/VBIAS pixel_3351/NB2 pixel_3351/AMP_IN pixel_3351/SF_IB
+ pixel_3351/PIX_OUT pixel_3351/CSA_VREF pixel
Xpixel_3340 pixel_3340/gring pixel_3340/VDD pixel_3340/GND pixel_3340/VREF pixel_3340/ROW_SEL
+ pixel_3340/NB1 pixel_3340/VBIAS pixel_3340/NB2 pixel_3340/AMP_IN pixel_3340/SF_IB
+ pixel_3340/PIX_OUT pixel_3340/CSA_VREF pixel
Xpixel_4063 pixel_4063/gring pixel_4063/VDD pixel_4063/GND pixel_4063/VREF pixel_4063/ROW_SEL
+ pixel_4063/NB1 pixel_4063/VBIAS pixel_4063/NB2 pixel_4063/AMP_IN pixel_4063/SF_IB
+ pixel_4063/PIX_OUT pixel_4063/CSA_VREF pixel
Xpixel_4074 pixel_4074/gring pixel_4074/VDD pixel_4074/GND pixel_4074/VREF pixel_4074/ROW_SEL
+ pixel_4074/NB1 pixel_4074/VBIAS pixel_4074/NB2 pixel_4074/AMP_IN pixel_4074/SF_IB
+ pixel_4074/PIX_OUT pixel_4074/CSA_VREF pixel
Xpixel_4085 pixel_4085/gring pixel_4085/VDD pixel_4085/GND pixel_4085/VREF pixel_4085/ROW_SEL
+ pixel_4085/NB1 pixel_4085/VBIAS pixel_4085/NB2 pixel_4085/AMP_IN pixel_4085/SF_IB
+ pixel_4085/PIX_OUT pixel_4085/CSA_VREF pixel
Xpixel_4096 pixel_4096/gring pixel_4096/VDD pixel_4096/GND pixel_4096/VREF pixel_4096/ROW_SEL
+ pixel_4096/NB1 pixel_4096/VBIAS pixel_4096/NB2 pixel_4096/AMP_IN pixel_4096/SF_IB
+ pixel_4096/PIX_OUT pixel_4096/CSA_VREF pixel
Xpixel_3384 pixel_3384/gring pixel_3384/VDD pixel_3384/GND pixel_3384/VREF pixel_3384/ROW_SEL
+ pixel_3384/NB1 pixel_3384/VBIAS pixel_3384/NB2 pixel_3384/AMP_IN pixel_3384/SF_IB
+ pixel_3384/PIX_OUT pixel_3384/CSA_VREF pixel
Xpixel_3373 pixel_3373/gring pixel_3373/VDD pixel_3373/GND pixel_3373/VREF pixel_3373/ROW_SEL
+ pixel_3373/NB1 pixel_3373/VBIAS pixel_3373/NB2 pixel_3373/AMP_IN pixel_3373/SF_IB
+ pixel_3373/PIX_OUT pixel_3373/CSA_VREF pixel
Xpixel_3362 pixel_3362/gring pixel_3362/VDD pixel_3362/GND pixel_3362/VREF pixel_3362/ROW_SEL
+ pixel_3362/NB1 pixel_3362/VBIAS pixel_3362/NB2 pixel_3362/AMP_IN pixel_3362/SF_IB
+ pixel_3362/PIX_OUT pixel_3362/CSA_VREF pixel
Xpixel_2672 pixel_2672/gring pixel_2672/VDD pixel_2672/GND pixel_2672/VREF pixel_2672/ROW_SEL
+ pixel_2672/NB1 pixel_2672/VBIAS pixel_2672/NB2 pixel_2672/AMP_IN pixel_2672/SF_IB
+ pixel_2672/PIX_OUT pixel_2672/CSA_VREF pixel
Xpixel_2661 pixel_2661/gring pixel_2661/VDD pixel_2661/GND pixel_2661/VREF pixel_2661/ROW_SEL
+ pixel_2661/NB1 pixel_2661/VBIAS pixel_2661/NB2 pixel_2661/AMP_IN pixel_2661/SF_IB
+ pixel_2661/PIX_OUT pixel_2661/CSA_VREF pixel
Xpixel_2650 pixel_2650/gring pixel_2650/VDD pixel_2650/GND pixel_2650/VREF pixel_2650/ROW_SEL
+ pixel_2650/NB1 pixel_2650/VBIAS pixel_2650/NB2 pixel_2650/AMP_IN pixel_2650/SF_IB
+ pixel_2650/PIX_OUT pixel_2650/CSA_VREF pixel
Xpixel_3395 pixel_3395/gring pixel_3395/VDD pixel_3395/GND pixel_3395/VREF pixel_3395/ROW_SEL
+ pixel_3395/NB1 pixel_3395/VBIAS pixel_3395/NB2 pixel_3395/AMP_IN pixel_3395/SF_IB
+ pixel_3395/PIX_OUT pixel_3395/CSA_VREF pixel
Xpixel_1971 pixel_1971/gring pixel_1971/VDD pixel_1971/GND pixel_1971/VREF pixel_1971/ROW_SEL
+ pixel_1971/NB1 pixel_1971/VBIAS pixel_1971/NB2 pixel_1971/AMP_IN pixel_1971/SF_IB
+ pixel_1971/PIX_OUT pixel_1971/CSA_VREF pixel
Xpixel_1960 pixel_1960/gring pixel_1960/VDD pixel_1960/GND pixel_1960/VREF pixel_1960/ROW_SEL
+ pixel_1960/NB1 pixel_1960/VBIAS pixel_1960/NB2 pixel_1960/AMP_IN pixel_1960/SF_IB
+ pixel_1960/PIX_OUT pixel_1960/CSA_VREF pixel
Xpixel_2694 pixel_2694/gring pixel_2694/VDD pixel_2694/GND pixel_2694/VREF pixel_2694/ROW_SEL
+ pixel_2694/NB1 pixel_2694/VBIAS pixel_2694/NB2 pixel_2694/AMP_IN pixel_2694/SF_IB
+ pixel_2694/PIX_OUT pixel_2694/CSA_VREF pixel
Xpixel_2683 pixel_2683/gring pixel_2683/VDD pixel_2683/GND pixel_2683/VREF pixel_2683/ROW_SEL
+ pixel_2683/NB1 pixel_2683/VBIAS pixel_2683/NB2 pixel_2683/AMP_IN pixel_2683/SF_IB
+ pixel_2683/PIX_OUT pixel_2683/CSA_VREF pixel
Xpixel_1993 pixel_1993/gring pixel_1993/VDD pixel_1993/GND pixel_1993/VREF pixel_1993/ROW_SEL
+ pixel_1993/NB1 pixel_1993/VBIAS pixel_1993/NB2 pixel_1993/AMP_IN pixel_1993/SF_IB
+ pixel_1993/PIX_OUT pixel_1993/CSA_VREF pixel
Xpixel_1982 pixel_1982/gring pixel_1982/VDD pixel_1982/GND pixel_1982/VREF pixel_1982/ROW_SEL
+ pixel_1982/NB1 pixel_1982/VBIAS pixel_1982/NB2 pixel_1982/AMP_IN pixel_1982/SF_IB
+ pixel_1982/PIX_OUT pixel_1982/CSA_VREF pixel
Xpixel_9019 pixel_9019/gring pixel_9019/VDD pixel_9019/GND pixel_9019/VREF pixel_9019/ROW_SEL
+ pixel_9019/NB1 pixel_9019/VBIAS pixel_9019/NB2 pixel_9019/AMP_IN pixel_9019/SF_IB
+ pixel_9019/PIX_OUT pixel_9019/CSA_VREF pixel
Xpixel_9008 pixel_9008/gring pixel_9008/VDD pixel_9008/GND pixel_9008/VREF pixel_9008/ROW_SEL
+ pixel_9008/NB1 pixel_9008/VBIAS pixel_9008/NB2 pixel_9008/AMP_IN pixel_9008/SF_IB
+ pixel_9008/PIX_OUT pixel_9008/CSA_VREF pixel
Xpixel_8307 pixel_8307/gring pixel_8307/VDD pixel_8307/GND pixel_8307/VREF pixel_8307/ROW_SEL
+ pixel_8307/NB1 pixel_8307/VBIAS pixel_8307/NB2 pixel_8307/AMP_IN pixel_8307/SF_IB
+ pixel_8307/PIX_OUT pixel_8307/CSA_VREF pixel
Xpixel_8318 pixel_8318/gring pixel_8318/VDD pixel_8318/GND pixel_8318/VREF pixel_8318/ROW_SEL
+ pixel_8318/NB1 pixel_8318/VBIAS pixel_8318/NB2 pixel_8318/AMP_IN pixel_8318/SF_IB
+ pixel_8318/PIX_OUT pixel_8318/CSA_VREF pixel
Xpixel_8329 pixel_8329/gring pixel_8329/VDD pixel_8329/GND pixel_8329/VREF pixel_8329/ROW_SEL
+ pixel_8329/NB1 pixel_8329/VBIAS pixel_8329/NB2 pixel_8329/AMP_IN pixel_8329/SF_IB
+ pixel_8329/PIX_OUT pixel_8329/CSA_VREF pixel
Xpixel_7606 pixel_7606/gring pixel_7606/VDD pixel_7606/GND pixel_7606/VREF pixel_7606/ROW_SEL
+ pixel_7606/NB1 pixel_7606/VBIAS pixel_7606/NB2 pixel_7606/AMP_IN pixel_7606/SF_IB
+ pixel_7606/PIX_OUT pixel_7606/CSA_VREF pixel
Xpixel_7617 pixel_7617/gring pixel_7617/VDD pixel_7617/GND pixel_7617/VREF pixel_7617/ROW_SEL
+ pixel_7617/NB1 pixel_7617/VBIAS pixel_7617/NB2 pixel_7617/AMP_IN pixel_7617/SF_IB
+ pixel_7617/PIX_OUT pixel_7617/CSA_VREF pixel
Xpixel_7628 pixel_7628/gring pixel_7628/VDD pixel_7628/GND pixel_7628/VREF pixel_7628/ROW_SEL
+ pixel_7628/NB1 pixel_7628/VBIAS pixel_7628/NB2 pixel_7628/AMP_IN pixel_7628/SF_IB
+ pixel_7628/PIX_OUT pixel_7628/CSA_VREF pixel
Xpixel_7639 pixel_7639/gring pixel_7639/VDD pixel_7639/GND pixel_7639/VREF pixel_7639/ROW_SEL
+ pixel_7639/NB1 pixel_7639/VBIAS pixel_7639/NB2 pixel_7639/AMP_IN pixel_7639/SF_IB
+ pixel_7639/PIX_OUT pixel_7639/CSA_VREF pixel
Xpixel_6905 pixel_6905/gring pixel_6905/VDD pixel_6905/GND pixel_6905/VREF pixel_6905/ROW_SEL
+ pixel_6905/NB1 pixel_6905/VBIAS pixel_6905/NB2 pixel_6905/AMP_IN pixel_6905/SF_IB
+ pixel_6905/PIX_OUT pixel_6905/CSA_VREF pixel
Xpixel_6916 pixel_6916/gring pixel_6916/VDD pixel_6916/GND pixel_6916/VREF pixel_6916/ROW_SEL
+ pixel_6916/NB1 pixel_6916/VBIAS pixel_6916/NB2 pixel_6916/AMP_IN pixel_6916/SF_IB
+ pixel_6916/PIX_OUT pixel_6916/CSA_VREF pixel
Xpixel_6927 pixel_6927/gring pixel_6927/VDD pixel_6927/GND pixel_6927/VREF pixel_6927/ROW_SEL
+ pixel_6927/NB1 pixel_6927/VBIAS pixel_6927/NB2 pixel_6927/AMP_IN pixel_6927/SF_IB
+ pixel_6927/PIX_OUT pixel_6927/CSA_VREF pixel
Xpixel_19 pixel_19/gring pixel_19/VDD pixel_19/GND pixel_19/VREF pixel_19/ROW_SEL
+ pixel_19/NB1 pixel_19/VBIAS pixel_19/NB2 pixel_19/AMP_IN pixel_19/SF_IB pixel_19/PIX_OUT
+ pixel_19/CSA_VREF pixel
Xpixel_6938 pixel_6938/gring pixel_6938/VDD pixel_6938/GND pixel_6938/VREF pixel_6938/ROW_SEL
+ pixel_6938/NB1 pixel_6938/VBIAS pixel_6938/NB2 pixel_6938/AMP_IN pixel_6938/SF_IB
+ pixel_6938/PIX_OUT pixel_6938/CSA_VREF pixel
Xpixel_6949 pixel_6949/gring pixel_6949/VDD pixel_6949/GND pixel_6949/VREF pixel_6949/ROW_SEL
+ pixel_6949/NB1 pixel_6949/VBIAS pixel_6949/NB2 pixel_6949/AMP_IN pixel_6949/SF_IB
+ pixel_6949/PIX_OUT pixel_6949/CSA_VREF pixel
Xpixel_1223 pixel_1223/gring pixel_1223/VDD pixel_1223/GND pixel_1223/VREF pixel_1223/ROW_SEL
+ pixel_1223/NB1 pixel_1223/VBIAS pixel_1223/NB2 pixel_1223/AMP_IN pixel_1223/SF_IB
+ pixel_1223/PIX_OUT pixel_1223/CSA_VREF pixel
Xpixel_1212 pixel_1212/gring pixel_1212/VDD pixel_1212/GND pixel_1212/VREF pixel_1212/ROW_SEL
+ pixel_1212/NB1 pixel_1212/VBIAS pixel_1212/NB2 pixel_1212/AMP_IN pixel_1212/SF_IB
+ pixel_1212/PIX_OUT pixel_1212/CSA_VREF pixel
Xpixel_1201 pixel_1201/gring pixel_1201/VDD pixel_1201/GND pixel_1201/VREF pixel_1201/ROW_SEL
+ pixel_1201/NB1 pixel_1201/VBIAS pixel_1201/NB2 pixel_1201/AMP_IN pixel_1201/SF_IB
+ pixel_1201/PIX_OUT pixel_1201/CSA_VREF pixel
Xpixel_1267 pixel_1267/gring pixel_1267/VDD pixel_1267/GND pixel_1267/VREF pixel_1267/ROW_SEL
+ pixel_1267/NB1 pixel_1267/VBIAS pixel_1267/NB2 pixel_1267/AMP_IN pixel_1267/SF_IB
+ pixel_1267/PIX_OUT pixel_1267/CSA_VREF pixel
Xpixel_1256 pixel_1256/gring pixel_1256/VDD pixel_1256/GND pixel_1256/VREF pixel_1256/ROW_SEL
+ pixel_1256/NB1 pixel_1256/VBIAS pixel_1256/NB2 pixel_1256/AMP_IN pixel_1256/SF_IB
+ pixel_1256/PIX_OUT pixel_1256/CSA_VREF pixel
Xpixel_1245 pixel_1245/gring pixel_1245/VDD pixel_1245/GND pixel_1245/VREF pixel_1245/ROW_SEL
+ pixel_1245/NB1 pixel_1245/VBIAS pixel_1245/NB2 pixel_1245/AMP_IN pixel_1245/SF_IB
+ pixel_1245/PIX_OUT pixel_1245/CSA_VREF pixel
Xpixel_1234 pixel_1234/gring pixel_1234/VDD pixel_1234/GND pixel_1234/VREF pixel_1234/ROW_SEL
+ pixel_1234/NB1 pixel_1234/VBIAS pixel_1234/NB2 pixel_1234/AMP_IN pixel_1234/SF_IB
+ pixel_1234/PIX_OUT pixel_1234/CSA_VREF pixel
Xpixel_1289 pixel_1289/gring pixel_1289/VDD pixel_1289/GND pixel_1289/VREF pixel_1289/ROW_SEL
+ pixel_1289/NB1 pixel_1289/VBIAS pixel_1289/NB2 pixel_1289/AMP_IN pixel_1289/SF_IB
+ pixel_1289/PIX_OUT pixel_1289/CSA_VREF pixel
Xpixel_1278 pixel_1278/gring pixel_1278/VDD pixel_1278/GND pixel_1278/VREF pixel_1278/ROW_SEL
+ pixel_1278/NB1 pixel_1278/VBIAS pixel_1278/NB2 pixel_1278/AMP_IN pixel_1278/SF_IB
+ pixel_1278/PIX_OUT pixel_1278/CSA_VREF pixel
Xpixel_9531 pixel_9531/gring pixel_9531/VDD pixel_9531/GND pixel_9531/VREF pixel_9531/ROW_SEL
+ pixel_9531/NB1 pixel_9531/VBIAS pixel_9531/NB2 pixel_9531/AMP_IN pixel_9531/SF_IB
+ pixel_9531/PIX_OUT pixel_9531/CSA_VREF pixel
Xpixel_9520 pixel_9520/gring pixel_9520/VDD pixel_9520/GND pixel_9520/VREF pixel_9520/ROW_SEL
+ pixel_9520/NB1 pixel_9520/VBIAS pixel_9520/NB2 pixel_9520/AMP_IN pixel_9520/SF_IB
+ pixel_9520/PIX_OUT pixel_9520/CSA_VREF pixel
Xpixel_8830 pixel_8830/gring pixel_8830/VDD pixel_8830/GND pixel_8830/VREF pixel_8830/ROW_SEL
+ pixel_8830/NB1 pixel_8830/VBIAS pixel_8830/NB2 pixel_8830/AMP_IN pixel_8830/SF_IB
+ pixel_8830/PIX_OUT pixel_8830/CSA_VREF pixel
Xpixel_9575 pixel_9575/gring pixel_9575/VDD pixel_9575/GND pixel_9575/VREF pixel_9575/ROW_SEL
+ pixel_9575/NB1 pixel_9575/VBIAS pixel_9575/NB2 pixel_9575/AMP_IN pixel_9575/SF_IB
+ pixel_9575/PIX_OUT pixel_9575/CSA_VREF pixel
Xpixel_9564 pixel_9564/gring pixel_9564/VDD pixel_9564/GND pixel_9564/VREF pixel_9564/ROW_SEL
+ pixel_9564/NB1 pixel_9564/VBIAS pixel_9564/NB2 pixel_9564/AMP_IN pixel_9564/SF_IB
+ pixel_9564/PIX_OUT pixel_9564/CSA_VREF pixel
Xpixel_9553 pixel_9553/gring pixel_9553/VDD pixel_9553/GND pixel_9553/VREF pixel_9553/ROW_SEL
+ pixel_9553/NB1 pixel_9553/VBIAS pixel_9553/NB2 pixel_9553/AMP_IN pixel_9553/SF_IB
+ pixel_9553/PIX_OUT pixel_9553/CSA_VREF pixel
Xpixel_9542 pixel_9542/gring pixel_9542/VDD pixel_9542/GND pixel_9542/VREF pixel_9542/ROW_SEL
+ pixel_9542/NB1 pixel_9542/VBIAS pixel_9542/NB2 pixel_9542/AMP_IN pixel_9542/SF_IB
+ pixel_9542/PIX_OUT pixel_9542/CSA_VREF pixel
Xpixel_8863 pixel_8863/gring pixel_8863/VDD pixel_8863/GND pixel_8863/VREF pixel_8863/ROW_SEL
+ pixel_8863/NB1 pixel_8863/VBIAS pixel_8863/NB2 pixel_8863/AMP_IN pixel_8863/SF_IB
+ pixel_8863/PIX_OUT pixel_8863/CSA_VREF pixel
Xpixel_8852 pixel_8852/gring pixel_8852/VDD pixel_8852/GND pixel_8852/VREF pixel_8852/ROW_SEL
+ pixel_8852/NB1 pixel_8852/VBIAS pixel_8852/NB2 pixel_8852/AMP_IN pixel_8852/SF_IB
+ pixel_8852/PIX_OUT pixel_8852/CSA_VREF pixel
Xpixel_8841 pixel_8841/gring pixel_8841/VDD pixel_8841/GND pixel_8841/VREF pixel_8841/ROW_SEL
+ pixel_8841/NB1 pixel_8841/VBIAS pixel_8841/NB2 pixel_8841/AMP_IN pixel_8841/SF_IB
+ pixel_8841/PIX_OUT pixel_8841/CSA_VREF pixel
Xpixel_9597 pixel_9597/gring pixel_9597/VDD pixel_9597/GND pixel_9597/VREF pixel_9597/ROW_SEL
+ pixel_9597/NB1 pixel_9597/VBIAS pixel_9597/NB2 pixel_9597/AMP_IN pixel_9597/SF_IB
+ pixel_9597/PIX_OUT pixel_9597/CSA_VREF pixel
Xpixel_9586 pixel_9586/gring pixel_9586/VDD pixel_9586/GND pixel_9586/VREF pixel_9586/ROW_SEL
+ pixel_9586/NB1 pixel_9586/VBIAS pixel_9586/NB2 pixel_9586/AMP_IN pixel_9586/SF_IB
+ pixel_9586/PIX_OUT pixel_9586/CSA_VREF pixel
Xpixel_8896 pixel_8896/gring pixel_8896/VDD pixel_8896/GND pixel_8896/VREF pixel_8896/ROW_SEL
+ pixel_8896/NB1 pixel_8896/VBIAS pixel_8896/NB2 pixel_8896/AMP_IN pixel_8896/SF_IB
+ pixel_8896/PIX_OUT pixel_8896/CSA_VREF pixel
Xpixel_8885 pixel_8885/gring pixel_8885/VDD pixel_8885/GND pixel_8885/VREF pixel_8885/ROW_SEL
+ pixel_8885/NB1 pixel_8885/VBIAS pixel_8885/NB2 pixel_8885/AMP_IN pixel_8885/SF_IB
+ pixel_8885/PIX_OUT pixel_8885/CSA_VREF pixel
Xpixel_8874 pixel_8874/gring pixel_8874/VDD pixel_8874/GND pixel_8874/VREF pixel_8874/ROW_SEL
+ pixel_8874/NB1 pixel_8874/VBIAS pixel_8874/NB2 pixel_8874/AMP_IN pixel_8874/SF_IB
+ pixel_8874/PIX_OUT pixel_8874/CSA_VREF pixel
Xpixel_3192 pixel_3192/gring pixel_3192/VDD pixel_3192/GND pixel_3192/VREF pixel_3192/ROW_SEL
+ pixel_3192/NB1 pixel_3192/VBIAS pixel_3192/NB2 pixel_3192/AMP_IN pixel_3192/SF_IB
+ pixel_3192/PIX_OUT pixel_3192/CSA_VREF pixel
Xpixel_3181 pixel_3181/gring pixel_3181/VDD pixel_3181/GND pixel_3181/VREF pixel_3181/ROW_SEL
+ pixel_3181/NB1 pixel_3181/VBIAS pixel_3181/NB2 pixel_3181/AMP_IN pixel_3181/SF_IB
+ pixel_3181/PIX_OUT pixel_3181/CSA_VREF pixel
Xpixel_3170 pixel_3170/gring pixel_3170/VDD pixel_3170/GND pixel_3170/VREF pixel_3170/ROW_SEL
+ pixel_3170/NB1 pixel_3170/VBIAS pixel_3170/NB2 pixel_3170/AMP_IN pixel_3170/SF_IB
+ pixel_3170/PIX_OUT pixel_3170/CSA_VREF pixel
Xpixel_2491 pixel_2491/gring pixel_2491/VDD pixel_2491/GND pixel_2491/VREF pixel_2491/ROW_SEL
+ pixel_2491/NB1 pixel_2491/VBIAS pixel_2491/NB2 pixel_2491/AMP_IN pixel_2491/SF_IB
+ pixel_2491/PIX_OUT pixel_2491/CSA_VREF pixel
Xpixel_2480 pixel_2480/gring pixel_2480/VDD pixel_2480/GND pixel_2480/VREF pixel_2480/ROW_SEL
+ pixel_2480/NB1 pixel_2480/VBIAS pixel_2480/NB2 pixel_2480/AMP_IN pixel_2480/SF_IB
+ pixel_2480/PIX_OUT pixel_2480/CSA_VREF pixel
Xpixel_1790 pixel_1790/gring pixel_1790/VDD pixel_1790/GND pixel_1790/VREF pixel_1790/ROW_SEL
+ pixel_1790/NB1 pixel_1790/VBIAS pixel_1790/NB2 pixel_1790/AMP_IN pixel_1790/SF_IB
+ pixel_1790/PIX_OUT pixel_1790/CSA_VREF pixel
Xpixel_805 pixel_805/gring pixel_805/VDD pixel_805/GND pixel_805/VREF pixel_805/ROW_SEL
+ pixel_805/NB1 pixel_805/VBIAS pixel_805/NB2 pixel_805/AMP_IN pixel_805/SF_IB pixel_805/PIX_OUT
+ pixel_805/CSA_VREF pixel
Xpixel_838 pixel_838/gring pixel_838/VDD pixel_838/GND pixel_838/VREF pixel_838/ROW_SEL
+ pixel_838/NB1 pixel_838/VBIAS pixel_838/NB2 pixel_838/AMP_IN pixel_838/SF_IB pixel_838/PIX_OUT
+ pixel_838/CSA_VREF pixel
Xpixel_827 pixel_827/gring pixel_827/VDD pixel_827/GND pixel_827/VREF pixel_827/ROW_SEL
+ pixel_827/NB1 pixel_827/VBIAS pixel_827/NB2 pixel_827/AMP_IN pixel_827/SF_IB pixel_827/PIX_OUT
+ pixel_827/CSA_VREF pixel
Xpixel_816 pixel_816/gring pixel_816/VDD pixel_816/GND pixel_816/VREF pixel_816/ROW_SEL
+ pixel_816/NB1 pixel_816/VBIAS pixel_816/NB2 pixel_816/AMP_IN pixel_816/SF_IB pixel_816/PIX_OUT
+ pixel_816/CSA_VREF pixel
Xpixel_849 pixel_849/gring pixel_849/VDD pixel_849/GND pixel_849/VREF pixel_849/ROW_SEL
+ pixel_849/NB1 pixel_849/VBIAS pixel_849/NB2 pixel_849/AMP_IN pixel_849/SF_IB pixel_849/PIX_OUT
+ pixel_849/CSA_VREF pixel
Xpixel_8104 pixel_8104/gring pixel_8104/VDD pixel_8104/GND pixel_8104/VREF pixel_8104/ROW_SEL
+ pixel_8104/NB1 pixel_8104/VBIAS pixel_8104/NB2 pixel_8104/AMP_IN pixel_8104/SF_IB
+ pixel_8104/PIX_OUT pixel_8104/CSA_VREF pixel
Xpixel_8115 pixel_8115/gring pixel_8115/VDD pixel_8115/GND pixel_8115/VREF pixel_8115/ROW_SEL
+ pixel_8115/NB1 pixel_8115/VBIAS pixel_8115/NB2 pixel_8115/AMP_IN pixel_8115/SF_IB
+ pixel_8115/PIX_OUT pixel_8115/CSA_VREF pixel
Xpixel_8126 pixel_8126/gring pixel_8126/VDD pixel_8126/GND pixel_8126/VREF pixel_8126/ROW_SEL
+ pixel_8126/NB1 pixel_8126/VBIAS pixel_8126/NB2 pixel_8126/AMP_IN pixel_8126/SF_IB
+ pixel_8126/PIX_OUT pixel_8126/CSA_VREF pixel
Xpixel_8137 pixel_8137/gring pixel_8137/VDD pixel_8137/GND pixel_8137/VREF pixel_8137/ROW_SEL
+ pixel_8137/NB1 pixel_8137/VBIAS pixel_8137/NB2 pixel_8137/AMP_IN pixel_8137/SF_IB
+ pixel_8137/PIX_OUT pixel_8137/CSA_VREF pixel
Xpixel_8148 pixel_8148/gring pixel_8148/VDD pixel_8148/GND pixel_8148/VREF pixel_8148/ROW_SEL
+ pixel_8148/NB1 pixel_8148/VBIAS pixel_8148/NB2 pixel_8148/AMP_IN pixel_8148/SF_IB
+ pixel_8148/PIX_OUT pixel_8148/CSA_VREF pixel
Xpixel_8159 pixel_8159/gring pixel_8159/VDD pixel_8159/GND pixel_8159/VREF pixel_8159/ROW_SEL
+ pixel_8159/NB1 pixel_8159/VBIAS pixel_8159/NB2 pixel_8159/AMP_IN pixel_8159/SF_IB
+ pixel_8159/PIX_OUT pixel_8159/CSA_VREF pixel
Xpixel_7403 pixel_7403/gring pixel_7403/VDD pixel_7403/GND pixel_7403/VREF pixel_7403/ROW_SEL
+ pixel_7403/NB1 pixel_7403/VBIAS pixel_7403/NB2 pixel_7403/AMP_IN pixel_7403/SF_IB
+ pixel_7403/PIX_OUT pixel_7403/CSA_VREF pixel
Xpixel_7414 pixel_7414/gring pixel_7414/VDD pixel_7414/GND pixel_7414/VREF pixel_7414/ROW_SEL
+ pixel_7414/NB1 pixel_7414/VBIAS pixel_7414/NB2 pixel_7414/AMP_IN pixel_7414/SF_IB
+ pixel_7414/PIX_OUT pixel_7414/CSA_VREF pixel
Xpixel_7425 pixel_7425/gring pixel_7425/VDD pixel_7425/GND pixel_7425/VREF pixel_7425/ROW_SEL
+ pixel_7425/NB1 pixel_7425/VBIAS pixel_7425/NB2 pixel_7425/AMP_IN pixel_7425/SF_IB
+ pixel_7425/PIX_OUT pixel_7425/CSA_VREF pixel
Xpixel_7436 pixel_7436/gring pixel_7436/VDD pixel_7436/GND pixel_7436/VREF pixel_7436/ROW_SEL
+ pixel_7436/NB1 pixel_7436/VBIAS pixel_7436/NB2 pixel_7436/AMP_IN pixel_7436/SF_IB
+ pixel_7436/PIX_OUT pixel_7436/CSA_VREF pixel
Xpixel_7447 pixel_7447/gring pixel_7447/VDD pixel_7447/GND pixel_7447/VREF pixel_7447/ROW_SEL
+ pixel_7447/NB1 pixel_7447/VBIAS pixel_7447/NB2 pixel_7447/AMP_IN pixel_7447/SF_IB
+ pixel_7447/PIX_OUT pixel_7447/CSA_VREF pixel
Xpixel_6702 pixel_6702/gring pixel_6702/VDD pixel_6702/GND pixel_6702/VREF pixel_6702/ROW_SEL
+ pixel_6702/NB1 pixel_6702/VBIAS pixel_6702/NB2 pixel_6702/AMP_IN pixel_6702/SF_IB
+ pixel_6702/PIX_OUT pixel_6702/CSA_VREF pixel
Xpixel_7458 pixel_7458/gring pixel_7458/VDD pixel_7458/GND pixel_7458/VREF pixel_7458/ROW_SEL
+ pixel_7458/NB1 pixel_7458/VBIAS pixel_7458/NB2 pixel_7458/AMP_IN pixel_7458/SF_IB
+ pixel_7458/PIX_OUT pixel_7458/CSA_VREF pixel
Xpixel_7469 pixel_7469/gring pixel_7469/VDD pixel_7469/GND pixel_7469/VREF pixel_7469/ROW_SEL
+ pixel_7469/NB1 pixel_7469/VBIAS pixel_7469/NB2 pixel_7469/AMP_IN pixel_7469/SF_IB
+ pixel_7469/PIX_OUT pixel_7469/CSA_VREF pixel
Xpixel_6713 pixel_6713/gring pixel_6713/VDD pixel_6713/GND pixel_6713/VREF pixel_6713/ROW_SEL
+ pixel_6713/NB1 pixel_6713/VBIAS pixel_6713/NB2 pixel_6713/AMP_IN pixel_6713/SF_IB
+ pixel_6713/PIX_OUT pixel_6713/CSA_VREF pixel
Xpixel_6724 pixel_6724/gring pixel_6724/VDD pixel_6724/GND pixel_6724/VREF pixel_6724/ROW_SEL
+ pixel_6724/NB1 pixel_6724/VBIAS pixel_6724/NB2 pixel_6724/AMP_IN pixel_6724/SF_IB
+ pixel_6724/PIX_OUT pixel_6724/CSA_VREF pixel
Xpixel_6735 pixel_6735/gring pixel_6735/VDD pixel_6735/GND pixel_6735/VREF pixel_6735/ROW_SEL
+ pixel_6735/NB1 pixel_6735/VBIAS pixel_6735/NB2 pixel_6735/AMP_IN pixel_6735/SF_IB
+ pixel_6735/PIX_OUT pixel_6735/CSA_VREF pixel
Xpixel_6746 pixel_6746/gring pixel_6746/VDD pixel_6746/GND pixel_6746/VREF pixel_6746/ROW_SEL
+ pixel_6746/NB1 pixel_6746/VBIAS pixel_6746/NB2 pixel_6746/AMP_IN pixel_6746/SF_IB
+ pixel_6746/PIX_OUT pixel_6746/CSA_VREF pixel
Xpixel_6757 pixel_6757/gring pixel_6757/VDD pixel_6757/GND pixel_6757/VREF pixel_6757/ROW_SEL
+ pixel_6757/NB1 pixel_6757/VBIAS pixel_6757/NB2 pixel_6757/AMP_IN pixel_6757/SF_IB
+ pixel_6757/PIX_OUT pixel_6757/CSA_VREF pixel
Xpixel_6768 pixel_6768/gring pixel_6768/VDD pixel_6768/GND pixel_6768/VREF pixel_6768/ROW_SEL
+ pixel_6768/NB1 pixel_6768/VBIAS pixel_6768/NB2 pixel_6768/AMP_IN pixel_6768/SF_IB
+ pixel_6768/PIX_OUT pixel_6768/CSA_VREF pixel
Xpixel_6779 pixel_6779/gring pixel_6779/VDD pixel_6779/GND pixel_6779/VREF pixel_6779/ROW_SEL
+ pixel_6779/NB1 pixel_6779/VBIAS pixel_6779/NB2 pixel_6779/AMP_IN pixel_6779/SF_IB
+ pixel_6779/PIX_OUT pixel_6779/CSA_VREF pixel
Xpixel_1042 pixel_1042/gring pixel_1042/VDD pixel_1042/GND pixel_1042/VREF pixel_1042/ROW_SEL
+ pixel_1042/NB1 pixel_1042/VBIAS pixel_1042/NB2 pixel_1042/AMP_IN pixel_1042/SF_IB
+ pixel_1042/PIX_OUT pixel_1042/CSA_VREF pixel
Xpixel_1031 pixel_1031/gring pixel_1031/VDD pixel_1031/GND pixel_1031/VREF pixel_1031/ROW_SEL
+ pixel_1031/NB1 pixel_1031/VBIAS pixel_1031/NB2 pixel_1031/AMP_IN pixel_1031/SF_IB
+ pixel_1031/PIX_OUT pixel_1031/CSA_VREF pixel
Xpixel_1020 pixel_1020/gring pixel_1020/VDD pixel_1020/GND pixel_1020/VREF pixel_1020/ROW_SEL
+ pixel_1020/NB1 pixel_1020/VBIAS pixel_1020/NB2 pixel_1020/AMP_IN pixel_1020/SF_IB
+ pixel_1020/PIX_OUT pixel_1020/CSA_VREF pixel
Xpixel_1075 pixel_1075/gring pixel_1075/VDD pixel_1075/GND pixel_1075/VREF pixel_1075/ROW_SEL
+ pixel_1075/NB1 pixel_1075/VBIAS pixel_1075/NB2 pixel_1075/AMP_IN pixel_1075/SF_IB
+ pixel_1075/PIX_OUT pixel_1075/CSA_VREF pixel
Xpixel_1064 pixel_1064/gring pixel_1064/VDD pixel_1064/GND pixel_1064/VREF pixel_1064/ROW_SEL
+ pixel_1064/NB1 pixel_1064/VBIAS pixel_1064/NB2 pixel_1064/AMP_IN pixel_1064/SF_IB
+ pixel_1064/PIX_OUT pixel_1064/CSA_VREF pixel
Xpixel_1053 pixel_1053/gring pixel_1053/VDD pixel_1053/GND pixel_1053/VREF pixel_1053/ROW_SEL
+ pixel_1053/NB1 pixel_1053/VBIAS pixel_1053/NB2 pixel_1053/AMP_IN pixel_1053/SF_IB
+ pixel_1053/PIX_OUT pixel_1053/CSA_VREF pixel
Xpixel_1097 pixel_1097/gring pixel_1097/VDD pixel_1097/GND pixel_1097/VREF pixel_1097/ROW_SEL
+ pixel_1097/NB1 pixel_1097/VBIAS pixel_1097/NB2 pixel_1097/AMP_IN pixel_1097/SF_IB
+ pixel_1097/PIX_OUT pixel_1097/CSA_VREF pixel
Xpixel_1086 pixel_1086/gring pixel_1086/VDD pixel_1086/GND pixel_1086/VREF pixel_1086/ROW_SEL
+ pixel_1086/NB1 pixel_1086/VBIAS pixel_1086/NB2 pixel_1086/AMP_IN pixel_1086/SF_IB
+ pixel_1086/PIX_OUT pixel_1086/CSA_VREF pixel
Xpixel_9350 pixel_9350/gring pixel_9350/VDD pixel_9350/GND pixel_9350/VREF pixel_9350/ROW_SEL
+ pixel_9350/NB1 pixel_9350/VBIAS pixel_9350/NB2 pixel_9350/AMP_IN pixel_9350/SF_IB
+ pixel_9350/PIX_OUT pixel_9350/CSA_VREF pixel
Xpixel_9383 pixel_9383/gring pixel_9383/VDD pixel_9383/GND pixel_9383/VREF pixel_9383/ROW_SEL
+ pixel_9383/NB1 pixel_9383/VBIAS pixel_9383/NB2 pixel_9383/AMP_IN pixel_9383/SF_IB
+ pixel_9383/PIX_OUT pixel_9383/CSA_VREF pixel
Xpixel_9372 pixel_9372/gring pixel_9372/VDD pixel_9372/GND pixel_9372/VREF pixel_9372/ROW_SEL
+ pixel_9372/NB1 pixel_9372/VBIAS pixel_9372/NB2 pixel_9372/AMP_IN pixel_9372/SF_IB
+ pixel_9372/PIX_OUT pixel_9372/CSA_VREF pixel
Xpixel_9361 pixel_9361/gring pixel_9361/VDD pixel_9361/GND pixel_9361/VREF pixel_9361/ROW_SEL
+ pixel_9361/NB1 pixel_9361/VBIAS pixel_9361/NB2 pixel_9361/AMP_IN pixel_9361/SF_IB
+ pixel_9361/PIX_OUT pixel_9361/CSA_VREF pixel
Xpixel_8671 pixel_8671/gring pixel_8671/VDD pixel_8671/GND pixel_8671/VREF pixel_8671/ROW_SEL
+ pixel_8671/NB1 pixel_8671/VBIAS pixel_8671/NB2 pixel_8671/AMP_IN pixel_8671/SF_IB
+ pixel_8671/PIX_OUT pixel_8671/CSA_VREF pixel
Xpixel_8660 pixel_8660/gring pixel_8660/VDD pixel_8660/GND pixel_8660/VREF pixel_8660/ROW_SEL
+ pixel_8660/NB1 pixel_8660/VBIAS pixel_8660/NB2 pixel_8660/AMP_IN pixel_8660/SF_IB
+ pixel_8660/PIX_OUT pixel_8660/CSA_VREF pixel
Xpixel_9394 pixel_9394/gring pixel_9394/VDD pixel_9394/GND pixel_9394/VREF pixel_9394/ROW_SEL
+ pixel_9394/NB1 pixel_9394/VBIAS pixel_9394/NB2 pixel_9394/AMP_IN pixel_9394/SF_IB
+ pixel_9394/PIX_OUT pixel_9394/CSA_VREF pixel
Xpixel_8693 pixel_8693/gring pixel_8693/VDD pixel_8693/GND pixel_8693/VREF pixel_8693/ROW_SEL
+ pixel_8693/NB1 pixel_8693/VBIAS pixel_8693/NB2 pixel_8693/AMP_IN pixel_8693/SF_IB
+ pixel_8693/PIX_OUT pixel_8693/CSA_VREF pixel
Xpixel_8682 pixel_8682/gring pixel_8682/VDD pixel_8682/GND pixel_8682/VREF pixel_8682/ROW_SEL
+ pixel_8682/NB1 pixel_8682/VBIAS pixel_8682/NB2 pixel_8682/AMP_IN pixel_8682/SF_IB
+ pixel_8682/PIX_OUT pixel_8682/CSA_VREF pixel
Xpixel_7970 pixel_7970/gring pixel_7970/VDD pixel_7970/GND pixel_7970/VREF pixel_7970/ROW_SEL
+ pixel_7970/NB1 pixel_7970/VBIAS pixel_7970/NB2 pixel_7970/AMP_IN pixel_7970/SF_IB
+ pixel_7970/PIX_OUT pixel_7970/CSA_VREF pixel
Xpixel_7981 pixel_7981/gring pixel_7981/VDD pixel_7981/GND pixel_7981/VREF pixel_7981/ROW_SEL
+ pixel_7981/NB1 pixel_7981/VBIAS pixel_7981/NB2 pixel_7981/AMP_IN pixel_7981/SF_IB
+ pixel_7981/PIX_OUT pixel_7981/CSA_VREF pixel
Xpixel_7992 pixel_7992/gring pixel_7992/VDD pixel_7992/GND pixel_7992/VREF pixel_7992/ROW_SEL
+ pixel_7992/NB1 pixel_7992/VBIAS pixel_7992/NB2 pixel_7992/AMP_IN pixel_7992/SF_IB
+ pixel_7992/PIX_OUT pixel_7992/CSA_VREF pixel
Xpixel_6009 pixel_6009/gring pixel_6009/VDD pixel_6009/GND pixel_6009/VREF pixel_6009/ROW_SEL
+ pixel_6009/NB1 pixel_6009/VBIAS pixel_6009/NB2 pixel_6009/AMP_IN pixel_6009/SF_IB
+ pixel_6009/PIX_OUT pixel_6009/CSA_VREF pixel
Xpixel_5308 pixel_5308/gring pixel_5308/VDD pixel_5308/GND pixel_5308/VREF pixel_5308/ROW_SEL
+ pixel_5308/NB1 pixel_5308/VBIAS pixel_5308/NB2 pixel_5308/AMP_IN pixel_5308/SF_IB
+ pixel_5308/PIX_OUT pixel_5308/CSA_VREF pixel
Xpixel_5319 pixel_5319/gring pixel_5319/VDD pixel_5319/GND pixel_5319/VREF pixel_5319/ROW_SEL
+ pixel_5319/NB1 pixel_5319/VBIAS pixel_5319/NB2 pixel_5319/AMP_IN pixel_5319/SF_IB
+ pixel_5319/PIX_OUT pixel_5319/CSA_VREF pixel
Xpixel_613 pixel_613/gring pixel_613/VDD pixel_613/GND pixel_613/VREF pixel_613/ROW_SEL
+ pixel_613/NB1 pixel_613/VBIAS pixel_613/NB2 pixel_613/AMP_IN pixel_613/SF_IB pixel_613/PIX_OUT
+ pixel_613/CSA_VREF pixel
Xpixel_602 pixel_602/gring pixel_602/VDD pixel_602/GND pixel_602/VREF pixel_602/ROW_SEL
+ pixel_602/NB1 pixel_602/VBIAS pixel_602/NB2 pixel_602/AMP_IN pixel_602/SF_IB pixel_602/PIX_OUT
+ pixel_602/CSA_VREF pixel
Xpixel_4607 pixel_4607/gring pixel_4607/VDD pixel_4607/GND pixel_4607/VREF pixel_4607/ROW_SEL
+ pixel_4607/NB1 pixel_4607/VBIAS pixel_4607/NB2 pixel_4607/AMP_IN pixel_4607/SF_IB
+ pixel_4607/PIX_OUT pixel_4607/CSA_VREF pixel
Xpixel_4618 pixel_4618/gring pixel_4618/VDD pixel_4618/GND pixel_4618/VREF pixel_4618/ROW_SEL
+ pixel_4618/NB1 pixel_4618/VBIAS pixel_4618/NB2 pixel_4618/AMP_IN pixel_4618/SF_IB
+ pixel_4618/PIX_OUT pixel_4618/CSA_VREF pixel
Xpixel_657 pixel_657/gring pixel_657/VDD pixel_657/GND pixel_657/VREF pixel_657/ROW_SEL
+ pixel_657/NB1 pixel_657/VBIAS pixel_657/NB2 pixel_657/AMP_IN pixel_657/SF_IB pixel_657/PIX_OUT
+ pixel_657/CSA_VREF pixel
Xpixel_646 pixel_646/gring pixel_646/VDD pixel_646/GND pixel_646/VREF pixel_646/ROW_SEL
+ pixel_646/NB1 pixel_646/VBIAS pixel_646/NB2 pixel_646/AMP_IN pixel_646/SF_IB pixel_646/PIX_OUT
+ pixel_646/CSA_VREF pixel
Xpixel_635 pixel_635/gring pixel_635/VDD pixel_635/GND pixel_635/VREF pixel_635/ROW_SEL
+ pixel_635/NB1 pixel_635/VBIAS pixel_635/NB2 pixel_635/AMP_IN pixel_635/SF_IB pixel_635/PIX_OUT
+ pixel_635/CSA_VREF pixel
Xpixel_624 pixel_624/gring pixel_624/VDD pixel_624/GND pixel_624/VREF pixel_624/ROW_SEL
+ pixel_624/NB1 pixel_624/VBIAS pixel_624/NB2 pixel_624/AMP_IN pixel_624/SF_IB pixel_624/PIX_OUT
+ pixel_624/CSA_VREF pixel
Xpixel_4629 pixel_4629/gring pixel_4629/VDD pixel_4629/GND pixel_4629/VREF pixel_4629/ROW_SEL
+ pixel_4629/NB1 pixel_4629/VBIAS pixel_4629/NB2 pixel_4629/AMP_IN pixel_4629/SF_IB
+ pixel_4629/PIX_OUT pixel_4629/CSA_VREF pixel
Xpixel_3906 pixel_3906/gring pixel_3906/VDD pixel_3906/GND pixel_3906/VREF pixel_3906/ROW_SEL
+ pixel_3906/NB1 pixel_3906/VBIAS pixel_3906/NB2 pixel_3906/AMP_IN pixel_3906/SF_IB
+ pixel_3906/PIX_OUT pixel_3906/CSA_VREF pixel
Xpixel_3917 pixel_3917/gring pixel_3917/VDD pixel_3917/GND pixel_3917/VREF pixel_3917/ROW_SEL
+ pixel_3917/NB1 pixel_3917/VBIAS pixel_3917/NB2 pixel_3917/AMP_IN pixel_3917/SF_IB
+ pixel_3917/PIX_OUT pixel_3917/CSA_VREF pixel
Xpixel_679 pixel_679/gring pixel_679/VDD pixel_679/GND pixel_679/VREF pixel_679/ROW_SEL
+ pixel_679/NB1 pixel_679/VBIAS pixel_679/NB2 pixel_679/AMP_IN pixel_679/SF_IB pixel_679/PIX_OUT
+ pixel_679/CSA_VREF pixel
Xpixel_668 pixel_668/gring pixel_668/VDD pixel_668/GND pixel_668/VREF pixel_668/ROW_SEL
+ pixel_668/NB1 pixel_668/VBIAS pixel_668/NB2 pixel_668/AMP_IN pixel_668/SF_IB pixel_668/PIX_OUT
+ pixel_668/CSA_VREF pixel
Xpixel_3928 pixel_3928/gring pixel_3928/VDD pixel_3928/GND pixel_3928/VREF pixel_3928/ROW_SEL
+ pixel_3928/NB1 pixel_3928/VBIAS pixel_3928/NB2 pixel_3928/AMP_IN pixel_3928/SF_IB
+ pixel_3928/PIX_OUT pixel_3928/CSA_VREF pixel
Xpixel_3939 pixel_3939/gring pixel_3939/VDD pixel_3939/GND pixel_3939/VREF pixel_3939/ROW_SEL
+ pixel_3939/NB1 pixel_3939/VBIAS pixel_3939/NB2 pixel_3939/AMP_IN pixel_3939/SF_IB
+ pixel_3939/PIX_OUT pixel_3939/CSA_VREF pixel
Xpixel_7200 pixel_7200/gring pixel_7200/VDD pixel_7200/GND pixel_7200/VREF pixel_7200/ROW_SEL
+ pixel_7200/NB1 pixel_7200/VBIAS pixel_7200/NB2 pixel_7200/AMP_IN pixel_7200/SF_IB
+ pixel_7200/PIX_OUT pixel_7200/CSA_VREF pixel
Xpixel_7211 pixel_7211/gring pixel_7211/VDD pixel_7211/GND pixel_7211/VREF pixel_7211/ROW_SEL
+ pixel_7211/NB1 pixel_7211/VBIAS pixel_7211/NB2 pixel_7211/AMP_IN pixel_7211/SF_IB
+ pixel_7211/PIX_OUT pixel_7211/CSA_VREF pixel
Xpixel_7222 pixel_7222/gring pixel_7222/VDD pixel_7222/GND pixel_7222/VREF pixel_7222/ROW_SEL
+ pixel_7222/NB1 pixel_7222/VBIAS pixel_7222/NB2 pixel_7222/AMP_IN pixel_7222/SF_IB
+ pixel_7222/PIX_OUT pixel_7222/CSA_VREF pixel
Xpixel_7233 pixel_7233/gring pixel_7233/VDD pixel_7233/GND pixel_7233/VREF pixel_7233/ROW_SEL
+ pixel_7233/NB1 pixel_7233/VBIAS pixel_7233/NB2 pixel_7233/AMP_IN pixel_7233/SF_IB
+ pixel_7233/PIX_OUT pixel_7233/CSA_VREF pixel
Xpixel_7244 pixel_7244/gring pixel_7244/VDD pixel_7244/GND pixel_7244/VREF pixel_7244/ROW_SEL
+ pixel_7244/NB1 pixel_7244/VBIAS pixel_7244/NB2 pixel_7244/AMP_IN pixel_7244/SF_IB
+ pixel_7244/PIX_OUT pixel_7244/CSA_VREF pixel
Xpixel_7255 pixel_7255/gring pixel_7255/VDD pixel_7255/GND pixel_7255/VREF pixel_7255/ROW_SEL
+ pixel_7255/NB1 pixel_7255/VBIAS pixel_7255/NB2 pixel_7255/AMP_IN pixel_7255/SF_IB
+ pixel_7255/PIX_OUT pixel_7255/CSA_VREF pixel
Xpixel_6510 pixel_6510/gring pixel_6510/VDD pixel_6510/GND pixel_6510/VREF pixel_6510/ROW_SEL
+ pixel_6510/NB1 pixel_6510/VBIAS pixel_6510/NB2 pixel_6510/AMP_IN pixel_6510/SF_IB
+ pixel_6510/PIX_OUT pixel_6510/CSA_VREF pixel
Xpixel_6521 pixel_6521/gring pixel_6521/VDD pixel_6521/GND pixel_6521/VREF pixel_6521/ROW_SEL
+ pixel_6521/NB1 pixel_6521/VBIAS pixel_6521/NB2 pixel_6521/AMP_IN pixel_6521/SF_IB
+ pixel_6521/PIX_OUT pixel_6521/CSA_VREF pixel
Xpixel_7266 pixel_7266/gring pixel_7266/VDD pixel_7266/GND pixel_7266/VREF pixel_7266/ROW_SEL
+ pixel_7266/NB1 pixel_7266/VBIAS pixel_7266/NB2 pixel_7266/AMP_IN pixel_7266/SF_IB
+ pixel_7266/PIX_OUT pixel_7266/CSA_VREF pixel
Xpixel_7277 pixel_7277/gring pixel_7277/VDD pixel_7277/GND pixel_7277/VREF pixel_7277/ROW_SEL
+ pixel_7277/NB1 pixel_7277/VBIAS pixel_7277/NB2 pixel_7277/AMP_IN pixel_7277/SF_IB
+ pixel_7277/PIX_OUT pixel_7277/CSA_VREF pixel
Xpixel_7288 pixel_7288/gring pixel_7288/VDD pixel_7288/GND pixel_7288/VREF pixel_7288/ROW_SEL
+ pixel_7288/NB1 pixel_7288/VBIAS pixel_7288/NB2 pixel_7288/AMP_IN pixel_7288/SF_IB
+ pixel_7288/PIX_OUT pixel_7288/CSA_VREF pixel
Xpixel_7299 pixel_7299/gring pixel_7299/VDD pixel_7299/GND pixel_7299/VREF pixel_7299/ROW_SEL
+ pixel_7299/NB1 pixel_7299/VBIAS pixel_7299/NB2 pixel_7299/AMP_IN pixel_7299/SF_IB
+ pixel_7299/PIX_OUT pixel_7299/CSA_VREF pixel
Xpixel_6532 pixel_6532/gring pixel_6532/VDD pixel_6532/GND pixel_6532/VREF pixel_6532/ROW_SEL
+ pixel_6532/NB1 pixel_6532/VBIAS pixel_6532/NB2 pixel_6532/AMP_IN pixel_6532/SF_IB
+ pixel_6532/PIX_OUT pixel_6532/CSA_VREF pixel
Xpixel_6543 pixel_6543/gring pixel_6543/VDD pixel_6543/GND pixel_6543/VREF pixel_6543/ROW_SEL
+ pixel_6543/NB1 pixel_6543/VBIAS pixel_6543/NB2 pixel_6543/AMP_IN pixel_6543/SF_IB
+ pixel_6543/PIX_OUT pixel_6543/CSA_VREF pixel
Xpixel_6554 pixel_6554/gring pixel_6554/VDD pixel_6554/GND pixel_6554/VREF pixel_6554/ROW_SEL
+ pixel_6554/NB1 pixel_6554/VBIAS pixel_6554/NB2 pixel_6554/AMP_IN pixel_6554/SF_IB
+ pixel_6554/PIX_OUT pixel_6554/CSA_VREF pixel
Xpixel_6565 pixel_6565/gring pixel_6565/VDD pixel_6565/GND pixel_6565/VREF pixel_6565/ROW_SEL
+ pixel_6565/NB1 pixel_6565/VBIAS pixel_6565/NB2 pixel_6565/AMP_IN pixel_6565/SF_IB
+ pixel_6565/PIX_OUT pixel_6565/CSA_VREF pixel
Xpixel_6576 pixel_6576/gring pixel_6576/VDD pixel_6576/GND pixel_6576/VREF pixel_6576/ROW_SEL
+ pixel_6576/NB1 pixel_6576/VBIAS pixel_6576/NB2 pixel_6576/AMP_IN pixel_6576/SF_IB
+ pixel_6576/PIX_OUT pixel_6576/CSA_VREF pixel
Xpixel_6587 pixel_6587/gring pixel_6587/VDD pixel_6587/GND pixel_6587/VREF pixel_6587/ROW_SEL
+ pixel_6587/NB1 pixel_6587/VBIAS pixel_6587/NB2 pixel_6587/AMP_IN pixel_6587/SF_IB
+ pixel_6587/PIX_OUT pixel_6587/CSA_VREF pixel
Xpixel_5820 pixel_5820/gring pixel_5820/VDD pixel_5820/GND pixel_5820/VREF pixel_5820/ROW_SEL
+ pixel_5820/NB1 pixel_5820/VBIAS pixel_5820/NB2 pixel_5820/AMP_IN pixel_5820/SF_IB
+ pixel_5820/PIX_OUT pixel_5820/CSA_VREF pixel
Xpixel_5831 pixel_5831/gring pixel_5831/VDD pixel_5831/GND pixel_5831/VREF pixel_5831/ROW_SEL
+ pixel_5831/NB1 pixel_5831/VBIAS pixel_5831/NB2 pixel_5831/AMP_IN pixel_5831/SF_IB
+ pixel_5831/PIX_OUT pixel_5831/CSA_VREF pixel
Xpixel_5842 pixel_5842/gring pixel_5842/VDD pixel_5842/GND pixel_5842/VREF pixel_5842/ROW_SEL
+ pixel_5842/NB1 pixel_5842/VBIAS pixel_5842/NB2 pixel_5842/AMP_IN pixel_5842/SF_IB
+ pixel_5842/PIX_OUT pixel_5842/CSA_VREF pixel
Xpixel_6598 pixel_6598/gring pixel_6598/VDD pixel_6598/GND pixel_6598/VREF pixel_6598/ROW_SEL
+ pixel_6598/NB1 pixel_6598/VBIAS pixel_6598/NB2 pixel_6598/AMP_IN pixel_6598/SF_IB
+ pixel_6598/PIX_OUT pixel_6598/CSA_VREF pixel
Xpixel_5853 pixel_5853/gring pixel_5853/VDD pixel_5853/GND pixel_5853/VREF pixel_5853/ROW_SEL
+ pixel_5853/NB1 pixel_5853/VBIAS pixel_5853/NB2 pixel_5853/AMP_IN pixel_5853/SF_IB
+ pixel_5853/PIX_OUT pixel_5853/CSA_VREF pixel
Xpixel_5864 pixel_5864/gring pixel_5864/VDD pixel_5864/GND pixel_5864/VREF pixel_5864/ROW_SEL
+ pixel_5864/NB1 pixel_5864/VBIAS pixel_5864/NB2 pixel_5864/AMP_IN pixel_5864/SF_IB
+ pixel_5864/PIX_OUT pixel_5864/CSA_VREF pixel
Xpixel_5875 pixel_5875/gring pixel_5875/VDD pixel_5875/GND pixel_5875/VREF pixel_5875/ROW_SEL
+ pixel_5875/NB1 pixel_5875/VBIAS pixel_5875/NB2 pixel_5875/AMP_IN pixel_5875/SF_IB
+ pixel_5875/PIX_OUT pixel_5875/CSA_VREF pixel
Xpixel_5886 pixel_5886/gring pixel_5886/VDD pixel_5886/GND pixel_5886/VREF pixel_5886/ROW_SEL
+ pixel_5886/NB1 pixel_5886/VBIAS pixel_5886/NB2 pixel_5886/AMP_IN pixel_5886/SF_IB
+ pixel_5886/PIX_OUT pixel_5886/CSA_VREF pixel
Xpixel_5897 pixel_5897/gring pixel_5897/VDD pixel_5897/GND pixel_5897/VREF pixel_5897/ROW_SEL
+ pixel_5897/NB1 pixel_5897/VBIAS pixel_5897/NB2 pixel_5897/AMP_IN pixel_5897/SF_IB
+ pixel_5897/PIX_OUT pixel_5897/CSA_VREF pixel
Xpixel_9191 pixel_9191/gring pixel_9191/VDD pixel_9191/GND pixel_9191/VREF pixel_9191/ROW_SEL
+ pixel_9191/NB1 pixel_9191/VBIAS pixel_9191/NB2 pixel_9191/AMP_IN pixel_9191/SF_IB
+ pixel_9191/PIX_OUT pixel_9191/CSA_VREF pixel
Xpixel_9180 pixel_9180/gring pixel_9180/VDD pixel_9180/GND pixel_9180/VREF pixel_9180/ROW_SEL
+ pixel_9180/NB1 pixel_9180/VBIAS pixel_9180/NB2 pixel_9180/AMP_IN pixel_9180/SF_IB
+ pixel_9180/PIX_OUT pixel_9180/CSA_VREF pixel
Xpixel_8490 pixel_8490/gring pixel_8490/VDD pixel_8490/GND pixel_8490/VREF pixel_8490/ROW_SEL
+ pixel_8490/NB1 pixel_8490/VBIAS pixel_8490/NB2 pixel_8490/AMP_IN pixel_8490/SF_IB
+ pixel_8490/PIX_OUT pixel_8490/CSA_VREF pixel
Xpixel_5105 pixel_5105/gring pixel_5105/VDD pixel_5105/GND pixel_5105/VREF pixel_5105/ROW_SEL
+ pixel_5105/NB1 pixel_5105/VBIAS pixel_5105/NB2 pixel_5105/AMP_IN pixel_5105/SF_IB
+ pixel_5105/PIX_OUT pixel_5105/CSA_VREF pixel
Xpixel_5116 pixel_5116/gring pixel_5116/VDD pixel_5116/GND pixel_5116/VREF pixel_5116/ROW_SEL
+ pixel_5116/NB1 pixel_5116/VBIAS pixel_5116/NB2 pixel_5116/AMP_IN pixel_5116/SF_IB
+ pixel_5116/PIX_OUT pixel_5116/CSA_VREF pixel
Xpixel_5127 pixel_5127/gring pixel_5127/VDD pixel_5127/GND pixel_5127/VREF pixel_5127/ROW_SEL
+ pixel_5127/NB1 pixel_5127/VBIAS pixel_5127/NB2 pixel_5127/AMP_IN pixel_5127/SF_IB
+ pixel_5127/PIX_OUT pixel_5127/CSA_VREF pixel
Xpixel_5138 pixel_5138/gring pixel_5138/VDD pixel_5138/GND pixel_5138/VREF pixel_5138/ROW_SEL
+ pixel_5138/NB1 pixel_5138/VBIAS pixel_5138/NB2 pixel_5138/AMP_IN pixel_5138/SF_IB
+ pixel_5138/PIX_OUT pixel_5138/CSA_VREF pixel
Xpixel_432 pixel_432/gring pixel_432/VDD pixel_432/GND pixel_432/VREF pixel_432/ROW_SEL
+ pixel_432/NB1 pixel_432/VBIAS pixel_432/NB2 pixel_432/AMP_IN pixel_432/SF_IB pixel_432/PIX_OUT
+ pixel_432/CSA_VREF pixel
Xpixel_421 pixel_421/gring pixel_421/VDD pixel_421/GND pixel_421/VREF pixel_421/ROW_SEL
+ pixel_421/NB1 pixel_421/VBIAS pixel_421/NB2 pixel_421/AMP_IN pixel_421/SF_IB pixel_421/PIX_OUT
+ pixel_421/CSA_VREF pixel
Xpixel_410 pixel_410/gring pixel_410/VDD pixel_410/GND pixel_410/VREF pixel_410/ROW_SEL
+ pixel_410/NB1 pixel_410/VBIAS pixel_410/NB2 pixel_410/AMP_IN pixel_410/SF_IB pixel_410/PIX_OUT
+ pixel_410/CSA_VREF pixel
Xpixel_5149 pixel_5149/gring pixel_5149/VDD pixel_5149/GND pixel_5149/VREF pixel_5149/ROW_SEL
+ pixel_5149/NB1 pixel_5149/VBIAS pixel_5149/NB2 pixel_5149/AMP_IN pixel_5149/SF_IB
+ pixel_5149/PIX_OUT pixel_5149/CSA_VREF pixel
Xpixel_4404 pixel_4404/gring pixel_4404/VDD pixel_4404/GND pixel_4404/VREF pixel_4404/ROW_SEL
+ pixel_4404/NB1 pixel_4404/VBIAS pixel_4404/NB2 pixel_4404/AMP_IN pixel_4404/SF_IB
+ pixel_4404/PIX_OUT pixel_4404/CSA_VREF pixel
Xpixel_4415 pixel_4415/gring pixel_4415/VDD pixel_4415/GND pixel_4415/VREF pixel_4415/ROW_SEL
+ pixel_4415/NB1 pixel_4415/VBIAS pixel_4415/NB2 pixel_4415/AMP_IN pixel_4415/SF_IB
+ pixel_4415/PIX_OUT pixel_4415/CSA_VREF pixel
Xpixel_4426 pixel_4426/gring pixel_4426/VDD pixel_4426/GND pixel_4426/VREF pixel_4426/ROW_SEL
+ pixel_4426/NB1 pixel_4426/VBIAS pixel_4426/NB2 pixel_4426/AMP_IN pixel_4426/SF_IB
+ pixel_4426/PIX_OUT pixel_4426/CSA_VREF pixel
Xpixel_465 pixel_465/gring pixel_465/VDD pixel_465/GND pixel_465/VREF pixel_465/ROW_SEL
+ pixel_465/NB1 pixel_465/VBIAS pixel_465/NB2 pixel_465/AMP_IN pixel_465/SF_IB pixel_465/PIX_OUT
+ pixel_465/CSA_VREF pixel
Xpixel_454 pixel_454/gring pixel_454/VDD pixel_454/GND pixel_454/VREF pixel_454/ROW_SEL
+ pixel_454/NB1 pixel_454/VBIAS pixel_454/NB2 pixel_454/AMP_IN pixel_454/SF_IB pixel_454/PIX_OUT
+ pixel_454/CSA_VREF pixel
Xpixel_443 pixel_443/gring pixel_443/VDD pixel_443/GND pixel_443/VREF pixel_443/ROW_SEL
+ pixel_443/NB1 pixel_443/VBIAS pixel_443/NB2 pixel_443/AMP_IN pixel_443/SF_IB pixel_443/PIX_OUT
+ pixel_443/CSA_VREF pixel
Xpixel_3725 pixel_3725/gring pixel_3725/VDD pixel_3725/GND pixel_3725/VREF pixel_3725/ROW_SEL
+ pixel_3725/NB1 pixel_3725/VBIAS pixel_3725/NB2 pixel_3725/AMP_IN pixel_3725/SF_IB
+ pixel_3725/PIX_OUT pixel_3725/CSA_VREF pixel
Xpixel_3714 pixel_3714/gring pixel_3714/VDD pixel_3714/GND pixel_3714/VREF pixel_3714/ROW_SEL
+ pixel_3714/NB1 pixel_3714/VBIAS pixel_3714/NB2 pixel_3714/AMP_IN pixel_3714/SF_IB
+ pixel_3714/PIX_OUT pixel_3714/CSA_VREF pixel
Xpixel_3703 pixel_3703/gring pixel_3703/VDD pixel_3703/GND pixel_3703/VREF pixel_3703/ROW_SEL
+ pixel_3703/NB1 pixel_3703/VBIAS pixel_3703/NB2 pixel_3703/AMP_IN pixel_3703/SF_IB
+ pixel_3703/PIX_OUT pixel_3703/CSA_VREF pixel
Xpixel_4437 pixel_4437/gring pixel_4437/VDD pixel_4437/GND pixel_4437/VREF pixel_4437/ROW_SEL
+ pixel_4437/NB1 pixel_4437/VBIAS pixel_4437/NB2 pixel_4437/AMP_IN pixel_4437/SF_IB
+ pixel_4437/PIX_OUT pixel_4437/CSA_VREF pixel
Xpixel_4448 pixel_4448/gring pixel_4448/VDD pixel_4448/GND pixel_4448/VREF pixel_4448/ROW_SEL
+ pixel_4448/NB1 pixel_4448/VBIAS pixel_4448/NB2 pixel_4448/AMP_IN pixel_4448/SF_IB
+ pixel_4448/PIX_OUT pixel_4448/CSA_VREF pixel
Xpixel_4459 pixel_4459/gring pixel_4459/VDD pixel_4459/GND pixel_4459/VREF pixel_4459/ROW_SEL
+ pixel_4459/NB1 pixel_4459/VBIAS pixel_4459/NB2 pixel_4459/AMP_IN pixel_4459/SF_IB
+ pixel_4459/PIX_OUT pixel_4459/CSA_VREF pixel
Xpixel_498 pixel_498/gring pixel_498/VDD pixel_498/GND pixel_498/VREF pixel_498/ROW_SEL
+ pixel_498/NB1 pixel_498/VBIAS pixel_498/NB2 pixel_498/AMP_IN pixel_498/SF_IB pixel_498/PIX_OUT
+ pixel_498/CSA_VREF pixel
Xpixel_487 pixel_487/gring pixel_487/VDD pixel_487/GND pixel_487/VREF pixel_487/ROW_SEL
+ pixel_487/NB1 pixel_487/VBIAS pixel_487/NB2 pixel_487/AMP_IN pixel_487/SF_IB pixel_487/PIX_OUT
+ pixel_487/CSA_VREF pixel
Xpixel_476 pixel_476/gring pixel_476/VDD pixel_476/GND pixel_476/VREF pixel_476/ROW_SEL
+ pixel_476/NB1 pixel_476/VBIAS pixel_476/NB2 pixel_476/AMP_IN pixel_476/SF_IB pixel_476/PIX_OUT
+ pixel_476/CSA_VREF pixel
Xpixel_3758 pixel_3758/gring pixel_3758/VDD pixel_3758/GND pixel_3758/VREF pixel_3758/ROW_SEL
+ pixel_3758/NB1 pixel_3758/VBIAS pixel_3758/NB2 pixel_3758/AMP_IN pixel_3758/SF_IB
+ pixel_3758/PIX_OUT pixel_3758/CSA_VREF pixel
Xpixel_3747 pixel_3747/gring pixel_3747/VDD pixel_3747/GND pixel_3747/VREF pixel_3747/ROW_SEL
+ pixel_3747/NB1 pixel_3747/VBIAS pixel_3747/NB2 pixel_3747/AMP_IN pixel_3747/SF_IB
+ pixel_3747/PIX_OUT pixel_3747/CSA_VREF pixel
Xpixel_3736 pixel_3736/gring pixel_3736/VDD pixel_3736/GND pixel_3736/VREF pixel_3736/ROW_SEL
+ pixel_3736/NB1 pixel_3736/VBIAS pixel_3736/NB2 pixel_3736/AMP_IN pixel_3736/SF_IB
+ pixel_3736/PIX_OUT pixel_3736/CSA_VREF pixel
Xpixel_3769 pixel_3769/gring pixel_3769/VDD pixel_3769/GND pixel_3769/VREF pixel_3769/ROW_SEL
+ pixel_3769/NB1 pixel_3769/VBIAS pixel_3769/NB2 pixel_3769/AMP_IN pixel_3769/SF_IB
+ pixel_3769/PIX_OUT pixel_3769/CSA_VREF pixel
Xpixel_7030 pixel_7030/gring pixel_7030/VDD pixel_7030/GND pixel_7030/VREF pixel_7030/ROW_SEL
+ pixel_7030/NB1 pixel_7030/VBIAS pixel_7030/NB2 pixel_7030/AMP_IN pixel_7030/SF_IB
+ pixel_7030/PIX_OUT pixel_7030/CSA_VREF pixel
Xpixel_7041 pixel_7041/gring pixel_7041/VDD pixel_7041/GND pixel_7041/VREF pixel_7041/ROW_SEL
+ pixel_7041/NB1 pixel_7041/VBIAS pixel_7041/NB2 pixel_7041/AMP_IN pixel_7041/SF_IB
+ pixel_7041/PIX_OUT pixel_7041/CSA_VREF pixel
Xpixel_7052 pixel_7052/gring pixel_7052/VDD pixel_7052/GND pixel_7052/VREF pixel_7052/ROW_SEL
+ pixel_7052/NB1 pixel_7052/VBIAS pixel_7052/NB2 pixel_7052/AMP_IN pixel_7052/SF_IB
+ pixel_7052/PIX_OUT pixel_7052/CSA_VREF pixel
Xpixel_7063 pixel_7063/gring pixel_7063/VDD pixel_7063/GND pixel_7063/VREF pixel_7063/ROW_SEL
+ pixel_7063/NB1 pixel_7063/VBIAS pixel_7063/NB2 pixel_7063/AMP_IN pixel_7063/SF_IB
+ pixel_7063/PIX_OUT pixel_7063/CSA_VREF pixel
Xpixel_7074 pixel_7074/gring pixel_7074/VDD pixel_7074/GND pixel_7074/VREF pixel_7074/ROW_SEL
+ pixel_7074/NB1 pixel_7074/VBIAS pixel_7074/NB2 pixel_7074/AMP_IN pixel_7074/SF_IB
+ pixel_7074/PIX_OUT pixel_7074/CSA_VREF pixel
Xpixel_7085 pixel_7085/gring pixel_7085/VDD pixel_7085/GND pixel_7085/VREF pixel_7085/ROW_SEL
+ pixel_7085/NB1 pixel_7085/VBIAS pixel_7085/NB2 pixel_7085/AMP_IN pixel_7085/SF_IB
+ pixel_7085/PIX_OUT pixel_7085/CSA_VREF pixel
Xpixel_7096 pixel_7096/gring pixel_7096/VDD pixel_7096/GND pixel_7096/VREF pixel_7096/ROW_SEL
+ pixel_7096/NB1 pixel_7096/VBIAS pixel_7096/NB2 pixel_7096/AMP_IN pixel_7096/SF_IB
+ pixel_7096/PIX_OUT pixel_7096/CSA_VREF pixel
Xpixel_6340 pixel_6340/gring pixel_6340/VDD pixel_6340/GND pixel_6340/VREF pixel_6340/ROW_SEL
+ pixel_6340/NB1 pixel_6340/VBIAS pixel_6340/NB2 pixel_6340/AMP_IN pixel_6340/SF_IB
+ pixel_6340/PIX_OUT pixel_6340/CSA_VREF pixel
Xpixel_6351 pixel_6351/gring pixel_6351/VDD pixel_6351/GND pixel_6351/VREF pixel_6351/ROW_SEL
+ pixel_6351/NB1 pixel_6351/VBIAS pixel_6351/NB2 pixel_6351/AMP_IN pixel_6351/SF_IB
+ pixel_6351/PIX_OUT pixel_6351/CSA_VREF pixel
Xpixel_6362 pixel_6362/gring pixel_6362/VDD pixel_6362/GND pixel_6362/VREF pixel_6362/ROW_SEL
+ pixel_6362/NB1 pixel_6362/VBIAS pixel_6362/NB2 pixel_6362/AMP_IN pixel_6362/SF_IB
+ pixel_6362/PIX_OUT pixel_6362/CSA_VREF pixel
Xpixel_6373 pixel_6373/gring pixel_6373/VDD pixel_6373/GND pixel_6373/VREF pixel_6373/ROW_SEL
+ pixel_6373/NB1 pixel_6373/VBIAS pixel_6373/NB2 pixel_6373/AMP_IN pixel_6373/SF_IB
+ pixel_6373/PIX_OUT pixel_6373/CSA_VREF pixel
Xpixel_6384 pixel_6384/gring pixel_6384/VDD pixel_6384/GND pixel_6384/VREF pixel_6384/ROW_SEL
+ pixel_6384/NB1 pixel_6384/VBIAS pixel_6384/NB2 pixel_6384/AMP_IN pixel_6384/SF_IB
+ pixel_6384/PIX_OUT pixel_6384/CSA_VREF pixel
Xpixel_6395 pixel_6395/gring pixel_6395/VDD pixel_6395/GND pixel_6395/VREF pixel_6395/ROW_SEL
+ pixel_6395/NB1 pixel_6395/VBIAS pixel_6395/NB2 pixel_6395/AMP_IN pixel_6395/SF_IB
+ pixel_6395/PIX_OUT pixel_6395/CSA_VREF pixel
Xpixel_5650 pixel_5650/gring pixel_5650/VDD pixel_5650/GND pixel_5650/VREF pixel_5650/ROW_SEL
+ pixel_5650/NB1 pixel_5650/VBIAS pixel_5650/NB2 pixel_5650/AMP_IN pixel_5650/SF_IB
+ pixel_5650/PIX_OUT pixel_5650/CSA_VREF pixel
Xpixel_5661 pixel_5661/gring pixel_5661/VDD pixel_5661/GND pixel_5661/VREF pixel_5661/ROW_SEL
+ pixel_5661/NB1 pixel_5661/VBIAS pixel_5661/NB2 pixel_5661/AMP_IN pixel_5661/SF_IB
+ pixel_5661/PIX_OUT pixel_5661/CSA_VREF pixel
Xpixel_5672 pixel_5672/gring pixel_5672/VDD pixel_5672/GND pixel_5672/VREF pixel_5672/ROW_SEL
+ pixel_5672/NB1 pixel_5672/VBIAS pixel_5672/NB2 pixel_5672/AMP_IN pixel_5672/SF_IB
+ pixel_5672/PIX_OUT pixel_5672/CSA_VREF pixel
Xpixel_5683 pixel_5683/gring pixel_5683/VDD pixel_5683/GND pixel_5683/VREF pixel_5683/ROW_SEL
+ pixel_5683/NB1 pixel_5683/VBIAS pixel_5683/NB2 pixel_5683/AMP_IN pixel_5683/SF_IB
+ pixel_5683/PIX_OUT pixel_5683/CSA_VREF pixel
Xpixel_5694 pixel_5694/gring pixel_5694/VDD pixel_5694/GND pixel_5694/VREF pixel_5694/ROW_SEL
+ pixel_5694/NB1 pixel_5694/VBIAS pixel_5694/NB2 pixel_5694/AMP_IN pixel_5694/SF_IB
+ pixel_5694/PIX_OUT pixel_5694/CSA_VREF pixel
Xpixel_4960 pixel_4960/gring pixel_4960/VDD pixel_4960/GND pixel_4960/VREF pixel_4960/ROW_SEL
+ pixel_4960/NB1 pixel_4960/VBIAS pixel_4960/NB2 pixel_4960/AMP_IN pixel_4960/SF_IB
+ pixel_4960/PIX_OUT pixel_4960/CSA_VREF pixel
Xpixel_4971 pixel_4971/gring pixel_4971/VDD pixel_4971/GND pixel_4971/VREF pixel_4971/ROW_SEL
+ pixel_4971/NB1 pixel_4971/VBIAS pixel_4971/NB2 pixel_4971/AMP_IN pixel_4971/SF_IB
+ pixel_4971/PIX_OUT pixel_4971/CSA_VREF pixel
Xpixel_4982 pixel_4982/gring pixel_4982/VDD pixel_4982/GND pixel_4982/VREF pixel_4982/ROW_SEL
+ pixel_4982/NB1 pixel_4982/VBIAS pixel_4982/NB2 pixel_4982/AMP_IN pixel_4982/SF_IB
+ pixel_4982/PIX_OUT pixel_4982/CSA_VREF pixel
Xpixel_4993 pixel_4993/gring pixel_4993/VDD pixel_4993/GND pixel_4993/VREF pixel_4993/ROW_SEL
+ pixel_4993/NB1 pixel_4993/VBIAS pixel_4993/NB2 pixel_4993/AMP_IN pixel_4993/SF_IB
+ pixel_4993/PIX_OUT pixel_4993/CSA_VREF pixel
Xpixel_2309 pixel_2309/gring pixel_2309/VDD pixel_2309/GND pixel_2309/VREF pixel_2309/ROW_SEL
+ pixel_2309/NB1 pixel_2309/VBIAS pixel_2309/NB2 pixel_2309/AMP_IN pixel_2309/SF_IB
+ pixel_2309/PIX_OUT pixel_2309/CSA_VREF pixel
Xpixel_1619 pixel_1619/gring pixel_1619/VDD pixel_1619/GND pixel_1619/VREF pixel_1619/ROW_SEL
+ pixel_1619/NB1 pixel_1619/VBIAS pixel_1619/NB2 pixel_1619/AMP_IN pixel_1619/SF_IB
+ pixel_1619/PIX_OUT pixel_1619/CSA_VREF pixel
Xpixel_1608 pixel_1608/gring pixel_1608/VDD pixel_1608/GND pixel_1608/VREF pixel_1608/ROW_SEL
+ pixel_1608/NB1 pixel_1608/VBIAS pixel_1608/NB2 pixel_1608/AMP_IN pixel_1608/SF_IB
+ pixel_1608/PIX_OUT pixel_1608/CSA_VREF pixel
Xpixel_9905 pixel_9905/gring pixel_9905/VDD pixel_9905/GND pixel_9905/VREF pixel_9905/ROW_SEL
+ pixel_9905/NB1 pixel_9905/VBIAS pixel_9905/NB2 pixel_9905/AMP_IN pixel_9905/SF_IB
+ pixel_9905/PIX_OUT pixel_9905/CSA_VREF pixel
Xpixel_9938 pixel_9938/gring pixel_9938/VDD pixel_9938/GND pixel_9938/VREF pixel_9938/ROW_SEL
+ pixel_9938/NB1 pixel_9938/VBIAS pixel_9938/NB2 pixel_9938/AMP_IN pixel_9938/SF_IB
+ pixel_9938/PIX_OUT pixel_9938/CSA_VREF pixel
Xpixel_9927 pixel_9927/gring pixel_9927/VDD pixel_9927/GND pixel_9927/VREF pixel_9927/ROW_SEL
+ pixel_9927/NB1 pixel_9927/VBIAS pixel_9927/NB2 pixel_9927/AMP_IN pixel_9927/SF_IB
+ pixel_9927/PIX_OUT pixel_9927/CSA_VREF pixel
Xpixel_9916 pixel_9916/gring pixel_9916/VDD pixel_9916/GND pixel_9916/VREF pixel_9916/ROW_SEL
+ pixel_9916/NB1 pixel_9916/VBIAS pixel_9916/NB2 pixel_9916/AMP_IN pixel_9916/SF_IB
+ pixel_9916/PIX_OUT pixel_9916/CSA_VREF pixel
Xpixel_9949 pixel_9949/gring pixel_9949/VDD pixel_9949/GND pixel_9949/VREF pixel_9949/ROW_SEL
+ pixel_9949/NB1 pixel_9949/VBIAS pixel_9949/NB2 pixel_9949/AMP_IN pixel_9949/SF_IB
+ pixel_9949/PIX_OUT pixel_9949/CSA_VREF pixel
Xpixel_4201 pixel_4201/gring pixel_4201/VDD pixel_4201/GND pixel_4201/VREF pixel_4201/ROW_SEL
+ pixel_4201/NB1 pixel_4201/VBIAS pixel_4201/NB2 pixel_4201/AMP_IN pixel_4201/SF_IB
+ pixel_4201/PIX_OUT pixel_4201/CSA_VREF pixel
Xpixel_240 pixel_240/gring pixel_240/VDD pixel_240/GND pixel_240/VREF pixel_240/ROW_SEL
+ pixel_240/NB1 pixel_240/VBIAS pixel_240/NB2 pixel_240/AMP_IN pixel_240/SF_IB pixel_240/PIX_OUT
+ pixel_240/CSA_VREF pixel
Xpixel_3500 pixel_3500/gring pixel_3500/VDD pixel_3500/GND pixel_3500/VREF pixel_3500/ROW_SEL
+ pixel_3500/NB1 pixel_3500/VBIAS pixel_3500/NB2 pixel_3500/AMP_IN pixel_3500/SF_IB
+ pixel_3500/PIX_OUT pixel_3500/CSA_VREF pixel
Xpixel_4212 pixel_4212/gring pixel_4212/VDD pixel_4212/GND pixel_4212/VREF pixel_4212/ROW_SEL
+ pixel_4212/NB1 pixel_4212/VBIAS pixel_4212/NB2 pixel_4212/AMP_IN pixel_4212/SF_IB
+ pixel_4212/PIX_OUT pixel_4212/CSA_VREF pixel
Xpixel_4223 pixel_4223/gring pixel_4223/VDD pixel_4223/GND pixel_4223/VREF pixel_4223/ROW_SEL
+ pixel_4223/NB1 pixel_4223/VBIAS pixel_4223/NB2 pixel_4223/AMP_IN pixel_4223/SF_IB
+ pixel_4223/PIX_OUT pixel_4223/CSA_VREF pixel
Xpixel_4234 pixel_4234/gring pixel_4234/VDD pixel_4234/GND pixel_4234/VREF pixel_4234/ROW_SEL
+ pixel_4234/NB1 pixel_4234/VBIAS pixel_4234/NB2 pixel_4234/AMP_IN pixel_4234/SF_IB
+ pixel_4234/PIX_OUT pixel_4234/CSA_VREF pixel
Xpixel_4245 pixel_4245/gring pixel_4245/VDD pixel_4245/GND pixel_4245/VREF pixel_4245/ROW_SEL
+ pixel_4245/NB1 pixel_4245/VBIAS pixel_4245/NB2 pixel_4245/AMP_IN pixel_4245/SF_IB
+ pixel_4245/PIX_OUT pixel_4245/CSA_VREF pixel
Xpixel_273 pixel_273/gring pixel_273/VDD pixel_273/GND pixel_273/VREF pixel_273/ROW_SEL
+ pixel_273/NB1 pixel_273/VBIAS pixel_273/NB2 pixel_273/AMP_IN pixel_273/SF_IB pixel_273/PIX_OUT
+ pixel_273/CSA_VREF pixel
Xpixel_262 pixel_262/gring pixel_262/VDD pixel_262/GND pixel_262/VREF pixel_262/ROW_SEL
+ pixel_262/NB1 pixel_262/VBIAS pixel_262/NB2 pixel_262/AMP_IN pixel_262/SF_IB pixel_262/PIX_OUT
+ pixel_262/CSA_VREF pixel
Xpixel_251 pixel_251/gring pixel_251/VDD pixel_251/GND pixel_251/VREF pixel_251/ROW_SEL
+ pixel_251/NB1 pixel_251/VBIAS pixel_251/NB2 pixel_251/AMP_IN pixel_251/SF_IB pixel_251/PIX_OUT
+ pixel_251/CSA_VREF pixel
Xpixel_3533 pixel_3533/gring pixel_3533/VDD pixel_3533/GND pixel_3533/VREF pixel_3533/ROW_SEL
+ pixel_3533/NB1 pixel_3533/VBIAS pixel_3533/NB2 pixel_3533/AMP_IN pixel_3533/SF_IB
+ pixel_3533/PIX_OUT pixel_3533/CSA_VREF pixel
Xpixel_3522 pixel_3522/gring pixel_3522/VDD pixel_3522/GND pixel_3522/VREF pixel_3522/ROW_SEL
+ pixel_3522/NB1 pixel_3522/VBIAS pixel_3522/NB2 pixel_3522/AMP_IN pixel_3522/SF_IB
+ pixel_3522/PIX_OUT pixel_3522/CSA_VREF pixel
Xpixel_3511 pixel_3511/gring pixel_3511/VDD pixel_3511/GND pixel_3511/VREF pixel_3511/ROW_SEL
+ pixel_3511/NB1 pixel_3511/VBIAS pixel_3511/NB2 pixel_3511/AMP_IN pixel_3511/SF_IB
+ pixel_3511/PIX_OUT pixel_3511/CSA_VREF pixel
Xpixel_4256 pixel_4256/gring pixel_4256/VDD pixel_4256/GND pixel_4256/VREF pixel_4256/ROW_SEL
+ pixel_4256/NB1 pixel_4256/VBIAS pixel_4256/NB2 pixel_4256/AMP_IN pixel_4256/SF_IB
+ pixel_4256/PIX_OUT pixel_4256/CSA_VREF pixel
Xpixel_4267 pixel_4267/gring pixel_4267/VDD pixel_4267/GND pixel_4267/VREF pixel_4267/ROW_SEL
+ pixel_4267/NB1 pixel_4267/VBIAS pixel_4267/NB2 pixel_4267/AMP_IN pixel_4267/SF_IB
+ pixel_4267/PIX_OUT pixel_4267/CSA_VREF pixel
Xpixel_4278 pixel_4278/gring pixel_4278/VDD pixel_4278/GND pixel_4278/VREF pixel_4278/ROW_SEL
+ pixel_4278/NB1 pixel_4278/VBIAS pixel_4278/NB2 pixel_4278/AMP_IN pixel_4278/SF_IB
+ pixel_4278/PIX_OUT pixel_4278/CSA_VREF pixel
Xpixel_295 pixel_295/gring pixel_295/VDD pixel_295/GND pixel_295/VREF pixel_295/ROW_SEL
+ pixel_295/NB1 pixel_295/VBIAS pixel_295/NB2 pixel_295/AMP_IN pixel_295/SF_IB pixel_295/PIX_OUT
+ pixel_295/CSA_VREF pixel
Xpixel_284 pixel_284/gring pixel_284/VDD pixel_284/GND pixel_284/VREF pixel_284/ROW_SEL
+ pixel_284/NB1 pixel_284/VBIAS pixel_284/NB2 pixel_284/AMP_IN pixel_284/SF_IB pixel_284/PIX_OUT
+ pixel_284/CSA_VREF pixel
Xpixel_2821 pixel_2821/gring pixel_2821/VDD pixel_2821/GND pixel_2821/VREF pixel_2821/ROW_SEL
+ pixel_2821/NB1 pixel_2821/VBIAS pixel_2821/NB2 pixel_2821/AMP_IN pixel_2821/SF_IB
+ pixel_2821/PIX_OUT pixel_2821/CSA_VREF pixel
Xpixel_2810 pixel_2810/gring pixel_2810/VDD pixel_2810/GND pixel_2810/VREF pixel_2810/ROW_SEL
+ pixel_2810/NB1 pixel_2810/VBIAS pixel_2810/NB2 pixel_2810/AMP_IN pixel_2810/SF_IB
+ pixel_2810/PIX_OUT pixel_2810/CSA_VREF pixel
Xpixel_3566 pixel_3566/gring pixel_3566/VDD pixel_3566/GND pixel_3566/VREF pixel_3566/ROW_SEL
+ pixel_3566/NB1 pixel_3566/VBIAS pixel_3566/NB2 pixel_3566/AMP_IN pixel_3566/SF_IB
+ pixel_3566/PIX_OUT pixel_3566/CSA_VREF pixel
Xpixel_3555 pixel_3555/gring pixel_3555/VDD pixel_3555/GND pixel_3555/VREF pixel_3555/ROW_SEL
+ pixel_3555/NB1 pixel_3555/VBIAS pixel_3555/NB2 pixel_3555/AMP_IN pixel_3555/SF_IB
+ pixel_3555/PIX_OUT pixel_3555/CSA_VREF pixel
Xpixel_3544 pixel_3544/gring pixel_3544/VDD pixel_3544/GND pixel_3544/VREF pixel_3544/ROW_SEL
+ pixel_3544/NB1 pixel_3544/VBIAS pixel_3544/NB2 pixel_3544/AMP_IN pixel_3544/SF_IB
+ pixel_3544/PIX_OUT pixel_3544/CSA_VREF pixel
Xpixel_4289 pixel_4289/gring pixel_4289/VDD pixel_4289/GND pixel_4289/VREF pixel_4289/ROW_SEL
+ pixel_4289/NB1 pixel_4289/VBIAS pixel_4289/NB2 pixel_4289/AMP_IN pixel_4289/SF_IB
+ pixel_4289/PIX_OUT pixel_4289/CSA_VREF pixel
Xpixel_2865 pixel_2865/gring pixel_2865/VDD pixel_2865/GND pixel_2865/VREF pixel_2865/ROW_SEL
+ pixel_2865/NB1 pixel_2865/VBIAS pixel_2865/NB2 pixel_2865/AMP_IN pixel_2865/SF_IB
+ pixel_2865/PIX_OUT pixel_2865/CSA_VREF pixel
Xpixel_2854 pixel_2854/gring pixel_2854/VDD pixel_2854/GND pixel_2854/VREF pixel_2854/ROW_SEL
+ pixel_2854/NB1 pixel_2854/VBIAS pixel_2854/NB2 pixel_2854/AMP_IN pixel_2854/SF_IB
+ pixel_2854/PIX_OUT pixel_2854/CSA_VREF pixel
Xpixel_2843 pixel_2843/gring pixel_2843/VDD pixel_2843/GND pixel_2843/VREF pixel_2843/ROW_SEL
+ pixel_2843/NB1 pixel_2843/VBIAS pixel_2843/NB2 pixel_2843/AMP_IN pixel_2843/SF_IB
+ pixel_2843/PIX_OUT pixel_2843/CSA_VREF pixel
Xpixel_2832 pixel_2832/gring pixel_2832/VDD pixel_2832/GND pixel_2832/VREF pixel_2832/ROW_SEL
+ pixel_2832/NB1 pixel_2832/VBIAS pixel_2832/NB2 pixel_2832/AMP_IN pixel_2832/SF_IB
+ pixel_2832/PIX_OUT pixel_2832/CSA_VREF pixel
Xpixel_3599 pixel_3599/gring pixel_3599/VDD pixel_3599/GND pixel_3599/VREF pixel_3599/ROW_SEL
+ pixel_3599/NB1 pixel_3599/VBIAS pixel_3599/NB2 pixel_3599/AMP_IN pixel_3599/SF_IB
+ pixel_3599/PIX_OUT pixel_3599/CSA_VREF pixel
Xpixel_3588 pixel_3588/gring pixel_3588/VDD pixel_3588/GND pixel_3588/VREF pixel_3588/ROW_SEL
+ pixel_3588/NB1 pixel_3588/VBIAS pixel_3588/NB2 pixel_3588/AMP_IN pixel_3588/SF_IB
+ pixel_3588/PIX_OUT pixel_3588/CSA_VREF pixel
Xpixel_3577 pixel_3577/gring pixel_3577/VDD pixel_3577/GND pixel_3577/VREF pixel_3577/ROW_SEL
+ pixel_3577/NB1 pixel_3577/VBIAS pixel_3577/NB2 pixel_3577/AMP_IN pixel_3577/SF_IB
+ pixel_3577/PIX_OUT pixel_3577/CSA_VREF pixel
Xpixel_2898 pixel_2898/gring pixel_2898/VDD pixel_2898/GND pixel_2898/VREF pixel_2898/ROW_SEL
+ pixel_2898/NB1 pixel_2898/VBIAS pixel_2898/NB2 pixel_2898/AMP_IN pixel_2898/SF_IB
+ pixel_2898/PIX_OUT pixel_2898/CSA_VREF pixel
Xpixel_2887 pixel_2887/gring pixel_2887/VDD pixel_2887/GND pixel_2887/VREF pixel_2887/ROW_SEL
+ pixel_2887/NB1 pixel_2887/VBIAS pixel_2887/NB2 pixel_2887/AMP_IN pixel_2887/SF_IB
+ pixel_2887/PIX_OUT pixel_2887/CSA_VREF pixel
Xpixel_2876 pixel_2876/gring pixel_2876/VDD pixel_2876/GND pixel_2876/VREF pixel_2876/ROW_SEL
+ pixel_2876/NB1 pixel_2876/VBIAS pixel_2876/NB2 pixel_2876/AMP_IN pixel_2876/SF_IB
+ pixel_2876/PIX_OUT pixel_2876/CSA_VREF pixel
Xpixel_6170 pixel_6170/gring pixel_6170/VDD pixel_6170/GND pixel_6170/VREF pixel_6170/ROW_SEL
+ pixel_6170/NB1 pixel_6170/VBIAS pixel_6170/NB2 pixel_6170/AMP_IN pixel_6170/SF_IB
+ pixel_6170/PIX_OUT pixel_6170/CSA_VREF pixel
Xpixel_6181 pixel_6181/gring pixel_6181/VDD pixel_6181/GND pixel_6181/VREF pixel_6181/ROW_SEL
+ pixel_6181/NB1 pixel_6181/VBIAS pixel_6181/NB2 pixel_6181/AMP_IN pixel_6181/SF_IB
+ pixel_6181/PIX_OUT pixel_6181/CSA_VREF pixel
Xpixel_6192 pixel_6192/gring pixel_6192/VDD pixel_6192/GND pixel_6192/VREF pixel_6192/ROW_SEL
+ pixel_6192/NB1 pixel_6192/VBIAS pixel_6192/NB2 pixel_6192/AMP_IN pixel_6192/SF_IB
+ pixel_6192/PIX_OUT pixel_6192/CSA_VREF pixel
Xpixel_5480 pixel_5480/gring pixel_5480/VDD pixel_5480/GND pixel_5480/VREF pixel_5480/ROW_SEL
+ pixel_5480/NB1 pixel_5480/VBIAS pixel_5480/NB2 pixel_5480/AMP_IN pixel_5480/SF_IB
+ pixel_5480/PIX_OUT pixel_5480/CSA_VREF pixel
Xpixel_5491 pixel_5491/gring pixel_5491/VDD pixel_5491/GND pixel_5491/VREF pixel_5491/ROW_SEL
+ pixel_5491/NB1 pixel_5491/VBIAS pixel_5491/NB2 pixel_5491/AMP_IN pixel_5491/SF_IB
+ pixel_5491/PIX_OUT pixel_5491/CSA_VREF pixel
Xpixel_4790 pixel_4790/gring pixel_4790/VDD pixel_4790/GND pixel_4790/VREF pixel_4790/ROW_SEL
+ pixel_4790/NB1 pixel_4790/VBIAS pixel_4790/NB2 pixel_4790/AMP_IN pixel_4790/SF_IB
+ pixel_4790/PIX_OUT pixel_4790/CSA_VREF pixel
Xpixel_2117 pixel_2117/gring pixel_2117/VDD pixel_2117/GND pixel_2117/VREF pixel_2117/ROW_SEL
+ pixel_2117/NB1 pixel_2117/VBIAS pixel_2117/NB2 pixel_2117/AMP_IN pixel_2117/SF_IB
+ pixel_2117/PIX_OUT pixel_2117/CSA_VREF pixel
Xpixel_2106 pixel_2106/gring pixel_2106/VDD pixel_2106/GND pixel_2106/VREF pixel_2106/ROW_SEL
+ pixel_2106/NB1 pixel_2106/VBIAS pixel_2106/NB2 pixel_2106/AMP_IN pixel_2106/SF_IB
+ pixel_2106/PIX_OUT pixel_2106/CSA_VREF pixel
Xpixel_1416 pixel_1416/gring pixel_1416/VDD pixel_1416/GND pixel_1416/VREF pixel_1416/ROW_SEL
+ pixel_1416/NB1 pixel_1416/VBIAS pixel_1416/NB2 pixel_1416/AMP_IN pixel_1416/SF_IB
+ pixel_1416/PIX_OUT pixel_1416/CSA_VREF pixel
Xpixel_1405 pixel_1405/gring pixel_1405/VDD pixel_1405/GND pixel_1405/VREF pixel_1405/ROW_SEL
+ pixel_1405/NB1 pixel_1405/VBIAS pixel_1405/NB2 pixel_1405/AMP_IN pixel_1405/SF_IB
+ pixel_1405/PIX_OUT pixel_1405/CSA_VREF pixel
Xpixel_2139 pixel_2139/gring pixel_2139/VDD pixel_2139/GND pixel_2139/VREF pixel_2139/ROW_SEL
+ pixel_2139/NB1 pixel_2139/VBIAS pixel_2139/NB2 pixel_2139/AMP_IN pixel_2139/SF_IB
+ pixel_2139/PIX_OUT pixel_2139/CSA_VREF pixel
Xpixel_2128 pixel_2128/gring pixel_2128/VDD pixel_2128/GND pixel_2128/VREF pixel_2128/ROW_SEL
+ pixel_2128/NB1 pixel_2128/VBIAS pixel_2128/NB2 pixel_2128/AMP_IN pixel_2128/SF_IB
+ pixel_2128/PIX_OUT pixel_2128/CSA_VREF pixel
Xpixel_1449 pixel_1449/gring pixel_1449/VDD pixel_1449/GND pixel_1449/VREF pixel_1449/ROW_SEL
+ pixel_1449/NB1 pixel_1449/VBIAS pixel_1449/NB2 pixel_1449/AMP_IN pixel_1449/SF_IB
+ pixel_1449/PIX_OUT pixel_1449/CSA_VREF pixel
Xpixel_1438 pixel_1438/gring pixel_1438/VDD pixel_1438/GND pixel_1438/VREF pixel_1438/ROW_SEL
+ pixel_1438/NB1 pixel_1438/VBIAS pixel_1438/NB2 pixel_1438/AMP_IN pixel_1438/SF_IB
+ pixel_1438/PIX_OUT pixel_1438/CSA_VREF pixel
Xpixel_1427 pixel_1427/gring pixel_1427/VDD pixel_1427/GND pixel_1427/VREF pixel_1427/ROW_SEL
+ pixel_1427/NB1 pixel_1427/VBIAS pixel_1427/NB2 pixel_1427/AMP_IN pixel_1427/SF_IB
+ pixel_1427/PIX_OUT pixel_1427/CSA_VREF pixel
Xpixel_9702 pixel_9702/gring pixel_9702/VDD pixel_9702/GND pixel_9702/VREF pixel_9702/ROW_SEL
+ pixel_9702/NB1 pixel_9702/VBIAS pixel_9702/NB2 pixel_9702/AMP_IN pixel_9702/SF_IB
+ pixel_9702/PIX_OUT pixel_9702/CSA_VREF pixel
Xpixel_9713 pixel_9713/gring pixel_9713/VDD pixel_9713/GND pixel_9713/VREF pixel_9713/ROW_SEL
+ pixel_9713/NB1 pixel_9713/VBIAS pixel_9713/NB2 pixel_9713/AMP_IN pixel_9713/SF_IB
+ pixel_9713/PIX_OUT pixel_9713/CSA_VREF pixel
Xpixel_9724 pixel_9724/gring pixel_9724/VDD pixel_9724/GND pixel_9724/VREF pixel_9724/ROW_SEL
+ pixel_9724/NB1 pixel_9724/VBIAS pixel_9724/NB2 pixel_9724/AMP_IN pixel_9724/SF_IB
+ pixel_9724/PIX_OUT pixel_9724/CSA_VREF pixel
Xpixel_9735 pixel_9735/gring pixel_9735/VDD pixel_9735/GND pixel_9735/VREF pixel_9735/ROW_SEL
+ pixel_9735/NB1 pixel_9735/VBIAS pixel_9735/NB2 pixel_9735/AMP_IN pixel_9735/SF_IB
+ pixel_9735/PIX_OUT pixel_9735/CSA_VREF pixel
Xpixel_9746 pixel_9746/gring pixel_9746/VDD pixel_9746/GND pixel_9746/VREF pixel_9746/ROW_SEL
+ pixel_9746/NB1 pixel_9746/VBIAS pixel_9746/NB2 pixel_9746/AMP_IN pixel_9746/SF_IB
+ pixel_9746/PIX_OUT pixel_9746/CSA_VREF pixel
Xpixel_9757 pixel_9757/gring pixel_9757/VDD pixel_9757/GND pixel_9757/VREF pixel_9757/ROW_SEL
+ pixel_9757/NB1 pixel_9757/VBIAS pixel_9757/NB2 pixel_9757/AMP_IN pixel_9757/SF_IB
+ pixel_9757/PIX_OUT pixel_9757/CSA_VREF pixel
Xpixel_9768 pixel_9768/gring pixel_9768/VDD pixel_9768/GND pixel_9768/VREF pixel_9768/ROW_SEL
+ pixel_9768/NB1 pixel_9768/VBIAS pixel_9768/NB2 pixel_9768/AMP_IN pixel_9768/SF_IB
+ pixel_9768/PIX_OUT pixel_9768/CSA_VREF pixel
Xpixel_9779 pixel_9779/gring pixel_9779/VDD pixel_9779/GND pixel_9779/VREF pixel_9779/ROW_SEL
+ pixel_9779/NB1 pixel_9779/VBIAS pixel_9779/NB2 pixel_9779/AMP_IN pixel_9779/SF_IB
+ pixel_9779/PIX_OUT pixel_9779/CSA_VREF pixel
Xpixel_4020 pixel_4020/gring pixel_4020/VDD pixel_4020/GND pixel_4020/VREF pixel_4020/ROW_SEL
+ pixel_4020/NB1 pixel_4020/VBIAS pixel_4020/NB2 pixel_4020/AMP_IN pixel_4020/SF_IB
+ pixel_4020/PIX_OUT pixel_4020/CSA_VREF pixel
Xpixel_4031 pixel_4031/gring pixel_4031/VDD pixel_4031/GND pixel_4031/VREF pixel_4031/ROW_SEL
+ pixel_4031/NB1 pixel_4031/VBIAS pixel_4031/NB2 pixel_4031/AMP_IN pixel_4031/SF_IB
+ pixel_4031/PIX_OUT pixel_4031/CSA_VREF pixel
Xpixel_4042 pixel_4042/gring pixel_4042/VDD pixel_4042/GND pixel_4042/VREF pixel_4042/ROW_SEL
+ pixel_4042/NB1 pixel_4042/VBIAS pixel_4042/NB2 pixel_4042/AMP_IN pixel_4042/SF_IB
+ pixel_4042/PIX_OUT pixel_4042/CSA_VREF pixel
Xpixel_4053 pixel_4053/gring pixel_4053/VDD pixel_4053/GND pixel_4053/VREF pixel_4053/ROW_SEL
+ pixel_4053/NB1 pixel_4053/VBIAS pixel_4053/NB2 pixel_4053/AMP_IN pixel_4053/SF_IB
+ pixel_4053/PIX_OUT pixel_4053/CSA_VREF pixel
Xpixel_3341 pixel_3341/gring pixel_3341/VDD pixel_3341/GND pixel_3341/VREF pixel_3341/ROW_SEL
+ pixel_3341/NB1 pixel_3341/VBIAS pixel_3341/NB2 pixel_3341/AMP_IN pixel_3341/SF_IB
+ pixel_3341/PIX_OUT pixel_3341/CSA_VREF pixel
Xpixel_3330 pixel_3330/gring pixel_3330/VDD pixel_3330/GND pixel_3330/VREF pixel_3330/ROW_SEL
+ pixel_3330/NB1 pixel_3330/VBIAS pixel_3330/NB2 pixel_3330/AMP_IN pixel_3330/SF_IB
+ pixel_3330/PIX_OUT pixel_3330/CSA_VREF pixel
Xpixel_4064 pixel_4064/gring pixel_4064/VDD pixel_4064/GND pixel_4064/VREF pixel_4064/ROW_SEL
+ pixel_4064/NB1 pixel_4064/VBIAS pixel_4064/NB2 pixel_4064/AMP_IN pixel_4064/SF_IB
+ pixel_4064/PIX_OUT pixel_4064/CSA_VREF pixel
Xpixel_4075 pixel_4075/gring pixel_4075/VDD pixel_4075/GND pixel_4075/VREF pixel_4075/ROW_SEL
+ pixel_4075/NB1 pixel_4075/VBIAS pixel_4075/NB2 pixel_4075/AMP_IN pixel_4075/SF_IB
+ pixel_4075/PIX_OUT pixel_4075/CSA_VREF pixel
Xpixel_4086 pixel_4086/gring pixel_4086/VDD pixel_4086/GND pixel_4086/VREF pixel_4086/ROW_SEL
+ pixel_4086/NB1 pixel_4086/VBIAS pixel_4086/NB2 pixel_4086/AMP_IN pixel_4086/SF_IB
+ pixel_4086/PIX_OUT pixel_4086/CSA_VREF pixel
Xpixel_2640 pixel_2640/gring pixel_2640/VDD pixel_2640/GND pixel_2640/VREF pixel_2640/ROW_SEL
+ pixel_2640/NB1 pixel_2640/VBIAS pixel_2640/NB2 pixel_2640/AMP_IN pixel_2640/SF_IB
+ pixel_2640/PIX_OUT pixel_2640/CSA_VREF pixel
Xpixel_3385 pixel_3385/gring pixel_3385/VDD pixel_3385/GND pixel_3385/VREF pixel_3385/ROW_SEL
+ pixel_3385/NB1 pixel_3385/VBIAS pixel_3385/NB2 pixel_3385/AMP_IN pixel_3385/SF_IB
+ pixel_3385/PIX_OUT pixel_3385/CSA_VREF pixel
Xpixel_3374 pixel_3374/gring pixel_3374/VDD pixel_3374/GND pixel_3374/VREF pixel_3374/ROW_SEL
+ pixel_3374/NB1 pixel_3374/VBIAS pixel_3374/NB2 pixel_3374/AMP_IN pixel_3374/SF_IB
+ pixel_3374/PIX_OUT pixel_3374/CSA_VREF pixel
Xpixel_3363 pixel_3363/gring pixel_3363/VDD pixel_3363/GND pixel_3363/VREF pixel_3363/ROW_SEL
+ pixel_3363/NB1 pixel_3363/VBIAS pixel_3363/NB2 pixel_3363/AMP_IN pixel_3363/SF_IB
+ pixel_3363/PIX_OUT pixel_3363/CSA_VREF pixel
Xpixel_3352 pixel_3352/gring pixel_3352/VDD pixel_3352/GND pixel_3352/VREF pixel_3352/ROW_SEL
+ pixel_3352/NB1 pixel_3352/VBIAS pixel_3352/NB2 pixel_3352/AMP_IN pixel_3352/SF_IB
+ pixel_3352/PIX_OUT pixel_3352/CSA_VREF pixel
Xpixel_4097 pixel_4097/gring pixel_4097/VDD pixel_4097/GND pixel_4097/VREF pixel_4097/ROW_SEL
+ pixel_4097/NB1 pixel_4097/VBIAS pixel_4097/NB2 pixel_4097/AMP_IN pixel_4097/SF_IB
+ pixel_4097/PIX_OUT pixel_4097/CSA_VREF pixel
Xpixel_2673 pixel_2673/gring pixel_2673/VDD pixel_2673/GND pixel_2673/VREF pixel_2673/ROW_SEL
+ pixel_2673/NB1 pixel_2673/VBIAS pixel_2673/NB2 pixel_2673/AMP_IN pixel_2673/SF_IB
+ pixel_2673/PIX_OUT pixel_2673/CSA_VREF pixel
Xpixel_2662 pixel_2662/gring pixel_2662/VDD pixel_2662/GND pixel_2662/VREF pixel_2662/ROW_SEL
+ pixel_2662/NB1 pixel_2662/VBIAS pixel_2662/NB2 pixel_2662/AMP_IN pixel_2662/SF_IB
+ pixel_2662/PIX_OUT pixel_2662/CSA_VREF pixel
Xpixel_2651 pixel_2651/gring pixel_2651/VDD pixel_2651/GND pixel_2651/VREF pixel_2651/ROW_SEL
+ pixel_2651/NB1 pixel_2651/VBIAS pixel_2651/NB2 pixel_2651/AMP_IN pixel_2651/SF_IB
+ pixel_2651/PIX_OUT pixel_2651/CSA_VREF pixel
Xpixel_3396 pixel_3396/gring pixel_3396/VDD pixel_3396/GND pixel_3396/VREF pixel_3396/ROW_SEL
+ pixel_3396/NB1 pixel_3396/VBIAS pixel_3396/NB2 pixel_3396/AMP_IN pixel_3396/SF_IB
+ pixel_3396/PIX_OUT pixel_3396/CSA_VREF pixel
Xpixel_1961 pixel_1961/gring pixel_1961/VDD pixel_1961/GND pixel_1961/VREF pixel_1961/ROW_SEL
+ pixel_1961/NB1 pixel_1961/VBIAS pixel_1961/NB2 pixel_1961/AMP_IN pixel_1961/SF_IB
+ pixel_1961/PIX_OUT pixel_1961/CSA_VREF pixel
Xpixel_1950 pixel_1950/gring pixel_1950/VDD pixel_1950/GND pixel_1950/VREF pixel_1950/ROW_SEL
+ pixel_1950/NB1 pixel_1950/VBIAS pixel_1950/NB2 pixel_1950/AMP_IN pixel_1950/SF_IB
+ pixel_1950/PIX_OUT pixel_1950/CSA_VREF pixel
Xpixel_2695 pixel_2695/gring pixel_2695/VDD pixel_2695/GND pixel_2695/VREF pixel_2695/ROW_SEL
+ pixel_2695/NB1 pixel_2695/VBIAS pixel_2695/NB2 pixel_2695/AMP_IN pixel_2695/SF_IB
+ pixel_2695/PIX_OUT pixel_2695/CSA_VREF pixel
Xpixel_2684 pixel_2684/gring pixel_2684/VDD pixel_2684/GND pixel_2684/VREF pixel_2684/ROW_SEL
+ pixel_2684/NB1 pixel_2684/VBIAS pixel_2684/NB2 pixel_2684/AMP_IN pixel_2684/SF_IB
+ pixel_2684/PIX_OUT pixel_2684/CSA_VREF pixel
Xpixel_1994 pixel_1994/gring pixel_1994/VDD pixel_1994/GND pixel_1994/VREF pixel_1994/ROW_SEL
+ pixel_1994/NB1 pixel_1994/VBIAS pixel_1994/NB2 pixel_1994/AMP_IN pixel_1994/SF_IB
+ pixel_1994/PIX_OUT pixel_1994/CSA_VREF pixel
Xpixel_1983 pixel_1983/gring pixel_1983/VDD pixel_1983/GND pixel_1983/VREF pixel_1983/ROW_SEL
+ pixel_1983/NB1 pixel_1983/VBIAS pixel_1983/NB2 pixel_1983/AMP_IN pixel_1983/SF_IB
+ pixel_1983/PIX_OUT pixel_1983/CSA_VREF pixel
Xpixel_1972 pixel_1972/gring pixel_1972/VDD pixel_1972/GND pixel_1972/VREF pixel_1972/ROW_SEL
+ pixel_1972/NB1 pixel_1972/VBIAS pixel_1972/NB2 pixel_1972/AMP_IN pixel_1972/SF_IB
+ pixel_1972/PIX_OUT pixel_1972/CSA_VREF pixel
Xpixel_9009 pixel_9009/gring pixel_9009/VDD pixel_9009/GND pixel_9009/VREF pixel_9009/ROW_SEL
+ pixel_9009/NB1 pixel_9009/VBIAS pixel_9009/NB2 pixel_9009/AMP_IN pixel_9009/SF_IB
+ pixel_9009/PIX_OUT pixel_9009/CSA_VREF pixel
Xpixel_8308 pixel_8308/gring pixel_8308/VDD pixel_8308/GND pixel_8308/VREF pixel_8308/ROW_SEL
+ pixel_8308/NB1 pixel_8308/VBIAS pixel_8308/NB2 pixel_8308/AMP_IN pixel_8308/SF_IB
+ pixel_8308/PIX_OUT pixel_8308/CSA_VREF pixel
Xpixel_8319 pixel_8319/gring pixel_8319/VDD pixel_8319/GND pixel_8319/VREF pixel_8319/ROW_SEL
+ pixel_8319/NB1 pixel_8319/VBIAS pixel_8319/NB2 pixel_8319/AMP_IN pixel_8319/SF_IB
+ pixel_8319/PIX_OUT pixel_8319/CSA_VREF pixel
Xpixel_7607 pixel_7607/gring pixel_7607/VDD pixel_7607/GND pixel_7607/VREF pixel_7607/ROW_SEL
+ pixel_7607/NB1 pixel_7607/VBIAS pixel_7607/NB2 pixel_7607/AMP_IN pixel_7607/SF_IB
+ pixel_7607/PIX_OUT pixel_7607/CSA_VREF pixel
Xpixel_7618 pixel_7618/gring pixel_7618/VDD pixel_7618/GND pixel_7618/VREF pixel_7618/ROW_SEL
+ pixel_7618/NB1 pixel_7618/VBIAS pixel_7618/NB2 pixel_7618/AMP_IN pixel_7618/SF_IB
+ pixel_7618/PIX_OUT pixel_7618/CSA_VREF pixel
Xpixel_7629 pixel_7629/gring pixel_7629/VDD pixel_7629/GND pixel_7629/VREF pixel_7629/ROW_SEL
+ pixel_7629/NB1 pixel_7629/VBIAS pixel_7629/NB2 pixel_7629/AMP_IN pixel_7629/SF_IB
+ pixel_7629/PIX_OUT pixel_7629/CSA_VREF pixel
Xpixel_6906 pixel_6906/gring pixel_6906/VDD pixel_6906/GND pixel_6906/VREF pixel_6906/ROW_SEL
+ pixel_6906/NB1 pixel_6906/VBIAS pixel_6906/NB2 pixel_6906/AMP_IN pixel_6906/SF_IB
+ pixel_6906/PIX_OUT pixel_6906/CSA_VREF pixel
Xpixel_6917 pixel_6917/gring pixel_6917/VDD pixel_6917/GND pixel_6917/VREF pixel_6917/ROW_SEL
+ pixel_6917/NB1 pixel_6917/VBIAS pixel_6917/NB2 pixel_6917/AMP_IN pixel_6917/SF_IB
+ pixel_6917/PIX_OUT pixel_6917/CSA_VREF pixel
Xpixel_6928 pixel_6928/gring pixel_6928/VDD pixel_6928/GND pixel_6928/VREF pixel_6928/ROW_SEL
+ pixel_6928/NB1 pixel_6928/VBIAS pixel_6928/NB2 pixel_6928/AMP_IN pixel_6928/SF_IB
+ pixel_6928/PIX_OUT pixel_6928/CSA_VREF pixel
Xpixel_6939 pixel_6939/gring pixel_6939/VDD pixel_6939/GND pixel_6939/VREF pixel_6939/ROW_SEL
+ pixel_6939/NB1 pixel_6939/VBIAS pixel_6939/NB2 pixel_6939/AMP_IN pixel_6939/SF_IB
+ pixel_6939/PIX_OUT pixel_6939/CSA_VREF pixel
Xpixel_1224 pixel_1224/gring pixel_1224/VDD pixel_1224/GND pixel_1224/VREF pixel_1224/ROW_SEL
+ pixel_1224/NB1 pixel_1224/VBIAS pixel_1224/NB2 pixel_1224/AMP_IN pixel_1224/SF_IB
+ pixel_1224/PIX_OUT pixel_1224/CSA_VREF pixel
Xpixel_1213 pixel_1213/gring pixel_1213/VDD pixel_1213/GND pixel_1213/VREF pixel_1213/ROW_SEL
+ pixel_1213/NB1 pixel_1213/VBIAS pixel_1213/NB2 pixel_1213/AMP_IN pixel_1213/SF_IB
+ pixel_1213/PIX_OUT pixel_1213/CSA_VREF pixel
Xpixel_1202 pixel_1202/gring pixel_1202/VDD pixel_1202/GND pixel_1202/VREF pixel_1202/ROW_SEL
+ pixel_1202/NB1 pixel_1202/VBIAS pixel_1202/NB2 pixel_1202/AMP_IN pixel_1202/SF_IB
+ pixel_1202/PIX_OUT pixel_1202/CSA_VREF pixel
Xpixel_1257 pixel_1257/gring pixel_1257/VDD pixel_1257/GND pixel_1257/VREF pixel_1257/ROW_SEL
+ pixel_1257/NB1 pixel_1257/VBIAS pixel_1257/NB2 pixel_1257/AMP_IN pixel_1257/SF_IB
+ pixel_1257/PIX_OUT pixel_1257/CSA_VREF pixel
Xpixel_1246 pixel_1246/gring pixel_1246/VDD pixel_1246/GND pixel_1246/VREF pixel_1246/ROW_SEL
+ pixel_1246/NB1 pixel_1246/VBIAS pixel_1246/NB2 pixel_1246/AMP_IN pixel_1246/SF_IB
+ pixel_1246/PIX_OUT pixel_1246/CSA_VREF pixel
Xpixel_1235 pixel_1235/gring pixel_1235/VDD pixel_1235/GND pixel_1235/VREF pixel_1235/ROW_SEL
+ pixel_1235/NB1 pixel_1235/VBIAS pixel_1235/NB2 pixel_1235/AMP_IN pixel_1235/SF_IB
+ pixel_1235/PIX_OUT pixel_1235/CSA_VREF pixel
Xpixel_1279 pixel_1279/gring pixel_1279/VDD pixel_1279/GND pixel_1279/VREF pixel_1279/ROW_SEL
+ pixel_1279/NB1 pixel_1279/VBIAS pixel_1279/NB2 pixel_1279/AMP_IN pixel_1279/SF_IB
+ pixel_1279/PIX_OUT pixel_1279/CSA_VREF pixel
Xpixel_1268 pixel_1268/gring pixel_1268/VDD pixel_1268/GND pixel_1268/VREF pixel_1268/ROW_SEL
+ pixel_1268/NB1 pixel_1268/VBIAS pixel_1268/NB2 pixel_1268/AMP_IN pixel_1268/SF_IB
+ pixel_1268/PIX_OUT pixel_1268/CSA_VREF pixel
Xpixel_9532 pixel_9532/gring pixel_9532/VDD pixel_9532/GND pixel_9532/VREF pixel_9532/ROW_SEL
+ pixel_9532/NB1 pixel_9532/VBIAS pixel_9532/NB2 pixel_9532/AMP_IN pixel_9532/SF_IB
+ pixel_9532/PIX_OUT pixel_9532/CSA_VREF pixel
Xpixel_9521 pixel_9521/gring pixel_9521/VDD pixel_9521/GND pixel_9521/VREF pixel_9521/ROW_SEL
+ pixel_9521/NB1 pixel_9521/VBIAS pixel_9521/NB2 pixel_9521/AMP_IN pixel_9521/SF_IB
+ pixel_9521/PIX_OUT pixel_9521/CSA_VREF pixel
Xpixel_9510 pixel_9510/gring pixel_9510/VDD pixel_9510/GND pixel_9510/VREF pixel_9510/ROW_SEL
+ pixel_9510/NB1 pixel_9510/VBIAS pixel_9510/NB2 pixel_9510/AMP_IN pixel_9510/SF_IB
+ pixel_9510/PIX_OUT pixel_9510/CSA_VREF pixel
Xpixel_8820 pixel_8820/gring pixel_8820/VDD pixel_8820/GND pixel_8820/VREF pixel_8820/ROW_SEL
+ pixel_8820/NB1 pixel_8820/VBIAS pixel_8820/NB2 pixel_8820/AMP_IN pixel_8820/SF_IB
+ pixel_8820/PIX_OUT pixel_8820/CSA_VREF pixel
Xpixel_9565 pixel_9565/gring pixel_9565/VDD pixel_9565/GND pixel_9565/VREF pixel_9565/ROW_SEL
+ pixel_9565/NB1 pixel_9565/VBIAS pixel_9565/NB2 pixel_9565/AMP_IN pixel_9565/SF_IB
+ pixel_9565/PIX_OUT pixel_9565/CSA_VREF pixel
Xpixel_9554 pixel_9554/gring pixel_9554/VDD pixel_9554/GND pixel_9554/VREF pixel_9554/ROW_SEL
+ pixel_9554/NB1 pixel_9554/VBIAS pixel_9554/NB2 pixel_9554/AMP_IN pixel_9554/SF_IB
+ pixel_9554/PIX_OUT pixel_9554/CSA_VREF pixel
Xpixel_9543 pixel_9543/gring pixel_9543/VDD pixel_9543/GND pixel_9543/VREF pixel_9543/ROW_SEL
+ pixel_9543/NB1 pixel_9543/VBIAS pixel_9543/NB2 pixel_9543/AMP_IN pixel_9543/SF_IB
+ pixel_9543/PIX_OUT pixel_9543/CSA_VREF pixel
Xpixel_8864 pixel_8864/gring pixel_8864/VDD pixel_8864/GND pixel_8864/VREF pixel_8864/ROW_SEL
+ pixel_8864/NB1 pixel_8864/VBIAS pixel_8864/NB2 pixel_8864/AMP_IN pixel_8864/SF_IB
+ pixel_8864/PIX_OUT pixel_8864/CSA_VREF pixel
Xpixel_8853 pixel_8853/gring pixel_8853/VDD pixel_8853/GND pixel_8853/VREF pixel_8853/ROW_SEL
+ pixel_8853/NB1 pixel_8853/VBIAS pixel_8853/NB2 pixel_8853/AMP_IN pixel_8853/SF_IB
+ pixel_8853/PIX_OUT pixel_8853/CSA_VREF pixel
Xpixel_8842 pixel_8842/gring pixel_8842/VDD pixel_8842/GND pixel_8842/VREF pixel_8842/ROW_SEL
+ pixel_8842/NB1 pixel_8842/VBIAS pixel_8842/NB2 pixel_8842/AMP_IN pixel_8842/SF_IB
+ pixel_8842/PIX_OUT pixel_8842/CSA_VREF pixel
Xpixel_8831 pixel_8831/gring pixel_8831/VDD pixel_8831/GND pixel_8831/VREF pixel_8831/ROW_SEL
+ pixel_8831/NB1 pixel_8831/VBIAS pixel_8831/NB2 pixel_8831/AMP_IN pixel_8831/SF_IB
+ pixel_8831/PIX_OUT pixel_8831/CSA_VREF pixel
Xpixel_9598 pixel_9598/gring pixel_9598/VDD pixel_9598/GND pixel_9598/VREF pixel_9598/ROW_SEL
+ pixel_9598/NB1 pixel_9598/VBIAS pixel_9598/NB2 pixel_9598/AMP_IN pixel_9598/SF_IB
+ pixel_9598/PIX_OUT pixel_9598/CSA_VREF pixel
Xpixel_9587 pixel_9587/gring pixel_9587/VDD pixel_9587/GND pixel_9587/VREF pixel_9587/ROW_SEL
+ pixel_9587/NB1 pixel_9587/VBIAS pixel_9587/NB2 pixel_9587/AMP_IN pixel_9587/SF_IB
+ pixel_9587/PIX_OUT pixel_9587/CSA_VREF pixel
Xpixel_9576 pixel_9576/gring pixel_9576/VDD pixel_9576/GND pixel_9576/VREF pixel_9576/ROW_SEL
+ pixel_9576/NB1 pixel_9576/VBIAS pixel_9576/NB2 pixel_9576/AMP_IN pixel_9576/SF_IB
+ pixel_9576/PIX_OUT pixel_9576/CSA_VREF pixel
Xpixel_8897 pixel_8897/gring pixel_8897/VDD pixel_8897/GND pixel_8897/VREF pixel_8897/ROW_SEL
+ pixel_8897/NB1 pixel_8897/VBIAS pixel_8897/NB2 pixel_8897/AMP_IN pixel_8897/SF_IB
+ pixel_8897/PIX_OUT pixel_8897/CSA_VREF pixel
Xpixel_8886 pixel_8886/gring pixel_8886/VDD pixel_8886/GND pixel_8886/VREF pixel_8886/ROW_SEL
+ pixel_8886/NB1 pixel_8886/VBIAS pixel_8886/NB2 pixel_8886/AMP_IN pixel_8886/SF_IB
+ pixel_8886/PIX_OUT pixel_8886/CSA_VREF pixel
Xpixel_8875 pixel_8875/gring pixel_8875/VDD pixel_8875/GND pixel_8875/VREF pixel_8875/ROW_SEL
+ pixel_8875/NB1 pixel_8875/VBIAS pixel_8875/NB2 pixel_8875/AMP_IN pixel_8875/SF_IB
+ pixel_8875/PIX_OUT pixel_8875/CSA_VREF pixel
Xpixel_3193 pixel_3193/gring pixel_3193/VDD pixel_3193/GND pixel_3193/VREF pixel_3193/ROW_SEL
+ pixel_3193/NB1 pixel_3193/VBIAS pixel_3193/NB2 pixel_3193/AMP_IN pixel_3193/SF_IB
+ pixel_3193/PIX_OUT pixel_3193/CSA_VREF pixel
Xpixel_3182 pixel_3182/gring pixel_3182/VDD pixel_3182/GND pixel_3182/VREF pixel_3182/ROW_SEL
+ pixel_3182/NB1 pixel_3182/VBIAS pixel_3182/NB2 pixel_3182/AMP_IN pixel_3182/SF_IB
+ pixel_3182/PIX_OUT pixel_3182/CSA_VREF pixel
Xpixel_3171 pixel_3171/gring pixel_3171/VDD pixel_3171/GND pixel_3171/VREF pixel_3171/ROW_SEL
+ pixel_3171/NB1 pixel_3171/VBIAS pixel_3171/NB2 pixel_3171/AMP_IN pixel_3171/SF_IB
+ pixel_3171/PIX_OUT pixel_3171/CSA_VREF pixel
Xpixel_3160 pixel_3160/gring pixel_3160/VDD pixel_3160/GND pixel_3160/VREF pixel_3160/ROW_SEL
+ pixel_3160/NB1 pixel_3160/VBIAS pixel_3160/NB2 pixel_3160/AMP_IN pixel_3160/SF_IB
+ pixel_3160/PIX_OUT pixel_3160/CSA_VREF pixel
Xpixel_2481 pixel_2481/gring pixel_2481/VDD pixel_2481/GND pixel_2481/VREF pixel_2481/ROW_SEL
+ pixel_2481/NB1 pixel_2481/VBIAS pixel_2481/NB2 pixel_2481/AMP_IN pixel_2481/SF_IB
+ pixel_2481/PIX_OUT pixel_2481/CSA_VREF pixel
Xpixel_2470 pixel_2470/gring pixel_2470/VDD pixel_2470/GND pixel_2470/VREF pixel_2470/ROW_SEL
+ pixel_2470/NB1 pixel_2470/VBIAS pixel_2470/NB2 pixel_2470/AMP_IN pixel_2470/SF_IB
+ pixel_2470/PIX_OUT pixel_2470/CSA_VREF pixel
Xpixel_1780 pixel_1780/gring pixel_1780/VDD pixel_1780/GND pixel_1780/VREF pixel_1780/ROW_SEL
+ pixel_1780/NB1 pixel_1780/VBIAS pixel_1780/NB2 pixel_1780/AMP_IN pixel_1780/SF_IB
+ pixel_1780/PIX_OUT pixel_1780/CSA_VREF pixel
Xpixel_2492 pixel_2492/gring pixel_2492/VDD pixel_2492/GND pixel_2492/VREF pixel_2492/ROW_SEL
+ pixel_2492/NB1 pixel_2492/VBIAS pixel_2492/NB2 pixel_2492/AMP_IN pixel_2492/SF_IB
+ pixel_2492/PIX_OUT pixel_2492/CSA_VREF pixel
Xpixel_1791 pixel_1791/gring pixel_1791/VDD pixel_1791/GND pixel_1791/VREF pixel_1791/ROW_SEL
+ pixel_1791/NB1 pixel_1791/VBIAS pixel_1791/NB2 pixel_1791/AMP_IN pixel_1791/SF_IB
+ pixel_1791/PIX_OUT pixel_1791/CSA_VREF pixel
Xpixel_806 pixel_806/gring pixel_806/VDD pixel_806/GND pixel_806/VREF pixel_806/ROW_SEL
+ pixel_806/NB1 pixel_806/VBIAS pixel_806/NB2 pixel_806/AMP_IN pixel_806/SF_IB pixel_806/PIX_OUT
+ pixel_806/CSA_VREF pixel
Xpixel_839 pixel_839/gring pixel_839/VDD pixel_839/GND pixel_839/VREF pixel_839/ROW_SEL
+ pixel_839/NB1 pixel_839/VBIAS pixel_839/NB2 pixel_839/AMP_IN pixel_839/SF_IB pixel_839/PIX_OUT
+ pixel_839/CSA_VREF pixel
Xpixel_828 pixel_828/gring pixel_828/VDD pixel_828/GND pixel_828/VREF pixel_828/ROW_SEL
+ pixel_828/NB1 pixel_828/VBIAS pixel_828/NB2 pixel_828/AMP_IN pixel_828/SF_IB pixel_828/PIX_OUT
+ pixel_828/CSA_VREF pixel
Xpixel_817 pixel_817/gring pixel_817/VDD pixel_817/GND pixel_817/VREF pixel_817/ROW_SEL
+ pixel_817/NB1 pixel_817/VBIAS pixel_817/NB2 pixel_817/AMP_IN pixel_817/SF_IB pixel_817/PIX_OUT
+ pixel_817/CSA_VREF pixel
Xpixel_8105 pixel_8105/gring pixel_8105/VDD pixel_8105/GND pixel_8105/VREF pixel_8105/ROW_SEL
+ pixel_8105/NB1 pixel_8105/VBIAS pixel_8105/NB2 pixel_8105/AMP_IN pixel_8105/SF_IB
+ pixel_8105/PIX_OUT pixel_8105/CSA_VREF pixel
Xpixel_8116 pixel_8116/gring pixel_8116/VDD pixel_8116/GND pixel_8116/VREF pixel_8116/ROW_SEL
+ pixel_8116/NB1 pixel_8116/VBIAS pixel_8116/NB2 pixel_8116/AMP_IN pixel_8116/SF_IB
+ pixel_8116/PIX_OUT pixel_8116/CSA_VREF pixel
Xpixel_8127 pixel_8127/gring pixel_8127/VDD pixel_8127/GND pixel_8127/VREF pixel_8127/ROW_SEL
+ pixel_8127/NB1 pixel_8127/VBIAS pixel_8127/NB2 pixel_8127/AMP_IN pixel_8127/SF_IB
+ pixel_8127/PIX_OUT pixel_8127/CSA_VREF pixel
Xpixel_8138 pixel_8138/gring pixel_8138/VDD pixel_8138/GND pixel_8138/VREF pixel_8138/ROW_SEL
+ pixel_8138/NB1 pixel_8138/VBIAS pixel_8138/NB2 pixel_8138/AMP_IN pixel_8138/SF_IB
+ pixel_8138/PIX_OUT pixel_8138/CSA_VREF pixel
Xpixel_8149 pixel_8149/gring pixel_8149/VDD pixel_8149/GND pixel_8149/VREF pixel_8149/ROW_SEL
+ pixel_8149/NB1 pixel_8149/VBIAS pixel_8149/NB2 pixel_8149/AMP_IN pixel_8149/SF_IB
+ pixel_8149/PIX_OUT pixel_8149/CSA_VREF pixel
Xpixel_7404 pixel_7404/gring pixel_7404/VDD pixel_7404/GND pixel_7404/VREF pixel_7404/ROW_SEL
+ pixel_7404/NB1 pixel_7404/VBIAS pixel_7404/NB2 pixel_7404/AMP_IN pixel_7404/SF_IB
+ pixel_7404/PIX_OUT pixel_7404/CSA_VREF pixel
Xpixel_7415 pixel_7415/gring pixel_7415/VDD pixel_7415/GND pixel_7415/VREF pixel_7415/ROW_SEL
+ pixel_7415/NB1 pixel_7415/VBIAS pixel_7415/NB2 pixel_7415/AMP_IN pixel_7415/SF_IB
+ pixel_7415/PIX_OUT pixel_7415/CSA_VREF pixel
Xpixel_7426 pixel_7426/gring pixel_7426/VDD pixel_7426/GND pixel_7426/VREF pixel_7426/ROW_SEL
+ pixel_7426/NB1 pixel_7426/VBIAS pixel_7426/NB2 pixel_7426/AMP_IN pixel_7426/SF_IB
+ pixel_7426/PIX_OUT pixel_7426/CSA_VREF pixel
Xpixel_7437 pixel_7437/gring pixel_7437/VDD pixel_7437/GND pixel_7437/VREF pixel_7437/ROW_SEL
+ pixel_7437/NB1 pixel_7437/VBIAS pixel_7437/NB2 pixel_7437/AMP_IN pixel_7437/SF_IB
+ pixel_7437/PIX_OUT pixel_7437/CSA_VREF pixel
Xpixel_7448 pixel_7448/gring pixel_7448/VDD pixel_7448/GND pixel_7448/VREF pixel_7448/ROW_SEL
+ pixel_7448/NB1 pixel_7448/VBIAS pixel_7448/NB2 pixel_7448/AMP_IN pixel_7448/SF_IB
+ pixel_7448/PIX_OUT pixel_7448/CSA_VREF pixel
Xpixel_6703 pixel_6703/gring pixel_6703/VDD pixel_6703/GND pixel_6703/VREF pixel_6703/ROW_SEL
+ pixel_6703/NB1 pixel_6703/VBIAS pixel_6703/NB2 pixel_6703/AMP_IN pixel_6703/SF_IB
+ pixel_6703/PIX_OUT pixel_6703/CSA_VREF pixel
Xpixel_7459 pixel_7459/gring pixel_7459/VDD pixel_7459/GND pixel_7459/VREF pixel_7459/ROW_SEL
+ pixel_7459/NB1 pixel_7459/VBIAS pixel_7459/NB2 pixel_7459/AMP_IN pixel_7459/SF_IB
+ pixel_7459/PIX_OUT pixel_7459/CSA_VREF pixel
Xpixel_6714 pixel_6714/gring pixel_6714/VDD pixel_6714/GND pixel_6714/VREF pixel_6714/ROW_SEL
+ pixel_6714/NB1 pixel_6714/VBIAS pixel_6714/NB2 pixel_6714/AMP_IN pixel_6714/SF_IB
+ pixel_6714/PIX_OUT pixel_6714/CSA_VREF pixel
Xpixel_6725 pixel_6725/gring pixel_6725/VDD pixel_6725/GND pixel_6725/VREF pixel_6725/ROW_SEL
+ pixel_6725/NB1 pixel_6725/VBIAS pixel_6725/NB2 pixel_6725/AMP_IN pixel_6725/SF_IB
+ pixel_6725/PIX_OUT pixel_6725/CSA_VREF pixel
Xpixel_6736 pixel_6736/gring pixel_6736/VDD pixel_6736/GND pixel_6736/VREF pixel_6736/ROW_SEL
+ pixel_6736/NB1 pixel_6736/VBIAS pixel_6736/NB2 pixel_6736/AMP_IN pixel_6736/SF_IB
+ pixel_6736/PIX_OUT pixel_6736/CSA_VREF pixel
Xpixel_6747 pixel_6747/gring pixel_6747/VDD pixel_6747/GND pixel_6747/VREF pixel_6747/ROW_SEL
+ pixel_6747/NB1 pixel_6747/VBIAS pixel_6747/NB2 pixel_6747/AMP_IN pixel_6747/SF_IB
+ pixel_6747/PIX_OUT pixel_6747/CSA_VREF pixel
Xpixel_6758 pixel_6758/gring pixel_6758/VDD pixel_6758/GND pixel_6758/VREF pixel_6758/ROW_SEL
+ pixel_6758/NB1 pixel_6758/VBIAS pixel_6758/NB2 pixel_6758/AMP_IN pixel_6758/SF_IB
+ pixel_6758/PIX_OUT pixel_6758/CSA_VREF pixel
Xpixel_6769 pixel_6769/gring pixel_6769/VDD pixel_6769/GND pixel_6769/VREF pixel_6769/ROW_SEL
+ pixel_6769/NB1 pixel_6769/VBIAS pixel_6769/NB2 pixel_6769/AMP_IN pixel_6769/SF_IB
+ pixel_6769/PIX_OUT pixel_6769/CSA_VREF pixel
Xpixel_1032 pixel_1032/gring pixel_1032/VDD pixel_1032/GND pixel_1032/VREF pixel_1032/ROW_SEL
+ pixel_1032/NB1 pixel_1032/VBIAS pixel_1032/NB2 pixel_1032/AMP_IN pixel_1032/SF_IB
+ pixel_1032/PIX_OUT pixel_1032/CSA_VREF pixel
Xpixel_1021 pixel_1021/gring pixel_1021/VDD pixel_1021/GND pixel_1021/VREF pixel_1021/ROW_SEL
+ pixel_1021/NB1 pixel_1021/VBIAS pixel_1021/NB2 pixel_1021/AMP_IN pixel_1021/SF_IB
+ pixel_1021/PIX_OUT pixel_1021/CSA_VREF pixel
Xpixel_1010 pixel_1010/gring pixel_1010/VDD pixel_1010/GND pixel_1010/VREF pixel_1010/ROW_SEL
+ pixel_1010/NB1 pixel_1010/VBIAS pixel_1010/NB2 pixel_1010/AMP_IN pixel_1010/SF_IB
+ pixel_1010/PIX_OUT pixel_1010/CSA_VREF pixel
Xpixel_1065 pixel_1065/gring pixel_1065/VDD pixel_1065/GND pixel_1065/VREF pixel_1065/ROW_SEL
+ pixel_1065/NB1 pixel_1065/VBIAS pixel_1065/NB2 pixel_1065/AMP_IN pixel_1065/SF_IB
+ pixel_1065/PIX_OUT pixel_1065/CSA_VREF pixel
Xpixel_1054 pixel_1054/gring pixel_1054/VDD pixel_1054/GND pixel_1054/VREF pixel_1054/ROW_SEL
+ pixel_1054/NB1 pixel_1054/VBIAS pixel_1054/NB2 pixel_1054/AMP_IN pixel_1054/SF_IB
+ pixel_1054/PIX_OUT pixel_1054/CSA_VREF pixel
Xpixel_1043 pixel_1043/gring pixel_1043/VDD pixel_1043/GND pixel_1043/VREF pixel_1043/ROW_SEL
+ pixel_1043/NB1 pixel_1043/VBIAS pixel_1043/NB2 pixel_1043/AMP_IN pixel_1043/SF_IB
+ pixel_1043/PIX_OUT pixel_1043/CSA_VREF pixel
Xpixel_1098 pixel_1098/gring pixel_1098/VDD pixel_1098/GND pixel_1098/VREF pixel_1098/ROW_SEL
+ pixel_1098/NB1 pixel_1098/VBIAS pixel_1098/NB2 pixel_1098/AMP_IN pixel_1098/SF_IB
+ pixel_1098/PIX_OUT pixel_1098/CSA_VREF pixel
Xpixel_1087 pixel_1087/gring pixel_1087/VDD pixel_1087/GND pixel_1087/VREF pixel_1087/ROW_SEL
+ pixel_1087/NB1 pixel_1087/VBIAS pixel_1087/NB2 pixel_1087/AMP_IN pixel_1087/SF_IB
+ pixel_1087/PIX_OUT pixel_1087/CSA_VREF pixel
Xpixel_1076 pixel_1076/gring pixel_1076/VDD pixel_1076/GND pixel_1076/VREF pixel_1076/ROW_SEL
+ pixel_1076/NB1 pixel_1076/VBIAS pixel_1076/NB2 pixel_1076/AMP_IN pixel_1076/SF_IB
+ pixel_1076/PIX_OUT pixel_1076/CSA_VREF pixel
Xpixel_9340 pixel_9340/gring pixel_9340/VDD pixel_9340/GND pixel_9340/VREF pixel_9340/ROW_SEL
+ pixel_9340/NB1 pixel_9340/VBIAS pixel_9340/NB2 pixel_9340/AMP_IN pixel_9340/SF_IB
+ pixel_9340/PIX_OUT pixel_9340/CSA_VREF pixel
Xpixel_9373 pixel_9373/gring pixel_9373/VDD pixel_9373/GND pixel_9373/VREF pixel_9373/ROW_SEL
+ pixel_9373/NB1 pixel_9373/VBIAS pixel_9373/NB2 pixel_9373/AMP_IN pixel_9373/SF_IB
+ pixel_9373/PIX_OUT pixel_9373/CSA_VREF pixel
Xpixel_9362 pixel_9362/gring pixel_9362/VDD pixel_9362/GND pixel_9362/VREF pixel_9362/ROW_SEL
+ pixel_9362/NB1 pixel_9362/VBIAS pixel_9362/NB2 pixel_9362/AMP_IN pixel_9362/SF_IB
+ pixel_9362/PIX_OUT pixel_9362/CSA_VREF pixel
Xpixel_9351 pixel_9351/gring pixel_9351/VDD pixel_9351/GND pixel_9351/VREF pixel_9351/ROW_SEL
+ pixel_9351/NB1 pixel_9351/VBIAS pixel_9351/NB2 pixel_9351/AMP_IN pixel_9351/SF_IB
+ pixel_9351/PIX_OUT pixel_9351/CSA_VREF pixel
Xpixel_8672 pixel_8672/gring pixel_8672/VDD pixel_8672/GND pixel_8672/VREF pixel_8672/ROW_SEL
+ pixel_8672/NB1 pixel_8672/VBIAS pixel_8672/NB2 pixel_8672/AMP_IN pixel_8672/SF_IB
+ pixel_8672/PIX_OUT pixel_8672/CSA_VREF pixel
Xpixel_8661 pixel_8661/gring pixel_8661/VDD pixel_8661/GND pixel_8661/VREF pixel_8661/ROW_SEL
+ pixel_8661/NB1 pixel_8661/VBIAS pixel_8661/NB2 pixel_8661/AMP_IN pixel_8661/SF_IB
+ pixel_8661/PIX_OUT pixel_8661/CSA_VREF pixel
Xpixel_8650 pixel_8650/gring pixel_8650/VDD pixel_8650/GND pixel_8650/VREF pixel_8650/ROW_SEL
+ pixel_8650/NB1 pixel_8650/VBIAS pixel_8650/NB2 pixel_8650/AMP_IN pixel_8650/SF_IB
+ pixel_8650/PIX_OUT pixel_8650/CSA_VREF pixel
Xpixel_9395 pixel_9395/gring pixel_9395/VDD pixel_9395/GND pixel_9395/VREF pixel_9395/ROW_SEL
+ pixel_9395/NB1 pixel_9395/VBIAS pixel_9395/NB2 pixel_9395/AMP_IN pixel_9395/SF_IB
+ pixel_9395/PIX_OUT pixel_9395/CSA_VREF pixel
Xpixel_9384 pixel_9384/gring pixel_9384/VDD pixel_9384/GND pixel_9384/VREF pixel_9384/ROW_SEL
+ pixel_9384/NB1 pixel_9384/VBIAS pixel_9384/NB2 pixel_9384/AMP_IN pixel_9384/SF_IB
+ pixel_9384/PIX_OUT pixel_9384/CSA_VREF pixel
Xpixel_8694 pixel_8694/gring pixel_8694/VDD pixel_8694/GND pixel_8694/VREF pixel_8694/ROW_SEL
+ pixel_8694/NB1 pixel_8694/VBIAS pixel_8694/NB2 pixel_8694/AMP_IN pixel_8694/SF_IB
+ pixel_8694/PIX_OUT pixel_8694/CSA_VREF pixel
Xpixel_8683 pixel_8683/gring pixel_8683/VDD pixel_8683/GND pixel_8683/VREF pixel_8683/ROW_SEL
+ pixel_8683/NB1 pixel_8683/VBIAS pixel_8683/NB2 pixel_8683/AMP_IN pixel_8683/SF_IB
+ pixel_8683/PIX_OUT pixel_8683/CSA_VREF pixel
Xpixel_7960 pixel_7960/gring pixel_7960/VDD pixel_7960/GND pixel_7960/VREF pixel_7960/ROW_SEL
+ pixel_7960/NB1 pixel_7960/VBIAS pixel_7960/NB2 pixel_7960/AMP_IN pixel_7960/SF_IB
+ pixel_7960/PIX_OUT pixel_7960/CSA_VREF pixel
Xpixel_7971 pixel_7971/gring pixel_7971/VDD pixel_7971/GND pixel_7971/VREF pixel_7971/ROW_SEL
+ pixel_7971/NB1 pixel_7971/VBIAS pixel_7971/NB2 pixel_7971/AMP_IN pixel_7971/SF_IB
+ pixel_7971/PIX_OUT pixel_7971/CSA_VREF pixel
Xpixel_7982 pixel_7982/gring pixel_7982/VDD pixel_7982/GND pixel_7982/VREF pixel_7982/ROW_SEL
+ pixel_7982/NB1 pixel_7982/VBIAS pixel_7982/NB2 pixel_7982/AMP_IN pixel_7982/SF_IB
+ pixel_7982/PIX_OUT pixel_7982/CSA_VREF pixel
Xpixel_7993 pixel_7993/gring pixel_7993/VDD pixel_7993/GND pixel_7993/VREF pixel_7993/ROW_SEL
+ pixel_7993/NB1 pixel_7993/VBIAS pixel_7993/NB2 pixel_7993/AMP_IN pixel_7993/SF_IB
+ pixel_7993/PIX_OUT pixel_7993/CSA_VREF pixel
Xpixel_5309 pixel_5309/gring pixel_5309/VDD pixel_5309/GND pixel_5309/VREF pixel_5309/ROW_SEL
+ pixel_5309/NB1 pixel_5309/VBIAS pixel_5309/NB2 pixel_5309/AMP_IN pixel_5309/SF_IB
+ pixel_5309/PIX_OUT pixel_5309/CSA_VREF pixel
Xpixel_614 pixel_614/gring pixel_614/VDD pixel_614/GND pixel_614/VREF pixel_614/ROW_SEL
+ pixel_614/NB1 pixel_614/VBIAS pixel_614/NB2 pixel_614/AMP_IN pixel_614/SF_IB pixel_614/PIX_OUT
+ pixel_614/CSA_VREF pixel
Xpixel_603 pixel_603/gring pixel_603/VDD pixel_603/GND pixel_603/VREF pixel_603/ROW_SEL
+ pixel_603/NB1 pixel_603/VBIAS pixel_603/NB2 pixel_603/AMP_IN pixel_603/SF_IB pixel_603/PIX_OUT
+ pixel_603/CSA_VREF pixel
Xpixel_4608 pixel_4608/gring pixel_4608/VDD pixel_4608/GND pixel_4608/VREF pixel_4608/ROW_SEL
+ pixel_4608/NB1 pixel_4608/VBIAS pixel_4608/NB2 pixel_4608/AMP_IN pixel_4608/SF_IB
+ pixel_4608/PIX_OUT pixel_4608/CSA_VREF pixel
Xpixel_4619 pixel_4619/gring pixel_4619/VDD pixel_4619/GND pixel_4619/VREF pixel_4619/ROW_SEL
+ pixel_4619/NB1 pixel_4619/VBIAS pixel_4619/NB2 pixel_4619/AMP_IN pixel_4619/SF_IB
+ pixel_4619/PIX_OUT pixel_4619/CSA_VREF pixel
Xpixel_647 pixel_647/gring pixel_647/VDD pixel_647/GND pixel_647/VREF pixel_647/ROW_SEL
+ pixel_647/NB1 pixel_647/VBIAS pixel_647/NB2 pixel_647/AMP_IN pixel_647/SF_IB pixel_647/PIX_OUT
+ pixel_647/CSA_VREF pixel
Xpixel_636 pixel_636/gring pixel_636/VDD pixel_636/GND pixel_636/VREF pixel_636/ROW_SEL
+ pixel_636/NB1 pixel_636/VBIAS pixel_636/NB2 pixel_636/AMP_IN pixel_636/SF_IB pixel_636/PIX_OUT
+ pixel_636/CSA_VREF pixel
Xpixel_625 pixel_625/gring pixel_625/VDD pixel_625/GND pixel_625/VREF pixel_625/ROW_SEL
+ pixel_625/NB1 pixel_625/VBIAS pixel_625/NB2 pixel_625/AMP_IN pixel_625/SF_IB pixel_625/PIX_OUT
+ pixel_625/CSA_VREF pixel
Xpixel_3907 pixel_3907/gring pixel_3907/VDD pixel_3907/GND pixel_3907/VREF pixel_3907/ROW_SEL
+ pixel_3907/NB1 pixel_3907/VBIAS pixel_3907/NB2 pixel_3907/AMP_IN pixel_3907/SF_IB
+ pixel_3907/PIX_OUT pixel_3907/CSA_VREF pixel
Xpixel_669 pixel_669/gring pixel_669/VDD pixel_669/GND pixel_669/VREF pixel_669/ROW_SEL
+ pixel_669/NB1 pixel_669/VBIAS pixel_669/NB2 pixel_669/AMP_IN pixel_669/SF_IB pixel_669/PIX_OUT
+ pixel_669/CSA_VREF pixel
Xpixel_658 pixel_658/gring pixel_658/VDD pixel_658/GND pixel_658/VREF pixel_658/ROW_SEL
+ pixel_658/NB1 pixel_658/VBIAS pixel_658/NB2 pixel_658/AMP_IN pixel_658/SF_IB pixel_658/PIX_OUT
+ pixel_658/CSA_VREF pixel
Xpixel_3918 pixel_3918/gring pixel_3918/VDD pixel_3918/GND pixel_3918/VREF pixel_3918/ROW_SEL
+ pixel_3918/NB1 pixel_3918/VBIAS pixel_3918/NB2 pixel_3918/AMP_IN pixel_3918/SF_IB
+ pixel_3918/PIX_OUT pixel_3918/CSA_VREF pixel
Xpixel_3929 pixel_3929/gring pixel_3929/VDD pixel_3929/GND pixel_3929/VREF pixel_3929/ROW_SEL
+ pixel_3929/NB1 pixel_3929/VBIAS pixel_3929/NB2 pixel_3929/AMP_IN pixel_3929/SF_IB
+ pixel_3929/PIX_OUT pixel_3929/CSA_VREF pixel
Xpixel_7201 pixel_7201/gring pixel_7201/VDD pixel_7201/GND pixel_7201/VREF pixel_7201/ROW_SEL
+ pixel_7201/NB1 pixel_7201/VBIAS pixel_7201/NB2 pixel_7201/AMP_IN pixel_7201/SF_IB
+ pixel_7201/PIX_OUT pixel_7201/CSA_VREF pixel
Xpixel_7212 pixel_7212/gring pixel_7212/VDD pixel_7212/GND pixel_7212/VREF pixel_7212/ROW_SEL
+ pixel_7212/NB1 pixel_7212/VBIAS pixel_7212/NB2 pixel_7212/AMP_IN pixel_7212/SF_IB
+ pixel_7212/PIX_OUT pixel_7212/CSA_VREF pixel
Xpixel_7223 pixel_7223/gring pixel_7223/VDD pixel_7223/GND pixel_7223/VREF pixel_7223/ROW_SEL
+ pixel_7223/NB1 pixel_7223/VBIAS pixel_7223/NB2 pixel_7223/AMP_IN pixel_7223/SF_IB
+ pixel_7223/PIX_OUT pixel_7223/CSA_VREF pixel
Xpixel_7234 pixel_7234/gring pixel_7234/VDD pixel_7234/GND pixel_7234/VREF pixel_7234/ROW_SEL
+ pixel_7234/NB1 pixel_7234/VBIAS pixel_7234/NB2 pixel_7234/AMP_IN pixel_7234/SF_IB
+ pixel_7234/PIX_OUT pixel_7234/CSA_VREF pixel
Xpixel_7245 pixel_7245/gring pixel_7245/VDD pixel_7245/GND pixel_7245/VREF pixel_7245/ROW_SEL
+ pixel_7245/NB1 pixel_7245/VBIAS pixel_7245/NB2 pixel_7245/AMP_IN pixel_7245/SF_IB
+ pixel_7245/PIX_OUT pixel_7245/CSA_VREF pixel
Xpixel_7256 pixel_7256/gring pixel_7256/VDD pixel_7256/GND pixel_7256/VREF pixel_7256/ROW_SEL
+ pixel_7256/NB1 pixel_7256/VBIAS pixel_7256/NB2 pixel_7256/AMP_IN pixel_7256/SF_IB
+ pixel_7256/PIX_OUT pixel_7256/CSA_VREF pixel
Xpixel_6500 pixel_6500/gring pixel_6500/VDD pixel_6500/GND pixel_6500/VREF pixel_6500/ROW_SEL
+ pixel_6500/NB1 pixel_6500/VBIAS pixel_6500/NB2 pixel_6500/AMP_IN pixel_6500/SF_IB
+ pixel_6500/PIX_OUT pixel_6500/CSA_VREF pixel
Xpixel_6511 pixel_6511/gring pixel_6511/VDD pixel_6511/GND pixel_6511/VREF pixel_6511/ROW_SEL
+ pixel_6511/NB1 pixel_6511/VBIAS pixel_6511/NB2 pixel_6511/AMP_IN pixel_6511/SF_IB
+ pixel_6511/PIX_OUT pixel_6511/CSA_VREF pixel
Xpixel_7267 pixel_7267/gring pixel_7267/VDD pixel_7267/GND pixel_7267/VREF pixel_7267/ROW_SEL
+ pixel_7267/NB1 pixel_7267/VBIAS pixel_7267/NB2 pixel_7267/AMP_IN pixel_7267/SF_IB
+ pixel_7267/PIX_OUT pixel_7267/CSA_VREF pixel
Xpixel_7278 pixel_7278/gring pixel_7278/VDD pixel_7278/GND pixel_7278/VREF pixel_7278/ROW_SEL
+ pixel_7278/NB1 pixel_7278/VBIAS pixel_7278/NB2 pixel_7278/AMP_IN pixel_7278/SF_IB
+ pixel_7278/PIX_OUT pixel_7278/CSA_VREF pixel
Xpixel_7289 pixel_7289/gring pixel_7289/VDD pixel_7289/GND pixel_7289/VREF pixel_7289/ROW_SEL
+ pixel_7289/NB1 pixel_7289/VBIAS pixel_7289/NB2 pixel_7289/AMP_IN pixel_7289/SF_IB
+ pixel_7289/PIX_OUT pixel_7289/CSA_VREF pixel
Xpixel_6522 pixel_6522/gring pixel_6522/VDD pixel_6522/GND pixel_6522/VREF pixel_6522/ROW_SEL
+ pixel_6522/NB1 pixel_6522/VBIAS pixel_6522/NB2 pixel_6522/AMP_IN pixel_6522/SF_IB
+ pixel_6522/PIX_OUT pixel_6522/CSA_VREF pixel
Xpixel_6533 pixel_6533/gring pixel_6533/VDD pixel_6533/GND pixel_6533/VREF pixel_6533/ROW_SEL
+ pixel_6533/NB1 pixel_6533/VBIAS pixel_6533/NB2 pixel_6533/AMP_IN pixel_6533/SF_IB
+ pixel_6533/PIX_OUT pixel_6533/CSA_VREF pixel
Xpixel_6544 pixel_6544/gring pixel_6544/VDD pixel_6544/GND pixel_6544/VREF pixel_6544/ROW_SEL
+ pixel_6544/NB1 pixel_6544/VBIAS pixel_6544/NB2 pixel_6544/AMP_IN pixel_6544/SF_IB
+ pixel_6544/PIX_OUT pixel_6544/CSA_VREF pixel
Xpixel_6555 pixel_6555/gring pixel_6555/VDD pixel_6555/GND pixel_6555/VREF pixel_6555/ROW_SEL
+ pixel_6555/NB1 pixel_6555/VBIAS pixel_6555/NB2 pixel_6555/AMP_IN pixel_6555/SF_IB
+ pixel_6555/PIX_OUT pixel_6555/CSA_VREF pixel
Xpixel_6566 pixel_6566/gring pixel_6566/VDD pixel_6566/GND pixel_6566/VREF pixel_6566/ROW_SEL
+ pixel_6566/NB1 pixel_6566/VBIAS pixel_6566/NB2 pixel_6566/AMP_IN pixel_6566/SF_IB
+ pixel_6566/PIX_OUT pixel_6566/CSA_VREF pixel
Xpixel_6577 pixel_6577/gring pixel_6577/VDD pixel_6577/GND pixel_6577/VREF pixel_6577/ROW_SEL
+ pixel_6577/NB1 pixel_6577/VBIAS pixel_6577/NB2 pixel_6577/AMP_IN pixel_6577/SF_IB
+ pixel_6577/PIX_OUT pixel_6577/CSA_VREF pixel
Xpixel_6588 pixel_6588/gring pixel_6588/VDD pixel_6588/GND pixel_6588/VREF pixel_6588/ROW_SEL
+ pixel_6588/NB1 pixel_6588/VBIAS pixel_6588/NB2 pixel_6588/AMP_IN pixel_6588/SF_IB
+ pixel_6588/PIX_OUT pixel_6588/CSA_VREF pixel
Xpixel_5810 pixel_5810/gring pixel_5810/VDD pixel_5810/GND pixel_5810/VREF pixel_5810/ROW_SEL
+ pixel_5810/NB1 pixel_5810/VBIAS pixel_5810/NB2 pixel_5810/AMP_IN pixel_5810/SF_IB
+ pixel_5810/PIX_OUT pixel_5810/CSA_VREF pixel
Xpixel_5821 pixel_5821/gring pixel_5821/VDD pixel_5821/GND pixel_5821/VREF pixel_5821/ROW_SEL
+ pixel_5821/NB1 pixel_5821/VBIAS pixel_5821/NB2 pixel_5821/AMP_IN pixel_5821/SF_IB
+ pixel_5821/PIX_OUT pixel_5821/CSA_VREF pixel
Xpixel_5832 pixel_5832/gring pixel_5832/VDD pixel_5832/GND pixel_5832/VREF pixel_5832/ROW_SEL
+ pixel_5832/NB1 pixel_5832/VBIAS pixel_5832/NB2 pixel_5832/AMP_IN pixel_5832/SF_IB
+ pixel_5832/PIX_OUT pixel_5832/CSA_VREF pixel
Xpixel_5843 pixel_5843/gring pixel_5843/VDD pixel_5843/GND pixel_5843/VREF pixel_5843/ROW_SEL
+ pixel_5843/NB1 pixel_5843/VBIAS pixel_5843/NB2 pixel_5843/AMP_IN pixel_5843/SF_IB
+ pixel_5843/PIX_OUT pixel_5843/CSA_VREF pixel
Xpixel_6599 pixel_6599/gring pixel_6599/VDD pixel_6599/GND pixel_6599/VREF pixel_6599/ROW_SEL
+ pixel_6599/NB1 pixel_6599/VBIAS pixel_6599/NB2 pixel_6599/AMP_IN pixel_6599/SF_IB
+ pixel_6599/PIX_OUT pixel_6599/CSA_VREF pixel
Xpixel_5854 pixel_5854/gring pixel_5854/VDD pixel_5854/GND pixel_5854/VREF pixel_5854/ROW_SEL
+ pixel_5854/NB1 pixel_5854/VBIAS pixel_5854/NB2 pixel_5854/AMP_IN pixel_5854/SF_IB
+ pixel_5854/PIX_OUT pixel_5854/CSA_VREF pixel
Xpixel_5865 pixel_5865/gring pixel_5865/VDD pixel_5865/GND pixel_5865/VREF pixel_5865/ROW_SEL
+ pixel_5865/NB1 pixel_5865/VBIAS pixel_5865/NB2 pixel_5865/AMP_IN pixel_5865/SF_IB
+ pixel_5865/PIX_OUT pixel_5865/CSA_VREF pixel
Xpixel_5876 pixel_5876/gring pixel_5876/VDD pixel_5876/GND pixel_5876/VREF pixel_5876/ROW_SEL
+ pixel_5876/NB1 pixel_5876/VBIAS pixel_5876/NB2 pixel_5876/AMP_IN pixel_5876/SF_IB
+ pixel_5876/PIX_OUT pixel_5876/CSA_VREF pixel
Xpixel_5887 pixel_5887/gring pixel_5887/VDD pixel_5887/GND pixel_5887/VREF pixel_5887/ROW_SEL
+ pixel_5887/NB1 pixel_5887/VBIAS pixel_5887/NB2 pixel_5887/AMP_IN pixel_5887/SF_IB
+ pixel_5887/PIX_OUT pixel_5887/CSA_VREF pixel
Xpixel_5898 pixel_5898/gring pixel_5898/VDD pixel_5898/GND pixel_5898/VREF pixel_5898/ROW_SEL
+ pixel_5898/NB1 pixel_5898/VBIAS pixel_5898/NB2 pixel_5898/AMP_IN pixel_5898/SF_IB
+ pixel_5898/PIX_OUT pixel_5898/CSA_VREF pixel
Xpixel_9192 pixel_9192/gring pixel_9192/VDD pixel_9192/GND pixel_9192/VREF pixel_9192/ROW_SEL
+ pixel_9192/NB1 pixel_9192/VBIAS pixel_9192/NB2 pixel_9192/AMP_IN pixel_9192/SF_IB
+ pixel_9192/PIX_OUT pixel_9192/CSA_VREF pixel
Xpixel_9181 pixel_9181/gring pixel_9181/VDD pixel_9181/GND pixel_9181/VREF pixel_9181/ROW_SEL
+ pixel_9181/NB1 pixel_9181/VBIAS pixel_9181/NB2 pixel_9181/AMP_IN pixel_9181/SF_IB
+ pixel_9181/PIX_OUT pixel_9181/CSA_VREF pixel
Xpixel_9170 pixel_9170/gring pixel_9170/VDD pixel_9170/GND pixel_9170/VREF pixel_9170/ROW_SEL
+ pixel_9170/NB1 pixel_9170/VBIAS pixel_9170/NB2 pixel_9170/AMP_IN pixel_9170/SF_IB
+ pixel_9170/PIX_OUT pixel_9170/CSA_VREF pixel
Xpixel_8480 pixel_8480/gring pixel_8480/VDD pixel_8480/GND pixel_8480/VREF pixel_8480/ROW_SEL
+ pixel_8480/NB1 pixel_8480/VBIAS pixel_8480/NB2 pixel_8480/AMP_IN pixel_8480/SF_IB
+ pixel_8480/PIX_OUT pixel_8480/CSA_VREF pixel
Xpixel_8491 pixel_8491/gring pixel_8491/VDD pixel_8491/GND pixel_8491/VREF pixel_8491/ROW_SEL
+ pixel_8491/NB1 pixel_8491/VBIAS pixel_8491/NB2 pixel_8491/AMP_IN pixel_8491/SF_IB
+ pixel_8491/PIX_OUT pixel_8491/CSA_VREF pixel
Xpixel_7790 pixel_7790/gring pixel_7790/VDD pixel_7790/GND pixel_7790/VREF pixel_7790/ROW_SEL
+ pixel_7790/NB1 pixel_7790/VBIAS pixel_7790/NB2 pixel_7790/AMP_IN pixel_7790/SF_IB
+ pixel_7790/PIX_OUT pixel_7790/CSA_VREF pixel
Xpixel_5106 pixel_5106/gring pixel_5106/VDD pixel_5106/GND pixel_5106/VREF pixel_5106/ROW_SEL
+ pixel_5106/NB1 pixel_5106/VBIAS pixel_5106/NB2 pixel_5106/AMP_IN pixel_5106/SF_IB
+ pixel_5106/PIX_OUT pixel_5106/CSA_VREF pixel
Xpixel_5117 pixel_5117/gring pixel_5117/VDD pixel_5117/GND pixel_5117/VREF pixel_5117/ROW_SEL
+ pixel_5117/NB1 pixel_5117/VBIAS pixel_5117/NB2 pixel_5117/AMP_IN pixel_5117/SF_IB
+ pixel_5117/PIX_OUT pixel_5117/CSA_VREF pixel
Xpixel_5128 pixel_5128/gring pixel_5128/VDD pixel_5128/GND pixel_5128/VREF pixel_5128/ROW_SEL
+ pixel_5128/NB1 pixel_5128/VBIAS pixel_5128/NB2 pixel_5128/AMP_IN pixel_5128/SF_IB
+ pixel_5128/PIX_OUT pixel_5128/CSA_VREF pixel
Xpixel_422 pixel_422/gring pixel_422/VDD pixel_422/GND pixel_422/VREF pixel_422/ROW_SEL
+ pixel_422/NB1 pixel_422/VBIAS pixel_422/NB2 pixel_422/AMP_IN pixel_422/SF_IB pixel_422/PIX_OUT
+ pixel_422/CSA_VREF pixel
Xpixel_411 pixel_411/gring pixel_411/VDD pixel_411/GND pixel_411/VREF pixel_411/ROW_SEL
+ pixel_411/NB1 pixel_411/VBIAS pixel_411/NB2 pixel_411/AMP_IN pixel_411/SF_IB pixel_411/PIX_OUT
+ pixel_411/CSA_VREF pixel
Xpixel_400 pixel_400/gring pixel_400/VDD pixel_400/GND pixel_400/VREF pixel_400/ROW_SEL
+ pixel_400/NB1 pixel_400/VBIAS pixel_400/NB2 pixel_400/AMP_IN pixel_400/SF_IB pixel_400/PIX_OUT
+ pixel_400/CSA_VREF pixel
Xpixel_5139 pixel_5139/gring pixel_5139/VDD pixel_5139/GND pixel_5139/VREF pixel_5139/ROW_SEL
+ pixel_5139/NB1 pixel_5139/VBIAS pixel_5139/NB2 pixel_5139/AMP_IN pixel_5139/SF_IB
+ pixel_5139/PIX_OUT pixel_5139/CSA_VREF pixel
Xpixel_4405 pixel_4405/gring pixel_4405/VDD pixel_4405/GND pixel_4405/VREF pixel_4405/ROW_SEL
+ pixel_4405/NB1 pixel_4405/VBIAS pixel_4405/NB2 pixel_4405/AMP_IN pixel_4405/SF_IB
+ pixel_4405/PIX_OUT pixel_4405/CSA_VREF pixel
Xpixel_4416 pixel_4416/gring pixel_4416/VDD pixel_4416/GND pixel_4416/VREF pixel_4416/ROW_SEL
+ pixel_4416/NB1 pixel_4416/VBIAS pixel_4416/NB2 pixel_4416/AMP_IN pixel_4416/SF_IB
+ pixel_4416/PIX_OUT pixel_4416/CSA_VREF pixel
Xpixel_4427 pixel_4427/gring pixel_4427/VDD pixel_4427/GND pixel_4427/VREF pixel_4427/ROW_SEL
+ pixel_4427/NB1 pixel_4427/VBIAS pixel_4427/NB2 pixel_4427/AMP_IN pixel_4427/SF_IB
+ pixel_4427/PIX_OUT pixel_4427/CSA_VREF pixel
Xpixel_455 pixel_455/gring pixel_455/VDD pixel_455/GND pixel_455/VREF pixel_455/ROW_SEL
+ pixel_455/NB1 pixel_455/VBIAS pixel_455/NB2 pixel_455/AMP_IN pixel_455/SF_IB pixel_455/PIX_OUT
+ pixel_455/CSA_VREF pixel
Xpixel_444 pixel_444/gring pixel_444/VDD pixel_444/GND pixel_444/VREF pixel_444/ROW_SEL
+ pixel_444/NB1 pixel_444/VBIAS pixel_444/NB2 pixel_444/AMP_IN pixel_444/SF_IB pixel_444/PIX_OUT
+ pixel_444/CSA_VREF pixel
Xpixel_433 pixel_433/gring pixel_433/VDD pixel_433/GND pixel_433/VREF pixel_433/ROW_SEL
+ pixel_433/NB1 pixel_433/VBIAS pixel_433/NB2 pixel_433/AMP_IN pixel_433/SF_IB pixel_433/PIX_OUT
+ pixel_433/CSA_VREF pixel
Xpixel_3715 pixel_3715/gring pixel_3715/VDD pixel_3715/GND pixel_3715/VREF pixel_3715/ROW_SEL
+ pixel_3715/NB1 pixel_3715/VBIAS pixel_3715/NB2 pixel_3715/AMP_IN pixel_3715/SF_IB
+ pixel_3715/PIX_OUT pixel_3715/CSA_VREF pixel
Xpixel_3704 pixel_3704/gring pixel_3704/VDD pixel_3704/GND pixel_3704/VREF pixel_3704/ROW_SEL
+ pixel_3704/NB1 pixel_3704/VBIAS pixel_3704/NB2 pixel_3704/AMP_IN pixel_3704/SF_IB
+ pixel_3704/PIX_OUT pixel_3704/CSA_VREF pixel
Xpixel_4438 pixel_4438/gring pixel_4438/VDD pixel_4438/GND pixel_4438/VREF pixel_4438/ROW_SEL
+ pixel_4438/NB1 pixel_4438/VBIAS pixel_4438/NB2 pixel_4438/AMP_IN pixel_4438/SF_IB
+ pixel_4438/PIX_OUT pixel_4438/CSA_VREF pixel
Xpixel_4449 pixel_4449/gring pixel_4449/VDD pixel_4449/GND pixel_4449/VREF pixel_4449/ROW_SEL
+ pixel_4449/NB1 pixel_4449/VBIAS pixel_4449/NB2 pixel_4449/AMP_IN pixel_4449/SF_IB
+ pixel_4449/PIX_OUT pixel_4449/CSA_VREF pixel
Xpixel_499 pixel_499/gring pixel_499/VDD pixel_499/GND pixel_499/VREF pixel_499/ROW_SEL
+ pixel_499/NB1 pixel_499/VBIAS pixel_499/NB2 pixel_499/AMP_IN pixel_499/SF_IB pixel_499/PIX_OUT
+ pixel_499/CSA_VREF pixel
Xpixel_488 pixel_488/gring pixel_488/VDD pixel_488/GND pixel_488/VREF pixel_488/ROW_SEL
+ pixel_488/NB1 pixel_488/VBIAS pixel_488/NB2 pixel_488/AMP_IN pixel_488/SF_IB pixel_488/PIX_OUT
+ pixel_488/CSA_VREF pixel
Xpixel_477 pixel_477/gring pixel_477/VDD pixel_477/GND pixel_477/VREF pixel_477/ROW_SEL
+ pixel_477/NB1 pixel_477/VBIAS pixel_477/NB2 pixel_477/AMP_IN pixel_477/SF_IB pixel_477/PIX_OUT
+ pixel_477/CSA_VREF pixel
Xpixel_466 pixel_466/gring pixel_466/VDD pixel_466/GND pixel_466/VREF pixel_466/ROW_SEL
+ pixel_466/NB1 pixel_466/VBIAS pixel_466/NB2 pixel_466/AMP_IN pixel_466/SF_IB pixel_466/PIX_OUT
+ pixel_466/CSA_VREF pixel
Xpixel_3759 pixel_3759/gring pixel_3759/VDD pixel_3759/GND pixel_3759/VREF pixel_3759/ROW_SEL
+ pixel_3759/NB1 pixel_3759/VBIAS pixel_3759/NB2 pixel_3759/AMP_IN pixel_3759/SF_IB
+ pixel_3759/PIX_OUT pixel_3759/CSA_VREF pixel
Xpixel_3748 pixel_3748/gring pixel_3748/VDD pixel_3748/GND pixel_3748/VREF pixel_3748/ROW_SEL
+ pixel_3748/NB1 pixel_3748/VBIAS pixel_3748/NB2 pixel_3748/AMP_IN pixel_3748/SF_IB
+ pixel_3748/PIX_OUT pixel_3748/CSA_VREF pixel
Xpixel_3737 pixel_3737/gring pixel_3737/VDD pixel_3737/GND pixel_3737/VREF pixel_3737/ROW_SEL
+ pixel_3737/NB1 pixel_3737/VBIAS pixel_3737/NB2 pixel_3737/AMP_IN pixel_3737/SF_IB
+ pixel_3737/PIX_OUT pixel_3737/CSA_VREF pixel
Xpixel_3726 pixel_3726/gring pixel_3726/VDD pixel_3726/GND pixel_3726/VREF pixel_3726/ROW_SEL
+ pixel_3726/NB1 pixel_3726/VBIAS pixel_3726/NB2 pixel_3726/AMP_IN pixel_3726/SF_IB
+ pixel_3726/PIX_OUT pixel_3726/CSA_VREF pixel
Xpixel_7020 pixel_7020/gring pixel_7020/VDD pixel_7020/GND pixel_7020/VREF pixel_7020/ROW_SEL
+ pixel_7020/NB1 pixel_7020/VBIAS pixel_7020/NB2 pixel_7020/AMP_IN pixel_7020/SF_IB
+ pixel_7020/PIX_OUT pixel_7020/CSA_VREF pixel
Xpixel_7031 pixel_7031/gring pixel_7031/VDD pixel_7031/GND pixel_7031/VREF pixel_7031/ROW_SEL
+ pixel_7031/NB1 pixel_7031/VBIAS pixel_7031/NB2 pixel_7031/AMP_IN pixel_7031/SF_IB
+ pixel_7031/PIX_OUT pixel_7031/CSA_VREF pixel
Xpixel_7042 pixel_7042/gring pixel_7042/VDD pixel_7042/GND pixel_7042/VREF pixel_7042/ROW_SEL
+ pixel_7042/NB1 pixel_7042/VBIAS pixel_7042/NB2 pixel_7042/AMP_IN pixel_7042/SF_IB
+ pixel_7042/PIX_OUT pixel_7042/CSA_VREF pixel
Xpixel_7053 pixel_7053/gring pixel_7053/VDD pixel_7053/GND pixel_7053/VREF pixel_7053/ROW_SEL
+ pixel_7053/NB1 pixel_7053/VBIAS pixel_7053/NB2 pixel_7053/AMP_IN pixel_7053/SF_IB
+ pixel_7053/PIX_OUT pixel_7053/CSA_VREF pixel
Xpixel_7064 pixel_7064/gring pixel_7064/VDD pixel_7064/GND pixel_7064/VREF pixel_7064/ROW_SEL
+ pixel_7064/NB1 pixel_7064/VBIAS pixel_7064/NB2 pixel_7064/AMP_IN pixel_7064/SF_IB
+ pixel_7064/PIX_OUT pixel_7064/CSA_VREF pixel
Xpixel_7075 pixel_7075/gring pixel_7075/VDD pixel_7075/GND pixel_7075/VREF pixel_7075/ROW_SEL
+ pixel_7075/NB1 pixel_7075/VBIAS pixel_7075/NB2 pixel_7075/AMP_IN pixel_7075/SF_IB
+ pixel_7075/PIX_OUT pixel_7075/CSA_VREF pixel
Xpixel_7086 pixel_7086/gring pixel_7086/VDD pixel_7086/GND pixel_7086/VREF pixel_7086/ROW_SEL
+ pixel_7086/NB1 pixel_7086/VBIAS pixel_7086/NB2 pixel_7086/AMP_IN pixel_7086/SF_IB
+ pixel_7086/PIX_OUT pixel_7086/CSA_VREF pixel
Xpixel_7097 pixel_7097/gring pixel_7097/VDD pixel_7097/GND pixel_7097/VREF pixel_7097/ROW_SEL
+ pixel_7097/NB1 pixel_7097/VBIAS pixel_7097/NB2 pixel_7097/AMP_IN pixel_7097/SF_IB
+ pixel_7097/PIX_OUT pixel_7097/CSA_VREF pixel
Xpixel_6330 pixel_6330/gring pixel_6330/VDD pixel_6330/GND pixel_6330/VREF pixel_6330/ROW_SEL
+ pixel_6330/NB1 pixel_6330/VBIAS pixel_6330/NB2 pixel_6330/AMP_IN pixel_6330/SF_IB
+ pixel_6330/PIX_OUT pixel_6330/CSA_VREF pixel
Xpixel_6341 pixel_6341/gring pixel_6341/VDD pixel_6341/GND pixel_6341/VREF pixel_6341/ROW_SEL
+ pixel_6341/NB1 pixel_6341/VBIAS pixel_6341/NB2 pixel_6341/AMP_IN pixel_6341/SF_IB
+ pixel_6341/PIX_OUT pixel_6341/CSA_VREF pixel
Xpixel_6352 pixel_6352/gring pixel_6352/VDD pixel_6352/GND pixel_6352/VREF pixel_6352/ROW_SEL
+ pixel_6352/NB1 pixel_6352/VBIAS pixel_6352/NB2 pixel_6352/AMP_IN pixel_6352/SF_IB
+ pixel_6352/PIX_OUT pixel_6352/CSA_VREF pixel
Xpixel_6363 pixel_6363/gring pixel_6363/VDD pixel_6363/GND pixel_6363/VREF pixel_6363/ROW_SEL
+ pixel_6363/NB1 pixel_6363/VBIAS pixel_6363/NB2 pixel_6363/AMP_IN pixel_6363/SF_IB
+ pixel_6363/PIX_OUT pixel_6363/CSA_VREF pixel
Xpixel_6374 pixel_6374/gring pixel_6374/VDD pixel_6374/GND pixel_6374/VREF pixel_6374/ROW_SEL
+ pixel_6374/NB1 pixel_6374/VBIAS pixel_6374/NB2 pixel_6374/AMP_IN pixel_6374/SF_IB
+ pixel_6374/PIX_OUT pixel_6374/CSA_VREF pixel
Xpixel_6385 pixel_6385/gring pixel_6385/VDD pixel_6385/GND pixel_6385/VREF pixel_6385/ROW_SEL
+ pixel_6385/NB1 pixel_6385/VBIAS pixel_6385/NB2 pixel_6385/AMP_IN pixel_6385/SF_IB
+ pixel_6385/PIX_OUT pixel_6385/CSA_VREF pixel
Xpixel_6396 pixel_6396/gring pixel_6396/VDD pixel_6396/GND pixel_6396/VREF pixel_6396/ROW_SEL
+ pixel_6396/NB1 pixel_6396/VBIAS pixel_6396/NB2 pixel_6396/AMP_IN pixel_6396/SF_IB
+ pixel_6396/PIX_OUT pixel_6396/CSA_VREF pixel
Xpixel_5640 pixel_5640/gring pixel_5640/VDD pixel_5640/GND pixel_5640/VREF pixel_5640/ROW_SEL
+ pixel_5640/NB1 pixel_5640/VBIAS pixel_5640/NB2 pixel_5640/AMP_IN pixel_5640/SF_IB
+ pixel_5640/PIX_OUT pixel_5640/CSA_VREF pixel
Xpixel_5651 pixel_5651/gring pixel_5651/VDD pixel_5651/GND pixel_5651/VREF pixel_5651/ROW_SEL
+ pixel_5651/NB1 pixel_5651/VBIAS pixel_5651/NB2 pixel_5651/AMP_IN pixel_5651/SF_IB
+ pixel_5651/PIX_OUT pixel_5651/CSA_VREF pixel
Xpixel_5662 pixel_5662/gring pixel_5662/VDD pixel_5662/GND pixel_5662/VREF pixel_5662/ROW_SEL
+ pixel_5662/NB1 pixel_5662/VBIAS pixel_5662/NB2 pixel_5662/AMP_IN pixel_5662/SF_IB
+ pixel_5662/PIX_OUT pixel_5662/CSA_VREF pixel
Xpixel_5673 pixel_5673/gring pixel_5673/VDD pixel_5673/GND pixel_5673/VREF pixel_5673/ROW_SEL
+ pixel_5673/NB1 pixel_5673/VBIAS pixel_5673/NB2 pixel_5673/AMP_IN pixel_5673/SF_IB
+ pixel_5673/PIX_OUT pixel_5673/CSA_VREF pixel
Xpixel_5684 pixel_5684/gring pixel_5684/VDD pixel_5684/GND pixel_5684/VREF pixel_5684/ROW_SEL
+ pixel_5684/NB1 pixel_5684/VBIAS pixel_5684/NB2 pixel_5684/AMP_IN pixel_5684/SF_IB
+ pixel_5684/PIX_OUT pixel_5684/CSA_VREF pixel
Xpixel_5695 pixel_5695/gring pixel_5695/VDD pixel_5695/GND pixel_5695/VREF pixel_5695/ROW_SEL
+ pixel_5695/NB1 pixel_5695/VBIAS pixel_5695/NB2 pixel_5695/AMP_IN pixel_5695/SF_IB
+ pixel_5695/PIX_OUT pixel_5695/CSA_VREF pixel
Xpixel_4950 pixel_4950/gring pixel_4950/VDD pixel_4950/GND pixel_4950/VREF pixel_4950/ROW_SEL
+ pixel_4950/NB1 pixel_4950/VBIAS pixel_4950/NB2 pixel_4950/AMP_IN pixel_4950/SF_IB
+ pixel_4950/PIX_OUT pixel_4950/CSA_VREF pixel
Xpixel_4961 pixel_4961/gring pixel_4961/VDD pixel_4961/GND pixel_4961/VREF pixel_4961/ROW_SEL
+ pixel_4961/NB1 pixel_4961/VBIAS pixel_4961/NB2 pixel_4961/AMP_IN pixel_4961/SF_IB
+ pixel_4961/PIX_OUT pixel_4961/CSA_VREF pixel
Xpixel_4972 pixel_4972/gring pixel_4972/VDD pixel_4972/GND pixel_4972/VREF pixel_4972/ROW_SEL
+ pixel_4972/NB1 pixel_4972/VBIAS pixel_4972/NB2 pixel_4972/AMP_IN pixel_4972/SF_IB
+ pixel_4972/PIX_OUT pixel_4972/CSA_VREF pixel
Xpixel_4983 pixel_4983/gring pixel_4983/VDD pixel_4983/GND pixel_4983/VREF pixel_4983/ROW_SEL
+ pixel_4983/NB1 pixel_4983/VBIAS pixel_4983/NB2 pixel_4983/AMP_IN pixel_4983/SF_IB
+ pixel_4983/PIX_OUT pixel_4983/CSA_VREF pixel
Xpixel_4994 pixel_4994/gring pixel_4994/VDD pixel_4994/GND pixel_4994/VREF pixel_4994/ROW_SEL
+ pixel_4994/NB1 pixel_4994/VBIAS pixel_4994/NB2 pixel_4994/AMP_IN pixel_4994/SF_IB
+ pixel_4994/PIX_OUT pixel_4994/CSA_VREF pixel
Xpixel_1609 pixel_1609/gring pixel_1609/VDD pixel_1609/GND pixel_1609/VREF pixel_1609/ROW_SEL
+ pixel_1609/NB1 pixel_1609/VBIAS pixel_1609/NB2 pixel_1609/AMP_IN pixel_1609/SF_IB
+ pixel_1609/PIX_OUT pixel_1609/CSA_VREF pixel
Xpixel_9906 pixel_9906/gring pixel_9906/VDD pixel_9906/GND pixel_9906/VREF pixel_9906/ROW_SEL
+ pixel_9906/NB1 pixel_9906/VBIAS pixel_9906/NB2 pixel_9906/AMP_IN pixel_9906/SF_IB
+ pixel_9906/PIX_OUT pixel_9906/CSA_VREF pixel
Xpixel_9939 pixel_9939/gring pixel_9939/VDD pixel_9939/GND pixel_9939/VREF pixel_9939/ROW_SEL
+ pixel_9939/NB1 pixel_9939/VBIAS pixel_9939/NB2 pixel_9939/AMP_IN pixel_9939/SF_IB
+ pixel_9939/PIX_OUT pixel_9939/CSA_VREF pixel
Xpixel_9928 pixel_9928/gring pixel_9928/VDD pixel_9928/GND pixel_9928/VREF pixel_9928/ROW_SEL
+ pixel_9928/NB1 pixel_9928/VBIAS pixel_9928/NB2 pixel_9928/AMP_IN pixel_9928/SF_IB
+ pixel_9928/PIX_OUT pixel_9928/CSA_VREF pixel
Xpixel_9917 pixel_9917/gring pixel_9917/VDD pixel_9917/GND pixel_9917/VREF pixel_9917/ROW_SEL
+ pixel_9917/NB1 pixel_9917/VBIAS pixel_9917/NB2 pixel_9917/AMP_IN pixel_9917/SF_IB
+ pixel_9917/PIX_OUT pixel_9917/CSA_VREF pixel
Xpixel_4202 pixel_4202/gring pixel_4202/VDD pixel_4202/GND pixel_4202/VREF pixel_4202/ROW_SEL
+ pixel_4202/NB1 pixel_4202/VBIAS pixel_4202/NB2 pixel_4202/AMP_IN pixel_4202/SF_IB
+ pixel_4202/PIX_OUT pixel_4202/CSA_VREF pixel
Xpixel_230 pixel_230/gring pixel_230/VDD pixel_230/GND pixel_230/VREF pixel_230/ROW_SEL
+ pixel_230/NB1 pixel_230/VBIAS pixel_230/NB2 pixel_230/AMP_IN pixel_230/SF_IB pixel_230/PIX_OUT
+ pixel_230/CSA_VREF pixel
Xpixel_4213 pixel_4213/gring pixel_4213/VDD pixel_4213/GND pixel_4213/VREF pixel_4213/ROW_SEL
+ pixel_4213/NB1 pixel_4213/VBIAS pixel_4213/NB2 pixel_4213/AMP_IN pixel_4213/SF_IB
+ pixel_4213/PIX_OUT pixel_4213/CSA_VREF pixel
Xpixel_4224 pixel_4224/gring pixel_4224/VDD pixel_4224/GND pixel_4224/VREF pixel_4224/ROW_SEL
+ pixel_4224/NB1 pixel_4224/VBIAS pixel_4224/NB2 pixel_4224/AMP_IN pixel_4224/SF_IB
+ pixel_4224/PIX_OUT pixel_4224/CSA_VREF pixel
Xpixel_4235 pixel_4235/gring pixel_4235/VDD pixel_4235/GND pixel_4235/VREF pixel_4235/ROW_SEL
+ pixel_4235/NB1 pixel_4235/VBIAS pixel_4235/NB2 pixel_4235/AMP_IN pixel_4235/SF_IB
+ pixel_4235/PIX_OUT pixel_4235/CSA_VREF pixel
Xpixel_274 pixel_274/gring pixel_274/VDD pixel_274/GND pixel_274/VREF pixel_274/ROW_SEL
+ pixel_274/NB1 pixel_274/VBIAS pixel_274/NB2 pixel_274/AMP_IN pixel_274/SF_IB pixel_274/PIX_OUT
+ pixel_274/CSA_VREF pixel
Xpixel_263 pixel_263/gring pixel_263/VDD pixel_263/GND pixel_263/VREF pixel_263/ROW_SEL
+ pixel_263/NB1 pixel_263/VBIAS pixel_263/NB2 pixel_263/AMP_IN pixel_263/SF_IB pixel_263/PIX_OUT
+ pixel_263/CSA_VREF pixel
Xpixel_252 pixel_252/gring pixel_252/VDD pixel_252/GND pixel_252/VREF pixel_252/ROW_SEL
+ pixel_252/NB1 pixel_252/VBIAS pixel_252/NB2 pixel_252/AMP_IN pixel_252/SF_IB pixel_252/PIX_OUT
+ pixel_252/CSA_VREF pixel
Xpixel_241 pixel_241/gring pixel_241/VDD pixel_241/GND pixel_241/VREF pixel_241/ROW_SEL
+ pixel_241/NB1 pixel_241/VBIAS pixel_241/NB2 pixel_241/AMP_IN pixel_241/SF_IB pixel_241/PIX_OUT
+ pixel_241/CSA_VREF pixel
Xpixel_3534 pixel_3534/gring pixel_3534/VDD pixel_3534/GND pixel_3534/VREF pixel_3534/ROW_SEL
+ pixel_3534/NB1 pixel_3534/VBIAS pixel_3534/NB2 pixel_3534/AMP_IN pixel_3534/SF_IB
+ pixel_3534/PIX_OUT pixel_3534/CSA_VREF pixel
Xpixel_3523 pixel_3523/gring pixel_3523/VDD pixel_3523/GND pixel_3523/VREF pixel_3523/ROW_SEL
+ pixel_3523/NB1 pixel_3523/VBIAS pixel_3523/NB2 pixel_3523/AMP_IN pixel_3523/SF_IB
+ pixel_3523/PIX_OUT pixel_3523/CSA_VREF pixel
Xpixel_3512 pixel_3512/gring pixel_3512/VDD pixel_3512/GND pixel_3512/VREF pixel_3512/ROW_SEL
+ pixel_3512/NB1 pixel_3512/VBIAS pixel_3512/NB2 pixel_3512/AMP_IN pixel_3512/SF_IB
+ pixel_3512/PIX_OUT pixel_3512/CSA_VREF pixel
Xpixel_3501 pixel_3501/gring pixel_3501/VDD pixel_3501/GND pixel_3501/VREF pixel_3501/ROW_SEL
+ pixel_3501/NB1 pixel_3501/VBIAS pixel_3501/NB2 pixel_3501/AMP_IN pixel_3501/SF_IB
+ pixel_3501/PIX_OUT pixel_3501/CSA_VREF pixel
Xpixel_4246 pixel_4246/gring pixel_4246/VDD pixel_4246/GND pixel_4246/VREF pixel_4246/ROW_SEL
+ pixel_4246/NB1 pixel_4246/VBIAS pixel_4246/NB2 pixel_4246/AMP_IN pixel_4246/SF_IB
+ pixel_4246/PIX_OUT pixel_4246/CSA_VREF pixel
Xpixel_4257 pixel_4257/gring pixel_4257/VDD pixel_4257/GND pixel_4257/VREF pixel_4257/ROW_SEL
+ pixel_4257/NB1 pixel_4257/VBIAS pixel_4257/NB2 pixel_4257/AMP_IN pixel_4257/SF_IB
+ pixel_4257/PIX_OUT pixel_4257/CSA_VREF pixel
Xpixel_4268 pixel_4268/gring pixel_4268/VDD pixel_4268/GND pixel_4268/VREF pixel_4268/ROW_SEL
+ pixel_4268/NB1 pixel_4268/VBIAS pixel_4268/NB2 pixel_4268/AMP_IN pixel_4268/SF_IB
+ pixel_4268/PIX_OUT pixel_4268/CSA_VREF pixel
Xpixel_296 pixel_296/gring pixel_296/VDD pixel_296/GND pixel_296/VREF pixel_296/ROW_SEL
+ pixel_296/NB1 pixel_296/VBIAS pixel_296/NB2 pixel_296/AMP_IN pixel_296/SF_IB pixel_296/PIX_OUT
+ pixel_296/CSA_VREF pixel
Xpixel_285 pixel_285/gring pixel_285/VDD pixel_285/GND pixel_285/VREF pixel_285/ROW_SEL
+ pixel_285/NB1 pixel_285/VBIAS pixel_285/NB2 pixel_285/AMP_IN pixel_285/SF_IB pixel_285/PIX_OUT
+ pixel_285/CSA_VREF pixel
Xpixel_2822 pixel_2822/gring pixel_2822/VDD pixel_2822/GND pixel_2822/VREF pixel_2822/ROW_SEL
+ pixel_2822/NB1 pixel_2822/VBIAS pixel_2822/NB2 pixel_2822/AMP_IN pixel_2822/SF_IB
+ pixel_2822/PIX_OUT pixel_2822/CSA_VREF pixel
Xpixel_2811 pixel_2811/gring pixel_2811/VDD pixel_2811/GND pixel_2811/VREF pixel_2811/ROW_SEL
+ pixel_2811/NB1 pixel_2811/VBIAS pixel_2811/NB2 pixel_2811/AMP_IN pixel_2811/SF_IB
+ pixel_2811/PIX_OUT pixel_2811/CSA_VREF pixel
Xpixel_2800 pixel_2800/gring pixel_2800/VDD pixel_2800/GND pixel_2800/VREF pixel_2800/ROW_SEL
+ pixel_2800/NB1 pixel_2800/VBIAS pixel_2800/NB2 pixel_2800/AMP_IN pixel_2800/SF_IB
+ pixel_2800/PIX_OUT pixel_2800/CSA_VREF pixel
Xpixel_3567 pixel_3567/gring pixel_3567/VDD pixel_3567/GND pixel_3567/VREF pixel_3567/ROW_SEL
+ pixel_3567/NB1 pixel_3567/VBIAS pixel_3567/NB2 pixel_3567/AMP_IN pixel_3567/SF_IB
+ pixel_3567/PIX_OUT pixel_3567/CSA_VREF pixel
Xpixel_3556 pixel_3556/gring pixel_3556/VDD pixel_3556/GND pixel_3556/VREF pixel_3556/ROW_SEL
+ pixel_3556/NB1 pixel_3556/VBIAS pixel_3556/NB2 pixel_3556/AMP_IN pixel_3556/SF_IB
+ pixel_3556/PIX_OUT pixel_3556/CSA_VREF pixel
Xpixel_3545 pixel_3545/gring pixel_3545/VDD pixel_3545/GND pixel_3545/VREF pixel_3545/ROW_SEL
+ pixel_3545/NB1 pixel_3545/VBIAS pixel_3545/NB2 pixel_3545/AMP_IN pixel_3545/SF_IB
+ pixel_3545/PIX_OUT pixel_3545/CSA_VREF pixel
Xpixel_4279 pixel_4279/gring pixel_4279/VDD pixel_4279/GND pixel_4279/VREF pixel_4279/ROW_SEL
+ pixel_4279/NB1 pixel_4279/VBIAS pixel_4279/NB2 pixel_4279/AMP_IN pixel_4279/SF_IB
+ pixel_4279/PIX_OUT pixel_4279/CSA_VREF pixel
Xpixel_2855 pixel_2855/gring pixel_2855/VDD pixel_2855/GND pixel_2855/VREF pixel_2855/ROW_SEL
+ pixel_2855/NB1 pixel_2855/VBIAS pixel_2855/NB2 pixel_2855/AMP_IN pixel_2855/SF_IB
+ pixel_2855/PIX_OUT pixel_2855/CSA_VREF pixel
Xpixel_2844 pixel_2844/gring pixel_2844/VDD pixel_2844/GND pixel_2844/VREF pixel_2844/ROW_SEL
+ pixel_2844/NB1 pixel_2844/VBIAS pixel_2844/NB2 pixel_2844/AMP_IN pixel_2844/SF_IB
+ pixel_2844/PIX_OUT pixel_2844/CSA_VREF pixel
Xpixel_2833 pixel_2833/gring pixel_2833/VDD pixel_2833/GND pixel_2833/VREF pixel_2833/ROW_SEL
+ pixel_2833/NB1 pixel_2833/VBIAS pixel_2833/NB2 pixel_2833/AMP_IN pixel_2833/SF_IB
+ pixel_2833/PIX_OUT pixel_2833/CSA_VREF pixel
Xpixel_3589 pixel_3589/gring pixel_3589/VDD pixel_3589/GND pixel_3589/VREF pixel_3589/ROW_SEL
+ pixel_3589/NB1 pixel_3589/VBIAS pixel_3589/NB2 pixel_3589/AMP_IN pixel_3589/SF_IB
+ pixel_3589/PIX_OUT pixel_3589/CSA_VREF pixel
Xpixel_3578 pixel_3578/gring pixel_3578/VDD pixel_3578/GND pixel_3578/VREF pixel_3578/ROW_SEL
+ pixel_3578/NB1 pixel_3578/VBIAS pixel_3578/NB2 pixel_3578/AMP_IN pixel_3578/SF_IB
+ pixel_3578/PIX_OUT pixel_3578/CSA_VREF pixel
Xpixel_2899 pixel_2899/gring pixel_2899/VDD pixel_2899/GND pixel_2899/VREF pixel_2899/ROW_SEL
+ pixel_2899/NB1 pixel_2899/VBIAS pixel_2899/NB2 pixel_2899/AMP_IN pixel_2899/SF_IB
+ pixel_2899/PIX_OUT pixel_2899/CSA_VREF pixel
Xpixel_2888 pixel_2888/gring pixel_2888/VDD pixel_2888/GND pixel_2888/VREF pixel_2888/ROW_SEL
+ pixel_2888/NB1 pixel_2888/VBIAS pixel_2888/NB2 pixel_2888/AMP_IN pixel_2888/SF_IB
+ pixel_2888/PIX_OUT pixel_2888/CSA_VREF pixel
Xpixel_2877 pixel_2877/gring pixel_2877/VDD pixel_2877/GND pixel_2877/VREF pixel_2877/ROW_SEL
+ pixel_2877/NB1 pixel_2877/VBIAS pixel_2877/NB2 pixel_2877/AMP_IN pixel_2877/SF_IB
+ pixel_2877/PIX_OUT pixel_2877/CSA_VREF pixel
Xpixel_2866 pixel_2866/gring pixel_2866/VDD pixel_2866/GND pixel_2866/VREF pixel_2866/ROW_SEL
+ pixel_2866/NB1 pixel_2866/VBIAS pixel_2866/NB2 pixel_2866/AMP_IN pixel_2866/SF_IB
+ pixel_2866/PIX_OUT pixel_2866/CSA_VREF pixel
Xpixel_6160 pixel_6160/gring pixel_6160/VDD pixel_6160/GND pixel_6160/VREF pixel_6160/ROW_SEL
+ pixel_6160/NB1 pixel_6160/VBIAS pixel_6160/NB2 pixel_6160/AMP_IN pixel_6160/SF_IB
+ pixel_6160/PIX_OUT pixel_6160/CSA_VREF pixel
Xpixel_6171 pixel_6171/gring pixel_6171/VDD pixel_6171/GND pixel_6171/VREF pixel_6171/ROW_SEL
+ pixel_6171/NB1 pixel_6171/VBIAS pixel_6171/NB2 pixel_6171/AMP_IN pixel_6171/SF_IB
+ pixel_6171/PIX_OUT pixel_6171/CSA_VREF pixel
Xpixel_6182 pixel_6182/gring pixel_6182/VDD pixel_6182/GND pixel_6182/VREF pixel_6182/ROW_SEL
+ pixel_6182/NB1 pixel_6182/VBIAS pixel_6182/NB2 pixel_6182/AMP_IN pixel_6182/SF_IB
+ pixel_6182/PIX_OUT pixel_6182/CSA_VREF pixel
Xpixel_6193 pixel_6193/gring pixel_6193/VDD pixel_6193/GND pixel_6193/VREF pixel_6193/ROW_SEL
+ pixel_6193/NB1 pixel_6193/VBIAS pixel_6193/NB2 pixel_6193/AMP_IN pixel_6193/SF_IB
+ pixel_6193/PIX_OUT pixel_6193/CSA_VREF pixel
Xpixel_5470 pixel_5470/gring pixel_5470/VDD pixel_5470/GND pixel_5470/VREF pixel_5470/ROW_SEL
+ pixel_5470/NB1 pixel_5470/VBIAS pixel_5470/NB2 pixel_5470/AMP_IN pixel_5470/SF_IB
+ pixel_5470/PIX_OUT pixel_5470/CSA_VREF pixel
Xpixel_5481 pixel_5481/gring pixel_5481/VDD pixel_5481/GND pixel_5481/VREF pixel_5481/ROW_SEL
+ pixel_5481/NB1 pixel_5481/VBIAS pixel_5481/NB2 pixel_5481/AMP_IN pixel_5481/SF_IB
+ pixel_5481/PIX_OUT pixel_5481/CSA_VREF pixel
Xpixel_5492 pixel_5492/gring pixel_5492/VDD pixel_5492/GND pixel_5492/VREF pixel_5492/ROW_SEL
+ pixel_5492/NB1 pixel_5492/VBIAS pixel_5492/NB2 pixel_5492/AMP_IN pixel_5492/SF_IB
+ pixel_5492/PIX_OUT pixel_5492/CSA_VREF pixel
Xpixel_4780 pixel_4780/gring pixel_4780/VDD pixel_4780/GND pixel_4780/VREF pixel_4780/ROW_SEL
+ pixel_4780/NB1 pixel_4780/VBIAS pixel_4780/NB2 pixel_4780/AMP_IN pixel_4780/SF_IB
+ pixel_4780/PIX_OUT pixel_4780/CSA_VREF pixel
Xpixel_4791 pixel_4791/gring pixel_4791/VDD pixel_4791/GND pixel_4791/VREF pixel_4791/ROW_SEL
+ pixel_4791/NB1 pixel_4791/VBIAS pixel_4791/NB2 pixel_4791/AMP_IN pixel_4791/SF_IB
+ pixel_4791/PIX_OUT pixel_4791/CSA_VREF pixel
Xpixel_2118 pixel_2118/gring pixel_2118/VDD pixel_2118/GND pixel_2118/VREF pixel_2118/ROW_SEL
+ pixel_2118/NB1 pixel_2118/VBIAS pixel_2118/NB2 pixel_2118/AMP_IN pixel_2118/SF_IB
+ pixel_2118/PIX_OUT pixel_2118/CSA_VREF pixel
Xpixel_2107 pixel_2107/gring pixel_2107/VDD pixel_2107/GND pixel_2107/VREF pixel_2107/ROW_SEL
+ pixel_2107/NB1 pixel_2107/VBIAS pixel_2107/NB2 pixel_2107/AMP_IN pixel_2107/SF_IB
+ pixel_2107/PIX_OUT pixel_2107/CSA_VREF pixel
Xpixel_1406 pixel_1406/gring pixel_1406/VDD pixel_1406/GND pixel_1406/VREF pixel_1406/ROW_SEL
+ pixel_1406/NB1 pixel_1406/VBIAS pixel_1406/NB2 pixel_1406/AMP_IN pixel_1406/SF_IB
+ pixel_1406/PIX_OUT pixel_1406/CSA_VREF pixel
Xpixel_2129 pixel_2129/gring pixel_2129/VDD pixel_2129/GND pixel_2129/VREF pixel_2129/ROW_SEL
+ pixel_2129/NB1 pixel_2129/VBIAS pixel_2129/NB2 pixel_2129/AMP_IN pixel_2129/SF_IB
+ pixel_2129/PIX_OUT pixel_2129/CSA_VREF pixel
Xpixel_1439 pixel_1439/gring pixel_1439/VDD pixel_1439/GND pixel_1439/VREF pixel_1439/ROW_SEL
+ pixel_1439/NB1 pixel_1439/VBIAS pixel_1439/NB2 pixel_1439/AMP_IN pixel_1439/SF_IB
+ pixel_1439/PIX_OUT pixel_1439/CSA_VREF pixel
Xpixel_1428 pixel_1428/gring pixel_1428/VDD pixel_1428/GND pixel_1428/VREF pixel_1428/ROW_SEL
+ pixel_1428/NB1 pixel_1428/VBIAS pixel_1428/NB2 pixel_1428/AMP_IN pixel_1428/SF_IB
+ pixel_1428/PIX_OUT pixel_1428/CSA_VREF pixel
Xpixel_1417 pixel_1417/gring pixel_1417/VDD pixel_1417/GND pixel_1417/VREF pixel_1417/ROW_SEL
+ pixel_1417/NB1 pixel_1417/VBIAS pixel_1417/NB2 pixel_1417/AMP_IN pixel_1417/SF_IB
+ pixel_1417/PIX_OUT pixel_1417/CSA_VREF pixel
Xpixel_9703 pixel_9703/gring pixel_9703/VDD pixel_9703/GND pixel_9703/VREF pixel_9703/ROW_SEL
+ pixel_9703/NB1 pixel_9703/VBIAS pixel_9703/NB2 pixel_9703/AMP_IN pixel_9703/SF_IB
+ pixel_9703/PIX_OUT pixel_9703/CSA_VREF pixel
Xpixel_9714 pixel_9714/gring pixel_9714/VDD pixel_9714/GND pixel_9714/VREF pixel_9714/ROW_SEL
+ pixel_9714/NB1 pixel_9714/VBIAS pixel_9714/NB2 pixel_9714/AMP_IN pixel_9714/SF_IB
+ pixel_9714/PIX_OUT pixel_9714/CSA_VREF pixel
Xpixel_9725 pixel_9725/gring pixel_9725/VDD pixel_9725/GND pixel_9725/VREF pixel_9725/ROW_SEL
+ pixel_9725/NB1 pixel_9725/VBIAS pixel_9725/NB2 pixel_9725/AMP_IN pixel_9725/SF_IB
+ pixel_9725/PIX_OUT pixel_9725/CSA_VREF pixel
Xpixel_9736 pixel_9736/gring pixel_9736/VDD pixel_9736/GND pixel_9736/VREF pixel_9736/ROW_SEL
+ pixel_9736/NB1 pixel_9736/VBIAS pixel_9736/NB2 pixel_9736/AMP_IN pixel_9736/SF_IB
+ pixel_9736/PIX_OUT pixel_9736/CSA_VREF pixel
Xpixel_9747 pixel_9747/gring pixel_9747/VDD pixel_9747/GND pixel_9747/VREF pixel_9747/ROW_SEL
+ pixel_9747/NB1 pixel_9747/VBIAS pixel_9747/NB2 pixel_9747/AMP_IN pixel_9747/SF_IB
+ pixel_9747/PIX_OUT pixel_9747/CSA_VREF pixel
Xpixel_9758 pixel_9758/gring pixel_9758/VDD pixel_9758/GND pixel_9758/VREF pixel_9758/ROW_SEL
+ pixel_9758/NB1 pixel_9758/VBIAS pixel_9758/NB2 pixel_9758/AMP_IN pixel_9758/SF_IB
+ pixel_9758/PIX_OUT pixel_9758/CSA_VREF pixel
Xpixel_9769 pixel_9769/gring pixel_9769/VDD pixel_9769/GND pixel_9769/VREF pixel_9769/ROW_SEL
+ pixel_9769/NB1 pixel_9769/VBIAS pixel_9769/NB2 pixel_9769/AMP_IN pixel_9769/SF_IB
+ pixel_9769/PIX_OUT pixel_9769/CSA_VREF pixel
Xpixel_4010 pixel_4010/gring pixel_4010/VDD pixel_4010/GND pixel_4010/VREF pixel_4010/ROW_SEL
+ pixel_4010/NB1 pixel_4010/VBIAS pixel_4010/NB2 pixel_4010/AMP_IN pixel_4010/SF_IB
+ pixel_4010/PIX_OUT pixel_4010/CSA_VREF pixel
Xpixel_4021 pixel_4021/gring pixel_4021/VDD pixel_4021/GND pixel_4021/VREF pixel_4021/ROW_SEL
+ pixel_4021/NB1 pixel_4021/VBIAS pixel_4021/NB2 pixel_4021/AMP_IN pixel_4021/SF_IB
+ pixel_4021/PIX_OUT pixel_4021/CSA_VREF pixel
Xpixel_4032 pixel_4032/gring pixel_4032/VDD pixel_4032/GND pixel_4032/VREF pixel_4032/ROW_SEL
+ pixel_4032/NB1 pixel_4032/VBIAS pixel_4032/NB2 pixel_4032/AMP_IN pixel_4032/SF_IB
+ pixel_4032/PIX_OUT pixel_4032/CSA_VREF pixel
Xpixel_4043 pixel_4043/gring pixel_4043/VDD pixel_4043/GND pixel_4043/VREF pixel_4043/ROW_SEL
+ pixel_4043/NB1 pixel_4043/VBIAS pixel_4043/NB2 pixel_4043/AMP_IN pixel_4043/SF_IB
+ pixel_4043/PIX_OUT pixel_4043/CSA_VREF pixel
Xpixel_3342 pixel_3342/gring pixel_3342/VDD pixel_3342/GND pixel_3342/VREF pixel_3342/ROW_SEL
+ pixel_3342/NB1 pixel_3342/VBIAS pixel_3342/NB2 pixel_3342/AMP_IN pixel_3342/SF_IB
+ pixel_3342/PIX_OUT pixel_3342/CSA_VREF pixel
Xpixel_3331 pixel_3331/gring pixel_3331/VDD pixel_3331/GND pixel_3331/VREF pixel_3331/ROW_SEL
+ pixel_3331/NB1 pixel_3331/VBIAS pixel_3331/NB2 pixel_3331/AMP_IN pixel_3331/SF_IB
+ pixel_3331/PIX_OUT pixel_3331/CSA_VREF pixel
Xpixel_3320 pixel_3320/gring pixel_3320/VDD pixel_3320/GND pixel_3320/VREF pixel_3320/ROW_SEL
+ pixel_3320/NB1 pixel_3320/VBIAS pixel_3320/NB2 pixel_3320/AMP_IN pixel_3320/SF_IB
+ pixel_3320/PIX_OUT pixel_3320/CSA_VREF pixel
Xpixel_4054 pixel_4054/gring pixel_4054/VDD pixel_4054/GND pixel_4054/VREF pixel_4054/ROW_SEL
+ pixel_4054/NB1 pixel_4054/VBIAS pixel_4054/NB2 pixel_4054/AMP_IN pixel_4054/SF_IB
+ pixel_4054/PIX_OUT pixel_4054/CSA_VREF pixel
Xpixel_4065 pixel_4065/gring pixel_4065/VDD pixel_4065/GND pixel_4065/VREF pixel_4065/ROW_SEL
+ pixel_4065/NB1 pixel_4065/VBIAS pixel_4065/NB2 pixel_4065/AMP_IN pixel_4065/SF_IB
+ pixel_4065/PIX_OUT pixel_4065/CSA_VREF pixel
Xpixel_4076 pixel_4076/gring pixel_4076/VDD pixel_4076/GND pixel_4076/VREF pixel_4076/ROW_SEL
+ pixel_4076/NB1 pixel_4076/VBIAS pixel_4076/NB2 pixel_4076/AMP_IN pixel_4076/SF_IB
+ pixel_4076/PIX_OUT pixel_4076/CSA_VREF pixel
Xpixel_4087 pixel_4087/gring pixel_4087/VDD pixel_4087/GND pixel_4087/VREF pixel_4087/ROW_SEL
+ pixel_4087/NB1 pixel_4087/VBIAS pixel_4087/NB2 pixel_4087/AMP_IN pixel_4087/SF_IB
+ pixel_4087/PIX_OUT pixel_4087/CSA_VREF pixel
Xpixel_2630 pixel_2630/gring pixel_2630/VDD pixel_2630/GND pixel_2630/VREF pixel_2630/ROW_SEL
+ pixel_2630/NB1 pixel_2630/VBIAS pixel_2630/NB2 pixel_2630/AMP_IN pixel_2630/SF_IB
+ pixel_2630/PIX_OUT pixel_2630/CSA_VREF pixel
Xpixel_3375 pixel_3375/gring pixel_3375/VDD pixel_3375/GND pixel_3375/VREF pixel_3375/ROW_SEL
+ pixel_3375/NB1 pixel_3375/VBIAS pixel_3375/NB2 pixel_3375/AMP_IN pixel_3375/SF_IB
+ pixel_3375/PIX_OUT pixel_3375/CSA_VREF pixel
Xpixel_3364 pixel_3364/gring pixel_3364/VDD pixel_3364/GND pixel_3364/VREF pixel_3364/ROW_SEL
+ pixel_3364/NB1 pixel_3364/VBIAS pixel_3364/NB2 pixel_3364/AMP_IN pixel_3364/SF_IB
+ pixel_3364/PIX_OUT pixel_3364/CSA_VREF pixel
Xpixel_3353 pixel_3353/gring pixel_3353/VDD pixel_3353/GND pixel_3353/VREF pixel_3353/ROW_SEL
+ pixel_3353/NB1 pixel_3353/VBIAS pixel_3353/NB2 pixel_3353/AMP_IN pixel_3353/SF_IB
+ pixel_3353/PIX_OUT pixel_3353/CSA_VREF pixel
Xpixel_4098 pixel_4098/gring pixel_4098/VDD pixel_4098/GND pixel_4098/VREF pixel_4098/ROW_SEL
+ pixel_4098/NB1 pixel_4098/VBIAS pixel_4098/NB2 pixel_4098/AMP_IN pixel_4098/SF_IB
+ pixel_4098/PIX_OUT pixel_4098/CSA_VREF pixel
Xpixel_2663 pixel_2663/gring pixel_2663/VDD pixel_2663/GND pixel_2663/VREF pixel_2663/ROW_SEL
+ pixel_2663/NB1 pixel_2663/VBIAS pixel_2663/NB2 pixel_2663/AMP_IN pixel_2663/SF_IB
+ pixel_2663/PIX_OUT pixel_2663/CSA_VREF pixel
Xpixel_2652 pixel_2652/gring pixel_2652/VDD pixel_2652/GND pixel_2652/VREF pixel_2652/ROW_SEL
+ pixel_2652/NB1 pixel_2652/VBIAS pixel_2652/NB2 pixel_2652/AMP_IN pixel_2652/SF_IB
+ pixel_2652/PIX_OUT pixel_2652/CSA_VREF pixel
Xpixel_2641 pixel_2641/gring pixel_2641/VDD pixel_2641/GND pixel_2641/VREF pixel_2641/ROW_SEL
+ pixel_2641/NB1 pixel_2641/VBIAS pixel_2641/NB2 pixel_2641/AMP_IN pixel_2641/SF_IB
+ pixel_2641/PIX_OUT pixel_2641/CSA_VREF pixel
Xpixel_3397 pixel_3397/gring pixel_3397/VDD pixel_3397/GND pixel_3397/VREF pixel_3397/ROW_SEL
+ pixel_3397/NB1 pixel_3397/VBIAS pixel_3397/NB2 pixel_3397/AMP_IN pixel_3397/SF_IB
+ pixel_3397/PIX_OUT pixel_3397/CSA_VREF pixel
Xpixel_3386 pixel_3386/gring pixel_3386/VDD pixel_3386/GND pixel_3386/VREF pixel_3386/ROW_SEL
+ pixel_3386/NB1 pixel_3386/VBIAS pixel_3386/NB2 pixel_3386/AMP_IN pixel_3386/SF_IB
+ pixel_3386/PIX_OUT pixel_3386/CSA_VREF pixel
Xpixel_1962 pixel_1962/gring pixel_1962/VDD pixel_1962/GND pixel_1962/VREF pixel_1962/ROW_SEL
+ pixel_1962/NB1 pixel_1962/VBIAS pixel_1962/NB2 pixel_1962/AMP_IN pixel_1962/SF_IB
+ pixel_1962/PIX_OUT pixel_1962/CSA_VREF pixel
Xpixel_1951 pixel_1951/gring pixel_1951/VDD pixel_1951/GND pixel_1951/VREF pixel_1951/ROW_SEL
+ pixel_1951/NB1 pixel_1951/VBIAS pixel_1951/NB2 pixel_1951/AMP_IN pixel_1951/SF_IB
+ pixel_1951/PIX_OUT pixel_1951/CSA_VREF pixel
Xpixel_1940 pixel_1940/gring pixel_1940/VDD pixel_1940/GND pixel_1940/VREF pixel_1940/ROW_SEL
+ pixel_1940/NB1 pixel_1940/VBIAS pixel_1940/NB2 pixel_1940/AMP_IN pixel_1940/SF_IB
+ pixel_1940/PIX_OUT pixel_1940/CSA_VREF pixel
Xpixel_2696 pixel_2696/gring pixel_2696/VDD pixel_2696/GND pixel_2696/VREF pixel_2696/ROW_SEL
+ pixel_2696/NB1 pixel_2696/VBIAS pixel_2696/NB2 pixel_2696/AMP_IN pixel_2696/SF_IB
+ pixel_2696/PIX_OUT pixel_2696/CSA_VREF pixel
Xpixel_2685 pixel_2685/gring pixel_2685/VDD pixel_2685/GND pixel_2685/VREF pixel_2685/ROW_SEL
+ pixel_2685/NB1 pixel_2685/VBIAS pixel_2685/NB2 pixel_2685/AMP_IN pixel_2685/SF_IB
+ pixel_2685/PIX_OUT pixel_2685/CSA_VREF pixel
Xpixel_2674 pixel_2674/gring pixel_2674/VDD pixel_2674/GND pixel_2674/VREF pixel_2674/ROW_SEL
+ pixel_2674/NB1 pixel_2674/VBIAS pixel_2674/NB2 pixel_2674/AMP_IN pixel_2674/SF_IB
+ pixel_2674/PIX_OUT pixel_2674/CSA_VREF pixel
Xpixel_1995 pixel_1995/gring pixel_1995/VDD pixel_1995/GND pixel_1995/VREF pixel_1995/ROW_SEL
+ pixel_1995/NB1 pixel_1995/VBIAS pixel_1995/NB2 pixel_1995/AMP_IN pixel_1995/SF_IB
+ pixel_1995/PIX_OUT pixel_1995/CSA_VREF pixel
Xpixel_1984 pixel_1984/gring pixel_1984/VDD pixel_1984/GND pixel_1984/VREF pixel_1984/ROW_SEL
+ pixel_1984/NB1 pixel_1984/VBIAS pixel_1984/NB2 pixel_1984/AMP_IN pixel_1984/SF_IB
+ pixel_1984/PIX_OUT pixel_1984/CSA_VREF pixel
Xpixel_1973 pixel_1973/gring pixel_1973/VDD pixel_1973/GND pixel_1973/VREF pixel_1973/ROW_SEL
+ pixel_1973/NB1 pixel_1973/VBIAS pixel_1973/NB2 pixel_1973/AMP_IN pixel_1973/SF_IB
+ pixel_1973/PIX_OUT pixel_1973/CSA_VREF pixel
Xpixel_8309 pixel_8309/gring pixel_8309/VDD pixel_8309/GND pixel_8309/VREF pixel_8309/ROW_SEL
+ pixel_8309/NB1 pixel_8309/VBIAS pixel_8309/NB2 pixel_8309/AMP_IN pixel_8309/SF_IB
+ pixel_8309/PIX_OUT pixel_8309/CSA_VREF pixel
Xpixel_7608 pixel_7608/gring pixel_7608/VDD pixel_7608/GND pixel_7608/VREF pixel_7608/ROW_SEL
+ pixel_7608/NB1 pixel_7608/VBIAS pixel_7608/NB2 pixel_7608/AMP_IN pixel_7608/SF_IB
+ pixel_7608/PIX_OUT pixel_7608/CSA_VREF pixel
Xpixel_7619 pixel_7619/gring pixel_7619/VDD pixel_7619/GND pixel_7619/VREF pixel_7619/ROW_SEL
+ pixel_7619/NB1 pixel_7619/VBIAS pixel_7619/NB2 pixel_7619/AMP_IN pixel_7619/SF_IB
+ pixel_7619/PIX_OUT pixel_7619/CSA_VREF pixel
Xpixel_6907 pixel_6907/gring pixel_6907/VDD pixel_6907/GND pixel_6907/VREF pixel_6907/ROW_SEL
+ pixel_6907/NB1 pixel_6907/VBIAS pixel_6907/NB2 pixel_6907/AMP_IN pixel_6907/SF_IB
+ pixel_6907/PIX_OUT pixel_6907/CSA_VREF pixel
Xpixel_6918 pixel_6918/gring pixel_6918/VDD pixel_6918/GND pixel_6918/VREF pixel_6918/ROW_SEL
+ pixel_6918/NB1 pixel_6918/VBIAS pixel_6918/NB2 pixel_6918/AMP_IN pixel_6918/SF_IB
+ pixel_6918/PIX_OUT pixel_6918/CSA_VREF pixel
Xpixel_6929 pixel_6929/gring pixel_6929/VDD pixel_6929/GND pixel_6929/VREF pixel_6929/ROW_SEL
+ pixel_6929/NB1 pixel_6929/VBIAS pixel_6929/NB2 pixel_6929/AMP_IN pixel_6929/SF_IB
+ pixel_6929/PIX_OUT pixel_6929/CSA_VREF pixel
Xpixel_1214 pixel_1214/gring pixel_1214/VDD pixel_1214/GND pixel_1214/VREF pixel_1214/ROW_SEL
+ pixel_1214/NB1 pixel_1214/VBIAS pixel_1214/NB2 pixel_1214/AMP_IN pixel_1214/SF_IB
+ pixel_1214/PIX_OUT pixel_1214/CSA_VREF pixel
Xpixel_1203 pixel_1203/gring pixel_1203/VDD pixel_1203/GND pixel_1203/VREF pixel_1203/ROW_SEL
+ pixel_1203/NB1 pixel_1203/VBIAS pixel_1203/NB2 pixel_1203/AMP_IN pixel_1203/SF_IB
+ pixel_1203/PIX_OUT pixel_1203/CSA_VREF pixel
Xpixel_1258 pixel_1258/gring pixel_1258/VDD pixel_1258/GND pixel_1258/VREF pixel_1258/ROW_SEL
+ pixel_1258/NB1 pixel_1258/VBIAS pixel_1258/NB2 pixel_1258/AMP_IN pixel_1258/SF_IB
+ pixel_1258/PIX_OUT pixel_1258/CSA_VREF pixel
Xpixel_1247 pixel_1247/gring pixel_1247/VDD pixel_1247/GND pixel_1247/VREF pixel_1247/ROW_SEL
+ pixel_1247/NB1 pixel_1247/VBIAS pixel_1247/NB2 pixel_1247/AMP_IN pixel_1247/SF_IB
+ pixel_1247/PIX_OUT pixel_1247/CSA_VREF pixel
Xpixel_1236 pixel_1236/gring pixel_1236/VDD pixel_1236/GND pixel_1236/VREF pixel_1236/ROW_SEL
+ pixel_1236/NB1 pixel_1236/VBIAS pixel_1236/NB2 pixel_1236/AMP_IN pixel_1236/SF_IB
+ pixel_1236/PIX_OUT pixel_1236/CSA_VREF pixel
Xpixel_1225 pixel_1225/gring pixel_1225/VDD pixel_1225/GND pixel_1225/VREF pixel_1225/ROW_SEL
+ pixel_1225/NB1 pixel_1225/VBIAS pixel_1225/NB2 pixel_1225/AMP_IN pixel_1225/SF_IB
+ pixel_1225/PIX_OUT pixel_1225/CSA_VREF pixel
Xpixel_1269 pixel_1269/gring pixel_1269/VDD pixel_1269/GND pixel_1269/VREF pixel_1269/ROW_SEL
+ pixel_1269/NB1 pixel_1269/VBIAS pixel_1269/NB2 pixel_1269/AMP_IN pixel_1269/SF_IB
+ pixel_1269/PIX_OUT pixel_1269/CSA_VREF pixel
Xpixel_9522 pixel_9522/gring pixel_9522/VDD pixel_9522/GND pixel_9522/VREF pixel_9522/ROW_SEL
+ pixel_9522/NB1 pixel_9522/VBIAS pixel_9522/NB2 pixel_9522/AMP_IN pixel_9522/SF_IB
+ pixel_9522/PIX_OUT pixel_9522/CSA_VREF pixel
Xpixel_9511 pixel_9511/gring pixel_9511/VDD pixel_9511/GND pixel_9511/VREF pixel_9511/ROW_SEL
+ pixel_9511/NB1 pixel_9511/VBIAS pixel_9511/NB2 pixel_9511/AMP_IN pixel_9511/SF_IB
+ pixel_9511/PIX_OUT pixel_9511/CSA_VREF pixel
Xpixel_9500 pixel_9500/gring pixel_9500/VDD pixel_9500/GND pixel_9500/VREF pixel_9500/ROW_SEL
+ pixel_9500/NB1 pixel_9500/VBIAS pixel_9500/NB2 pixel_9500/AMP_IN pixel_9500/SF_IB
+ pixel_9500/PIX_OUT pixel_9500/CSA_VREF pixel
Xpixel_8821 pixel_8821/gring pixel_8821/VDD pixel_8821/GND pixel_8821/VREF pixel_8821/ROW_SEL
+ pixel_8821/NB1 pixel_8821/VBIAS pixel_8821/NB2 pixel_8821/AMP_IN pixel_8821/SF_IB
+ pixel_8821/PIX_OUT pixel_8821/CSA_VREF pixel
Xpixel_8810 pixel_8810/gring pixel_8810/VDD pixel_8810/GND pixel_8810/VREF pixel_8810/ROW_SEL
+ pixel_8810/NB1 pixel_8810/VBIAS pixel_8810/NB2 pixel_8810/AMP_IN pixel_8810/SF_IB
+ pixel_8810/PIX_OUT pixel_8810/CSA_VREF pixel
Xpixel_9566 pixel_9566/gring pixel_9566/VDD pixel_9566/GND pixel_9566/VREF pixel_9566/ROW_SEL
+ pixel_9566/NB1 pixel_9566/VBIAS pixel_9566/NB2 pixel_9566/AMP_IN pixel_9566/SF_IB
+ pixel_9566/PIX_OUT pixel_9566/CSA_VREF pixel
Xpixel_9555 pixel_9555/gring pixel_9555/VDD pixel_9555/GND pixel_9555/VREF pixel_9555/ROW_SEL
+ pixel_9555/NB1 pixel_9555/VBIAS pixel_9555/NB2 pixel_9555/AMP_IN pixel_9555/SF_IB
+ pixel_9555/PIX_OUT pixel_9555/CSA_VREF pixel
Xpixel_9544 pixel_9544/gring pixel_9544/VDD pixel_9544/GND pixel_9544/VREF pixel_9544/ROW_SEL
+ pixel_9544/NB1 pixel_9544/VBIAS pixel_9544/NB2 pixel_9544/AMP_IN pixel_9544/SF_IB
+ pixel_9544/PIX_OUT pixel_9544/CSA_VREF pixel
Xpixel_9533 pixel_9533/gring pixel_9533/VDD pixel_9533/GND pixel_9533/VREF pixel_9533/ROW_SEL
+ pixel_9533/NB1 pixel_9533/VBIAS pixel_9533/NB2 pixel_9533/AMP_IN pixel_9533/SF_IB
+ pixel_9533/PIX_OUT pixel_9533/CSA_VREF pixel
Xpixel_8854 pixel_8854/gring pixel_8854/VDD pixel_8854/GND pixel_8854/VREF pixel_8854/ROW_SEL
+ pixel_8854/NB1 pixel_8854/VBIAS pixel_8854/NB2 pixel_8854/AMP_IN pixel_8854/SF_IB
+ pixel_8854/PIX_OUT pixel_8854/CSA_VREF pixel
Xpixel_8843 pixel_8843/gring pixel_8843/VDD pixel_8843/GND pixel_8843/VREF pixel_8843/ROW_SEL
+ pixel_8843/NB1 pixel_8843/VBIAS pixel_8843/NB2 pixel_8843/AMP_IN pixel_8843/SF_IB
+ pixel_8843/PIX_OUT pixel_8843/CSA_VREF pixel
Xpixel_8832 pixel_8832/gring pixel_8832/VDD pixel_8832/GND pixel_8832/VREF pixel_8832/ROW_SEL
+ pixel_8832/NB1 pixel_8832/VBIAS pixel_8832/NB2 pixel_8832/AMP_IN pixel_8832/SF_IB
+ pixel_8832/PIX_OUT pixel_8832/CSA_VREF pixel
Xpixel_9599 pixel_9599/gring pixel_9599/VDD pixel_9599/GND pixel_9599/VREF pixel_9599/ROW_SEL
+ pixel_9599/NB1 pixel_9599/VBIAS pixel_9599/NB2 pixel_9599/AMP_IN pixel_9599/SF_IB
+ pixel_9599/PIX_OUT pixel_9599/CSA_VREF pixel
Xpixel_9588 pixel_9588/gring pixel_9588/VDD pixel_9588/GND pixel_9588/VREF pixel_9588/ROW_SEL
+ pixel_9588/NB1 pixel_9588/VBIAS pixel_9588/NB2 pixel_9588/AMP_IN pixel_9588/SF_IB
+ pixel_9588/PIX_OUT pixel_9588/CSA_VREF pixel
Xpixel_9577 pixel_9577/gring pixel_9577/VDD pixel_9577/GND pixel_9577/VREF pixel_9577/ROW_SEL
+ pixel_9577/NB1 pixel_9577/VBIAS pixel_9577/NB2 pixel_9577/AMP_IN pixel_9577/SF_IB
+ pixel_9577/PIX_OUT pixel_9577/CSA_VREF pixel
Xpixel_8887 pixel_8887/gring pixel_8887/VDD pixel_8887/GND pixel_8887/VREF pixel_8887/ROW_SEL
+ pixel_8887/NB1 pixel_8887/VBIAS pixel_8887/NB2 pixel_8887/AMP_IN pixel_8887/SF_IB
+ pixel_8887/PIX_OUT pixel_8887/CSA_VREF pixel
Xpixel_8876 pixel_8876/gring pixel_8876/VDD pixel_8876/GND pixel_8876/VREF pixel_8876/ROW_SEL
+ pixel_8876/NB1 pixel_8876/VBIAS pixel_8876/NB2 pixel_8876/AMP_IN pixel_8876/SF_IB
+ pixel_8876/PIX_OUT pixel_8876/CSA_VREF pixel
Xpixel_8865 pixel_8865/gring pixel_8865/VDD pixel_8865/GND pixel_8865/VREF pixel_8865/ROW_SEL
+ pixel_8865/NB1 pixel_8865/VBIAS pixel_8865/NB2 pixel_8865/AMP_IN pixel_8865/SF_IB
+ pixel_8865/PIX_OUT pixel_8865/CSA_VREF pixel
Xpixel_8898 pixel_8898/gring pixel_8898/VDD pixel_8898/GND pixel_8898/VREF pixel_8898/ROW_SEL
+ pixel_8898/NB1 pixel_8898/VBIAS pixel_8898/NB2 pixel_8898/AMP_IN pixel_8898/SF_IB
+ pixel_8898/PIX_OUT pixel_8898/CSA_VREF pixel
Xpixel_3150 pixel_3150/gring pixel_3150/VDD pixel_3150/GND pixel_3150/VREF pixel_3150/ROW_SEL
+ pixel_3150/NB1 pixel_3150/VBIAS pixel_3150/NB2 pixel_3150/AMP_IN pixel_3150/SF_IB
+ pixel_3150/PIX_OUT pixel_3150/CSA_VREF pixel
Xpixel_3183 pixel_3183/gring pixel_3183/VDD pixel_3183/GND pixel_3183/VREF pixel_3183/ROW_SEL
+ pixel_3183/NB1 pixel_3183/VBIAS pixel_3183/NB2 pixel_3183/AMP_IN pixel_3183/SF_IB
+ pixel_3183/PIX_OUT pixel_3183/CSA_VREF pixel
Xpixel_3172 pixel_3172/gring pixel_3172/VDD pixel_3172/GND pixel_3172/VREF pixel_3172/ROW_SEL
+ pixel_3172/NB1 pixel_3172/VBIAS pixel_3172/NB2 pixel_3172/AMP_IN pixel_3172/SF_IB
+ pixel_3172/PIX_OUT pixel_3172/CSA_VREF pixel
Xpixel_3161 pixel_3161/gring pixel_3161/VDD pixel_3161/GND pixel_3161/VREF pixel_3161/ROW_SEL
+ pixel_3161/NB1 pixel_3161/VBIAS pixel_3161/NB2 pixel_3161/AMP_IN pixel_3161/SF_IB
+ pixel_3161/PIX_OUT pixel_3161/CSA_VREF pixel
Xpixel_2482 pixel_2482/gring pixel_2482/VDD pixel_2482/GND pixel_2482/VREF pixel_2482/ROW_SEL
+ pixel_2482/NB1 pixel_2482/VBIAS pixel_2482/NB2 pixel_2482/AMP_IN pixel_2482/SF_IB
+ pixel_2482/PIX_OUT pixel_2482/CSA_VREF pixel
Xpixel_2471 pixel_2471/gring pixel_2471/VDD pixel_2471/GND pixel_2471/VREF pixel_2471/ROW_SEL
+ pixel_2471/NB1 pixel_2471/VBIAS pixel_2471/NB2 pixel_2471/AMP_IN pixel_2471/SF_IB
+ pixel_2471/PIX_OUT pixel_2471/CSA_VREF pixel
Xpixel_2460 pixel_2460/gring pixel_2460/VDD pixel_2460/GND pixel_2460/VREF pixel_2460/ROW_SEL
+ pixel_2460/NB1 pixel_2460/VBIAS pixel_2460/NB2 pixel_2460/AMP_IN pixel_2460/SF_IB
+ pixel_2460/PIX_OUT pixel_2460/CSA_VREF pixel
Xpixel_3194 pixel_3194/gring pixel_3194/VDD pixel_3194/GND pixel_3194/VREF pixel_3194/ROW_SEL
+ pixel_3194/NB1 pixel_3194/VBIAS pixel_3194/NB2 pixel_3194/AMP_IN pixel_3194/SF_IB
+ pixel_3194/PIX_OUT pixel_3194/CSA_VREF pixel
Xpixel_1770 pixel_1770/gring pixel_1770/VDD pixel_1770/GND pixel_1770/VREF pixel_1770/ROW_SEL
+ pixel_1770/NB1 pixel_1770/VBIAS pixel_1770/NB2 pixel_1770/AMP_IN pixel_1770/SF_IB
+ pixel_1770/PIX_OUT pixel_1770/CSA_VREF pixel
Xpixel_2493 pixel_2493/gring pixel_2493/VDD pixel_2493/GND pixel_2493/VREF pixel_2493/ROW_SEL
+ pixel_2493/NB1 pixel_2493/VBIAS pixel_2493/NB2 pixel_2493/AMP_IN pixel_2493/SF_IB
+ pixel_2493/PIX_OUT pixel_2493/CSA_VREF pixel
Xpixel_1792 pixel_1792/gring pixel_1792/VDD pixel_1792/GND pixel_1792/VREF pixel_1792/ROW_SEL
+ pixel_1792/NB1 pixel_1792/VBIAS pixel_1792/NB2 pixel_1792/AMP_IN pixel_1792/SF_IB
+ pixel_1792/PIX_OUT pixel_1792/CSA_VREF pixel
Xpixel_1781 pixel_1781/gring pixel_1781/VDD pixel_1781/GND pixel_1781/VREF pixel_1781/ROW_SEL
+ pixel_1781/NB1 pixel_1781/VBIAS pixel_1781/NB2 pixel_1781/AMP_IN pixel_1781/SF_IB
+ pixel_1781/PIX_OUT pixel_1781/CSA_VREF pixel
Xpixel_829 pixel_829/gring pixel_829/VDD pixel_829/GND pixel_829/VREF pixel_829/ROW_SEL
+ pixel_829/NB1 pixel_829/VBIAS pixel_829/NB2 pixel_829/AMP_IN pixel_829/SF_IB pixel_829/PIX_OUT
+ pixel_829/CSA_VREF pixel
Xpixel_818 pixel_818/gring pixel_818/VDD pixel_818/GND pixel_818/VREF pixel_818/ROW_SEL
+ pixel_818/NB1 pixel_818/VBIAS pixel_818/NB2 pixel_818/AMP_IN pixel_818/SF_IB pixel_818/PIX_OUT
+ pixel_818/CSA_VREF pixel
Xpixel_807 pixel_807/gring pixel_807/VDD pixel_807/GND pixel_807/VREF pixel_807/ROW_SEL
+ pixel_807/NB1 pixel_807/VBIAS pixel_807/NB2 pixel_807/AMP_IN pixel_807/SF_IB pixel_807/PIX_OUT
+ pixel_807/CSA_VREF pixel
Xpixel_8106 pixel_8106/gring pixel_8106/VDD pixel_8106/GND pixel_8106/VREF pixel_8106/ROW_SEL
+ pixel_8106/NB1 pixel_8106/VBIAS pixel_8106/NB2 pixel_8106/AMP_IN pixel_8106/SF_IB
+ pixel_8106/PIX_OUT pixel_8106/CSA_VREF pixel
Xpixel_8117 pixel_8117/gring pixel_8117/VDD pixel_8117/GND pixel_8117/VREF pixel_8117/ROW_SEL
+ pixel_8117/NB1 pixel_8117/VBIAS pixel_8117/NB2 pixel_8117/AMP_IN pixel_8117/SF_IB
+ pixel_8117/PIX_OUT pixel_8117/CSA_VREF pixel
Xpixel_8128 pixel_8128/gring pixel_8128/VDD pixel_8128/GND pixel_8128/VREF pixel_8128/ROW_SEL
+ pixel_8128/NB1 pixel_8128/VBIAS pixel_8128/NB2 pixel_8128/AMP_IN pixel_8128/SF_IB
+ pixel_8128/PIX_OUT pixel_8128/CSA_VREF pixel
Xpixel_8139 pixel_8139/gring pixel_8139/VDD pixel_8139/GND pixel_8139/VREF pixel_8139/ROW_SEL
+ pixel_8139/NB1 pixel_8139/VBIAS pixel_8139/NB2 pixel_8139/AMP_IN pixel_8139/SF_IB
+ pixel_8139/PIX_OUT pixel_8139/CSA_VREF pixel
Xpixel_7405 pixel_7405/gring pixel_7405/VDD pixel_7405/GND pixel_7405/VREF pixel_7405/ROW_SEL
+ pixel_7405/NB1 pixel_7405/VBIAS pixel_7405/NB2 pixel_7405/AMP_IN pixel_7405/SF_IB
+ pixel_7405/PIX_OUT pixel_7405/CSA_VREF pixel
Xpixel_7416 pixel_7416/gring pixel_7416/VDD pixel_7416/GND pixel_7416/VREF pixel_7416/ROW_SEL
+ pixel_7416/NB1 pixel_7416/VBIAS pixel_7416/NB2 pixel_7416/AMP_IN pixel_7416/SF_IB
+ pixel_7416/PIX_OUT pixel_7416/CSA_VREF pixel
Xpixel_7427 pixel_7427/gring pixel_7427/VDD pixel_7427/GND pixel_7427/VREF pixel_7427/ROW_SEL
+ pixel_7427/NB1 pixel_7427/VBIAS pixel_7427/NB2 pixel_7427/AMP_IN pixel_7427/SF_IB
+ pixel_7427/PIX_OUT pixel_7427/CSA_VREF pixel
Xpixel_7438 pixel_7438/gring pixel_7438/VDD pixel_7438/GND pixel_7438/VREF pixel_7438/ROW_SEL
+ pixel_7438/NB1 pixel_7438/VBIAS pixel_7438/NB2 pixel_7438/AMP_IN pixel_7438/SF_IB
+ pixel_7438/PIX_OUT pixel_7438/CSA_VREF pixel
Xpixel_7449 pixel_7449/gring pixel_7449/VDD pixel_7449/GND pixel_7449/VREF pixel_7449/ROW_SEL
+ pixel_7449/NB1 pixel_7449/VBIAS pixel_7449/NB2 pixel_7449/AMP_IN pixel_7449/SF_IB
+ pixel_7449/PIX_OUT pixel_7449/CSA_VREF pixel
Xpixel_6704 pixel_6704/gring pixel_6704/VDD pixel_6704/GND pixel_6704/VREF pixel_6704/ROW_SEL
+ pixel_6704/NB1 pixel_6704/VBIAS pixel_6704/NB2 pixel_6704/AMP_IN pixel_6704/SF_IB
+ pixel_6704/PIX_OUT pixel_6704/CSA_VREF pixel
Xpixel_6715 pixel_6715/gring pixel_6715/VDD pixel_6715/GND pixel_6715/VREF pixel_6715/ROW_SEL
+ pixel_6715/NB1 pixel_6715/VBIAS pixel_6715/NB2 pixel_6715/AMP_IN pixel_6715/SF_IB
+ pixel_6715/PIX_OUT pixel_6715/CSA_VREF pixel
Xpixel_6726 pixel_6726/gring pixel_6726/VDD pixel_6726/GND pixel_6726/VREF pixel_6726/ROW_SEL
+ pixel_6726/NB1 pixel_6726/VBIAS pixel_6726/NB2 pixel_6726/AMP_IN pixel_6726/SF_IB
+ pixel_6726/PIX_OUT pixel_6726/CSA_VREF pixel
Xpixel_6737 pixel_6737/gring pixel_6737/VDD pixel_6737/GND pixel_6737/VREF pixel_6737/ROW_SEL
+ pixel_6737/NB1 pixel_6737/VBIAS pixel_6737/NB2 pixel_6737/AMP_IN pixel_6737/SF_IB
+ pixel_6737/PIX_OUT pixel_6737/CSA_VREF pixel
Xpixel_6748 pixel_6748/gring pixel_6748/VDD pixel_6748/GND pixel_6748/VREF pixel_6748/ROW_SEL
+ pixel_6748/NB1 pixel_6748/VBIAS pixel_6748/NB2 pixel_6748/AMP_IN pixel_6748/SF_IB
+ pixel_6748/PIX_OUT pixel_6748/CSA_VREF pixel
Xpixel_6759 pixel_6759/gring pixel_6759/VDD pixel_6759/GND pixel_6759/VREF pixel_6759/ROW_SEL
+ pixel_6759/NB1 pixel_6759/VBIAS pixel_6759/NB2 pixel_6759/AMP_IN pixel_6759/SF_IB
+ pixel_6759/PIX_OUT pixel_6759/CSA_VREF pixel
Xpixel_1033 pixel_1033/gring pixel_1033/VDD pixel_1033/GND pixel_1033/VREF pixel_1033/ROW_SEL
+ pixel_1033/NB1 pixel_1033/VBIAS pixel_1033/NB2 pixel_1033/AMP_IN pixel_1033/SF_IB
+ pixel_1033/PIX_OUT pixel_1033/CSA_VREF pixel
Xpixel_1022 pixel_1022/gring pixel_1022/VDD pixel_1022/GND pixel_1022/VREF pixel_1022/ROW_SEL
+ pixel_1022/NB1 pixel_1022/VBIAS pixel_1022/NB2 pixel_1022/AMP_IN pixel_1022/SF_IB
+ pixel_1022/PIX_OUT pixel_1022/CSA_VREF pixel
Xpixel_1011 pixel_1011/gring pixel_1011/VDD pixel_1011/GND pixel_1011/VREF pixel_1011/ROW_SEL
+ pixel_1011/NB1 pixel_1011/VBIAS pixel_1011/NB2 pixel_1011/AMP_IN pixel_1011/SF_IB
+ pixel_1011/PIX_OUT pixel_1011/CSA_VREF pixel
Xpixel_1000 pixel_1000/gring pixel_1000/VDD pixel_1000/GND pixel_1000/VREF pixel_1000/ROW_SEL
+ pixel_1000/NB1 pixel_1000/VBIAS pixel_1000/NB2 pixel_1000/AMP_IN pixel_1000/SF_IB
+ pixel_1000/PIX_OUT pixel_1000/CSA_VREF pixel
Xpixel_1066 pixel_1066/gring pixel_1066/VDD pixel_1066/GND pixel_1066/VREF pixel_1066/ROW_SEL
+ pixel_1066/NB1 pixel_1066/VBIAS pixel_1066/NB2 pixel_1066/AMP_IN pixel_1066/SF_IB
+ pixel_1066/PIX_OUT pixel_1066/CSA_VREF pixel
Xpixel_1055 pixel_1055/gring pixel_1055/VDD pixel_1055/GND pixel_1055/VREF pixel_1055/ROW_SEL
+ pixel_1055/NB1 pixel_1055/VBIAS pixel_1055/NB2 pixel_1055/AMP_IN pixel_1055/SF_IB
+ pixel_1055/PIX_OUT pixel_1055/CSA_VREF pixel
Xpixel_1044 pixel_1044/gring pixel_1044/VDD pixel_1044/GND pixel_1044/VREF pixel_1044/ROW_SEL
+ pixel_1044/NB1 pixel_1044/VBIAS pixel_1044/NB2 pixel_1044/AMP_IN pixel_1044/SF_IB
+ pixel_1044/PIX_OUT pixel_1044/CSA_VREF pixel
Xpixel_1099 pixel_1099/gring pixel_1099/VDD pixel_1099/GND pixel_1099/VREF pixel_1099/ROW_SEL
+ pixel_1099/NB1 pixel_1099/VBIAS pixel_1099/NB2 pixel_1099/AMP_IN pixel_1099/SF_IB
+ pixel_1099/PIX_OUT pixel_1099/CSA_VREF pixel
Xpixel_1088 pixel_1088/gring pixel_1088/VDD pixel_1088/GND pixel_1088/VREF pixel_1088/ROW_SEL
+ pixel_1088/NB1 pixel_1088/VBIAS pixel_1088/NB2 pixel_1088/AMP_IN pixel_1088/SF_IB
+ pixel_1088/PIX_OUT pixel_1088/CSA_VREF pixel
Xpixel_1077 pixel_1077/gring pixel_1077/VDD pixel_1077/GND pixel_1077/VREF pixel_1077/ROW_SEL
+ pixel_1077/NB1 pixel_1077/VBIAS pixel_1077/NB2 pixel_1077/AMP_IN pixel_1077/SF_IB
+ pixel_1077/PIX_OUT pixel_1077/CSA_VREF pixel
Xpixel_9341 pixel_9341/gring pixel_9341/VDD pixel_9341/GND pixel_9341/VREF pixel_9341/ROW_SEL
+ pixel_9341/NB1 pixel_9341/VBIAS pixel_9341/NB2 pixel_9341/AMP_IN pixel_9341/SF_IB
+ pixel_9341/PIX_OUT pixel_9341/CSA_VREF pixel
Xpixel_9330 pixel_9330/gring pixel_9330/VDD pixel_9330/GND pixel_9330/VREF pixel_9330/ROW_SEL
+ pixel_9330/NB1 pixel_9330/VBIAS pixel_9330/NB2 pixel_9330/AMP_IN pixel_9330/SF_IB
+ pixel_9330/PIX_OUT pixel_9330/CSA_VREF pixel
Xpixel_9374 pixel_9374/gring pixel_9374/VDD pixel_9374/GND pixel_9374/VREF pixel_9374/ROW_SEL
+ pixel_9374/NB1 pixel_9374/VBIAS pixel_9374/NB2 pixel_9374/AMP_IN pixel_9374/SF_IB
+ pixel_9374/PIX_OUT pixel_9374/CSA_VREF pixel
Xpixel_9363 pixel_9363/gring pixel_9363/VDD pixel_9363/GND pixel_9363/VREF pixel_9363/ROW_SEL
+ pixel_9363/NB1 pixel_9363/VBIAS pixel_9363/NB2 pixel_9363/AMP_IN pixel_9363/SF_IB
+ pixel_9363/PIX_OUT pixel_9363/CSA_VREF pixel
Xpixel_9352 pixel_9352/gring pixel_9352/VDD pixel_9352/GND pixel_9352/VREF pixel_9352/ROW_SEL
+ pixel_9352/NB1 pixel_9352/VBIAS pixel_9352/NB2 pixel_9352/AMP_IN pixel_9352/SF_IB
+ pixel_9352/PIX_OUT pixel_9352/CSA_VREF pixel
Xpixel_8662 pixel_8662/gring pixel_8662/VDD pixel_8662/GND pixel_8662/VREF pixel_8662/ROW_SEL
+ pixel_8662/NB1 pixel_8662/VBIAS pixel_8662/NB2 pixel_8662/AMP_IN pixel_8662/SF_IB
+ pixel_8662/PIX_OUT pixel_8662/CSA_VREF pixel
Xpixel_8651 pixel_8651/gring pixel_8651/VDD pixel_8651/GND pixel_8651/VREF pixel_8651/ROW_SEL
+ pixel_8651/NB1 pixel_8651/VBIAS pixel_8651/NB2 pixel_8651/AMP_IN pixel_8651/SF_IB
+ pixel_8651/PIX_OUT pixel_8651/CSA_VREF pixel
Xpixel_8640 pixel_8640/gring pixel_8640/VDD pixel_8640/GND pixel_8640/VREF pixel_8640/ROW_SEL
+ pixel_8640/NB1 pixel_8640/VBIAS pixel_8640/NB2 pixel_8640/AMP_IN pixel_8640/SF_IB
+ pixel_8640/PIX_OUT pixel_8640/CSA_VREF pixel
Xpixel_9396 pixel_9396/gring pixel_9396/VDD pixel_9396/GND pixel_9396/VREF pixel_9396/ROW_SEL
+ pixel_9396/NB1 pixel_9396/VBIAS pixel_9396/NB2 pixel_9396/AMP_IN pixel_9396/SF_IB
+ pixel_9396/PIX_OUT pixel_9396/CSA_VREF pixel
Xpixel_9385 pixel_9385/gring pixel_9385/VDD pixel_9385/GND pixel_9385/VREF pixel_9385/ROW_SEL
+ pixel_9385/NB1 pixel_9385/VBIAS pixel_9385/NB2 pixel_9385/AMP_IN pixel_9385/SF_IB
+ pixel_9385/PIX_OUT pixel_9385/CSA_VREF pixel
Xpixel_8695 pixel_8695/gring pixel_8695/VDD pixel_8695/GND pixel_8695/VREF pixel_8695/ROW_SEL
+ pixel_8695/NB1 pixel_8695/VBIAS pixel_8695/NB2 pixel_8695/AMP_IN pixel_8695/SF_IB
+ pixel_8695/PIX_OUT pixel_8695/CSA_VREF pixel
Xpixel_8684 pixel_8684/gring pixel_8684/VDD pixel_8684/GND pixel_8684/VREF pixel_8684/ROW_SEL
+ pixel_8684/NB1 pixel_8684/VBIAS pixel_8684/NB2 pixel_8684/AMP_IN pixel_8684/SF_IB
+ pixel_8684/PIX_OUT pixel_8684/CSA_VREF pixel
Xpixel_8673 pixel_8673/gring pixel_8673/VDD pixel_8673/GND pixel_8673/VREF pixel_8673/ROW_SEL
+ pixel_8673/NB1 pixel_8673/VBIAS pixel_8673/NB2 pixel_8673/AMP_IN pixel_8673/SF_IB
+ pixel_8673/PIX_OUT pixel_8673/CSA_VREF pixel
Xpixel_7950 pixel_7950/gring pixel_7950/VDD pixel_7950/GND pixel_7950/VREF pixel_7950/ROW_SEL
+ pixel_7950/NB1 pixel_7950/VBIAS pixel_7950/NB2 pixel_7950/AMP_IN pixel_7950/SF_IB
+ pixel_7950/PIX_OUT pixel_7950/CSA_VREF pixel
Xpixel_7961 pixel_7961/gring pixel_7961/VDD pixel_7961/GND pixel_7961/VREF pixel_7961/ROW_SEL
+ pixel_7961/NB1 pixel_7961/VBIAS pixel_7961/NB2 pixel_7961/AMP_IN pixel_7961/SF_IB
+ pixel_7961/PIX_OUT pixel_7961/CSA_VREF pixel
Xpixel_7972 pixel_7972/gring pixel_7972/VDD pixel_7972/GND pixel_7972/VREF pixel_7972/ROW_SEL
+ pixel_7972/NB1 pixel_7972/VBIAS pixel_7972/NB2 pixel_7972/AMP_IN pixel_7972/SF_IB
+ pixel_7972/PIX_OUT pixel_7972/CSA_VREF pixel
Xpixel_7983 pixel_7983/gring pixel_7983/VDD pixel_7983/GND pixel_7983/VREF pixel_7983/ROW_SEL
+ pixel_7983/NB1 pixel_7983/VBIAS pixel_7983/NB2 pixel_7983/AMP_IN pixel_7983/SF_IB
+ pixel_7983/PIX_OUT pixel_7983/CSA_VREF pixel
Xpixel_7994 pixel_7994/gring pixel_7994/VDD pixel_7994/GND pixel_7994/VREF pixel_7994/ROW_SEL
+ pixel_7994/NB1 pixel_7994/VBIAS pixel_7994/NB2 pixel_7994/AMP_IN pixel_7994/SF_IB
+ pixel_7994/PIX_OUT pixel_7994/CSA_VREF pixel
Xpixel_2290 pixel_2290/gring pixel_2290/VDD pixel_2290/GND pixel_2290/VREF pixel_2290/ROW_SEL
+ pixel_2290/NB1 pixel_2290/VBIAS pixel_2290/NB2 pixel_2290/AMP_IN pixel_2290/SF_IB
+ pixel_2290/PIX_OUT pixel_2290/CSA_VREF pixel
Xpixel_604 pixel_604/gring pixel_604/VDD pixel_604/GND pixel_604/VREF pixel_604/ROW_SEL
+ pixel_604/NB1 pixel_604/VBIAS pixel_604/NB2 pixel_604/AMP_IN pixel_604/SF_IB pixel_604/PIX_OUT
+ pixel_604/CSA_VREF pixel
Xpixel_4609 pixel_4609/gring pixel_4609/VDD pixel_4609/GND pixel_4609/VREF pixel_4609/ROW_SEL
+ pixel_4609/NB1 pixel_4609/VBIAS pixel_4609/NB2 pixel_4609/AMP_IN pixel_4609/SF_IB
+ pixel_4609/PIX_OUT pixel_4609/CSA_VREF pixel
Xpixel_648 pixel_648/gring pixel_648/VDD pixel_648/GND pixel_648/VREF pixel_648/ROW_SEL
+ pixel_648/NB1 pixel_648/VBIAS pixel_648/NB2 pixel_648/AMP_IN pixel_648/SF_IB pixel_648/PIX_OUT
+ pixel_648/CSA_VREF pixel
Xpixel_637 pixel_637/gring pixel_637/VDD pixel_637/GND pixel_637/VREF pixel_637/ROW_SEL
+ pixel_637/NB1 pixel_637/VBIAS pixel_637/NB2 pixel_637/AMP_IN pixel_637/SF_IB pixel_637/PIX_OUT
+ pixel_637/CSA_VREF pixel
Xpixel_626 pixel_626/gring pixel_626/VDD pixel_626/GND pixel_626/VREF pixel_626/ROW_SEL
+ pixel_626/NB1 pixel_626/VBIAS pixel_626/NB2 pixel_626/AMP_IN pixel_626/SF_IB pixel_626/PIX_OUT
+ pixel_626/CSA_VREF pixel
Xpixel_615 pixel_615/gring pixel_615/VDD pixel_615/GND pixel_615/VREF pixel_615/ROW_SEL
+ pixel_615/NB1 pixel_615/VBIAS pixel_615/NB2 pixel_615/AMP_IN pixel_615/SF_IB pixel_615/PIX_OUT
+ pixel_615/CSA_VREF pixel
Xpixel_3908 pixel_3908/gring pixel_3908/VDD pixel_3908/GND pixel_3908/VREF pixel_3908/ROW_SEL
+ pixel_3908/NB1 pixel_3908/VBIAS pixel_3908/NB2 pixel_3908/AMP_IN pixel_3908/SF_IB
+ pixel_3908/PIX_OUT pixel_3908/CSA_VREF pixel
Xpixel_659 pixel_659/gring pixel_659/VDD pixel_659/GND pixel_659/VREF pixel_659/ROW_SEL
+ pixel_659/NB1 pixel_659/VBIAS pixel_659/NB2 pixel_659/AMP_IN pixel_659/SF_IB pixel_659/PIX_OUT
+ pixel_659/CSA_VREF pixel
Xpixel_3919 pixel_3919/gring pixel_3919/VDD pixel_3919/GND pixel_3919/VREF pixel_3919/ROW_SEL
+ pixel_3919/NB1 pixel_3919/VBIAS pixel_3919/NB2 pixel_3919/AMP_IN pixel_3919/SF_IB
+ pixel_3919/PIX_OUT pixel_3919/CSA_VREF pixel
Xpixel_7202 pixel_7202/gring pixel_7202/VDD pixel_7202/GND pixel_7202/VREF pixel_7202/ROW_SEL
+ pixel_7202/NB1 pixel_7202/VBIAS pixel_7202/NB2 pixel_7202/AMP_IN pixel_7202/SF_IB
+ pixel_7202/PIX_OUT pixel_7202/CSA_VREF pixel
Xpixel_7213 pixel_7213/gring pixel_7213/VDD pixel_7213/GND pixel_7213/VREF pixel_7213/ROW_SEL
+ pixel_7213/NB1 pixel_7213/VBIAS pixel_7213/NB2 pixel_7213/AMP_IN pixel_7213/SF_IB
+ pixel_7213/PIX_OUT pixel_7213/CSA_VREF pixel
Xpixel_7224 pixel_7224/gring pixel_7224/VDD pixel_7224/GND pixel_7224/VREF pixel_7224/ROW_SEL
+ pixel_7224/NB1 pixel_7224/VBIAS pixel_7224/NB2 pixel_7224/AMP_IN pixel_7224/SF_IB
+ pixel_7224/PIX_OUT pixel_7224/CSA_VREF pixel
Xpixel_7235 pixel_7235/gring pixel_7235/VDD pixel_7235/GND pixel_7235/VREF pixel_7235/ROW_SEL
+ pixel_7235/NB1 pixel_7235/VBIAS pixel_7235/NB2 pixel_7235/AMP_IN pixel_7235/SF_IB
+ pixel_7235/PIX_OUT pixel_7235/CSA_VREF pixel
Xpixel_7246 pixel_7246/gring pixel_7246/VDD pixel_7246/GND pixel_7246/VREF pixel_7246/ROW_SEL
+ pixel_7246/NB1 pixel_7246/VBIAS pixel_7246/NB2 pixel_7246/AMP_IN pixel_7246/SF_IB
+ pixel_7246/PIX_OUT pixel_7246/CSA_VREF pixel
Xpixel_6501 pixel_6501/gring pixel_6501/VDD pixel_6501/GND pixel_6501/VREF pixel_6501/ROW_SEL
+ pixel_6501/NB1 pixel_6501/VBIAS pixel_6501/NB2 pixel_6501/AMP_IN pixel_6501/SF_IB
+ pixel_6501/PIX_OUT pixel_6501/CSA_VREF pixel
Xpixel_6512 pixel_6512/gring pixel_6512/VDD pixel_6512/GND pixel_6512/VREF pixel_6512/ROW_SEL
+ pixel_6512/NB1 pixel_6512/VBIAS pixel_6512/NB2 pixel_6512/AMP_IN pixel_6512/SF_IB
+ pixel_6512/PIX_OUT pixel_6512/CSA_VREF pixel
Xpixel_7257 pixel_7257/gring pixel_7257/VDD pixel_7257/GND pixel_7257/VREF pixel_7257/ROW_SEL
+ pixel_7257/NB1 pixel_7257/VBIAS pixel_7257/NB2 pixel_7257/AMP_IN pixel_7257/SF_IB
+ pixel_7257/PIX_OUT pixel_7257/CSA_VREF pixel
Xpixel_7268 pixel_7268/gring pixel_7268/VDD pixel_7268/GND pixel_7268/VREF pixel_7268/ROW_SEL
+ pixel_7268/NB1 pixel_7268/VBIAS pixel_7268/NB2 pixel_7268/AMP_IN pixel_7268/SF_IB
+ pixel_7268/PIX_OUT pixel_7268/CSA_VREF pixel
Xpixel_7279 pixel_7279/gring pixel_7279/VDD pixel_7279/GND pixel_7279/VREF pixel_7279/ROW_SEL
+ pixel_7279/NB1 pixel_7279/VBIAS pixel_7279/NB2 pixel_7279/AMP_IN pixel_7279/SF_IB
+ pixel_7279/PIX_OUT pixel_7279/CSA_VREF pixel
Xpixel_6523 pixel_6523/gring pixel_6523/VDD pixel_6523/GND pixel_6523/VREF pixel_6523/ROW_SEL
+ pixel_6523/NB1 pixel_6523/VBIAS pixel_6523/NB2 pixel_6523/AMP_IN pixel_6523/SF_IB
+ pixel_6523/PIX_OUT pixel_6523/CSA_VREF pixel
Xpixel_6534 pixel_6534/gring pixel_6534/VDD pixel_6534/GND pixel_6534/VREF pixel_6534/ROW_SEL
+ pixel_6534/NB1 pixel_6534/VBIAS pixel_6534/NB2 pixel_6534/AMP_IN pixel_6534/SF_IB
+ pixel_6534/PIX_OUT pixel_6534/CSA_VREF pixel
Xpixel_6545 pixel_6545/gring pixel_6545/VDD pixel_6545/GND pixel_6545/VREF pixel_6545/ROW_SEL
+ pixel_6545/NB1 pixel_6545/VBIAS pixel_6545/NB2 pixel_6545/AMP_IN pixel_6545/SF_IB
+ pixel_6545/PIX_OUT pixel_6545/CSA_VREF pixel
Xpixel_5800 pixel_5800/gring pixel_5800/VDD pixel_5800/GND pixel_5800/VREF pixel_5800/ROW_SEL
+ pixel_5800/NB1 pixel_5800/VBIAS pixel_5800/NB2 pixel_5800/AMP_IN pixel_5800/SF_IB
+ pixel_5800/PIX_OUT pixel_5800/CSA_VREF pixel
Xpixel_6556 pixel_6556/gring pixel_6556/VDD pixel_6556/GND pixel_6556/VREF pixel_6556/ROW_SEL
+ pixel_6556/NB1 pixel_6556/VBIAS pixel_6556/NB2 pixel_6556/AMP_IN pixel_6556/SF_IB
+ pixel_6556/PIX_OUT pixel_6556/CSA_VREF pixel
Xpixel_6567 pixel_6567/gring pixel_6567/VDD pixel_6567/GND pixel_6567/VREF pixel_6567/ROW_SEL
+ pixel_6567/NB1 pixel_6567/VBIAS pixel_6567/NB2 pixel_6567/AMP_IN pixel_6567/SF_IB
+ pixel_6567/PIX_OUT pixel_6567/CSA_VREF pixel
Xpixel_6578 pixel_6578/gring pixel_6578/VDD pixel_6578/GND pixel_6578/VREF pixel_6578/ROW_SEL
+ pixel_6578/NB1 pixel_6578/VBIAS pixel_6578/NB2 pixel_6578/AMP_IN pixel_6578/SF_IB
+ pixel_6578/PIX_OUT pixel_6578/CSA_VREF pixel
Xpixel_5811 pixel_5811/gring pixel_5811/VDD pixel_5811/GND pixel_5811/VREF pixel_5811/ROW_SEL
+ pixel_5811/NB1 pixel_5811/VBIAS pixel_5811/NB2 pixel_5811/AMP_IN pixel_5811/SF_IB
+ pixel_5811/PIX_OUT pixel_5811/CSA_VREF pixel
Xpixel_5822 pixel_5822/gring pixel_5822/VDD pixel_5822/GND pixel_5822/VREF pixel_5822/ROW_SEL
+ pixel_5822/NB1 pixel_5822/VBIAS pixel_5822/NB2 pixel_5822/AMP_IN pixel_5822/SF_IB
+ pixel_5822/PIX_OUT pixel_5822/CSA_VREF pixel
Xpixel_5833 pixel_5833/gring pixel_5833/VDD pixel_5833/GND pixel_5833/VREF pixel_5833/ROW_SEL
+ pixel_5833/NB1 pixel_5833/VBIAS pixel_5833/NB2 pixel_5833/AMP_IN pixel_5833/SF_IB
+ pixel_5833/PIX_OUT pixel_5833/CSA_VREF pixel
Xpixel_6589 pixel_6589/gring pixel_6589/VDD pixel_6589/GND pixel_6589/VREF pixel_6589/ROW_SEL
+ pixel_6589/NB1 pixel_6589/VBIAS pixel_6589/NB2 pixel_6589/AMP_IN pixel_6589/SF_IB
+ pixel_6589/PIX_OUT pixel_6589/CSA_VREF pixel
Xpixel_5844 pixel_5844/gring pixel_5844/VDD pixel_5844/GND pixel_5844/VREF pixel_5844/ROW_SEL
+ pixel_5844/NB1 pixel_5844/VBIAS pixel_5844/NB2 pixel_5844/AMP_IN pixel_5844/SF_IB
+ pixel_5844/PIX_OUT pixel_5844/CSA_VREF pixel
Xpixel_5855 pixel_5855/gring pixel_5855/VDD pixel_5855/GND pixel_5855/VREF pixel_5855/ROW_SEL
+ pixel_5855/NB1 pixel_5855/VBIAS pixel_5855/NB2 pixel_5855/AMP_IN pixel_5855/SF_IB
+ pixel_5855/PIX_OUT pixel_5855/CSA_VREF pixel
Xpixel_5866 pixel_5866/gring pixel_5866/VDD pixel_5866/GND pixel_5866/VREF pixel_5866/ROW_SEL
+ pixel_5866/NB1 pixel_5866/VBIAS pixel_5866/NB2 pixel_5866/AMP_IN pixel_5866/SF_IB
+ pixel_5866/PIX_OUT pixel_5866/CSA_VREF pixel
Xpixel_5877 pixel_5877/gring pixel_5877/VDD pixel_5877/GND pixel_5877/VREF pixel_5877/ROW_SEL
+ pixel_5877/NB1 pixel_5877/VBIAS pixel_5877/NB2 pixel_5877/AMP_IN pixel_5877/SF_IB
+ pixel_5877/PIX_OUT pixel_5877/CSA_VREF pixel
Xpixel_5888 pixel_5888/gring pixel_5888/VDD pixel_5888/GND pixel_5888/VREF pixel_5888/ROW_SEL
+ pixel_5888/NB1 pixel_5888/VBIAS pixel_5888/NB2 pixel_5888/AMP_IN pixel_5888/SF_IB
+ pixel_5888/PIX_OUT pixel_5888/CSA_VREF pixel
Xpixel_5899 pixel_5899/gring pixel_5899/VDD pixel_5899/GND pixel_5899/VREF pixel_5899/ROW_SEL
+ pixel_5899/NB1 pixel_5899/VBIAS pixel_5899/NB2 pixel_5899/AMP_IN pixel_5899/SF_IB
+ pixel_5899/PIX_OUT pixel_5899/CSA_VREF pixel
Xpixel_9182 pixel_9182/gring pixel_9182/VDD pixel_9182/GND pixel_9182/VREF pixel_9182/ROW_SEL
+ pixel_9182/NB1 pixel_9182/VBIAS pixel_9182/NB2 pixel_9182/AMP_IN pixel_9182/SF_IB
+ pixel_9182/PIX_OUT pixel_9182/CSA_VREF pixel
Xpixel_9171 pixel_9171/gring pixel_9171/VDD pixel_9171/GND pixel_9171/VREF pixel_9171/ROW_SEL
+ pixel_9171/NB1 pixel_9171/VBIAS pixel_9171/NB2 pixel_9171/AMP_IN pixel_9171/SF_IB
+ pixel_9171/PIX_OUT pixel_9171/CSA_VREF pixel
Xpixel_9160 pixel_9160/gring pixel_9160/VDD pixel_9160/GND pixel_9160/VREF pixel_9160/ROW_SEL
+ pixel_9160/NB1 pixel_9160/VBIAS pixel_9160/NB2 pixel_9160/AMP_IN pixel_9160/SF_IB
+ pixel_9160/PIX_OUT pixel_9160/CSA_VREF pixel
Xpixel_9193 pixel_9193/gring pixel_9193/VDD pixel_9193/GND pixel_9193/VREF pixel_9193/ROW_SEL
+ pixel_9193/NB1 pixel_9193/VBIAS pixel_9193/NB2 pixel_9193/AMP_IN pixel_9193/SF_IB
+ pixel_9193/PIX_OUT pixel_9193/CSA_VREF pixel
Xpixel_8470 pixel_8470/gring pixel_8470/VDD pixel_8470/GND pixel_8470/VREF pixel_8470/ROW_SEL
+ pixel_8470/NB1 pixel_8470/VBIAS pixel_8470/NB2 pixel_8470/AMP_IN pixel_8470/SF_IB
+ pixel_8470/PIX_OUT pixel_8470/CSA_VREF pixel
Xpixel_8481 pixel_8481/gring pixel_8481/VDD pixel_8481/GND pixel_8481/VREF pixel_8481/ROW_SEL
+ pixel_8481/NB1 pixel_8481/VBIAS pixel_8481/NB2 pixel_8481/AMP_IN pixel_8481/SF_IB
+ pixel_8481/PIX_OUT pixel_8481/CSA_VREF pixel
Xpixel_8492 pixel_8492/gring pixel_8492/VDD pixel_8492/GND pixel_8492/VREF pixel_8492/ROW_SEL
+ pixel_8492/NB1 pixel_8492/VBIAS pixel_8492/NB2 pixel_8492/AMP_IN pixel_8492/SF_IB
+ pixel_8492/PIX_OUT pixel_8492/CSA_VREF pixel
Xpixel_7780 pixel_7780/gring pixel_7780/VDD pixel_7780/GND pixel_7780/VREF pixel_7780/ROW_SEL
+ pixel_7780/NB1 pixel_7780/VBIAS pixel_7780/NB2 pixel_7780/AMP_IN pixel_7780/SF_IB
+ pixel_7780/PIX_OUT pixel_7780/CSA_VREF pixel
Xpixel_7791 pixel_7791/gring pixel_7791/VDD pixel_7791/GND pixel_7791/VREF pixel_7791/ROW_SEL
+ pixel_7791/NB1 pixel_7791/VBIAS pixel_7791/NB2 pixel_7791/AMP_IN pixel_7791/SF_IB
+ pixel_7791/PIX_OUT pixel_7791/CSA_VREF pixel
Xpixel_5107 pixel_5107/gring pixel_5107/VDD pixel_5107/GND pixel_5107/VREF pixel_5107/ROW_SEL
+ pixel_5107/NB1 pixel_5107/VBIAS pixel_5107/NB2 pixel_5107/AMP_IN pixel_5107/SF_IB
+ pixel_5107/PIX_OUT pixel_5107/CSA_VREF pixel
Xpixel_5118 pixel_5118/gring pixel_5118/VDD pixel_5118/GND pixel_5118/VREF pixel_5118/ROW_SEL
+ pixel_5118/NB1 pixel_5118/VBIAS pixel_5118/NB2 pixel_5118/AMP_IN pixel_5118/SF_IB
+ pixel_5118/PIX_OUT pixel_5118/CSA_VREF pixel
Xpixel_5129 pixel_5129/gring pixel_5129/VDD pixel_5129/GND pixel_5129/VREF pixel_5129/ROW_SEL
+ pixel_5129/NB1 pixel_5129/VBIAS pixel_5129/NB2 pixel_5129/AMP_IN pixel_5129/SF_IB
+ pixel_5129/PIX_OUT pixel_5129/CSA_VREF pixel
Xpixel_423 pixel_423/gring pixel_423/VDD pixel_423/GND pixel_423/VREF pixel_423/ROW_SEL
+ pixel_423/NB1 pixel_423/VBIAS pixel_423/NB2 pixel_423/AMP_IN pixel_423/SF_IB pixel_423/PIX_OUT
+ pixel_423/CSA_VREF pixel
Xpixel_412 pixel_412/gring pixel_412/VDD pixel_412/GND pixel_412/VREF pixel_412/ROW_SEL
+ pixel_412/NB1 pixel_412/VBIAS pixel_412/NB2 pixel_412/AMP_IN pixel_412/SF_IB pixel_412/PIX_OUT
+ pixel_412/CSA_VREF pixel
Xpixel_401 pixel_401/gring pixel_401/VDD pixel_401/GND pixel_401/VREF pixel_401/ROW_SEL
+ pixel_401/NB1 pixel_401/VBIAS pixel_401/NB2 pixel_401/AMP_IN pixel_401/SF_IB pixel_401/PIX_OUT
+ pixel_401/CSA_VREF pixel
Xpixel_4406 pixel_4406/gring pixel_4406/VDD pixel_4406/GND pixel_4406/VREF pixel_4406/ROW_SEL
+ pixel_4406/NB1 pixel_4406/VBIAS pixel_4406/NB2 pixel_4406/AMP_IN pixel_4406/SF_IB
+ pixel_4406/PIX_OUT pixel_4406/CSA_VREF pixel
Xpixel_4417 pixel_4417/gring pixel_4417/VDD pixel_4417/GND pixel_4417/VREF pixel_4417/ROW_SEL
+ pixel_4417/NB1 pixel_4417/VBIAS pixel_4417/NB2 pixel_4417/AMP_IN pixel_4417/SF_IB
+ pixel_4417/PIX_OUT pixel_4417/CSA_VREF pixel
Xpixel_456 pixel_456/gring pixel_456/VDD pixel_456/GND pixel_456/VREF pixel_456/ROW_SEL
+ pixel_456/NB1 pixel_456/VBIAS pixel_456/NB2 pixel_456/AMP_IN pixel_456/SF_IB pixel_456/PIX_OUT
+ pixel_456/CSA_VREF pixel
Xpixel_445 pixel_445/gring pixel_445/VDD pixel_445/GND pixel_445/VREF pixel_445/ROW_SEL
+ pixel_445/NB1 pixel_445/VBIAS pixel_445/NB2 pixel_445/AMP_IN pixel_445/SF_IB pixel_445/PIX_OUT
+ pixel_445/CSA_VREF pixel
Xpixel_434 pixel_434/gring pixel_434/VDD pixel_434/GND pixel_434/VREF pixel_434/ROW_SEL
+ pixel_434/NB1 pixel_434/VBIAS pixel_434/NB2 pixel_434/AMP_IN pixel_434/SF_IB pixel_434/PIX_OUT
+ pixel_434/CSA_VREF pixel
Xpixel_3716 pixel_3716/gring pixel_3716/VDD pixel_3716/GND pixel_3716/VREF pixel_3716/ROW_SEL
+ pixel_3716/NB1 pixel_3716/VBIAS pixel_3716/NB2 pixel_3716/AMP_IN pixel_3716/SF_IB
+ pixel_3716/PIX_OUT pixel_3716/CSA_VREF pixel
Xpixel_3705 pixel_3705/gring pixel_3705/VDD pixel_3705/GND pixel_3705/VREF pixel_3705/ROW_SEL
+ pixel_3705/NB1 pixel_3705/VBIAS pixel_3705/NB2 pixel_3705/AMP_IN pixel_3705/SF_IB
+ pixel_3705/PIX_OUT pixel_3705/CSA_VREF pixel
Xpixel_4428 pixel_4428/gring pixel_4428/VDD pixel_4428/GND pixel_4428/VREF pixel_4428/ROW_SEL
+ pixel_4428/NB1 pixel_4428/VBIAS pixel_4428/NB2 pixel_4428/AMP_IN pixel_4428/SF_IB
+ pixel_4428/PIX_OUT pixel_4428/CSA_VREF pixel
Xpixel_4439 pixel_4439/gring pixel_4439/VDD pixel_4439/GND pixel_4439/VREF pixel_4439/ROW_SEL
+ pixel_4439/NB1 pixel_4439/VBIAS pixel_4439/NB2 pixel_4439/AMP_IN pixel_4439/SF_IB
+ pixel_4439/PIX_OUT pixel_4439/CSA_VREF pixel
Xpixel_489 pixel_489/gring pixel_489/VDD pixel_489/GND pixel_489/VREF pixel_489/ROW_SEL
+ pixel_489/NB1 pixel_489/VBIAS pixel_489/NB2 pixel_489/AMP_IN pixel_489/SF_IB pixel_489/PIX_OUT
+ pixel_489/CSA_VREF pixel
Xpixel_478 pixel_478/gring pixel_478/VDD pixel_478/GND pixel_478/VREF pixel_478/ROW_SEL
+ pixel_478/NB1 pixel_478/VBIAS pixel_478/NB2 pixel_478/AMP_IN pixel_478/SF_IB pixel_478/PIX_OUT
+ pixel_478/CSA_VREF pixel
Xpixel_467 pixel_467/gring pixel_467/VDD pixel_467/GND pixel_467/VREF pixel_467/ROW_SEL
+ pixel_467/NB1 pixel_467/VBIAS pixel_467/NB2 pixel_467/AMP_IN pixel_467/SF_IB pixel_467/PIX_OUT
+ pixel_467/CSA_VREF pixel
Xpixel_3749 pixel_3749/gring pixel_3749/VDD pixel_3749/GND pixel_3749/VREF pixel_3749/ROW_SEL
+ pixel_3749/NB1 pixel_3749/VBIAS pixel_3749/NB2 pixel_3749/AMP_IN pixel_3749/SF_IB
+ pixel_3749/PIX_OUT pixel_3749/CSA_VREF pixel
Xpixel_3738 pixel_3738/gring pixel_3738/VDD pixel_3738/GND pixel_3738/VREF pixel_3738/ROW_SEL
+ pixel_3738/NB1 pixel_3738/VBIAS pixel_3738/NB2 pixel_3738/AMP_IN pixel_3738/SF_IB
+ pixel_3738/PIX_OUT pixel_3738/CSA_VREF pixel
Xpixel_3727 pixel_3727/gring pixel_3727/VDD pixel_3727/GND pixel_3727/VREF pixel_3727/ROW_SEL
+ pixel_3727/NB1 pixel_3727/VBIAS pixel_3727/NB2 pixel_3727/AMP_IN pixel_3727/SF_IB
+ pixel_3727/PIX_OUT pixel_3727/CSA_VREF pixel
Xpixel_7010 pixel_7010/gring pixel_7010/VDD pixel_7010/GND pixel_7010/VREF pixel_7010/ROW_SEL
+ pixel_7010/NB1 pixel_7010/VBIAS pixel_7010/NB2 pixel_7010/AMP_IN pixel_7010/SF_IB
+ pixel_7010/PIX_OUT pixel_7010/CSA_VREF pixel
Xpixel_7021 pixel_7021/gring pixel_7021/VDD pixel_7021/GND pixel_7021/VREF pixel_7021/ROW_SEL
+ pixel_7021/NB1 pixel_7021/VBIAS pixel_7021/NB2 pixel_7021/AMP_IN pixel_7021/SF_IB
+ pixel_7021/PIX_OUT pixel_7021/CSA_VREF pixel
Xpixel_7032 pixel_7032/gring pixel_7032/VDD pixel_7032/GND pixel_7032/VREF pixel_7032/ROW_SEL
+ pixel_7032/NB1 pixel_7032/VBIAS pixel_7032/NB2 pixel_7032/AMP_IN pixel_7032/SF_IB
+ pixel_7032/PIX_OUT pixel_7032/CSA_VREF pixel
Xpixel_7043 pixel_7043/gring pixel_7043/VDD pixel_7043/GND pixel_7043/VREF pixel_7043/ROW_SEL
+ pixel_7043/NB1 pixel_7043/VBIAS pixel_7043/NB2 pixel_7043/AMP_IN pixel_7043/SF_IB
+ pixel_7043/PIX_OUT pixel_7043/CSA_VREF pixel
Xpixel_7054 pixel_7054/gring pixel_7054/VDD pixel_7054/GND pixel_7054/VREF pixel_7054/ROW_SEL
+ pixel_7054/NB1 pixel_7054/VBIAS pixel_7054/NB2 pixel_7054/AMP_IN pixel_7054/SF_IB
+ pixel_7054/PIX_OUT pixel_7054/CSA_VREF pixel
Xpixel_7065 pixel_7065/gring pixel_7065/VDD pixel_7065/GND pixel_7065/VREF pixel_7065/ROW_SEL
+ pixel_7065/NB1 pixel_7065/VBIAS pixel_7065/NB2 pixel_7065/AMP_IN pixel_7065/SF_IB
+ pixel_7065/PIX_OUT pixel_7065/CSA_VREF pixel
Xpixel_6320 pixel_6320/gring pixel_6320/VDD pixel_6320/GND pixel_6320/VREF pixel_6320/ROW_SEL
+ pixel_6320/NB1 pixel_6320/VBIAS pixel_6320/NB2 pixel_6320/AMP_IN pixel_6320/SF_IB
+ pixel_6320/PIX_OUT pixel_6320/CSA_VREF pixel
Xpixel_7076 pixel_7076/gring pixel_7076/VDD pixel_7076/GND pixel_7076/VREF pixel_7076/ROW_SEL
+ pixel_7076/NB1 pixel_7076/VBIAS pixel_7076/NB2 pixel_7076/AMP_IN pixel_7076/SF_IB
+ pixel_7076/PIX_OUT pixel_7076/CSA_VREF pixel
Xpixel_7087 pixel_7087/gring pixel_7087/VDD pixel_7087/GND pixel_7087/VREF pixel_7087/ROW_SEL
+ pixel_7087/NB1 pixel_7087/VBIAS pixel_7087/NB2 pixel_7087/AMP_IN pixel_7087/SF_IB
+ pixel_7087/PIX_OUT pixel_7087/CSA_VREF pixel
Xpixel_7098 pixel_7098/gring pixel_7098/VDD pixel_7098/GND pixel_7098/VREF pixel_7098/ROW_SEL
+ pixel_7098/NB1 pixel_7098/VBIAS pixel_7098/NB2 pixel_7098/AMP_IN pixel_7098/SF_IB
+ pixel_7098/PIX_OUT pixel_7098/CSA_VREF pixel
Xpixel_6331 pixel_6331/gring pixel_6331/VDD pixel_6331/GND pixel_6331/VREF pixel_6331/ROW_SEL
+ pixel_6331/NB1 pixel_6331/VBIAS pixel_6331/NB2 pixel_6331/AMP_IN pixel_6331/SF_IB
+ pixel_6331/PIX_OUT pixel_6331/CSA_VREF pixel
Xpixel_6342 pixel_6342/gring pixel_6342/VDD pixel_6342/GND pixel_6342/VREF pixel_6342/ROW_SEL
+ pixel_6342/NB1 pixel_6342/VBIAS pixel_6342/NB2 pixel_6342/AMP_IN pixel_6342/SF_IB
+ pixel_6342/PIX_OUT pixel_6342/CSA_VREF pixel
Xpixel_6353 pixel_6353/gring pixel_6353/VDD pixel_6353/GND pixel_6353/VREF pixel_6353/ROW_SEL
+ pixel_6353/NB1 pixel_6353/VBIAS pixel_6353/NB2 pixel_6353/AMP_IN pixel_6353/SF_IB
+ pixel_6353/PIX_OUT pixel_6353/CSA_VREF pixel
Xpixel_6364 pixel_6364/gring pixel_6364/VDD pixel_6364/GND pixel_6364/VREF pixel_6364/ROW_SEL
+ pixel_6364/NB1 pixel_6364/VBIAS pixel_6364/NB2 pixel_6364/AMP_IN pixel_6364/SF_IB
+ pixel_6364/PIX_OUT pixel_6364/CSA_VREF pixel
Xpixel_6375 pixel_6375/gring pixel_6375/VDD pixel_6375/GND pixel_6375/VREF pixel_6375/ROW_SEL
+ pixel_6375/NB1 pixel_6375/VBIAS pixel_6375/NB2 pixel_6375/AMP_IN pixel_6375/SF_IB
+ pixel_6375/PIX_OUT pixel_6375/CSA_VREF pixel
Xpixel_6386 pixel_6386/gring pixel_6386/VDD pixel_6386/GND pixel_6386/VREF pixel_6386/ROW_SEL
+ pixel_6386/NB1 pixel_6386/VBIAS pixel_6386/NB2 pixel_6386/AMP_IN pixel_6386/SF_IB
+ pixel_6386/PIX_OUT pixel_6386/CSA_VREF pixel
Xpixel_5630 pixel_5630/gring pixel_5630/VDD pixel_5630/GND pixel_5630/VREF pixel_5630/ROW_SEL
+ pixel_5630/NB1 pixel_5630/VBIAS pixel_5630/NB2 pixel_5630/AMP_IN pixel_5630/SF_IB
+ pixel_5630/PIX_OUT pixel_5630/CSA_VREF pixel
Xpixel_5641 pixel_5641/gring pixel_5641/VDD pixel_5641/GND pixel_5641/VREF pixel_5641/ROW_SEL
+ pixel_5641/NB1 pixel_5641/VBIAS pixel_5641/NB2 pixel_5641/AMP_IN pixel_5641/SF_IB
+ pixel_5641/PIX_OUT pixel_5641/CSA_VREF pixel
Xpixel_6397 pixel_6397/gring pixel_6397/VDD pixel_6397/GND pixel_6397/VREF pixel_6397/ROW_SEL
+ pixel_6397/NB1 pixel_6397/VBIAS pixel_6397/NB2 pixel_6397/AMP_IN pixel_6397/SF_IB
+ pixel_6397/PIX_OUT pixel_6397/CSA_VREF pixel
Xpixel_5652 pixel_5652/gring pixel_5652/VDD pixel_5652/GND pixel_5652/VREF pixel_5652/ROW_SEL
+ pixel_5652/NB1 pixel_5652/VBIAS pixel_5652/NB2 pixel_5652/AMP_IN pixel_5652/SF_IB
+ pixel_5652/PIX_OUT pixel_5652/CSA_VREF pixel
Xpixel_5663 pixel_5663/gring pixel_5663/VDD pixel_5663/GND pixel_5663/VREF pixel_5663/ROW_SEL
+ pixel_5663/NB1 pixel_5663/VBIAS pixel_5663/NB2 pixel_5663/AMP_IN pixel_5663/SF_IB
+ pixel_5663/PIX_OUT pixel_5663/CSA_VREF pixel
Xpixel_5674 pixel_5674/gring pixel_5674/VDD pixel_5674/GND pixel_5674/VREF pixel_5674/ROW_SEL
+ pixel_5674/NB1 pixel_5674/VBIAS pixel_5674/NB2 pixel_5674/AMP_IN pixel_5674/SF_IB
+ pixel_5674/PIX_OUT pixel_5674/CSA_VREF pixel
Xpixel_5685 pixel_5685/gring pixel_5685/VDD pixel_5685/GND pixel_5685/VREF pixel_5685/ROW_SEL
+ pixel_5685/NB1 pixel_5685/VBIAS pixel_5685/NB2 pixel_5685/AMP_IN pixel_5685/SF_IB
+ pixel_5685/PIX_OUT pixel_5685/CSA_VREF pixel
Xpixel_4940 pixel_4940/gring pixel_4940/VDD pixel_4940/GND pixel_4940/VREF pixel_4940/ROW_SEL
+ pixel_4940/NB1 pixel_4940/VBIAS pixel_4940/NB2 pixel_4940/AMP_IN pixel_4940/SF_IB
+ pixel_4940/PIX_OUT pixel_4940/CSA_VREF pixel
Xpixel_5696 pixel_5696/gring pixel_5696/VDD pixel_5696/GND pixel_5696/VREF pixel_5696/ROW_SEL
+ pixel_5696/NB1 pixel_5696/VBIAS pixel_5696/NB2 pixel_5696/AMP_IN pixel_5696/SF_IB
+ pixel_5696/PIX_OUT pixel_5696/CSA_VREF pixel
Xpixel_4951 pixel_4951/gring pixel_4951/VDD pixel_4951/GND pixel_4951/VREF pixel_4951/ROW_SEL
+ pixel_4951/NB1 pixel_4951/VBIAS pixel_4951/NB2 pixel_4951/AMP_IN pixel_4951/SF_IB
+ pixel_4951/PIX_OUT pixel_4951/CSA_VREF pixel
Xpixel_4962 pixel_4962/gring pixel_4962/VDD pixel_4962/GND pixel_4962/VREF pixel_4962/ROW_SEL
+ pixel_4962/NB1 pixel_4962/VBIAS pixel_4962/NB2 pixel_4962/AMP_IN pixel_4962/SF_IB
+ pixel_4962/PIX_OUT pixel_4962/CSA_VREF pixel
Xpixel_4973 pixel_4973/gring pixel_4973/VDD pixel_4973/GND pixel_4973/VREF pixel_4973/ROW_SEL
+ pixel_4973/NB1 pixel_4973/VBIAS pixel_4973/NB2 pixel_4973/AMP_IN pixel_4973/SF_IB
+ pixel_4973/PIX_OUT pixel_4973/CSA_VREF pixel
Xpixel_990 pixel_990/gring pixel_990/VDD pixel_990/GND pixel_990/VREF pixel_990/ROW_SEL
+ pixel_990/NB1 pixel_990/VBIAS pixel_990/NB2 pixel_990/AMP_IN pixel_990/SF_IB pixel_990/PIX_OUT
+ pixel_990/CSA_VREF pixel
Xpixel_4984 pixel_4984/gring pixel_4984/VDD pixel_4984/GND pixel_4984/VREF pixel_4984/ROW_SEL
+ pixel_4984/NB1 pixel_4984/VBIAS pixel_4984/NB2 pixel_4984/AMP_IN pixel_4984/SF_IB
+ pixel_4984/PIX_OUT pixel_4984/CSA_VREF pixel
Xpixel_4995 pixel_4995/gring pixel_4995/VDD pixel_4995/GND pixel_4995/VREF pixel_4995/ROW_SEL
+ pixel_4995/NB1 pixel_4995/VBIAS pixel_4995/NB2 pixel_4995/AMP_IN pixel_4995/SF_IB
+ pixel_4995/PIX_OUT pixel_4995/CSA_VREF pixel
Xpixel_9929 pixel_9929/gring pixel_9929/VDD pixel_9929/GND pixel_9929/VREF pixel_9929/ROW_SEL
+ pixel_9929/NB1 pixel_9929/VBIAS pixel_9929/NB2 pixel_9929/AMP_IN pixel_9929/SF_IB
+ pixel_9929/PIX_OUT pixel_9929/CSA_VREF pixel
Xpixel_9918 pixel_9918/gring pixel_9918/VDD pixel_9918/GND pixel_9918/VREF pixel_9918/ROW_SEL
+ pixel_9918/NB1 pixel_9918/VBIAS pixel_9918/NB2 pixel_9918/AMP_IN pixel_9918/SF_IB
+ pixel_9918/PIX_OUT pixel_9918/CSA_VREF pixel
Xpixel_9907 pixel_9907/gring pixel_9907/VDD pixel_9907/GND pixel_9907/VREF pixel_9907/ROW_SEL
+ pixel_9907/NB1 pixel_9907/VBIAS pixel_9907/NB2 pixel_9907/AMP_IN pixel_9907/SF_IB
+ pixel_9907/PIX_OUT pixel_9907/CSA_VREF pixel
Xpixel_231 pixel_231/gring pixel_231/VDD pixel_231/GND pixel_231/VREF pixel_231/ROW_SEL
+ pixel_231/NB1 pixel_231/VBIAS pixel_231/NB2 pixel_231/AMP_IN pixel_231/SF_IB pixel_231/PIX_OUT
+ pixel_231/CSA_VREF pixel
Xpixel_220 pixel_220/gring pixel_220/VDD pixel_220/GND pixel_220/VREF pixel_220/ROW_SEL
+ pixel_220/NB1 pixel_220/VBIAS pixel_220/NB2 pixel_220/AMP_IN pixel_220/SF_IB pixel_220/PIX_OUT
+ pixel_220/CSA_VREF pixel
Xpixel_4203 pixel_4203/gring pixel_4203/VDD pixel_4203/GND pixel_4203/VREF pixel_4203/ROW_SEL
+ pixel_4203/NB1 pixel_4203/VBIAS pixel_4203/NB2 pixel_4203/AMP_IN pixel_4203/SF_IB
+ pixel_4203/PIX_OUT pixel_4203/CSA_VREF pixel
Xpixel_4214 pixel_4214/gring pixel_4214/VDD pixel_4214/GND pixel_4214/VREF pixel_4214/ROW_SEL
+ pixel_4214/NB1 pixel_4214/VBIAS pixel_4214/NB2 pixel_4214/AMP_IN pixel_4214/SF_IB
+ pixel_4214/PIX_OUT pixel_4214/CSA_VREF pixel
Xpixel_4225 pixel_4225/gring pixel_4225/VDD pixel_4225/GND pixel_4225/VREF pixel_4225/ROW_SEL
+ pixel_4225/NB1 pixel_4225/VBIAS pixel_4225/NB2 pixel_4225/AMP_IN pixel_4225/SF_IB
+ pixel_4225/PIX_OUT pixel_4225/CSA_VREF pixel
Xpixel_4236 pixel_4236/gring pixel_4236/VDD pixel_4236/GND pixel_4236/VREF pixel_4236/ROW_SEL
+ pixel_4236/NB1 pixel_4236/VBIAS pixel_4236/NB2 pixel_4236/AMP_IN pixel_4236/SF_IB
+ pixel_4236/PIX_OUT pixel_4236/CSA_VREF pixel
Xpixel_264 pixel_264/gring pixel_264/VDD pixel_264/GND pixel_264/VREF pixel_264/ROW_SEL
+ pixel_264/NB1 pixel_264/VBIAS pixel_264/NB2 pixel_264/AMP_IN pixel_264/SF_IB pixel_264/PIX_OUT
+ pixel_264/CSA_VREF pixel
Xpixel_253 pixel_253/gring pixel_253/VDD pixel_253/GND pixel_253/VREF pixel_253/ROW_SEL
+ pixel_253/NB1 pixel_253/VBIAS pixel_253/NB2 pixel_253/AMP_IN pixel_253/SF_IB pixel_253/PIX_OUT
+ pixel_253/CSA_VREF pixel
Xpixel_242 pixel_242/gring pixel_242/VDD pixel_242/GND pixel_242/VREF pixel_242/ROW_SEL
+ pixel_242/NB1 pixel_242/VBIAS pixel_242/NB2 pixel_242/AMP_IN pixel_242/SF_IB pixel_242/PIX_OUT
+ pixel_242/CSA_VREF pixel
Xpixel_3524 pixel_3524/gring pixel_3524/VDD pixel_3524/GND pixel_3524/VREF pixel_3524/ROW_SEL
+ pixel_3524/NB1 pixel_3524/VBIAS pixel_3524/NB2 pixel_3524/AMP_IN pixel_3524/SF_IB
+ pixel_3524/PIX_OUT pixel_3524/CSA_VREF pixel
Xpixel_3513 pixel_3513/gring pixel_3513/VDD pixel_3513/GND pixel_3513/VREF pixel_3513/ROW_SEL
+ pixel_3513/NB1 pixel_3513/VBIAS pixel_3513/NB2 pixel_3513/AMP_IN pixel_3513/SF_IB
+ pixel_3513/PIX_OUT pixel_3513/CSA_VREF pixel
Xpixel_3502 pixel_3502/gring pixel_3502/VDD pixel_3502/GND pixel_3502/VREF pixel_3502/ROW_SEL
+ pixel_3502/NB1 pixel_3502/VBIAS pixel_3502/NB2 pixel_3502/AMP_IN pixel_3502/SF_IB
+ pixel_3502/PIX_OUT pixel_3502/CSA_VREF pixel
Xpixel_4247 pixel_4247/gring pixel_4247/VDD pixel_4247/GND pixel_4247/VREF pixel_4247/ROW_SEL
+ pixel_4247/NB1 pixel_4247/VBIAS pixel_4247/NB2 pixel_4247/AMP_IN pixel_4247/SF_IB
+ pixel_4247/PIX_OUT pixel_4247/CSA_VREF pixel
Xpixel_4258 pixel_4258/gring pixel_4258/VDD pixel_4258/GND pixel_4258/VREF pixel_4258/ROW_SEL
+ pixel_4258/NB1 pixel_4258/VBIAS pixel_4258/NB2 pixel_4258/AMP_IN pixel_4258/SF_IB
+ pixel_4258/PIX_OUT pixel_4258/CSA_VREF pixel
Xpixel_4269 pixel_4269/gring pixel_4269/VDD pixel_4269/GND pixel_4269/VREF pixel_4269/ROW_SEL
+ pixel_4269/NB1 pixel_4269/VBIAS pixel_4269/NB2 pixel_4269/AMP_IN pixel_4269/SF_IB
+ pixel_4269/PIX_OUT pixel_4269/CSA_VREF pixel
Xpixel_297 pixel_297/gring pixel_297/VDD pixel_297/GND pixel_297/VREF pixel_297/ROW_SEL
+ pixel_297/NB1 pixel_297/VBIAS pixel_297/NB2 pixel_297/AMP_IN pixel_297/SF_IB pixel_297/PIX_OUT
+ pixel_297/CSA_VREF pixel
Xpixel_286 pixel_286/gring pixel_286/VDD pixel_286/GND pixel_286/VREF pixel_286/ROW_SEL
+ pixel_286/NB1 pixel_286/VBIAS pixel_286/NB2 pixel_286/AMP_IN pixel_286/SF_IB pixel_286/PIX_OUT
+ pixel_286/CSA_VREF pixel
Xpixel_275 pixel_275/gring pixel_275/VDD pixel_275/GND pixel_275/VREF pixel_275/ROW_SEL
+ pixel_275/NB1 pixel_275/VBIAS pixel_275/NB2 pixel_275/AMP_IN pixel_275/SF_IB pixel_275/PIX_OUT
+ pixel_275/CSA_VREF pixel
Xpixel_2812 pixel_2812/gring pixel_2812/VDD pixel_2812/GND pixel_2812/VREF pixel_2812/ROW_SEL
+ pixel_2812/NB1 pixel_2812/VBIAS pixel_2812/NB2 pixel_2812/AMP_IN pixel_2812/SF_IB
+ pixel_2812/PIX_OUT pixel_2812/CSA_VREF pixel
Xpixel_2801 pixel_2801/gring pixel_2801/VDD pixel_2801/GND pixel_2801/VREF pixel_2801/ROW_SEL
+ pixel_2801/NB1 pixel_2801/VBIAS pixel_2801/NB2 pixel_2801/AMP_IN pixel_2801/SF_IB
+ pixel_2801/PIX_OUT pixel_2801/CSA_VREF pixel
Xpixel_3557 pixel_3557/gring pixel_3557/VDD pixel_3557/GND pixel_3557/VREF pixel_3557/ROW_SEL
+ pixel_3557/NB1 pixel_3557/VBIAS pixel_3557/NB2 pixel_3557/AMP_IN pixel_3557/SF_IB
+ pixel_3557/PIX_OUT pixel_3557/CSA_VREF pixel
Xpixel_3546 pixel_3546/gring pixel_3546/VDD pixel_3546/GND pixel_3546/VREF pixel_3546/ROW_SEL
+ pixel_3546/NB1 pixel_3546/VBIAS pixel_3546/NB2 pixel_3546/AMP_IN pixel_3546/SF_IB
+ pixel_3546/PIX_OUT pixel_3546/CSA_VREF pixel
Xpixel_3535 pixel_3535/gring pixel_3535/VDD pixel_3535/GND pixel_3535/VREF pixel_3535/ROW_SEL
+ pixel_3535/NB1 pixel_3535/VBIAS pixel_3535/NB2 pixel_3535/AMP_IN pixel_3535/SF_IB
+ pixel_3535/PIX_OUT pixel_3535/CSA_VREF pixel
Xpixel_2856 pixel_2856/gring pixel_2856/VDD pixel_2856/GND pixel_2856/VREF pixel_2856/ROW_SEL
+ pixel_2856/NB1 pixel_2856/VBIAS pixel_2856/NB2 pixel_2856/AMP_IN pixel_2856/SF_IB
+ pixel_2856/PIX_OUT pixel_2856/CSA_VREF pixel
Xpixel_2845 pixel_2845/gring pixel_2845/VDD pixel_2845/GND pixel_2845/VREF pixel_2845/ROW_SEL
+ pixel_2845/NB1 pixel_2845/VBIAS pixel_2845/NB2 pixel_2845/AMP_IN pixel_2845/SF_IB
+ pixel_2845/PIX_OUT pixel_2845/CSA_VREF pixel
Xpixel_2834 pixel_2834/gring pixel_2834/VDD pixel_2834/GND pixel_2834/VREF pixel_2834/ROW_SEL
+ pixel_2834/NB1 pixel_2834/VBIAS pixel_2834/NB2 pixel_2834/AMP_IN pixel_2834/SF_IB
+ pixel_2834/PIX_OUT pixel_2834/CSA_VREF pixel
Xpixel_2823 pixel_2823/gring pixel_2823/VDD pixel_2823/GND pixel_2823/VREF pixel_2823/ROW_SEL
+ pixel_2823/NB1 pixel_2823/VBIAS pixel_2823/NB2 pixel_2823/AMP_IN pixel_2823/SF_IB
+ pixel_2823/PIX_OUT pixel_2823/CSA_VREF pixel
Xpixel_3579 pixel_3579/gring pixel_3579/VDD pixel_3579/GND pixel_3579/VREF pixel_3579/ROW_SEL
+ pixel_3579/NB1 pixel_3579/VBIAS pixel_3579/NB2 pixel_3579/AMP_IN pixel_3579/SF_IB
+ pixel_3579/PIX_OUT pixel_3579/CSA_VREF pixel
Xpixel_3568 pixel_3568/gring pixel_3568/VDD pixel_3568/GND pixel_3568/VREF pixel_3568/ROW_SEL
+ pixel_3568/NB1 pixel_3568/VBIAS pixel_3568/NB2 pixel_3568/AMP_IN pixel_3568/SF_IB
+ pixel_3568/PIX_OUT pixel_3568/CSA_VREF pixel
Xpixel_2889 pixel_2889/gring pixel_2889/VDD pixel_2889/GND pixel_2889/VREF pixel_2889/ROW_SEL
+ pixel_2889/NB1 pixel_2889/VBIAS pixel_2889/NB2 pixel_2889/AMP_IN pixel_2889/SF_IB
+ pixel_2889/PIX_OUT pixel_2889/CSA_VREF pixel
Xpixel_2878 pixel_2878/gring pixel_2878/VDD pixel_2878/GND pixel_2878/VREF pixel_2878/ROW_SEL
+ pixel_2878/NB1 pixel_2878/VBIAS pixel_2878/NB2 pixel_2878/AMP_IN pixel_2878/SF_IB
+ pixel_2878/PIX_OUT pixel_2878/CSA_VREF pixel
Xpixel_2867 pixel_2867/gring pixel_2867/VDD pixel_2867/GND pixel_2867/VREF pixel_2867/ROW_SEL
+ pixel_2867/NB1 pixel_2867/VBIAS pixel_2867/NB2 pixel_2867/AMP_IN pixel_2867/SF_IB
+ pixel_2867/PIX_OUT pixel_2867/CSA_VREF pixel
Xpixel_6150 pixel_6150/gring pixel_6150/VDD pixel_6150/GND pixel_6150/VREF pixel_6150/ROW_SEL
+ pixel_6150/NB1 pixel_6150/VBIAS pixel_6150/NB2 pixel_6150/AMP_IN pixel_6150/SF_IB
+ pixel_6150/PIX_OUT pixel_6150/CSA_VREF pixel
Xpixel_6161 pixel_6161/gring pixel_6161/VDD pixel_6161/GND pixel_6161/VREF pixel_6161/ROW_SEL
+ pixel_6161/NB1 pixel_6161/VBIAS pixel_6161/NB2 pixel_6161/AMP_IN pixel_6161/SF_IB
+ pixel_6161/PIX_OUT pixel_6161/CSA_VREF pixel
Xpixel_6172 pixel_6172/gring pixel_6172/VDD pixel_6172/GND pixel_6172/VREF pixel_6172/ROW_SEL
+ pixel_6172/NB1 pixel_6172/VBIAS pixel_6172/NB2 pixel_6172/AMP_IN pixel_6172/SF_IB
+ pixel_6172/PIX_OUT pixel_6172/CSA_VREF pixel
Xpixel_6183 pixel_6183/gring pixel_6183/VDD pixel_6183/GND pixel_6183/VREF pixel_6183/ROW_SEL
+ pixel_6183/NB1 pixel_6183/VBIAS pixel_6183/NB2 pixel_6183/AMP_IN pixel_6183/SF_IB
+ pixel_6183/PIX_OUT pixel_6183/CSA_VREF pixel
Xpixel_6194 pixel_6194/gring pixel_6194/VDD pixel_6194/GND pixel_6194/VREF pixel_6194/ROW_SEL
+ pixel_6194/NB1 pixel_6194/VBIAS pixel_6194/NB2 pixel_6194/AMP_IN pixel_6194/SF_IB
+ pixel_6194/PIX_OUT pixel_6194/CSA_VREF pixel
Xpixel_5460 pixel_5460/gring pixel_5460/VDD pixel_5460/GND pixel_5460/VREF pixel_5460/ROW_SEL
+ pixel_5460/NB1 pixel_5460/VBIAS pixel_5460/NB2 pixel_5460/AMP_IN pixel_5460/SF_IB
+ pixel_5460/PIX_OUT pixel_5460/CSA_VREF pixel
Xpixel_5471 pixel_5471/gring pixel_5471/VDD pixel_5471/GND pixel_5471/VREF pixel_5471/ROW_SEL
+ pixel_5471/NB1 pixel_5471/VBIAS pixel_5471/NB2 pixel_5471/AMP_IN pixel_5471/SF_IB
+ pixel_5471/PIX_OUT pixel_5471/CSA_VREF pixel
Xpixel_5482 pixel_5482/gring pixel_5482/VDD pixel_5482/GND pixel_5482/VREF pixel_5482/ROW_SEL
+ pixel_5482/NB1 pixel_5482/VBIAS pixel_5482/NB2 pixel_5482/AMP_IN pixel_5482/SF_IB
+ pixel_5482/PIX_OUT pixel_5482/CSA_VREF pixel
Xpixel_5493 pixel_5493/gring pixel_5493/VDD pixel_5493/GND pixel_5493/VREF pixel_5493/ROW_SEL
+ pixel_5493/NB1 pixel_5493/VBIAS pixel_5493/NB2 pixel_5493/AMP_IN pixel_5493/SF_IB
+ pixel_5493/PIX_OUT pixel_5493/CSA_VREF pixel
Xpixel_4770 pixel_4770/gring pixel_4770/VDD pixel_4770/GND pixel_4770/VREF pixel_4770/ROW_SEL
+ pixel_4770/NB1 pixel_4770/VBIAS pixel_4770/NB2 pixel_4770/AMP_IN pixel_4770/SF_IB
+ pixel_4770/PIX_OUT pixel_4770/CSA_VREF pixel
Xpixel_4781 pixel_4781/gring pixel_4781/VDD pixel_4781/GND pixel_4781/VREF pixel_4781/ROW_SEL
+ pixel_4781/NB1 pixel_4781/VBIAS pixel_4781/NB2 pixel_4781/AMP_IN pixel_4781/SF_IB
+ pixel_4781/PIX_OUT pixel_4781/CSA_VREF pixel
Xpixel_4792 pixel_4792/gring pixel_4792/VDD pixel_4792/GND pixel_4792/VREF pixel_4792/ROW_SEL
+ pixel_4792/NB1 pixel_4792/VBIAS pixel_4792/NB2 pixel_4792/AMP_IN pixel_4792/SF_IB
+ pixel_4792/PIX_OUT pixel_4792/CSA_VREF pixel
Xpixel_2108 pixel_2108/gring pixel_2108/VDD pixel_2108/GND pixel_2108/VREF pixel_2108/ROW_SEL
+ pixel_2108/NB1 pixel_2108/VBIAS pixel_2108/NB2 pixel_2108/AMP_IN pixel_2108/SF_IB
+ pixel_2108/PIX_OUT pixel_2108/CSA_VREF pixel
Xpixel_1407 pixel_1407/gring pixel_1407/VDD pixel_1407/GND pixel_1407/VREF pixel_1407/ROW_SEL
+ pixel_1407/NB1 pixel_1407/VBIAS pixel_1407/NB2 pixel_1407/AMP_IN pixel_1407/SF_IB
+ pixel_1407/PIX_OUT pixel_1407/CSA_VREF pixel
Xpixel_2119 pixel_2119/gring pixel_2119/VDD pixel_2119/GND pixel_2119/VREF pixel_2119/ROW_SEL
+ pixel_2119/NB1 pixel_2119/VBIAS pixel_2119/NB2 pixel_2119/AMP_IN pixel_2119/SF_IB
+ pixel_2119/PIX_OUT pixel_2119/CSA_VREF pixel
Xpixel_1429 pixel_1429/gring pixel_1429/VDD pixel_1429/GND pixel_1429/VREF pixel_1429/ROW_SEL
+ pixel_1429/NB1 pixel_1429/VBIAS pixel_1429/NB2 pixel_1429/AMP_IN pixel_1429/SF_IB
+ pixel_1429/PIX_OUT pixel_1429/CSA_VREF pixel
Xpixel_1418 pixel_1418/gring pixel_1418/VDD pixel_1418/GND pixel_1418/VREF pixel_1418/ROW_SEL
+ pixel_1418/NB1 pixel_1418/VBIAS pixel_1418/NB2 pixel_1418/AMP_IN pixel_1418/SF_IB
+ pixel_1418/PIX_OUT pixel_1418/CSA_VREF pixel
Xpixel_9704 pixel_9704/gring pixel_9704/VDD pixel_9704/GND pixel_9704/VREF pixel_9704/ROW_SEL
+ pixel_9704/NB1 pixel_9704/VBIAS pixel_9704/NB2 pixel_9704/AMP_IN pixel_9704/SF_IB
+ pixel_9704/PIX_OUT pixel_9704/CSA_VREF pixel
Xpixel_9715 pixel_9715/gring pixel_9715/VDD pixel_9715/GND pixel_9715/VREF pixel_9715/ROW_SEL
+ pixel_9715/NB1 pixel_9715/VBIAS pixel_9715/NB2 pixel_9715/AMP_IN pixel_9715/SF_IB
+ pixel_9715/PIX_OUT pixel_9715/CSA_VREF pixel
Xpixel_9726 pixel_9726/gring pixel_9726/VDD pixel_9726/GND pixel_9726/VREF pixel_9726/ROW_SEL
+ pixel_9726/NB1 pixel_9726/VBIAS pixel_9726/NB2 pixel_9726/AMP_IN pixel_9726/SF_IB
+ pixel_9726/PIX_OUT pixel_9726/CSA_VREF pixel
Xpixel_9737 pixel_9737/gring pixel_9737/VDD pixel_9737/GND pixel_9737/VREF pixel_9737/ROW_SEL
+ pixel_9737/NB1 pixel_9737/VBIAS pixel_9737/NB2 pixel_9737/AMP_IN pixel_9737/SF_IB
+ pixel_9737/PIX_OUT pixel_9737/CSA_VREF pixel
Xpixel_9748 pixel_9748/gring pixel_9748/VDD pixel_9748/GND pixel_9748/VREF pixel_9748/ROW_SEL
+ pixel_9748/NB1 pixel_9748/VBIAS pixel_9748/NB2 pixel_9748/AMP_IN pixel_9748/SF_IB
+ pixel_9748/PIX_OUT pixel_9748/CSA_VREF pixel
Xpixel_9759 pixel_9759/gring pixel_9759/VDD pixel_9759/GND pixel_9759/VREF pixel_9759/ROW_SEL
+ pixel_9759/NB1 pixel_9759/VBIAS pixel_9759/NB2 pixel_9759/AMP_IN pixel_9759/SF_IB
+ pixel_9759/PIX_OUT pixel_9759/CSA_VREF pixel
Xpixel_4000 pixel_4000/gring pixel_4000/VDD pixel_4000/GND pixel_4000/VREF pixel_4000/ROW_SEL
+ pixel_4000/NB1 pixel_4000/VBIAS pixel_4000/NB2 pixel_4000/AMP_IN pixel_4000/SF_IB
+ pixel_4000/PIX_OUT pixel_4000/CSA_VREF pixel
Xpixel_4011 pixel_4011/gring pixel_4011/VDD pixel_4011/GND pixel_4011/VREF pixel_4011/ROW_SEL
+ pixel_4011/NB1 pixel_4011/VBIAS pixel_4011/NB2 pixel_4011/AMP_IN pixel_4011/SF_IB
+ pixel_4011/PIX_OUT pixel_4011/CSA_VREF pixel
Xpixel_4022 pixel_4022/gring pixel_4022/VDD pixel_4022/GND pixel_4022/VREF pixel_4022/ROW_SEL
+ pixel_4022/NB1 pixel_4022/VBIAS pixel_4022/NB2 pixel_4022/AMP_IN pixel_4022/SF_IB
+ pixel_4022/PIX_OUT pixel_4022/CSA_VREF pixel
Xpixel_4033 pixel_4033/gring pixel_4033/VDD pixel_4033/GND pixel_4033/VREF pixel_4033/ROW_SEL
+ pixel_4033/NB1 pixel_4033/VBIAS pixel_4033/NB2 pixel_4033/AMP_IN pixel_4033/SF_IB
+ pixel_4033/PIX_OUT pixel_4033/CSA_VREF pixel
Xpixel_4044 pixel_4044/gring pixel_4044/VDD pixel_4044/GND pixel_4044/VREF pixel_4044/ROW_SEL
+ pixel_4044/NB1 pixel_4044/VBIAS pixel_4044/NB2 pixel_4044/AMP_IN pixel_4044/SF_IB
+ pixel_4044/PIX_OUT pixel_4044/CSA_VREF pixel
Xpixel_3332 pixel_3332/gring pixel_3332/VDD pixel_3332/GND pixel_3332/VREF pixel_3332/ROW_SEL
+ pixel_3332/NB1 pixel_3332/VBIAS pixel_3332/NB2 pixel_3332/AMP_IN pixel_3332/SF_IB
+ pixel_3332/PIX_OUT pixel_3332/CSA_VREF pixel
Xpixel_3321 pixel_3321/gring pixel_3321/VDD pixel_3321/GND pixel_3321/VREF pixel_3321/ROW_SEL
+ pixel_3321/NB1 pixel_3321/VBIAS pixel_3321/NB2 pixel_3321/AMP_IN pixel_3321/SF_IB
+ pixel_3321/PIX_OUT pixel_3321/CSA_VREF pixel
Xpixel_3310 pixel_3310/gring pixel_3310/VDD pixel_3310/GND pixel_3310/VREF pixel_3310/ROW_SEL
+ pixel_3310/NB1 pixel_3310/VBIAS pixel_3310/NB2 pixel_3310/AMP_IN pixel_3310/SF_IB
+ pixel_3310/PIX_OUT pixel_3310/CSA_VREF pixel
Xpixel_4055 pixel_4055/gring pixel_4055/VDD pixel_4055/GND pixel_4055/VREF pixel_4055/ROW_SEL
+ pixel_4055/NB1 pixel_4055/VBIAS pixel_4055/NB2 pixel_4055/AMP_IN pixel_4055/SF_IB
+ pixel_4055/PIX_OUT pixel_4055/CSA_VREF pixel
Xpixel_4066 pixel_4066/gring pixel_4066/VDD pixel_4066/GND pixel_4066/VREF pixel_4066/ROW_SEL
+ pixel_4066/NB1 pixel_4066/VBIAS pixel_4066/NB2 pixel_4066/AMP_IN pixel_4066/SF_IB
+ pixel_4066/PIX_OUT pixel_4066/CSA_VREF pixel
Xpixel_4077 pixel_4077/gring pixel_4077/VDD pixel_4077/GND pixel_4077/VREF pixel_4077/ROW_SEL
+ pixel_4077/NB1 pixel_4077/VBIAS pixel_4077/NB2 pixel_4077/AMP_IN pixel_4077/SF_IB
+ pixel_4077/PIX_OUT pixel_4077/CSA_VREF pixel
Xpixel_2631 pixel_2631/gring pixel_2631/VDD pixel_2631/GND pixel_2631/VREF pixel_2631/ROW_SEL
+ pixel_2631/NB1 pixel_2631/VBIAS pixel_2631/NB2 pixel_2631/AMP_IN pixel_2631/SF_IB
+ pixel_2631/PIX_OUT pixel_2631/CSA_VREF pixel
Xpixel_2620 pixel_2620/gring pixel_2620/VDD pixel_2620/GND pixel_2620/VREF pixel_2620/ROW_SEL
+ pixel_2620/NB1 pixel_2620/VBIAS pixel_2620/NB2 pixel_2620/AMP_IN pixel_2620/SF_IB
+ pixel_2620/PIX_OUT pixel_2620/CSA_VREF pixel
Xpixel_3376 pixel_3376/gring pixel_3376/VDD pixel_3376/GND pixel_3376/VREF pixel_3376/ROW_SEL
+ pixel_3376/NB1 pixel_3376/VBIAS pixel_3376/NB2 pixel_3376/AMP_IN pixel_3376/SF_IB
+ pixel_3376/PIX_OUT pixel_3376/CSA_VREF pixel
Xpixel_3365 pixel_3365/gring pixel_3365/VDD pixel_3365/GND pixel_3365/VREF pixel_3365/ROW_SEL
+ pixel_3365/NB1 pixel_3365/VBIAS pixel_3365/NB2 pixel_3365/AMP_IN pixel_3365/SF_IB
+ pixel_3365/PIX_OUT pixel_3365/CSA_VREF pixel
Xpixel_3354 pixel_3354/gring pixel_3354/VDD pixel_3354/GND pixel_3354/VREF pixel_3354/ROW_SEL
+ pixel_3354/NB1 pixel_3354/VBIAS pixel_3354/NB2 pixel_3354/AMP_IN pixel_3354/SF_IB
+ pixel_3354/PIX_OUT pixel_3354/CSA_VREF pixel
Xpixel_3343 pixel_3343/gring pixel_3343/VDD pixel_3343/GND pixel_3343/VREF pixel_3343/ROW_SEL
+ pixel_3343/NB1 pixel_3343/VBIAS pixel_3343/NB2 pixel_3343/AMP_IN pixel_3343/SF_IB
+ pixel_3343/PIX_OUT pixel_3343/CSA_VREF pixel
Xpixel_4088 pixel_4088/gring pixel_4088/VDD pixel_4088/GND pixel_4088/VREF pixel_4088/ROW_SEL
+ pixel_4088/NB1 pixel_4088/VBIAS pixel_4088/NB2 pixel_4088/AMP_IN pixel_4088/SF_IB
+ pixel_4088/PIX_OUT pixel_4088/CSA_VREF pixel
Xpixel_4099 pixel_4099/gring pixel_4099/VDD pixel_4099/GND pixel_4099/VREF pixel_4099/ROW_SEL
+ pixel_4099/NB1 pixel_4099/VBIAS pixel_4099/NB2 pixel_4099/AMP_IN pixel_4099/SF_IB
+ pixel_4099/PIX_OUT pixel_4099/CSA_VREF pixel
Xpixel_2664 pixel_2664/gring pixel_2664/VDD pixel_2664/GND pixel_2664/VREF pixel_2664/ROW_SEL
+ pixel_2664/NB1 pixel_2664/VBIAS pixel_2664/NB2 pixel_2664/AMP_IN pixel_2664/SF_IB
+ pixel_2664/PIX_OUT pixel_2664/CSA_VREF pixel
Xpixel_2653 pixel_2653/gring pixel_2653/VDD pixel_2653/GND pixel_2653/VREF pixel_2653/ROW_SEL
+ pixel_2653/NB1 pixel_2653/VBIAS pixel_2653/NB2 pixel_2653/AMP_IN pixel_2653/SF_IB
+ pixel_2653/PIX_OUT pixel_2653/CSA_VREF pixel
Xpixel_2642 pixel_2642/gring pixel_2642/VDD pixel_2642/GND pixel_2642/VREF pixel_2642/ROW_SEL
+ pixel_2642/NB1 pixel_2642/VBIAS pixel_2642/NB2 pixel_2642/AMP_IN pixel_2642/SF_IB
+ pixel_2642/PIX_OUT pixel_2642/CSA_VREF pixel
Xpixel_3398 pixel_3398/gring pixel_3398/VDD pixel_3398/GND pixel_3398/VREF pixel_3398/ROW_SEL
+ pixel_3398/NB1 pixel_3398/VBIAS pixel_3398/NB2 pixel_3398/AMP_IN pixel_3398/SF_IB
+ pixel_3398/PIX_OUT pixel_3398/CSA_VREF pixel
Xpixel_3387 pixel_3387/gring pixel_3387/VDD pixel_3387/GND pixel_3387/VREF pixel_3387/ROW_SEL
+ pixel_3387/NB1 pixel_3387/VBIAS pixel_3387/NB2 pixel_3387/AMP_IN pixel_3387/SF_IB
+ pixel_3387/PIX_OUT pixel_3387/CSA_VREF pixel
Xpixel_1952 pixel_1952/gring pixel_1952/VDD pixel_1952/GND pixel_1952/VREF pixel_1952/ROW_SEL
+ pixel_1952/NB1 pixel_1952/VBIAS pixel_1952/NB2 pixel_1952/AMP_IN pixel_1952/SF_IB
+ pixel_1952/PIX_OUT pixel_1952/CSA_VREF pixel
Xpixel_1941 pixel_1941/gring pixel_1941/VDD pixel_1941/GND pixel_1941/VREF pixel_1941/ROW_SEL
+ pixel_1941/NB1 pixel_1941/VBIAS pixel_1941/NB2 pixel_1941/AMP_IN pixel_1941/SF_IB
+ pixel_1941/PIX_OUT pixel_1941/CSA_VREF pixel
Xpixel_1930 pixel_1930/gring pixel_1930/VDD pixel_1930/GND pixel_1930/VREF pixel_1930/ROW_SEL
+ pixel_1930/NB1 pixel_1930/VBIAS pixel_1930/NB2 pixel_1930/AMP_IN pixel_1930/SF_IB
+ pixel_1930/PIX_OUT pixel_1930/CSA_VREF pixel
Xpixel_2697 pixel_2697/gring pixel_2697/VDD pixel_2697/GND pixel_2697/VREF pixel_2697/ROW_SEL
+ pixel_2697/NB1 pixel_2697/VBIAS pixel_2697/NB2 pixel_2697/AMP_IN pixel_2697/SF_IB
+ pixel_2697/PIX_OUT pixel_2697/CSA_VREF pixel
Xpixel_2686 pixel_2686/gring pixel_2686/VDD pixel_2686/GND pixel_2686/VREF pixel_2686/ROW_SEL
+ pixel_2686/NB1 pixel_2686/VBIAS pixel_2686/NB2 pixel_2686/AMP_IN pixel_2686/SF_IB
+ pixel_2686/PIX_OUT pixel_2686/CSA_VREF pixel
Xpixel_2675 pixel_2675/gring pixel_2675/VDD pixel_2675/GND pixel_2675/VREF pixel_2675/ROW_SEL
+ pixel_2675/NB1 pixel_2675/VBIAS pixel_2675/NB2 pixel_2675/AMP_IN pixel_2675/SF_IB
+ pixel_2675/PIX_OUT pixel_2675/CSA_VREF pixel
Xpixel_1996 pixel_1996/gring pixel_1996/VDD pixel_1996/GND pixel_1996/VREF pixel_1996/ROW_SEL
+ pixel_1996/NB1 pixel_1996/VBIAS pixel_1996/NB2 pixel_1996/AMP_IN pixel_1996/SF_IB
+ pixel_1996/PIX_OUT pixel_1996/CSA_VREF pixel
Xpixel_1985 pixel_1985/gring pixel_1985/VDD pixel_1985/GND pixel_1985/VREF pixel_1985/ROW_SEL
+ pixel_1985/NB1 pixel_1985/VBIAS pixel_1985/NB2 pixel_1985/AMP_IN pixel_1985/SF_IB
+ pixel_1985/PIX_OUT pixel_1985/CSA_VREF pixel
Xpixel_1974 pixel_1974/gring pixel_1974/VDD pixel_1974/GND pixel_1974/VREF pixel_1974/ROW_SEL
+ pixel_1974/NB1 pixel_1974/VBIAS pixel_1974/NB2 pixel_1974/AMP_IN pixel_1974/SF_IB
+ pixel_1974/PIX_OUT pixel_1974/CSA_VREF pixel
Xpixel_1963 pixel_1963/gring pixel_1963/VDD pixel_1963/GND pixel_1963/VREF pixel_1963/ROW_SEL
+ pixel_1963/NB1 pixel_1963/VBIAS pixel_1963/NB2 pixel_1963/AMP_IN pixel_1963/SF_IB
+ pixel_1963/PIX_OUT pixel_1963/CSA_VREF pixel
Xpixel_5290 pixel_5290/gring pixel_5290/VDD pixel_5290/GND pixel_5290/VREF pixel_5290/ROW_SEL
+ pixel_5290/NB1 pixel_5290/VBIAS pixel_5290/NB2 pixel_5290/AMP_IN pixel_5290/SF_IB
+ pixel_5290/PIX_OUT pixel_5290/CSA_VREF pixel
Xpixel_7609 pixel_7609/gring pixel_7609/VDD pixel_7609/GND pixel_7609/VREF pixel_7609/ROW_SEL
+ pixel_7609/NB1 pixel_7609/VBIAS pixel_7609/NB2 pixel_7609/AMP_IN pixel_7609/SF_IB
+ pixel_7609/PIX_OUT pixel_7609/CSA_VREF pixel
Xpixel_6908 pixel_6908/gring pixel_6908/VDD pixel_6908/GND pixel_6908/VREF pixel_6908/ROW_SEL
+ pixel_6908/NB1 pixel_6908/VBIAS pixel_6908/NB2 pixel_6908/AMP_IN pixel_6908/SF_IB
+ pixel_6908/PIX_OUT pixel_6908/CSA_VREF pixel
Xpixel_6919 pixel_6919/gring pixel_6919/VDD pixel_6919/GND pixel_6919/VREF pixel_6919/ROW_SEL
+ pixel_6919/NB1 pixel_6919/VBIAS pixel_6919/NB2 pixel_6919/AMP_IN pixel_6919/SF_IB
+ pixel_6919/PIX_OUT pixel_6919/CSA_VREF pixel
Xpixel_1215 pixel_1215/gring pixel_1215/VDD pixel_1215/GND pixel_1215/VREF pixel_1215/ROW_SEL
+ pixel_1215/NB1 pixel_1215/VBIAS pixel_1215/NB2 pixel_1215/AMP_IN pixel_1215/SF_IB
+ pixel_1215/PIX_OUT pixel_1215/CSA_VREF pixel
Xpixel_1204 pixel_1204/gring pixel_1204/VDD pixel_1204/GND pixel_1204/VREF pixel_1204/ROW_SEL
+ pixel_1204/NB1 pixel_1204/VBIAS pixel_1204/NB2 pixel_1204/AMP_IN pixel_1204/SF_IB
+ pixel_1204/PIX_OUT pixel_1204/CSA_VREF pixel
Xpixel_1248 pixel_1248/gring pixel_1248/VDD pixel_1248/GND pixel_1248/VREF pixel_1248/ROW_SEL
+ pixel_1248/NB1 pixel_1248/VBIAS pixel_1248/NB2 pixel_1248/AMP_IN pixel_1248/SF_IB
+ pixel_1248/PIX_OUT pixel_1248/CSA_VREF pixel
Xpixel_1237 pixel_1237/gring pixel_1237/VDD pixel_1237/GND pixel_1237/VREF pixel_1237/ROW_SEL
+ pixel_1237/NB1 pixel_1237/VBIAS pixel_1237/NB2 pixel_1237/AMP_IN pixel_1237/SF_IB
+ pixel_1237/PIX_OUT pixel_1237/CSA_VREF pixel
Xpixel_1226 pixel_1226/gring pixel_1226/VDD pixel_1226/GND pixel_1226/VREF pixel_1226/ROW_SEL
+ pixel_1226/NB1 pixel_1226/VBIAS pixel_1226/NB2 pixel_1226/AMP_IN pixel_1226/SF_IB
+ pixel_1226/PIX_OUT pixel_1226/CSA_VREF pixel
Xpixel_1259 pixel_1259/gring pixel_1259/VDD pixel_1259/GND pixel_1259/VREF pixel_1259/ROW_SEL
+ pixel_1259/NB1 pixel_1259/VBIAS pixel_1259/NB2 pixel_1259/AMP_IN pixel_1259/SF_IB
+ pixel_1259/PIX_OUT pixel_1259/CSA_VREF pixel
Xpixel_9523 pixel_9523/gring pixel_9523/VDD pixel_9523/GND pixel_9523/VREF pixel_9523/ROW_SEL
+ pixel_9523/NB1 pixel_9523/VBIAS pixel_9523/NB2 pixel_9523/AMP_IN pixel_9523/SF_IB
+ pixel_9523/PIX_OUT pixel_9523/CSA_VREF pixel
Xpixel_9512 pixel_9512/gring pixel_9512/VDD pixel_9512/GND pixel_9512/VREF pixel_9512/ROW_SEL
+ pixel_9512/NB1 pixel_9512/VBIAS pixel_9512/NB2 pixel_9512/AMP_IN pixel_9512/SF_IB
+ pixel_9512/PIX_OUT pixel_9512/CSA_VREF pixel
Xpixel_9501 pixel_9501/gring pixel_9501/VDD pixel_9501/GND pixel_9501/VREF pixel_9501/ROW_SEL
+ pixel_9501/NB1 pixel_9501/VBIAS pixel_9501/NB2 pixel_9501/AMP_IN pixel_9501/SF_IB
+ pixel_9501/PIX_OUT pixel_9501/CSA_VREF pixel
Xpixel_8811 pixel_8811/gring pixel_8811/VDD pixel_8811/GND pixel_8811/VREF pixel_8811/ROW_SEL
+ pixel_8811/NB1 pixel_8811/VBIAS pixel_8811/NB2 pixel_8811/AMP_IN pixel_8811/SF_IB
+ pixel_8811/PIX_OUT pixel_8811/CSA_VREF pixel
Xpixel_8800 pixel_8800/gring pixel_8800/VDD pixel_8800/GND pixel_8800/VREF pixel_8800/ROW_SEL
+ pixel_8800/NB1 pixel_8800/VBIAS pixel_8800/NB2 pixel_8800/AMP_IN pixel_8800/SF_IB
+ pixel_8800/PIX_OUT pixel_8800/CSA_VREF pixel
Xpixel_9556 pixel_9556/gring pixel_9556/VDD pixel_9556/GND pixel_9556/VREF pixel_9556/ROW_SEL
+ pixel_9556/NB1 pixel_9556/VBIAS pixel_9556/NB2 pixel_9556/AMP_IN pixel_9556/SF_IB
+ pixel_9556/PIX_OUT pixel_9556/CSA_VREF pixel
Xpixel_9545 pixel_9545/gring pixel_9545/VDD pixel_9545/GND pixel_9545/VREF pixel_9545/ROW_SEL
+ pixel_9545/NB1 pixel_9545/VBIAS pixel_9545/NB2 pixel_9545/AMP_IN pixel_9545/SF_IB
+ pixel_9545/PIX_OUT pixel_9545/CSA_VREF pixel
Xpixel_9534 pixel_9534/gring pixel_9534/VDD pixel_9534/GND pixel_9534/VREF pixel_9534/ROW_SEL
+ pixel_9534/NB1 pixel_9534/VBIAS pixel_9534/NB2 pixel_9534/AMP_IN pixel_9534/SF_IB
+ pixel_9534/PIX_OUT pixel_9534/CSA_VREF pixel
Xpixel_8855 pixel_8855/gring pixel_8855/VDD pixel_8855/GND pixel_8855/VREF pixel_8855/ROW_SEL
+ pixel_8855/NB1 pixel_8855/VBIAS pixel_8855/NB2 pixel_8855/AMP_IN pixel_8855/SF_IB
+ pixel_8855/PIX_OUT pixel_8855/CSA_VREF pixel
Xpixel_8844 pixel_8844/gring pixel_8844/VDD pixel_8844/GND pixel_8844/VREF pixel_8844/ROW_SEL
+ pixel_8844/NB1 pixel_8844/VBIAS pixel_8844/NB2 pixel_8844/AMP_IN pixel_8844/SF_IB
+ pixel_8844/PIX_OUT pixel_8844/CSA_VREF pixel
Xpixel_8833 pixel_8833/gring pixel_8833/VDD pixel_8833/GND pixel_8833/VREF pixel_8833/ROW_SEL
+ pixel_8833/NB1 pixel_8833/VBIAS pixel_8833/NB2 pixel_8833/AMP_IN pixel_8833/SF_IB
+ pixel_8833/PIX_OUT pixel_8833/CSA_VREF pixel
Xpixel_8822 pixel_8822/gring pixel_8822/VDD pixel_8822/GND pixel_8822/VREF pixel_8822/ROW_SEL
+ pixel_8822/NB1 pixel_8822/VBIAS pixel_8822/NB2 pixel_8822/AMP_IN pixel_8822/SF_IB
+ pixel_8822/PIX_OUT pixel_8822/CSA_VREF pixel
Xpixel_9589 pixel_9589/gring pixel_9589/VDD pixel_9589/GND pixel_9589/VREF pixel_9589/ROW_SEL
+ pixel_9589/NB1 pixel_9589/VBIAS pixel_9589/NB2 pixel_9589/AMP_IN pixel_9589/SF_IB
+ pixel_9589/PIX_OUT pixel_9589/CSA_VREF pixel
Xpixel_9578 pixel_9578/gring pixel_9578/VDD pixel_9578/GND pixel_9578/VREF pixel_9578/ROW_SEL
+ pixel_9578/NB1 pixel_9578/VBIAS pixel_9578/NB2 pixel_9578/AMP_IN pixel_9578/SF_IB
+ pixel_9578/PIX_OUT pixel_9578/CSA_VREF pixel
Xpixel_9567 pixel_9567/gring pixel_9567/VDD pixel_9567/GND pixel_9567/VREF pixel_9567/ROW_SEL
+ pixel_9567/NB1 pixel_9567/VBIAS pixel_9567/NB2 pixel_9567/AMP_IN pixel_9567/SF_IB
+ pixel_9567/PIX_OUT pixel_9567/CSA_VREF pixel
Xpixel_8888 pixel_8888/gring pixel_8888/VDD pixel_8888/GND pixel_8888/VREF pixel_8888/ROW_SEL
+ pixel_8888/NB1 pixel_8888/VBIAS pixel_8888/NB2 pixel_8888/AMP_IN pixel_8888/SF_IB
+ pixel_8888/PIX_OUT pixel_8888/CSA_VREF pixel
Xpixel_8877 pixel_8877/gring pixel_8877/VDD pixel_8877/GND pixel_8877/VREF pixel_8877/ROW_SEL
+ pixel_8877/NB1 pixel_8877/VBIAS pixel_8877/NB2 pixel_8877/AMP_IN pixel_8877/SF_IB
+ pixel_8877/PIX_OUT pixel_8877/CSA_VREF pixel
Xpixel_8866 pixel_8866/gring pixel_8866/VDD pixel_8866/GND pixel_8866/VREF pixel_8866/ROW_SEL
+ pixel_8866/NB1 pixel_8866/VBIAS pixel_8866/NB2 pixel_8866/AMP_IN pixel_8866/SF_IB
+ pixel_8866/PIX_OUT pixel_8866/CSA_VREF pixel
Xpixel_8899 pixel_8899/gring pixel_8899/VDD pixel_8899/GND pixel_8899/VREF pixel_8899/ROW_SEL
+ pixel_8899/NB1 pixel_8899/VBIAS pixel_8899/NB2 pixel_8899/AMP_IN pixel_8899/SF_IB
+ pixel_8899/PIX_OUT pixel_8899/CSA_VREF pixel
Xpixel_3140 pixel_3140/gring pixel_3140/VDD pixel_3140/GND pixel_3140/VREF pixel_3140/ROW_SEL
+ pixel_3140/NB1 pixel_3140/VBIAS pixel_3140/NB2 pixel_3140/AMP_IN pixel_3140/SF_IB
+ pixel_3140/PIX_OUT pixel_3140/CSA_VREF pixel
Xpixel_3184 pixel_3184/gring pixel_3184/VDD pixel_3184/GND pixel_3184/VREF pixel_3184/ROW_SEL
+ pixel_3184/NB1 pixel_3184/VBIAS pixel_3184/NB2 pixel_3184/AMP_IN pixel_3184/SF_IB
+ pixel_3184/PIX_OUT pixel_3184/CSA_VREF pixel
Xpixel_3173 pixel_3173/gring pixel_3173/VDD pixel_3173/GND pixel_3173/VREF pixel_3173/ROW_SEL
+ pixel_3173/NB1 pixel_3173/VBIAS pixel_3173/NB2 pixel_3173/AMP_IN pixel_3173/SF_IB
+ pixel_3173/PIX_OUT pixel_3173/CSA_VREF pixel
Xpixel_3162 pixel_3162/gring pixel_3162/VDD pixel_3162/GND pixel_3162/VREF pixel_3162/ROW_SEL
+ pixel_3162/NB1 pixel_3162/VBIAS pixel_3162/NB2 pixel_3162/AMP_IN pixel_3162/SF_IB
+ pixel_3162/PIX_OUT pixel_3162/CSA_VREF pixel
Xpixel_3151 pixel_3151/gring pixel_3151/VDD pixel_3151/GND pixel_3151/VREF pixel_3151/ROW_SEL
+ pixel_3151/NB1 pixel_3151/VBIAS pixel_3151/NB2 pixel_3151/AMP_IN pixel_3151/SF_IB
+ pixel_3151/PIX_OUT pixel_3151/CSA_VREF pixel
Xpixel_2472 pixel_2472/gring pixel_2472/VDD pixel_2472/GND pixel_2472/VREF pixel_2472/ROW_SEL
+ pixel_2472/NB1 pixel_2472/VBIAS pixel_2472/NB2 pixel_2472/AMP_IN pixel_2472/SF_IB
+ pixel_2472/PIX_OUT pixel_2472/CSA_VREF pixel
Xpixel_2461 pixel_2461/gring pixel_2461/VDD pixel_2461/GND pixel_2461/VREF pixel_2461/ROW_SEL
+ pixel_2461/NB1 pixel_2461/VBIAS pixel_2461/NB2 pixel_2461/AMP_IN pixel_2461/SF_IB
+ pixel_2461/PIX_OUT pixel_2461/CSA_VREF pixel
Xpixel_2450 pixel_2450/gring pixel_2450/VDD pixel_2450/GND pixel_2450/VREF pixel_2450/ROW_SEL
+ pixel_2450/NB1 pixel_2450/VBIAS pixel_2450/NB2 pixel_2450/AMP_IN pixel_2450/SF_IB
+ pixel_2450/PIX_OUT pixel_2450/CSA_VREF pixel
Xpixel_3195 pixel_3195/gring pixel_3195/VDD pixel_3195/GND pixel_3195/VREF pixel_3195/ROW_SEL
+ pixel_3195/NB1 pixel_3195/VBIAS pixel_3195/NB2 pixel_3195/AMP_IN pixel_3195/SF_IB
+ pixel_3195/PIX_OUT pixel_3195/CSA_VREF pixel
Xpixel_1771 pixel_1771/gring pixel_1771/VDD pixel_1771/GND pixel_1771/VREF pixel_1771/ROW_SEL
+ pixel_1771/NB1 pixel_1771/VBIAS pixel_1771/NB2 pixel_1771/AMP_IN pixel_1771/SF_IB
+ pixel_1771/PIX_OUT pixel_1771/CSA_VREF pixel
Xpixel_1760 pixel_1760/gring pixel_1760/VDD pixel_1760/GND pixel_1760/VREF pixel_1760/ROW_SEL
+ pixel_1760/NB1 pixel_1760/VBIAS pixel_1760/NB2 pixel_1760/AMP_IN pixel_1760/SF_IB
+ pixel_1760/PIX_OUT pixel_1760/CSA_VREF pixel
Xpixel_2494 pixel_2494/gring pixel_2494/VDD pixel_2494/GND pixel_2494/VREF pixel_2494/ROW_SEL
+ pixel_2494/NB1 pixel_2494/VBIAS pixel_2494/NB2 pixel_2494/AMP_IN pixel_2494/SF_IB
+ pixel_2494/PIX_OUT pixel_2494/CSA_VREF pixel
Xpixel_2483 pixel_2483/gring pixel_2483/VDD pixel_2483/GND pixel_2483/VREF pixel_2483/ROW_SEL
+ pixel_2483/NB1 pixel_2483/VBIAS pixel_2483/NB2 pixel_2483/AMP_IN pixel_2483/SF_IB
+ pixel_2483/PIX_OUT pixel_2483/CSA_VREF pixel
Xpixel_1793 pixel_1793/gring pixel_1793/VDD pixel_1793/GND pixel_1793/VREF pixel_1793/ROW_SEL
+ pixel_1793/NB1 pixel_1793/VBIAS pixel_1793/NB2 pixel_1793/AMP_IN pixel_1793/SF_IB
+ pixel_1793/PIX_OUT pixel_1793/CSA_VREF pixel
Xpixel_1782 pixel_1782/gring pixel_1782/VDD pixel_1782/GND pixel_1782/VREF pixel_1782/ROW_SEL
+ pixel_1782/NB1 pixel_1782/VBIAS pixel_1782/NB2 pixel_1782/AMP_IN pixel_1782/SF_IB
+ pixel_1782/PIX_OUT pixel_1782/CSA_VREF pixel
Xpixel_819 pixel_819/gring pixel_819/VDD pixel_819/GND pixel_819/VREF pixel_819/ROW_SEL
+ pixel_819/NB1 pixel_819/VBIAS pixel_819/NB2 pixel_819/AMP_IN pixel_819/SF_IB pixel_819/PIX_OUT
+ pixel_819/CSA_VREF pixel
Xpixel_808 pixel_808/gring pixel_808/VDD pixel_808/GND pixel_808/VREF pixel_808/ROW_SEL
+ pixel_808/NB1 pixel_808/VBIAS pixel_808/NB2 pixel_808/AMP_IN pixel_808/SF_IB pixel_808/PIX_OUT
+ pixel_808/CSA_VREF pixel
Xpixel_8107 pixel_8107/gring pixel_8107/VDD pixel_8107/GND pixel_8107/VREF pixel_8107/ROW_SEL
+ pixel_8107/NB1 pixel_8107/VBIAS pixel_8107/NB2 pixel_8107/AMP_IN pixel_8107/SF_IB
+ pixel_8107/PIX_OUT pixel_8107/CSA_VREF pixel
Xpixel_8118 pixel_8118/gring pixel_8118/VDD pixel_8118/GND pixel_8118/VREF pixel_8118/ROW_SEL
+ pixel_8118/NB1 pixel_8118/VBIAS pixel_8118/NB2 pixel_8118/AMP_IN pixel_8118/SF_IB
+ pixel_8118/PIX_OUT pixel_8118/CSA_VREF pixel
Xpixel_8129 pixel_8129/gring pixel_8129/VDD pixel_8129/GND pixel_8129/VREF pixel_8129/ROW_SEL
+ pixel_8129/NB1 pixel_8129/VBIAS pixel_8129/NB2 pixel_8129/AMP_IN pixel_8129/SF_IB
+ pixel_8129/PIX_OUT pixel_8129/CSA_VREF pixel
Xpixel_7406 pixel_7406/gring pixel_7406/VDD pixel_7406/GND pixel_7406/VREF pixel_7406/ROW_SEL
+ pixel_7406/NB1 pixel_7406/VBIAS pixel_7406/NB2 pixel_7406/AMP_IN pixel_7406/SF_IB
+ pixel_7406/PIX_OUT pixel_7406/CSA_VREF pixel
Xpixel_7417 pixel_7417/gring pixel_7417/VDD pixel_7417/GND pixel_7417/VREF pixel_7417/ROW_SEL
+ pixel_7417/NB1 pixel_7417/VBIAS pixel_7417/NB2 pixel_7417/AMP_IN pixel_7417/SF_IB
+ pixel_7417/PIX_OUT pixel_7417/CSA_VREF pixel
Xpixel_7428 pixel_7428/gring pixel_7428/VDD pixel_7428/GND pixel_7428/VREF pixel_7428/ROW_SEL
+ pixel_7428/NB1 pixel_7428/VBIAS pixel_7428/NB2 pixel_7428/AMP_IN pixel_7428/SF_IB
+ pixel_7428/PIX_OUT pixel_7428/CSA_VREF pixel
Xpixel_7439 pixel_7439/gring pixel_7439/VDD pixel_7439/GND pixel_7439/VREF pixel_7439/ROW_SEL
+ pixel_7439/NB1 pixel_7439/VBIAS pixel_7439/NB2 pixel_7439/AMP_IN pixel_7439/SF_IB
+ pixel_7439/PIX_OUT pixel_7439/CSA_VREF pixel
Xpixel_6705 pixel_6705/gring pixel_6705/VDD pixel_6705/GND pixel_6705/VREF pixel_6705/ROW_SEL
+ pixel_6705/NB1 pixel_6705/VBIAS pixel_6705/NB2 pixel_6705/AMP_IN pixel_6705/SF_IB
+ pixel_6705/PIX_OUT pixel_6705/CSA_VREF pixel
Xpixel_6716 pixel_6716/gring pixel_6716/VDD pixel_6716/GND pixel_6716/VREF pixel_6716/ROW_SEL
+ pixel_6716/NB1 pixel_6716/VBIAS pixel_6716/NB2 pixel_6716/AMP_IN pixel_6716/SF_IB
+ pixel_6716/PIX_OUT pixel_6716/CSA_VREF pixel
Xpixel_6727 pixel_6727/gring pixel_6727/VDD pixel_6727/GND pixel_6727/VREF pixel_6727/ROW_SEL
+ pixel_6727/NB1 pixel_6727/VBIAS pixel_6727/NB2 pixel_6727/AMP_IN pixel_6727/SF_IB
+ pixel_6727/PIX_OUT pixel_6727/CSA_VREF pixel
Xpixel_6738 pixel_6738/gring pixel_6738/VDD pixel_6738/GND pixel_6738/VREF pixel_6738/ROW_SEL
+ pixel_6738/NB1 pixel_6738/VBIAS pixel_6738/NB2 pixel_6738/AMP_IN pixel_6738/SF_IB
+ pixel_6738/PIX_OUT pixel_6738/CSA_VREF pixel
Xpixel_6749 pixel_6749/gring pixel_6749/VDD pixel_6749/GND pixel_6749/VREF pixel_6749/ROW_SEL
+ pixel_6749/NB1 pixel_6749/VBIAS pixel_6749/NB2 pixel_6749/AMP_IN pixel_6749/SF_IB
+ pixel_6749/PIX_OUT pixel_6749/CSA_VREF pixel
Xpixel_1023 pixel_1023/gring pixel_1023/VDD pixel_1023/GND pixel_1023/VREF pixel_1023/ROW_SEL
+ pixel_1023/NB1 pixel_1023/VBIAS pixel_1023/NB2 pixel_1023/AMP_IN pixel_1023/SF_IB
+ pixel_1023/PIX_OUT pixel_1023/CSA_VREF pixel
Xpixel_1012 pixel_1012/gring pixel_1012/VDD pixel_1012/GND pixel_1012/VREF pixel_1012/ROW_SEL
+ pixel_1012/NB1 pixel_1012/VBIAS pixel_1012/NB2 pixel_1012/AMP_IN pixel_1012/SF_IB
+ pixel_1012/PIX_OUT pixel_1012/CSA_VREF pixel
Xpixel_1001 pixel_1001/gring pixel_1001/VDD pixel_1001/GND pixel_1001/VREF pixel_1001/ROW_SEL
+ pixel_1001/NB1 pixel_1001/VBIAS pixel_1001/NB2 pixel_1001/AMP_IN pixel_1001/SF_IB
+ pixel_1001/PIX_OUT pixel_1001/CSA_VREF pixel
Xpixel_1056 pixel_1056/gring pixel_1056/VDD pixel_1056/GND pixel_1056/VREF pixel_1056/ROW_SEL
+ pixel_1056/NB1 pixel_1056/VBIAS pixel_1056/NB2 pixel_1056/AMP_IN pixel_1056/SF_IB
+ pixel_1056/PIX_OUT pixel_1056/CSA_VREF pixel
Xpixel_1045 pixel_1045/gring pixel_1045/VDD pixel_1045/GND pixel_1045/VREF pixel_1045/ROW_SEL
+ pixel_1045/NB1 pixel_1045/VBIAS pixel_1045/NB2 pixel_1045/AMP_IN pixel_1045/SF_IB
+ pixel_1045/PIX_OUT pixel_1045/CSA_VREF pixel
Xpixel_1034 pixel_1034/gring pixel_1034/VDD pixel_1034/GND pixel_1034/VREF pixel_1034/ROW_SEL
+ pixel_1034/NB1 pixel_1034/VBIAS pixel_1034/NB2 pixel_1034/AMP_IN pixel_1034/SF_IB
+ pixel_1034/PIX_OUT pixel_1034/CSA_VREF pixel
Xpixel_1089 pixel_1089/gring pixel_1089/VDD pixel_1089/GND pixel_1089/VREF pixel_1089/ROW_SEL
+ pixel_1089/NB1 pixel_1089/VBIAS pixel_1089/NB2 pixel_1089/AMP_IN pixel_1089/SF_IB
+ pixel_1089/PIX_OUT pixel_1089/CSA_VREF pixel
Xpixel_1078 pixel_1078/gring pixel_1078/VDD pixel_1078/GND pixel_1078/VREF pixel_1078/ROW_SEL
+ pixel_1078/NB1 pixel_1078/VBIAS pixel_1078/NB2 pixel_1078/AMP_IN pixel_1078/SF_IB
+ pixel_1078/PIX_OUT pixel_1078/CSA_VREF pixel
Xpixel_1067 pixel_1067/gring pixel_1067/VDD pixel_1067/GND pixel_1067/VREF pixel_1067/ROW_SEL
+ pixel_1067/NB1 pixel_1067/VBIAS pixel_1067/NB2 pixel_1067/AMP_IN pixel_1067/SF_IB
+ pixel_1067/PIX_OUT pixel_1067/CSA_VREF pixel
Xpixel_9331 pixel_9331/gring pixel_9331/VDD pixel_9331/GND pixel_9331/VREF pixel_9331/ROW_SEL
+ pixel_9331/NB1 pixel_9331/VBIAS pixel_9331/NB2 pixel_9331/AMP_IN pixel_9331/SF_IB
+ pixel_9331/PIX_OUT pixel_9331/CSA_VREF pixel
Xpixel_9320 pixel_9320/gring pixel_9320/VDD pixel_9320/GND pixel_9320/VREF pixel_9320/ROW_SEL
+ pixel_9320/NB1 pixel_9320/VBIAS pixel_9320/NB2 pixel_9320/AMP_IN pixel_9320/SF_IB
+ pixel_9320/PIX_OUT pixel_9320/CSA_VREF pixel
Xpixel_9364 pixel_9364/gring pixel_9364/VDD pixel_9364/GND pixel_9364/VREF pixel_9364/ROW_SEL
+ pixel_9364/NB1 pixel_9364/VBIAS pixel_9364/NB2 pixel_9364/AMP_IN pixel_9364/SF_IB
+ pixel_9364/PIX_OUT pixel_9364/CSA_VREF pixel
Xpixel_9353 pixel_9353/gring pixel_9353/VDD pixel_9353/GND pixel_9353/VREF pixel_9353/ROW_SEL
+ pixel_9353/NB1 pixel_9353/VBIAS pixel_9353/NB2 pixel_9353/AMP_IN pixel_9353/SF_IB
+ pixel_9353/PIX_OUT pixel_9353/CSA_VREF pixel
Xpixel_9342 pixel_9342/gring pixel_9342/VDD pixel_9342/GND pixel_9342/VREF pixel_9342/ROW_SEL
+ pixel_9342/NB1 pixel_9342/VBIAS pixel_9342/NB2 pixel_9342/AMP_IN pixel_9342/SF_IB
+ pixel_9342/PIX_OUT pixel_9342/CSA_VREF pixel
Xpixel_8663 pixel_8663/gring pixel_8663/VDD pixel_8663/GND pixel_8663/VREF pixel_8663/ROW_SEL
+ pixel_8663/NB1 pixel_8663/VBIAS pixel_8663/NB2 pixel_8663/AMP_IN pixel_8663/SF_IB
+ pixel_8663/PIX_OUT pixel_8663/CSA_VREF pixel
Xpixel_8652 pixel_8652/gring pixel_8652/VDD pixel_8652/GND pixel_8652/VREF pixel_8652/ROW_SEL
+ pixel_8652/NB1 pixel_8652/VBIAS pixel_8652/NB2 pixel_8652/AMP_IN pixel_8652/SF_IB
+ pixel_8652/PIX_OUT pixel_8652/CSA_VREF pixel
Xpixel_8641 pixel_8641/gring pixel_8641/VDD pixel_8641/GND pixel_8641/VREF pixel_8641/ROW_SEL
+ pixel_8641/NB1 pixel_8641/VBIAS pixel_8641/NB2 pixel_8641/AMP_IN pixel_8641/SF_IB
+ pixel_8641/PIX_OUT pixel_8641/CSA_VREF pixel
Xpixel_8630 pixel_8630/gring pixel_8630/VDD pixel_8630/GND pixel_8630/VREF pixel_8630/ROW_SEL
+ pixel_8630/NB1 pixel_8630/VBIAS pixel_8630/NB2 pixel_8630/AMP_IN pixel_8630/SF_IB
+ pixel_8630/PIX_OUT pixel_8630/CSA_VREF pixel
Xpixel_9397 pixel_9397/gring pixel_9397/VDD pixel_9397/GND pixel_9397/VREF pixel_9397/ROW_SEL
+ pixel_9397/NB1 pixel_9397/VBIAS pixel_9397/NB2 pixel_9397/AMP_IN pixel_9397/SF_IB
+ pixel_9397/PIX_OUT pixel_9397/CSA_VREF pixel
Xpixel_9386 pixel_9386/gring pixel_9386/VDD pixel_9386/GND pixel_9386/VREF pixel_9386/ROW_SEL
+ pixel_9386/NB1 pixel_9386/VBIAS pixel_9386/NB2 pixel_9386/AMP_IN pixel_9386/SF_IB
+ pixel_9386/PIX_OUT pixel_9386/CSA_VREF pixel
Xpixel_9375 pixel_9375/gring pixel_9375/VDD pixel_9375/GND pixel_9375/VREF pixel_9375/ROW_SEL
+ pixel_9375/NB1 pixel_9375/VBIAS pixel_9375/NB2 pixel_9375/AMP_IN pixel_9375/SF_IB
+ pixel_9375/PIX_OUT pixel_9375/CSA_VREF pixel
Xpixel_8696 pixel_8696/gring pixel_8696/VDD pixel_8696/GND pixel_8696/VREF pixel_8696/ROW_SEL
+ pixel_8696/NB1 pixel_8696/VBIAS pixel_8696/NB2 pixel_8696/AMP_IN pixel_8696/SF_IB
+ pixel_8696/PIX_OUT pixel_8696/CSA_VREF pixel
Xpixel_8685 pixel_8685/gring pixel_8685/VDD pixel_8685/GND pixel_8685/VREF pixel_8685/ROW_SEL
+ pixel_8685/NB1 pixel_8685/VBIAS pixel_8685/NB2 pixel_8685/AMP_IN pixel_8685/SF_IB
+ pixel_8685/PIX_OUT pixel_8685/CSA_VREF pixel
Xpixel_8674 pixel_8674/gring pixel_8674/VDD pixel_8674/GND pixel_8674/VREF pixel_8674/ROW_SEL
+ pixel_8674/NB1 pixel_8674/VBIAS pixel_8674/NB2 pixel_8674/AMP_IN pixel_8674/SF_IB
+ pixel_8674/PIX_OUT pixel_8674/CSA_VREF pixel
Xpixel_7940 pixel_7940/gring pixel_7940/VDD pixel_7940/GND pixel_7940/VREF pixel_7940/ROW_SEL
+ pixel_7940/NB1 pixel_7940/VBIAS pixel_7940/NB2 pixel_7940/AMP_IN pixel_7940/SF_IB
+ pixel_7940/PIX_OUT pixel_7940/CSA_VREF pixel
Xpixel_7951 pixel_7951/gring pixel_7951/VDD pixel_7951/GND pixel_7951/VREF pixel_7951/ROW_SEL
+ pixel_7951/NB1 pixel_7951/VBIAS pixel_7951/NB2 pixel_7951/AMP_IN pixel_7951/SF_IB
+ pixel_7951/PIX_OUT pixel_7951/CSA_VREF pixel
Xpixel_7962 pixel_7962/gring pixel_7962/VDD pixel_7962/GND pixel_7962/VREF pixel_7962/ROW_SEL
+ pixel_7962/NB1 pixel_7962/VBIAS pixel_7962/NB2 pixel_7962/AMP_IN pixel_7962/SF_IB
+ pixel_7962/PIX_OUT pixel_7962/CSA_VREF pixel
Xpixel_7973 pixel_7973/gring pixel_7973/VDD pixel_7973/GND pixel_7973/VREF pixel_7973/ROW_SEL
+ pixel_7973/NB1 pixel_7973/VBIAS pixel_7973/NB2 pixel_7973/AMP_IN pixel_7973/SF_IB
+ pixel_7973/PIX_OUT pixel_7973/CSA_VREF pixel
Xpixel_7984 pixel_7984/gring pixel_7984/VDD pixel_7984/GND pixel_7984/VREF pixel_7984/ROW_SEL
+ pixel_7984/NB1 pixel_7984/VBIAS pixel_7984/NB2 pixel_7984/AMP_IN pixel_7984/SF_IB
+ pixel_7984/PIX_OUT pixel_7984/CSA_VREF pixel
Xpixel_7995 pixel_7995/gring pixel_7995/VDD pixel_7995/GND pixel_7995/VREF pixel_7995/ROW_SEL
+ pixel_7995/NB1 pixel_7995/VBIAS pixel_7995/NB2 pixel_7995/AMP_IN pixel_7995/SF_IB
+ pixel_7995/PIX_OUT pixel_7995/CSA_VREF pixel
Xpixel_2280 pixel_2280/gring pixel_2280/VDD pixel_2280/GND pixel_2280/VREF pixel_2280/ROW_SEL
+ pixel_2280/NB1 pixel_2280/VBIAS pixel_2280/NB2 pixel_2280/AMP_IN pixel_2280/SF_IB
+ pixel_2280/PIX_OUT pixel_2280/CSA_VREF pixel
Xpixel_2291 pixel_2291/gring pixel_2291/VDD pixel_2291/GND pixel_2291/VREF pixel_2291/ROW_SEL
+ pixel_2291/NB1 pixel_2291/VBIAS pixel_2291/NB2 pixel_2291/AMP_IN pixel_2291/SF_IB
+ pixel_2291/PIX_OUT pixel_2291/CSA_VREF pixel
Xpixel_1590 pixel_1590/gring pixel_1590/VDD pixel_1590/GND pixel_1590/VREF pixel_1590/ROW_SEL
+ pixel_1590/NB1 pixel_1590/VBIAS pixel_1590/NB2 pixel_1590/AMP_IN pixel_1590/SF_IB
+ pixel_1590/PIX_OUT pixel_1590/CSA_VREF pixel
Xpixel_605 pixel_605/gring pixel_605/VDD pixel_605/GND pixel_605/VREF pixel_605/ROW_SEL
+ pixel_605/NB1 pixel_605/VBIAS pixel_605/NB2 pixel_605/AMP_IN pixel_605/SF_IB pixel_605/PIX_OUT
+ pixel_605/CSA_VREF pixel
Xpixel_638 pixel_638/gring pixel_638/VDD pixel_638/GND pixel_638/VREF pixel_638/ROW_SEL
+ pixel_638/NB1 pixel_638/VBIAS pixel_638/NB2 pixel_638/AMP_IN pixel_638/SF_IB pixel_638/PIX_OUT
+ pixel_638/CSA_VREF pixel
Xpixel_627 pixel_627/gring pixel_627/VDD pixel_627/GND pixel_627/VREF pixel_627/ROW_SEL
+ pixel_627/NB1 pixel_627/VBIAS pixel_627/NB2 pixel_627/AMP_IN pixel_627/SF_IB pixel_627/PIX_OUT
+ pixel_627/CSA_VREF pixel
Xpixel_616 pixel_616/gring pixel_616/VDD pixel_616/GND pixel_616/VREF pixel_616/ROW_SEL
+ pixel_616/NB1 pixel_616/VBIAS pixel_616/NB2 pixel_616/AMP_IN pixel_616/SF_IB pixel_616/PIX_OUT
+ pixel_616/CSA_VREF pixel
Xpixel_649 pixel_649/gring pixel_649/VDD pixel_649/GND pixel_649/VREF pixel_649/ROW_SEL
+ pixel_649/NB1 pixel_649/VBIAS pixel_649/NB2 pixel_649/AMP_IN pixel_649/SF_IB pixel_649/PIX_OUT
+ pixel_649/CSA_VREF pixel
Xpixel_3909 pixel_3909/gring pixel_3909/VDD pixel_3909/GND pixel_3909/VREF pixel_3909/ROW_SEL
+ pixel_3909/NB1 pixel_3909/VBIAS pixel_3909/NB2 pixel_3909/AMP_IN pixel_3909/SF_IB
+ pixel_3909/PIX_OUT pixel_3909/CSA_VREF pixel
Xpixel_7203 pixel_7203/gring pixel_7203/VDD pixel_7203/GND pixel_7203/VREF pixel_7203/ROW_SEL
+ pixel_7203/NB1 pixel_7203/VBIAS pixel_7203/NB2 pixel_7203/AMP_IN pixel_7203/SF_IB
+ pixel_7203/PIX_OUT pixel_7203/CSA_VREF pixel
Xpixel_7214 pixel_7214/gring pixel_7214/VDD pixel_7214/GND pixel_7214/VREF pixel_7214/ROW_SEL
+ pixel_7214/NB1 pixel_7214/VBIAS pixel_7214/NB2 pixel_7214/AMP_IN pixel_7214/SF_IB
+ pixel_7214/PIX_OUT pixel_7214/CSA_VREF pixel
Xpixel_7225 pixel_7225/gring pixel_7225/VDD pixel_7225/GND pixel_7225/VREF pixel_7225/ROW_SEL
+ pixel_7225/NB1 pixel_7225/VBIAS pixel_7225/NB2 pixel_7225/AMP_IN pixel_7225/SF_IB
+ pixel_7225/PIX_OUT pixel_7225/CSA_VREF pixel
Xpixel_7236 pixel_7236/gring pixel_7236/VDD pixel_7236/GND pixel_7236/VREF pixel_7236/ROW_SEL
+ pixel_7236/NB1 pixel_7236/VBIAS pixel_7236/NB2 pixel_7236/AMP_IN pixel_7236/SF_IB
+ pixel_7236/PIX_OUT pixel_7236/CSA_VREF pixel
Xpixel_7247 pixel_7247/gring pixel_7247/VDD pixel_7247/GND pixel_7247/VREF pixel_7247/ROW_SEL
+ pixel_7247/NB1 pixel_7247/VBIAS pixel_7247/NB2 pixel_7247/AMP_IN pixel_7247/SF_IB
+ pixel_7247/PIX_OUT pixel_7247/CSA_VREF pixel
Xpixel_6502 pixel_6502/gring pixel_6502/VDD pixel_6502/GND pixel_6502/VREF pixel_6502/ROW_SEL
+ pixel_6502/NB1 pixel_6502/VBIAS pixel_6502/NB2 pixel_6502/AMP_IN pixel_6502/SF_IB
+ pixel_6502/PIX_OUT pixel_6502/CSA_VREF pixel
Xpixel_7258 pixel_7258/gring pixel_7258/VDD pixel_7258/GND pixel_7258/VREF pixel_7258/ROW_SEL
+ pixel_7258/NB1 pixel_7258/VBIAS pixel_7258/NB2 pixel_7258/AMP_IN pixel_7258/SF_IB
+ pixel_7258/PIX_OUT pixel_7258/CSA_VREF pixel
Xpixel_7269 pixel_7269/gring pixel_7269/VDD pixel_7269/GND pixel_7269/VREF pixel_7269/ROW_SEL
+ pixel_7269/NB1 pixel_7269/VBIAS pixel_7269/NB2 pixel_7269/AMP_IN pixel_7269/SF_IB
+ pixel_7269/PIX_OUT pixel_7269/CSA_VREF pixel
Xpixel_6513 pixel_6513/gring pixel_6513/VDD pixel_6513/GND pixel_6513/VREF pixel_6513/ROW_SEL
+ pixel_6513/NB1 pixel_6513/VBIAS pixel_6513/NB2 pixel_6513/AMP_IN pixel_6513/SF_IB
+ pixel_6513/PIX_OUT pixel_6513/CSA_VREF pixel
Xpixel_6524 pixel_6524/gring pixel_6524/VDD pixel_6524/GND pixel_6524/VREF pixel_6524/ROW_SEL
+ pixel_6524/NB1 pixel_6524/VBIAS pixel_6524/NB2 pixel_6524/AMP_IN pixel_6524/SF_IB
+ pixel_6524/PIX_OUT pixel_6524/CSA_VREF pixel
Xpixel_6535 pixel_6535/gring pixel_6535/VDD pixel_6535/GND pixel_6535/VREF pixel_6535/ROW_SEL
+ pixel_6535/NB1 pixel_6535/VBIAS pixel_6535/NB2 pixel_6535/AMP_IN pixel_6535/SF_IB
+ pixel_6535/PIX_OUT pixel_6535/CSA_VREF pixel
Xpixel_6546 pixel_6546/gring pixel_6546/VDD pixel_6546/GND pixel_6546/VREF pixel_6546/ROW_SEL
+ pixel_6546/NB1 pixel_6546/VBIAS pixel_6546/NB2 pixel_6546/AMP_IN pixel_6546/SF_IB
+ pixel_6546/PIX_OUT pixel_6546/CSA_VREF pixel
Xpixel_6557 pixel_6557/gring pixel_6557/VDD pixel_6557/GND pixel_6557/VREF pixel_6557/ROW_SEL
+ pixel_6557/NB1 pixel_6557/VBIAS pixel_6557/NB2 pixel_6557/AMP_IN pixel_6557/SF_IB
+ pixel_6557/PIX_OUT pixel_6557/CSA_VREF pixel
Xpixel_6568 pixel_6568/gring pixel_6568/VDD pixel_6568/GND pixel_6568/VREF pixel_6568/ROW_SEL
+ pixel_6568/NB1 pixel_6568/VBIAS pixel_6568/NB2 pixel_6568/AMP_IN pixel_6568/SF_IB
+ pixel_6568/PIX_OUT pixel_6568/CSA_VREF pixel
Xpixel_6579 pixel_6579/gring pixel_6579/VDD pixel_6579/GND pixel_6579/VREF pixel_6579/ROW_SEL
+ pixel_6579/NB1 pixel_6579/VBIAS pixel_6579/NB2 pixel_6579/AMP_IN pixel_6579/SF_IB
+ pixel_6579/PIX_OUT pixel_6579/CSA_VREF pixel
Xpixel_5801 pixel_5801/gring pixel_5801/VDD pixel_5801/GND pixel_5801/VREF pixel_5801/ROW_SEL
+ pixel_5801/NB1 pixel_5801/VBIAS pixel_5801/NB2 pixel_5801/AMP_IN pixel_5801/SF_IB
+ pixel_5801/PIX_OUT pixel_5801/CSA_VREF pixel
Xpixel_5812 pixel_5812/gring pixel_5812/VDD pixel_5812/GND pixel_5812/VREF pixel_5812/ROW_SEL
+ pixel_5812/NB1 pixel_5812/VBIAS pixel_5812/NB2 pixel_5812/AMP_IN pixel_5812/SF_IB
+ pixel_5812/PIX_OUT pixel_5812/CSA_VREF pixel
Xpixel_5823 pixel_5823/gring pixel_5823/VDD pixel_5823/GND pixel_5823/VREF pixel_5823/ROW_SEL
+ pixel_5823/NB1 pixel_5823/VBIAS pixel_5823/NB2 pixel_5823/AMP_IN pixel_5823/SF_IB
+ pixel_5823/PIX_OUT pixel_5823/CSA_VREF pixel
Xpixel_5834 pixel_5834/gring pixel_5834/VDD pixel_5834/GND pixel_5834/VREF pixel_5834/ROW_SEL
+ pixel_5834/NB1 pixel_5834/VBIAS pixel_5834/NB2 pixel_5834/AMP_IN pixel_5834/SF_IB
+ pixel_5834/PIX_OUT pixel_5834/CSA_VREF pixel
Xpixel_5845 pixel_5845/gring pixel_5845/VDD pixel_5845/GND pixel_5845/VREF pixel_5845/ROW_SEL
+ pixel_5845/NB1 pixel_5845/VBIAS pixel_5845/NB2 pixel_5845/AMP_IN pixel_5845/SF_IB
+ pixel_5845/PIX_OUT pixel_5845/CSA_VREF pixel
Xpixel_5856 pixel_5856/gring pixel_5856/VDD pixel_5856/GND pixel_5856/VREF pixel_5856/ROW_SEL
+ pixel_5856/NB1 pixel_5856/VBIAS pixel_5856/NB2 pixel_5856/AMP_IN pixel_5856/SF_IB
+ pixel_5856/PIX_OUT pixel_5856/CSA_VREF pixel
Xpixel_5867 pixel_5867/gring pixel_5867/VDD pixel_5867/GND pixel_5867/VREF pixel_5867/ROW_SEL
+ pixel_5867/NB1 pixel_5867/VBIAS pixel_5867/NB2 pixel_5867/AMP_IN pixel_5867/SF_IB
+ pixel_5867/PIX_OUT pixel_5867/CSA_VREF pixel
Xpixel_5878 pixel_5878/gring pixel_5878/VDD pixel_5878/GND pixel_5878/VREF pixel_5878/ROW_SEL
+ pixel_5878/NB1 pixel_5878/VBIAS pixel_5878/NB2 pixel_5878/AMP_IN pixel_5878/SF_IB
+ pixel_5878/PIX_OUT pixel_5878/CSA_VREF pixel
Xpixel_5889 pixel_5889/gring pixel_5889/VDD pixel_5889/GND pixel_5889/VREF pixel_5889/ROW_SEL
+ pixel_5889/NB1 pixel_5889/VBIAS pixel_5889/NB2 pixel_5889/AMP_IN pixel_5889/SF_IB
+ pixel_5889/PIX_OUT pixel_5889/CSA_VREF pixel
Xpixel_9183 pixel_9183/gring pixel_9183/VDD pixel_9183/GND pixel_9183/VREF pixel_9183/ROW_SEL
+ pixel_9183/NB1 pixel_9183/VBIAS pixel_9183/NB2 pixel_9183/AMP_IN pixel_9183/SF_IB
+ pixel_9183/PIX_OUT pixel_9183/CSA_VREF pixel
Xpixel_9172 pixel_9172/gring pixel_9172/VDD pixel_9172/GND pixel_9172/VREF pixel_9172/ROW_SEL
+ pixel_9172/NB1 pixel_9172/VBIAS pixel_9172/NB2 pixel_9172/AMP_IN pixel_9172/SF_IB
+ pixel_9172/PIX_OUT pixel_9172/CSA_VREF pixel
Xpixel_9161 pixel_9161/gring pixel_9161/VDD pixel_9161/GND pixel_9161/VREF pixel_9161/ROW_SEL
+ pixel_9161/NB1 pixel_9161/VBIAS pixel_9161/NB2 pixel_9161/AMP_IN pixel_9161/SF_IB
+ pixel_9161/PIX_OUT pixel_9161/CSA_VREF pixel
Xpixel_9150 pixel_9150/gring pixel_9150/VDD pixel_9150/GND pixel_9150/VREF pixel_9150/ROW_SEL
+ pixel_9150/NB1 pixel_9150/VBIAS pixel_9150/NB2 pixel_9150/AMP_IN pixel_9150/SF_IB
+ pixel_9150/PIX_OUT pixel_9150/CSA_VREF pixel
Xpixel_9194 pixel_9194/gring pixel_9194/VDD pixel_9194/GND pixel_9194/VREF pixel_9194/ROW_SEL
+ pixel_9194/NB1 pixel_9194/VBIAS pixel_9194/NB2 pixel_9194/AMP_IN pixel_9194/SF_IB
+ pixel_9194/PIX_OUT pixel_9194/CSA_VREF pixel
Xpixel_8460 pixel_8460/gring pixel_8460/VDD pixel_8460/GND pixel_8460/VREF pixel_8460/ROW_SEL
+ pixel_8460/NB1 pixel_8460/VBIAS pixel_8460/NB2 pixel_8460/AMP_IN pixel_8460/SF_IB
+ pixel_8460/PIX_OUT pixel_8460/CSA_VREF pixel
Xpixel_8471 pixel_8471/gring pixel_8471/VDD pixel_8471/GND pixel_8471/VREF pixel_8471/ROW_SEL
+ pixel_8471/NB1 pixel_8471/VBIAS pixel_8471/NB2 pixel_8471/AMP_IN pixel_8471/SF_IB
+ pixel_8471/PIX_OUT pixel_8471/CSA_VREF pixel
Xpixel_8482 pixel_8482/gring pixel_8482/VDD pixel_8482/GND pixel_8482/VREF pixel_8482/ROW_SEL
+ pixel_8482/NB1 pixel_8482/VBIAS pixel_8482/NB2 pixel_8482/AMP_IN pixel_8482/SF_IB
+ pixel_8482/PIX_OUT pixel_8482/CSA_VREF pixel
Xpixel_8493 pixel_8493/gring pixel_8493/VDD pixel_8493/GND pixel_8493/VREF pixel_8493/ROW_SEL
+ pixel_8493/NB1 pixel_8493/VBIAS pixel_8493/NB2 pixel_8493/AMP_IN pixel_8493/SF_IB
+ pixel_8493/PIX_OUT pixel_8493/CSA_VREF pixel
Xpixel_7770 pixel_7770/gring pixel_7770/VDD pixel_7770/GND pixel_7770/VREF pixel_7770/ROW_SEL
+ pixel_7770/NB1 pixel_7770/VBIAS pixel_7770/NB2 pixel_7770/AMP_IN pixel_7770/SF_IB
+ pixel_7770/PIX_OUT pixel_7770/CSA_VREF pixel
Xpixel_7781 pixel_7781/gring pixel_7781/VDD pixel_7781/GND pixel_7781/VREF pixel_7781/ROW_SEL
+ pixel_7781/NB1 pixel_7781/VBIAS pixel_7781/NB2 pixel_7781/AMP_IN pixel_7781/SF_IB
+ pixel_7781/PIX_OUT pixel_7781/CSA_VREF pixel
Xpixel_7792 pixel_7792/gring pixel_7792/VDD pixel_7792/GND pixel_7792/VREF pixel_7792/ROW_SEL
+ pixel_7792/NB1 pixel_7792/VBIAS pixel_7792/NB2 pixel_7792/AMP_IN pixel_7792/SF_IB
+ pixel_7792/PIX_OUT pixel_7792/CSA_VREF pixel
Xpixel_5108 pixel_5108/gring pixel_5108/VDD pixel_5108/GND pixel_5108/VREF pixel_5108/ROW_SEL
+ pixel_5108/NB1 pixel_5108/VBIAS pixel_5108/NB2 pixel_5108/AMP_IN pixel_5108/SF_IB
+ pixel_5108/PIX_OUT pixel_5108/CSA_VREF pixel
Xpixel_5119 pixel_5119/gring pixel_5119/VDD pixel_5119/GND pixel_5119/VREF pixel_5119/ROW_SEL
+ pixel_5119/NB1 pixel_5119/VBIAS pixel_5119/NB2 pixel_5119/AMP_IN pixel_5119/SF_IB
+ pixel_5119/PIX_OUT pixel_5119/CSA_VREF pixel
Xpixel_413 pixel_413/gring pixel_413/VDD pixel_413/GND pixel_413/VREF pixel_413/ROW_SEL
+ pixel_413/NB1 pixel_413/VBIAS pixel_413/NB2 pixel_413/AMP_IN pixel_413/SF_IB pixel_413/PIX_OUT
+ pixel_413/CSA_VREF pixel
Xpixel_402 pixel_402/gring pixel_402/VDD pixel_402/GND pixel_402/VREF pixel_402/ROW_SEL
+ pixel_402/NB1 pixel_402/VBIAS pixel_402/NB2 pixel_402/AMP_IN pixel_402/SF_IB pixel_402/PIX_OUT
+ pixel_402/CSA_VREF pixel
Xpixel_4407 pixel_4407/gring pixel_4407/VDD pixel_4407/GND pixel_4407/VREF pixel_4407/ROW_SEL
+ pixel_4407/NB1 pixel_4407/VBIAS pixel_4407/NB2 pixel_4407/AMP_IN pixel_4407/SF_IB
+ pixel_4407/PIX_OUT pixel_4407/CSA_VREF pixel
Xpixel_4418 pixel_4418/gring pixel_4418/VDD pixel_4418/GND pixel_4418/VREF pixel_4418/ROW_SEL
+ pixel_4418/NB1 pixel_4418/VBIAS pixel_4418/NB2 pixel_4418/AMP_IN pixel_4418/SF_IB
+ pixel_4418/PIX_OUT pixel_4418/CSA_VREF pixel
Xpixel_446 pixel_446/gring pixel_446/VDD pixel_446/GND pixel_446/VREF pixel_446/ROW_SEL
+ pixel_446/NB1 pixel_446/VBIAS pixel_446/NB2 pixel_446/AMP_IN pixel_446/SF_IB pixel_446/PIX_OUT
+ pixel_446/CSA_VREF pixel
Xpixel_435 pixel_435/gring pixel_435/VDD pixel_435/GND pixel_435/VREF pixel_435/ROW_SEL
+ pixel_435/NB1 pixel_435/VBIAS pixel_435/NB2 pixel_435/AMP_IN pixel_435/SF_IB pixel_435/PIX_OUT
+ pixel_435/CSA_VREF pixel
Xpixel_424 pixel_424/gring pixel_424/VDD pixel_424/GND pixel_424/VREF pixel_424/ROW_SEL
+ pixel_424/NB1 pixel_424/VBIAS pixel_424/NB2 pixel_424/AMP_IN pixel_424/SF_IB pixel_424/PIX_OUT
+ pixel_424/CSA_VREF pixel
Xpixel_3706 pixel_3706/gring pixel_3706/VDD pixel_3706/GND pixel_3706/VREF pixel_3706/ROW_SEL
+ pixel_3706/NB1 pixel_3706/VBIAS pixel_3706/NB2 pixel_3706/AMP_IN pixel_3706/SF_IB
+ pixel_3706/PIX_OUT pixel_3706/CSA_VREF pixel
Xpixel_4429 pixel_4429/gring pixel_4429/VDD pixel_4429/GND pixel_4429/VREF pixel_4429/ROW_SEL
+ pixel_4429/NB1 pixel_4429/VBIAS pixel_4429/NB2 pixel_4429/AMP_IN pixel_4429/SF_IB
+ pixel_4429/PIX_OUT pixel_4429/CSA_VREF pixel
Xpixel_479 pixel_479/gring pixel_479/VDD pixel_479/GND pixel_479/VREF pixel_479/ROW_SEL
+ pixel_479/NB1 pixel_479/VBIAS pixel_479/NB2 pixel_479/AMP_IN pixel_479/SF_IB pixel_479/PIX_OUT
+ pixel_479/CSA_VREF pixel
Xpixel_468 pixel_468/gring pixel_468/VDD pixel_468/GND pixel_468/VREF pixel_468/ROW_SEL
+ pixel_468/NB1 pixel_468/VBIAS pixel_468/NB2 pixel_468/AMP_IN pixel_468/SF_IB pixel_468/PIX_OUT
+ pixel_468/CSA_VREF pixel
Xpixel_457 pixel_457/gring pixel_457/VDD pixel_457/GND pixel_457/VREF pixel_457/ROW_SEL
+ pixel_457/NB1 pixel_457/VBIAS pixel_457/NB2 pixel_457/AMP_IN pixel_457/SF_IB pixel_457/PIX_OUT
+ pixel_457/CSA_VREF pixel
Xpixel_3739 pixel_3739/gring pixel_3739/VDD pixel_3739/GND pixel_3739/VREF pixel_3739/ROW_SEL
+ pixel_3739/NB1 pixel_3739/VBIAS pixel_3739/NB2 pixel_3739/AMP_IN pixel_3739/SF_IB
+ pixel_3739/PIX_OUT pixel_3739/CSA_VREF pixel
Xpixel_3728 pixel_3728/gring pixel_3728/VDD pixel_3728/GND pixel_3728/VREF pixel_3728/ROW_SEL
+ pixel_3728/NB1 pixel_3728/VBIAS pixel_3728/NB2 pixel_3728/AMP_IN pixel_3728/SF_IB
+ pixel_3728/PIX_OUT pixel_3728/CSA_VREF pixel
Xpixel_3717 pixel_3717/gring pixel_3717/VDD pixel_3717/GND pixel_3717/VREF pixel_3717/ROW_SEL
+ pixel_3717/NB1 pixel_3717/VBIAS pixel_3717/NB2 pixel_3717/AMP_IN pixel_3717/SF_IB
+ pixel_3717/PIX_OUT pixel_3717/CSA_VREF pixel
Xpixel_7000 pixel_7000/gring pixel_7000/VDD pixel_7000/GND pixel_7000/VREF pixel_7000/ROW_SEL
+ pixel_7000/NB1 pixel_7000/VBIAS pixel_7000/NB2 pixel_7000/AMP_IN pixel_7000/SF_IB
+ pixel_7000/PIX_OUT pixel_7000/CSA_VREF pixel
Xpixel_7011 pixel_7011/gring pixel_7011/VDD pixel_7011/GND pixel_7011/VREF pixel_7011/ROW_SEL
+ pixel_7011/NB1 pixel_7011/VBIAS pixel_7011/NB2 pixel_7011/AMP_IN pixel_7011/SF_IB
+ pixel_7011/PIX_OUT pixel_7011/CSA_VREF pixel
Xpixel_7022 pixel_7022/gring pixel_7022/VDD pixel_7022/GND pixel_7022/VREF pixel_7022/ROW_SEL
+ pixel_7022/NB1 pixel_7022/VBIAS pixel_7022/NB2 pixel_7022/AMP_IN pixel_7022/SF_IB
+ pixel_7022/PIX_OUT pixel_7022/CSA_VREF pixel
Xpixel_7033 pixel_7033/gring pixel_7033/VDD pixel_7033/GND pixel_7033/VREF pixel_7033/ROW_SEL
+ pixel_7033/NB1 pixel_7033/VBIAS pixel_7033/NB2 pixel_7033/AMP_IN pixel_7033/SF_IB
+ pixel_7033/PIX_OUT pixel_7033/CSA_VREF pixel
Xpixel_7044 pixel_7044/gring pixel_7044/VDD pixel_7044/GND pixel_7044/VREF pixel_7044/ROW_SEL
+ pixel_7044/NB1 pixel_7044/VBIAS pixel_7044/NB2 pixel_7044/AMP_IN pixel_7044/SF_IB
+ pixel_7044/PIX_OUT pixel_7044/CSA_VREF pixel
Xpixel_7055 pixel_7055/gring pixel_7055/VDD pixel_7055/GND pixel_7055/VREF pixel_7055/ROW_SEL
+ pixel_7055/NB1 pixel_7055/VBIAS pixel_7055/NB2 pixel_7055/AMP_IN pixel_7055/SF_IB
+ pixel_7055/PIX_OUT pixel_7055/CSA_VREF pixel
Xpixel_6310 pixel_6310/gring pixel_6310/VDD pixel_6310/GND pixel_6310/VREF pixel_6310/ROW_SEL
+ pixel_6310/NB1 pixel_6310/VBIAS pixel_6310/NB2 pixel_6310/AMP_IN pixel_6310/SF_IB
+ pixel_6310/PIX_OUT pixel_6310/CSA_VREF pixel
Xpixel_7066 pixel_7066/gring pixel_7066/VDD pixel_7066/GND pixel_7066/VREF pixel_7066/ROW_SEL
+ pixel_7066/NB1 pixel_7066/VBIAS pixel_7066/NB2 pixel_7066/AMP_IN pixel_7066/SF_IB
+ pixel_7066/PIX_OUT pixel_7066/CSA_VREF pixel
Xpixel_7077 pixel_7077/gring pixel_7077/VDD pixel_7077/GND pixel_7077/VREF pixel_7077/ROW_SEL
+ pixel_7077/NB1 pixel_7077/VBIAS pixel_7077/NB2 pixel_7077/AMP_IN pixel_7077/SF_IB
+ pixel_7077/PIX_OUT pixel_7077/CSA_VREF pixel
Xpixel_7088 pixel_7088/gring pixel_7088/VDD pixel_7088/GND pixel_7088/VREF pixel_7088/ROW_SEL
+ pixel_7088/NB1 pixel_7088/VBIAS pixel_7088/NB2 pixel_7088/AMP_IN pixel_7088/SF_IB
+ pixel_7088/PIX_OUT pixel_7088/CSA_VREF pixel
Xpixel_6321 pixel_6321/gring pixel_6321/VDD pixel_6321/GND pixel_6321/VREF pixel_6321/ROW_SEL
+ pixel_6321/NB1 pixel_6321/VBIAS pixel_6321/NB2 pixel_6321/AMP_IN pixel_6321/SF_IB
+ pixel_6321/PIX_OUT pixel_6321/CSA_VREF pixel
Xpixel_6332 pixel_6332/gring pixel_6332/VDD pixel_6332/GND pixel_6332/VREF pixel_6332/ROW_SEL
+ pixel_6332/NB1 pixel_6332/VBIAS pixel_6332/NB2 pixel_6332/AMP_IN pixel_6332/SF_IB
+ pixel_6332/PIX_OUT pixel_6332/CSA_VREF pixel
Xpixel_6343 pixel_6343/gring pixel_6343/VDD pixel_6343/GND pixel_6343/VREF pixel_6343/ROW_SEL
+ pixel_6343/NB1 pixel_6343/VBIAS pixel_6343/NB2 pixel_6343/AMP_IN pixel_6343/SF_IB
+ pixel_6343/PIX_OUT pixel_6343/CSA_VREF pixel
Xpixel_6354 pixel_6354/gring pixel_6354/VDD pixel_6354/GND pixel_6354/VREF pixel_6354/ROW_SEL
+ pixel_6354/NB1 pixel_6354/VBIAS pixel_6354/NB2 pixel_6354/AMP_IN pixel_6354/SF_IB
+ pixel_6354/PIX_OUT pixel_6354/CSA_VREF pixel
Xpixel_7099 pixel_7099/gring pixel_7099/VDD pixel_7099/GND pixel_7099/VREF pixel_7099/ROW_SEL
+ pixel_7099/NB1 pixel_7099/VBIAS pixel_7099/NB2 pixel_7099/AMP_IN pixel_7099/SF_IB
+ pixel_7099/PIX_OUT pixel_7099/CSA_VREF pixel
Xpixel_6365 pixel_6365/gring pixel_6365/VDD pixel_6365/GND pixel_6365/VREF pixel_6365/ROW_SEL
+ pixel_6365/NB1 pixel_6365/VBIAS pixel_6365/NB2 pixel_6365/AMP_IN pixel_6365/SF_IB
+ pixel_6365/PIX_OUT pixel_6365/CSA_VREF pixel
Xpixel_6376 pixel_6376/gring pixel_6376/VDD pixel_6376/GND pixel_6376/VREF pixel_6376/ROW_SEL
+ pixel_6376/NB1 pixel_6376/VBIAS pixel_6376/NB2 pixel_6376/AMP_IN pixel_6376/SF_IB
+ pixel_6376/PIX_OUT pixel_6376/CSA_VREF pixel
Xpixel_6387 pixel_6387/gring pixel_6387/VDD pixel_6387/GND pixel_6387/VREF pixel_6387/ROW_SEL
+ pixel_6387/NB1 pixel_6387/VBIAS pixel_6387/NB2 pixel_6387/AMP_IN pixel_6387/SF_IB
+ pixel_6387/PIX_OUT pixel_6387/CSA_VREF pixel
Xpixel_5620 pixel_5620/gring pixel_5620/VDD pixel_5620/GND pixel_5620/VREF pixel_5620/ROW_SEL
+ pixel_5620/NB1 pixel_5620/VBIAS pixel_5620/NB2 pixel_5620/AMP_IN pixel_5620/SF_IB
+ pixel_5620/PIX_OUT pixel_5620/CSA_VREF pixel
Xpixel_5631 pixel_5631/gring pixel_5631/VDD pixel_5631/GND pixel_5631/VREF pixel_5631/ROW_SEL
+ pixel_5631/NB1 pixel_5631/VBIAS pixel_5631/NB2 pixel_5631/AMP_IN pixel_5631/SF_IB
+ pixel_5631/PIX_OUT pixel_5631/CSA_VREF pixel
Xpixel_5642 pixel_5642/gring pixel_5642/VDD pixel_5642/GND pixel_5642/VREF pixel_5642/ROW_SEL
+ pixel_5642/NB1 pixel_5642/VBIAS pixel_5642/NB2 pixel_5642/AMP_IN pixel_5642/SF_IB
+ pixel_5642/PIX_OUT pixel_5642/CSA_VREF pixel
Xpixel_6398 pixel_6398/gring pixel_6398/VDD pixel_6398/GND pixel_6398/VREF pixel_6398/ROW_SEL
+ pixel_6398/NB1 pixel_6398/VBIAS pixel_6398/NB2 pixel_6398/AMP_IN pixel_6398/SF_IB
+ pixel_6398/PIX_OUT pixel_6398/CSA_VREF pixel
Xpixel_5653 pixel_5653/gring pixel_5653/VDD pixel_5653/GND pixel_5653/VREF pixel_5653/ROW_SEL
+ pixel_5653/NB1 pixel_5653/VBIAS pixel_5653/NB2 pixel_5653/AMP_IN pixel_5653/SF_IB
+ pixel_5653/PIX_OUT pixel_5653/CSA_VREF pixel
Xpixel_5664 pixel_5664/gring pixel_5664/VDD pixel_5664/GND pixel_5664/VREF pixel_5664/ROW_SEL
+ pixel_5664/NB1 pixel_5664/VBIAS pixel_5664/NB2 pixel_5664/AMP_IN pixel_5664/SF_IB
+ pixel_5664/PIX_OUT pixel_5664/CSA_VREF pixel
Xpixel_5675 pixel_5675/gring pixel_5675/VDD pixel_5675/GND pixel_5675/VREF pixel_5675/ROW_SEL
+ pixel_5675/NB1 pixel_5675/VBIAS pixel_5675/NB2 pixel_5675/AMP_IN pixel_5675/SF_IB
+ pixel_5675/PIX_OUT pixel_5675/CSA_VREF pixel
Xpixel_4930 pixel_4930/gring pixel_4930/VDD pixel_4930/GND pixel_4930/VREF pixel_4930/ROW_SEL
+ pixel_4930/NB1 pixel_4930/VBIAS pixel_4930/NB2 pixel_4930/AMP_IN pixel_4930/SF_IB
+ pixel_4930/PIX_OUT pixel_4930/CSA_VREF pixel
Xpixel_5686 pixel_5686/gring pixel_5686/VDD pixel_5686/GND pixel_5686/VREF pixel_5686/ROW_SEL
+ pixel_5686/NB1 pixel_5686/VBIAS pixel_5686/NB2 pixel_5686/AMP_IN pixel_5686/SF_IB
+ pixel_5686/PIX_OUT pixel_5686/CSA_VREF pixel
Xpixel_5697 pixel_5697/gring pixel_5697/VDD pixel_5697/GND pixel_5697/VREF pixel_5697/ROW_SEL
+ pixel_5697/NB1 pixel_5697/VBIAS pixel_5697/NB2 pixel_5697/AMP_IN pixel_5697/SF_IB
+ pixel_5697/PIX_OUT pixel_5697/CSA_VREF pixel
Xpixel_4941 pixel_4941/gring pixel_4941/VDD pixel_4941/GND pixel_4941/VREF pixel_4941/ROW_SEL
+ pixel_4941/NB1 pixel_4941/VBIAS pixel_4941/NB2 pixel_4941/AMP_IN pixel_4941/SF_IB
+ pixel_4941/PIX_OUT pixel_4941/CSA_VREF pixel
Xpixel_4952 pixel_4952/gring pixel_4952/VDD pixel_4952/GND pixel_4952/VREF pixel_4952/ROW_SEL
+ pixel_4952/NB1 pixel_4952/VBIAS pixel_4952/NB2 pixel_4952/AMP_IN pixel_4952/SF_IB
+ pixel_4952/PIX_OUT pixel_4952/CSA_VREF pixel
Xpixel_4963 pixel_4963/gring pixel_4963/VDD pixel_4963/GND pixel_4963/VREF pixel_4963/ROW_SEL
+ pixel_4963/NB1 pixel_4963/VBIAS pixel_4963/NB2 pixel_4963/AMP_IN pixel_4963/SF_IB
+ pixel_4963/PIX_OUT pixel_4963/CSA_VREF pixel
Xpixel_4974 pixel_4974/gring pixel_4974/VDD pixel_4974/GND pixel_4974/VREF pixel_4974/ROW_SEL
+ pixel_4974/NB1 pixel_4974/VBIAS pixel_4974/NB2 pixel_4974/AMP_IN pixel_4974/SF_IB
+ pixel_4974/PIX_OUT pixel_4974/CSA_VREF pixel
Xpixel_991 pixel_991/gring pixel_991/VDD pixel_991/GND pixel_991/VREF pixel_991/ROW_SEL
+ pixel_991/NB1 pixel_991/VBIAS pixel_991/NB2 pixel_991/AMP_IN pixel_991/SF_IB pixel_991/PIX_OUT
+ pixel_991/CSA_VREF pixel
Xpixel_980 pixel_980/gring pixel_980/VDD pixel_980/GND pixel_980/VREF pixel_980/ROW_SEL
+ pixel_980/NB1 pixel_980/VBIAS pixel_980/NB2 pixel_980/AMP_IN pixel_980/SF_IB pixel_980/PIX_OUT
+ pixel_980/CSA_VREF pixel
Xpixel_4985 pixel_4985/gring pixel_4985/VDD pixel_4985/GND pixel_4985/VREF pixel_4985/ROW_SEL
+ pixel_4985/NB1 pixel_4985/VBIAS pixel_4985/NB2 pixel_4985/AMP_IN pixel_4985/SF_IB
+ pixel_4985/PIX_OUT pixel_4985/CSA_VREF pixel
Xpixel_4996 pixel_4996/gring pixel_4996/VDD pixel_4996/GND pixel_4996/VREF pixel_4996/ROW_SEL
+ pixel_4996/NB1 pixel_4996/VBIAS pixel_4996/NB2 pixel_4996/AMP_IN pixel_4996/SF_IB
+ pixel_4996/PIX_OUT pixel_4996/CSA_VREF pixel
Xpixel_8290 pixel_8290/gring pixel_8290/VDD pixel_8290/GND pixel_8290/VREF pixel_8290/ROW_SEL
+ pixel_8290/NB1 pixel_8290/VBIAS pixel_8290/NB2 pixel_8290/AMP_IN pixel_8290/SF_IB
+ pixel_8290/PIX_OUT pixel_8290/CSA_VREF pixel
Xpixel_9919 pixel_9919/gring pixel_9919/VDD pixel_9919/GND pixel_9919/VREF pixel_9919/ROW_SEL
+ pixel_9919/NB1 pixel_9919/VBIAS pixel_9919/NB2 pixel_9919/AMP_IN pixel_9919/SF_IB
+ pixel_9919/PIX_OUT pixel_9919/CSA_VREF pixel
Xpixel_9908 pixel_9908/gring pixel_9908/VDD pixel_9908/GND pixel_9908/VREF pixel_9908/ROW_SEL
+ pixel_9908/NB1 pixel_9908/VBIAS pixel_9908/NB2 pixel_9908/AMP_IN pixel_9908/SF_IB
+ pixel_9908/PIX_OUT pixel_9908/CSA_VREF pixel
Xpixel_221 pixel_221/gring pixel_221/VDD pixel_221/GND pixel_221/VREF pixel_221/ROW_SEL
+ pixel_221/NB1 pixel_221/VBIAS pixel_221/NB2 pixel_221/AMP_IN pixel_221/SF_IB pixel_221/PIX_OUT
+ pixel_221/CSA_VREF pixel
Xpixel_210 pixel_210/gring pixel_210/VDD pixel_210/GND pixel_210/VREF pixel_210/ROW_SEL
+ pixel_210/NB1 pixel_210/VBIAS pixel_210/NB2 pixel_210/AMP_IN pixel_210/SF_IB pixel_210/PIX_OUT
+ pixel_210/CSA_VREF pixel
Xpixel_4204 pixel_4204/gring pixel_4204/VDD pixel_4204/GND pixel_4204/VREF pixel_4204/ROW_SEL
+ pixel_4204/NB1 pixel_4204/VBIAS pixel_4204/NB2 pixel_4204/AMP_IN pixel_4204/SF_IB
+ pixel_4204/PIX_OUT pixel_4204/CSA_VREF pixel
Xpixel_4215 pixel_4215/gring pixel_4215/VDD pixel_4215/GND pixel_4215/VREF pixel_4215/ROW_SEL
+ pixel_4215/NB1 pixel_4215/VBIAS pixel_4215/NB2 pixel_4215/AMP_IN pixel_4215/SF_IB
+ pixel_4215/PIX_OUT pixel_4215/CSA_VREF pixel
Xpixel_4226 pixel_4226/gring pixel_4226/VDD pixel_4226/GND pixel_4226/VREF pixel_4226/ROW_SEL
+ pixel_4226/NB1 pixel_4226/VBIAS pixel_4226/NB2 pixel_4226/AMP_IN pixel_4226/SF_IB
+ pixel_4226/PIX_OUT pixel_4226/CSA_VREF pixel
Xpixel_265 pixel_265/gring pixel_265/VDD pixel_265/GND pixel_265/VREF pixel_265/ROW_SEL
+ pixel_265/NB1 pixel_265/VBIAS pixel_265/NB2 pixel_265/AMP_IN pixel_265/SF_IB pixel_265/PIX_OUT
+ pixel_265/CSA_VREF pixel
Xpixel_254 pixel_254/gring pixel_254/VDD pixel_254/GND pixel_254/VREF pixel_254/ROW_SEL
+ pixel_254/NB1 pixel_254/VBIAS pixel_254/NB2 pixel_254/AMP_IN pixel_254/SF_IB pixel_254/PIX_OUT
+ pixel_254/CSA_VREF pixel
Xpixel_243 pixel_243/gring pixel_243/VDD pixel_243/GND pixel_243/VREF pixel_243/ROW_SEL
+ pixel_243/NB1 pixel_243/VBIAS pixel_243/NB2 pixel_243/AMP_IN pixel_243/SF_IB pixel_243/PIX_OUT
+ pixel_243/CSA_VREF pixel
Xpixel_232 pixel_232/gring pixel_232/VDD pixel_232/GND pixel_232/VREF pixel_232/ROW_SEL
+ pixel_232/NB1 pixel_232/VBIAS pixel_232/NB2 pixel_232/AMP_IN pixel_232/SF_IB pixel_232/PIX_OUT
+ pixel_232/CSA_VREF pixel
Xpixel_3525 pixel_3525/gring pixel_3525/VDD pixel_3525/GND pixel_3525/VREF pixel_3525/ROW_SEL
+ pixel_3525/NB1 pixel_3525/VBIAS pixel_3525/NB2 pixel_3525/AMP_IN pixel_3525/SF_IB
+ pixel_3525/PIX_OUT pixel_3525/CSA_VREF pixel
Xpixel_3514 pixel_3514/gring pixel_3514/VDD pixel_3514/GND pixel_3514/VREF pixel_3514/ROW_SEL
+ pixel_3514/NB1 pixel_3514/VBIAS pixel_3514/NB2 pixel_3514/AMP_IN pixel_3514/SF_IB
+ pixel_3514/PIX_OUT pixel_3514/CSA_VREF pixel
Xpixel_3503 pixel_3503/gring pixel_3503/VDD pixel_3503/GND pixel_3503/VREF pixel_3503/ROW_SEL
+ pixel_3503/NB1 pixel_3503/VBIAS pixel_3503/NB2 pixel_3503/AMP_IN pixel_3503/SF_IB
+ pixel_3503/PIX_OUT pixel_3503/CSA_VREF pixel
Xpixel_4237 pixel_4237/gring pixel_4237/VDD pixel_4237/GND pixel_4237/VREF pixel_4237/ROW_SEL
+ pixel_4237/NB1 pixel_4237/VBIAS pixel_4237/NB2 pixel_4237/AMP_IN pixel_4237/SF_IB
+ pixel_4237/PIX_OUT pixel_4237/CSA_VREF pixel
Xpixel_4248 pixel_4248/gring pixel_4248/VDD pixel_4248/GND pixel_4248/VREF pixel_4248/ROW_SEL
+ pixel_4248/NB1 pixel_4248/VBIAS pixel_4248/NB2 pixel_4248/AMP_IN pixel_4248/SF_IB
+ pixel_4248/PIX_OUT pixel_4248/CSA_VREF pixel
Xpixel_4259 pixel_4259/gring pixel_4259/VDD pixel_4259/GND pixel_4259/VREF pixel_4259/ROW_SEL
+ pixel_4259/NB1 pixel_4259/VBIAS pixel_4259/NB2 pixel_4259/AMP_IN pixel_4259/SF_IB
+ pixel_4259/PIX_OUT pixel_4259/CSA_VREF pixel
Xpixel_298 pixel_298/gring pixel_298/VDD pixel_298/GND pixel_298/VREF pixel_298/ROW_SEL
+ pixel_298/NB1 pixel_298/VBIAS pixel_298/NB2 pixel_298/AMP_IN pixel_298/SF_IB pixel_298/PIX_OUT
+ pixel_298/CSA_VREF pixel
Xpixel_287 pixel_287/gring pixel_287/VDD pixel_287/GND pixel_287/VREF pixel_287/ROW_SEL
+ pixel_287/NB1 pixel_287/VBIAS pixel_287/NB2 pixel_287/AMP_IN pixel_287/SF_IB pixel_287/PIX_OUT
+ pixel_287/CSA_VREF pixel
Xpixel_276 pixel_276/gring pixel_276/VDD pixel_276/GND pixel_276/VREF pixel_276/ROW_SEL
+ pixel_276/NB1 pixel_276/VBIAS pixel_276/NB2 pixel_276/AMP_IN pixel_276/SF_IB pixel_276/PIX_OUT
+ pixel_276/CSA_VREF pixel
Xpixel_2813 pixel_2813/gring pixel_2813/VDD pixel_2813/GND pixel_2813/VREF pixel_2813/ROW_SEL
+ pixel_2813/NB1 pixel_2813/VBIAS pixel_2813/NB2 pixel_2813/AMP_IN pixel_2813/SF_IB
+ pixel_2813/PIX_OUT pixel_2813/CSA_VREF pixel
Xpixel_2802 pixel_2802/gring pixel_2802/VDD pixel_2802/GND pixel_2802/VREF pixel_2802/ROW_SEL
+ pixel_2802/NB1 pixel_2802/VBIAS pixel_2802/NB2 pixel_2802/AMP_IN pixel_2802/SF_IB
+ pixel_2802/PIX_OUT pixel_2802/CSA_VREF pixel
Xpixel_3558 pixel_3558/gring pixel_3558/VDD pixel_3558/GND pixel_3558/VREF pixel_3558/ROW_SEL
+ pixel_3558/NB1 pixel_3558/VBIAS pixel_3558/NB2 pixel_3558/AMP_IN pixel_3558/SF_IB
+ pixel_3558/PIX_OUT pixel_3558/CSA_VREF pixel
Xpixel_3547 pixel_3547/gring pixel_3547/VDD pixel_3547/GND pixel_3547/VREF pixel_3547/ROW_SEL
+ pixel_3547/NB1 pixel_3547/VBIAS pixel_3547/NB2 pixel_3547/AMP_IN pixel_3547/SF_IB
+ pixel_3547/PIX_OUT pixel_3547/CSA_VREF pixel
Xpixel_3536 pixel_3536/gring pixel_3536/VDD pixel_3536/GND pixel_3536/VREF pixel_3536/ROW_SEL
+ pixel_3536/NB1 pixel_3536/VBIAS pixel_3536/NB2 pixel_3536/AMP_IN pixel_3536/SF_IB
+ pixel_3536/PIX_OUT pixel_3536/CSA_VREF pixel
Xpixel_2846 pixel_2846/gring pixel_2846/VDD pixel_2846/GND pixel_2846/VREF pixel_2846/ROW_SEL
+ pixel_2846/NB1 pixel_2846/VBIAS pixel_2846/NB2 pixel_2846/AMP_IN pixel_2846/SF_IB
+ pixel_2846/PIX_OUT pixel_2846/CSA_VREF pixel
Xpixel_2835 pixel_2835/gring pixel_2835/VDD pixel_2835/GND pixel_2835/VREF pixel_2835/ROW_SEL
+ pixel_2835/NB1 pixel_2835/VBIAS pixel_2835/NB2 pixel_2835/AMP_IN pixel_2835/SF_IB
+ pixel_2835/PIX_OUT pixel_2835/CSA_VREF pixel
Xpixel_2824 pixel_2824/gring pixel_2824/VDD pixel_2824/GND pixel_2824/VREF pixel_2824/ROW_SEL
+ pixel_2824/NB1 pixel_2824/VBIAS pixel_2824/NB2 pixel_2824/AMP_IN pixel_2824/SF_IB
+ pixel_2824/PIX_OUT pixel_2824/CSA_VREF pixel
Xpixel_3569 pixel_3569/gring pixel_3569/VDD pixel_3569/GND pixel_3569/VREF pixel_3569/ROW_SEL
+ pixel_3569/NB1 pixel_3569/VBIAS pixel_3569/NB2 pixel_3569/AMP_IN pixel_3569/SF_IB
+ pixel_3569/PIX_OUT pixel_3569/CSA_VREF pixel
Xpixel_2879 pixel_2879/gring pixel_2879/VDD pixel_2879/GND pixel_2879/VREF pixel_2879/ROW_SEL
+ pixel_2879/NB1 pixel_2879/VBIAS pixel_2879/NB2 pixel_2879/AMP_IN pixel_2879/SF_IB
+ pixel_2879/PIX_OUT pixel_2879/CSA_VREF pixel
Xpixel_2868 pixel_2868/gring pixel_2868/VDD pixel_2868/GND pixel_2868/VREF pixel_2868/ROW_SEL
+ pixel_2868/NB1 pixel_2868/VBIAS pixel_2868/NB2 pixel_2868/AMP_IN pixel_2868/SF_IB
+ pixel_2868/PIX_OUT pixel_2868/CSA_VREF pixel
Xpixel_2857 pixel_2857/gring pixel_2857/VDD pixel_2857/GND pixel_2857/VREF pixel_2857/ROW_SEL
+ pixel_2857/NB1 pixel_2857/VBIAS pixel_2857/NB2 pixel_2857/AMP_IN pixel_2857/SF_IB
+ pixel_2857/PIX_OUT pixel_2857/CSA_VREF pixel
Xpixel_6140 pixel_6140/gring pixel_6140/VDD pixel_6140/GND pixel_6140/VREF pixel_6140/ROW_SEL
+ pixel_6140/NB1 pixel_6140/VBIAS pixel_6140/NB2 pixel_6140/AMP_IN pixel_6140/SF_IB
+ pixel_6140/PIX_OUT pixel_6140/CSA_VREF pixel
Xpixel_6151 pixel_6151/gring pixel_6151/VDD pixel_6151/GND pixel_6151/VREF pixel_6151/ROW_SEL
+ pixel_6151/NB1 pixel_6151/VBIAS pixel_6151/NB2 pixel_6151/AMP_IN pixel_6151/SF_IB
+ pixel_6151/PIX_OUT pixel_6151/CSA_VREF pixel
Xpixel_6162 pixel_6162/gring pixel_6162/VDD pixel_6162/GND pixel_6162/VREF pixel_6162/ROW_SEL
+ pixel_6162/NB1 pixel_6162/VBIAS pixel_6162/NB2 pixel_6162/AMP_IN pixel_6162/SF_IB
+ pixel_6162/PIX_OUT pixel_6162/CSA_VREF pixel
Xpixel_6173 pixel_6173/gring pixel_6173/VDD pixel_6173/GND pixel_6173/VREF pixel_6173/ROW_SEL
+ pixel_6173/NB1 pixel_6173/VBIAS pixel_6173/NB2 pixel_6173/AMP_IN pixel_6173/SF_IB
+ pixel_6173/PIX_OUT pixel_6173/CSA_VREF pixel
Xpixel_6184 pixel_6184/gring pixel_6184/VDD pixel_6184/GND pixel_6184/VREF pixel_6184/ROW_SEL
+ pixel_6184/NB1 pixel_6184/VBIAS pixel_6184/NB2 pixel_6184/AMP_IN pixel_6184/SF_IB
+ pixel_6184/PIX_OUT pixel_6184/CSA_VREF pixel
Xpixel_6195 pixel_6195/gring pixel_6195/VDD pixel_6195/GND pixel_6195/VREF pixel_6195/ROW_SEL
+ pixel_6195/NB1 pixel_6195/VBIAS pixel_6195/NB2 pixel_6195/AMP_IN pixel_6195/SF_IB
+ pixel_6195/PIX_OUT pixel_6195/CSA_VREF pixel
Xpixel_5450 pixel_5450/gring pixel_5450/VDD pixel_5450/GND pixel_5450/VREF pixel_5450/ROW_SEL
+ pixel_5450/NB1 pixel_5450/VBIAS pixel_5450/NB2 pixel_5450/AMP_IN pixel_5450/SF_IB
+ pixel_5450/PIX_OUT pixel_5450/CSA_VREF pixel
Xpixel_5461 pixel_5461/gring pixel_5461/VDD pixel_5461/GND pixel_5461/VREF pixel_5461/ROW_SEL
+ pixel_5461/NB1 pixel_5461/VBIAS pixel_5461/NB2 pixel_5461/AMP_IN pixel_5461/SF_IB
+ pixel_5461/PIX_OUT pixel_5461/CSA_VREF pixel
Xpixel_5472 pixel_5472/gring pixel_5472/VDD pixel_5472/GND pixel_5472/VREF pixel_5472/ROW_SEL
+ pixel_5472/NB1 pixel_5472/VBIAS pixel_5472/NB2 pixel_5472/AMP_IN pixel_5472/SF_IB
+ pixel_5472/PIX_OUT pixel_5472/CSA_VREF pixel
Xpixel_5483 pixel_5483/gring pixel_5483/VDD pixel_5483/GND pixel_5483/VREF pixel_5483/ROW_SEL
+ pixel_5483/NB1 pixel_5483/VBIAS pixel_5483/NB2 pixel_5483/AMP_IN pixel_5483/SF_IB
+ pixel_5483/PIX_OUT pixel_5483/CSA_VREF pixel
Xpixel_5494 pixel_5494/gring pixel_5494/VDD pixel_5494/GND pixel_5494/VREF pixel_5494/ROW_SEL
+ pixel_5494/NB1 pixel_5494/VBIAS pixel_5494/NB2 pixel_5494/AMP_IN pixel_5494/SF_IB
+ pixel_5494/PIX_OUT pixel_5494/CSA_VREF pixel
Xpixel_4760 pixel_4760/gring pixel_4760/VDD pixel_4760/GND pixel_4760/VREF pixel_4760/ROW_SEL
+ pixel_4760/NB1 pixel_4760/VBIAS pixel_4760/NB2 pixel_4760/AMP_IN pixel_4760/SF_IB
+ pixel_4760/PIX_OUT pixel_4760/CSA_VREF pixel
Xpixel_4771 pixel_4771/gring pixel_4771/VDD pixel_4771/GND pixel_4771/VREF pixel_4771/ROW_SEL
+ pixel_4771/NB1 pixel_4771/VBIAS pixel_4771/NB2 pixel_4771/AMP_IN pixel_4771/SF_IB
+ pixel_4771/PIX_OUT pixel_4771/CSA_VREF pixel
Xpixel_4782 pixel_4782/gring pixel_4782/VDD pixel_4782/GND pixel_4782/VREF pixel_4782/ROW_SEL
+ pixel_4782/NB1 pixel_4782/VBIAS pixel_4782/NB2 pixel_4782/AMP_IN pixel_4782/SF_IB
+ pixel_4782/PIX_OUT pixel_4782/CSA_VREF pixel
Xpixel_4793 pixel_4793/gring pixel_4793/VDD pixel_4793/GND pixel_4793/VREF pixel_4793/ROW_SEL
+ pixel_4793/NB1 pixel_4793/VBIAS pixel_4793/NB2 pixel_4793/AMP_IN pixel_4793/SF_IB
+ pixel_4793/PIX_OUT pixel_4793/CSA_VREF pixel
Xpixel_2109 pixel_2109/gring pixel_2109/VDD pixel_2109/GND pixel_2109/VREF pixel_2109/ROW_SEL
+ pixel_2109/NB1 pixel_2109/VBIAS pixel_2109/NB2 pixel_2109/AMP_IN pixel_2109/SF_IB
+ pixel_2109/PIX_OUT pixel_2109/CSA_VREF pixel
Xpixel_1419 pixel_1419/gring pixel_1419/VDD pixel_1419/GND pixel_1419/VREF pixel_1419/ROW_SEL
+ pixel_1419/NB1 pixel_1419/VBIAS pixel_1419/NB2 pixel_1419/AMP_IN pixel_1419/SF_IB
+ pixel_1419/PIX_OUT pixel_1419/CSA_VREF pixel
Xpixel_1408 pixel_1408/gring pixel_1408/VDD pixel_1408/GND pixel_1408/VREF pixel_1408/ROW_SEL
+ pixel_1408/NB1 pixel_1408/VBIAS pixel_1408/NB2 pixel_1408/AMP_IN pixel_1408/SF_IB
+ pixel_1408/PIX_OUT pixel_1408/CSA_VREF pixel
Xpixel_9705 pixel_9705/gring pixel_9705/VDD pixel_9705/GND pixel_9705/VREF pixel_9705/ROW_SEL
+ pixel_9705/NB1 pixel_9705/VBIAS pixel_9705/NB2 pixel_9705/AMP_IN pixel_9705/SF_IB
+ pixel_9705/PIX_OUT pixel_9705/CSA_VREF pixel
Xpixel_9716 pixel_9716/gring pixel_9716/VDD pixel_9716/GND pixel_9716/VREF pixel_9716/ROW_SEL
+ pixel_9716/NB1 pixel_9716/VBIAS pixel_9716/NB2 pixel_9716/AMP_IN pixel_9716/SF_IB
+ pixel_9716/PIX_OUT pixel_9716/CSA_VREF pixel
Xpixel_9727 pixel_9727/gring pixel_9727/VDD pixel_9727/GND pixel_9727/VREF pixel_9727/ROW_SEL
+ pixel_9727/NB1 pixel_9727/VBIAS pixel_9727/NB2 pixel_9727/AMP_IN pixel_9727/SF_IB
+ pixel_9727/PIX_OUT pixel_9727/CSA_VREF pixel
Xpixel_9738 pixel_9738/gring pixel_9738/VDD pixel_9738/GND pixel_9738/VREF pixel_9738/ROW_SEL
+ pixel_9738/NB1 pixel_9738/VBIAS pixel_9738/NB2 pixel_9738/AMP_IN pixel_9738/SF_IB
+ pixel_9738/PIX_OUT pixel_9738/CSA_VREF pixel
Xpixel_9749 pixel_9749/gring pixel_9749/VDD pixel_9749/GND pixel_9749/VREF pixel_9749/ROW_SEL
+ pixel_9749/NB1 pixel_9749/VBIAS pixel_9749/NB2 pixel_9749/AMP_IN pixel_9749/SF_IB
+ pixel_9749/PIX_OUT pixel_9749/CSA_VREF pixel
Xpixel_4001 pixel_4001/gring pixel_4001/VDD pixel_4001/GND pixel_4001/VREF pixel_4001/ROW_SEL
+ pixel_4001/NB1 pixel_4001/VBIAS pixel_4001/NB2 pixel_4001/AMP_IN pixel_4001/SF_IB
+ pixel_4001/PIX_OUT pixel_4001/CSA_VREF pixel
Xpixel_4012 pixel_4012/gring pixel_4012/VDD pixel_4012/GND pixel_4012/VREF pixel_4012/ROW_SEL
+ pixel_4012/NB1 pixel_4012/VBIAS pixel_4012/NB2 pixel_4012/AMP_IN pixel_4012/SF_IB
+ pixel_4012/PIX_OUT pixel_4012/CSA_VREF pixel
Xpixel_4023 pixel_4023/gring pixel_4023/VDD pixel_4023/GND pixel_4023/VREF pixel_4023/ROW_SEL
+ pixel_4023/NB1 pixel_4023/VBIAS pixel_4023/NB2 pixel_4023/AMP_IN pixel_4023/SF_IB
+ pixel_4023/PIX_OUT pixel_4023/CSA_VREF pixel
Xpixel_4034 pixel_4034/gring pixel_4034/VDD pixel_4034/GND pixel_4034/VREF pixel_4034/ROW_SEL
+ pixel_4034/NB1 pixel_4034/VBIAS pixel_4034/NB2 pixel_4034/AMP_IN pixel_4034/SF_IB
+ pixel_4034/PIX_OUT pixel_4034/CSA_VREF pixel
Xpixel_3333 pixel_3333/gring pixel_3333/VDD pixel_3333/GND pixel_3333/VREF pixel_3333/ROW_SEL
+ pixel_3333/NB1 pixel_3333/VBIAS pixel_3333/NB2 pixel_3333/AMP_IN pixel_3333/SF_IB
+ pixel_3333/PIX_OUT pixel_3333/CSA_VREF pixel
Xpixel_3322 pixel_3322/gring pixel_3322/VDD pixel_3322/GND pixel_3322/VREF pixel_3322/ROW_SEL
+ pixel_3322/NB1 pixel_3322/VBIAS pixel_3322/NB2 pixel_3322/AMP_IN pixel_3322/SF_IB
+ pixel_3322/PIX_OUT pixel_3322/CSA_VREF pixel
Xpixel_3311 pixel_3311/gring pixel_3311/VDD pixel_3311/GND pixel_3311/VREF pixel_3311/ROW_SEL
+ pixel_3311/NB1 pixel_3311/VBIAS pixel_3311/NB2 pixel_3311/AMP_IN pixel_3311/SF_IB
+ pixel_3311/PIX_OUT pixel_3311/CSA_VREF pixel
Xpixel_3300 pixel_3300/gring pixel_3300/VDD pixel_3300/GND pixel_3300/VREF pixel_3300/ROW_SEL
+ pixel_3300/NB1 pixel_3300/VBIAS pixel_3300/NB2 pixel_3300/AMP_IN pixel_3300/SF_IB
+ pixel_3300/PIX_OUT pixel_3300/CSA_VREF pixel
Xpixel_4045 pixel_4045/gring pixel_4045/VDD pixel_4045/GND pixel_4045/VREF pixel_4045/ROW_SEL
+ pixel_4045/NB1 pixel_4045/VBIAS pixel_4045/NB2 pixel_4045/AMP_IN pixel_4045/SF_IB
+ pixel_4045/PIX_OUT pixel_4045/CSA_VREF pixel
Xpixel_4056 pixel_4056/gring pixel_4056/VDD pixel_4056/GND pixel_4056/VREF pixel_4056/ROW_SEL
+ pixel_4056/NB1 pixel_4056/VBIAS pixel_4056/NB2 pixel_4056/AMP_IN pixel_4056/SF_IB
+ pixel_4056/PIX_OUT pixel_4056/CSA_VREF pixel
Xpixel_4067 pixel_4067/gring pixel_4067/VDD pixel_4067/GND pixel_4067/VREF pixel_4067/ROW_SEL
+ pixel_4067/NB1 pixel_4067/VBIAS pixel_4067/NB2 pixel_4067/AMP_IN pixel_4067/SF_IB
+ pixel_4067/PIX_OUT pixel_4067/CSA_VREF pixel
Xpixel_4078 pixel_4078/gring pixel_4078/VDD pixel_4078/GND pixel_4078/VREF pixel_4078/ROW_SEL
+ pixel_4078/NB1 pixel_4078/VBIAS pixel_4078/NB2 pixel_4078/AMP_IN pixel_4078/SF_IB
+ pixel_4078/PIX_OUT pixel_4078/CSA_VREF pixel
Xpixel_2621 pixel_2621/gring pixel_2621/VDD pixel_2621/GND pixel_2621/VREF pixel_2621/ROW_SEL
+ pixel_2621/NB1 pixel_2621/VBIAS pixel_2621/NB2 pixel_2621/AMP_IN pixel_2621/SF_IB
+ pixel_2621/PIX_OUT pixel_2621/CSA_VREF pixel
Xpixel_2610 pixel_2610/gring pixel_2610/VDD pixel_2610/GND pixel_2610/VREF pixel_2610/ROW_SEL
+ pixel_2610/NB1 pixel_2610/VBIAS pixel_2610/NB2 pixel_2610/AMP_IN pixel_2610/SF_IB
+ pixel_2610/PIX_OUT pixel_2610/CSA_VREF pixel
Xpixel_3366 pixel_3366/gring pixel_3366/VDD pixel_3366/GND pixel_3366/VREF pixel_3366/ROW_SEL
+ pixel_3366/NB1 pixel_3366/VBIAS pixel_3366/NB2 pixel_3366/AMP_IN pixel_3366/SF_IB
+ pixel_3366/PIX_OUT pixel_3366/CSA_VREF pixel
Xpixel_3355 pixel_3355/gring pixel_3355/VDD pixel_3355/GND pixel_3355/VREF pixel_3355/ROW_SEL
+ pixel_3355/NB1 pixel_3355/VBIAS pixel_3355/NB2 pixel_3355/AMP_IN pixel_3355/SF_IB
+ pixel_3355/PIX_OUT pixel_3355/CSA_VREF pixel
Xpixel_3344 pixel_3344/gring pixel_3344/VDD pixel_3344/GND pixel_3344/VREF pixel_3344/ROW_SEL
+ pixel_3344/NB1 pixel_3344/VBIAS pixel_3344/NB2 pixel_3344/AMP_IN pixel_3344/SF_IB
+ pixel_3344/PIX_OUT pixel_3344/CSA_VREF pixel
Xpixel_4089 pixel_4089/gring pixel_4089/VDD pixel_4089/GND pixel_4089/VREF pixel_4089/ROW_SEL
+ pixel_4089/NB1 pixel_4089/VBIAS pixel_4089/NB2 pixel_4089/AMP_IN pixel_4089/SF_IB
+ pixel_4089/PIX_OUT pixel_4089/CSA_VREF pixel
Xpixel_1920 pixel_1920/gring pixel_1920/VDD pixel_1920/GND pixel_1920/VREF pixel_1920/ROW_SEL
+ pixel_1920/NB1 pixel_1920/VBIAS pixel_1920/NB2 pixel_1920/AMP_IN pixel_1920/SF_IB
+ pixel_1920/PIX_OUT pixel_1920/CSA_VREF pixel
Xpixel_2654 pixel_2654/gring pixel_2654/VDD pixel_2654/GND pixel_2654/VREF pixel_2654/ROW_SEL
+ pixel_2654/NB1 pixel_2654/VBIAS pixel_2654/NB2 pixel_2654/AMP_IN pixel_2654/SF_IB
+ pixel_2654/PIX_OUT pixel_2654/CSA_VREF pixel
Xpixel_2643 pixel_2643/gring pixel_2643/VDD pixel_2643/GND pixel_2643/VREF pixel_2643/ROW_SEL
+ pixel_2643/NB1 pixel_2643/VBIAS pixel_2643/NB2 pixel_2643/AMP_IN pixel_2643/SF_IB
+ pixel_2643/PIX_OUT pixel_2643/CSA_VREF pixel
Xpixel_2632 pixel_2632/gring pixel_2632/VDD pixel_2632/GND pixel_2632/VREF pixel_2632/ROW_SEL
+ pixel_2632/NB1 pixel_2632/VBIAS pixel_2632/NB2 pixel_2632/AMP_IN pixel_2632/SF_IB
+ pixel_2632/PIX_OUT pixel_2632/CSA_VREF pixel
Xpixel_3399 pixel_3399/gring pixel_3399/VDD pixel_3399/GND pixel_3399/VREF pixel_3399/ROW_SEL
+ pixel_3399/NB1 pixel_3399/VBIAS pixel_3399/NB2 pixel_3399/AMP_IN pixel_3399/SF_IB
+ pixel_3399/PIX_OUT pixel_3399/CSA_VREF pixel
Xpixel_3388 pixel_3388/gring pixel_3388/VDD pixel_3388/GND pixel_3388/VREF pixel_3388/ROW_SEL
+ pixel_3388/NB1 pixel_3388/VBIAS pixel_3388/NB2 pixel_3388/AMP_IN pixel_3388/SF_IB
+ pixel_3388/PIX_OUT pixel_3388/CSA_VREF pixel
Xpixel_3377 pixel_3377/gring pixel_3377/VDD pixel_3377/GND pixel_3377/VREF pixel_3377/ROW_SEL
+ pixel_3377/NB1 pixel_3377/VBIAS pixel_3377/NB2 pixel_3377/AMP_IN pixel_3377/SF_IB
+ pixel_3377/PIX_OUT pixel_3377/CSA_VREF pixel
Xpixel_1953 pixel_1953/gring pixel_1953/VDD pixel_1953/GND pixel_1953/VREF pixel_1953/ROW_SEL
+ pixel_1953/NB1 pixel_1953/VBIAS pixel_1953/NB2 pixel_1953/AMP_IN pixel_1953/SF_IB
+ pixel_1953/PIX_OUT pixel_1953/CSA_VREF pixel
Xpixel_1942 pixel_1942/gring pixel_1942/VDD pixel_1942/GND pixel_1942/VREF pixel_1942/ROW_SEL
+ pixel_1942/NB1 pixel_1942/VBIAS pixel_1942/NB2 pixel_1942/AMP_IN pixel_1942/SF_IB
+ pixel_1942/PIX_OUT pixel_1942/CSA_VREF pixel
Xpixel_1931 pixel_1931/gring pixel_1931/VDD pixel_1931/GND pixel_1931/VREF pixel_1931/ROW_SEL
+ pixel_1931/NB1 pixel_1931/VBIAS pixel_1931/NB2 pixel_1931/AMP_IN pixel_1931/SF_IB
+ pixel_1931/PIX_OUT pixel_1931/CSA_VREF pixel
Xpixel_2698 pixel_2698/gring pixel_2698/VDD pixel_2698/GND pixel_2698/VREF pixel_2698/ROW_SEL
+ pixel_2698/NB1 pixel_2698/VBIAS pixel_2698/NB2 pixel_2698/AMP_IN pixel_2698/SF_IB
+ pixel_2698/PIX_OUT pixel_2698/CSA_VREF pixel
Xpixel_2687 pixel_2687/gring pixel_2687/VDD pixel_2687/GND pixel_2687/VREF pixel_2687/ROW_SEL
+ pixel_2687/NB1 pixel_2687/VBIAS pixel_2687/NB2 pixel_2687/AMP_IN pixel_2687/SF_IB
+ pixel_2687/PIX_OUT pixel_2687/CSA_VREF pixel
Xpixel_2676 pixel_2676/gring pixel_2676/VDD pixel_2676/GND pixel_2676/VREF pixel_2676/ROW_SEL
+ pixel_2676/NB1 pixel_2676/VBIAS pixel_2676/NB2 pixel_2676/AMP_IN pixel_2676/SF_IB
+ pixel_2676/PIX_OUT pixel_2676/CSA_VREF pixel
Xpixel_2665 pixel_2665/gring pixel_2665/VDD pixel_2665/GND pixel_2665/VREF pixel_2665/ROW_SEL
+ pixel_2665/NB1 pixel_2665/VBIAS pixel_2665/NB2 pixel_2665/AMP_IN pixel_2665/SF_IB
+ pixel_2665/PIX_OUT pixel_2665/CSA_VREF pixel
Xpixel_1986 pixel_1986/gring pixel_1986/VDD pixel_1986/GND pixel_1986/VREF pixel_1986/ROW_SEL
+ pixel_1986/NB1 pixel_1986/VBIAS pixel_1986/NB2 pixel_1986/AMP_IN pixel_1986/SF_IB
+ pixel_1986/PIX_OUT pixel_1986/CSA_VREF pixel
Xpixel_1975 pixel_1975/gring pixel_1975/VDD pixel_1975/GND pixel_1975/VREF pixel_1975/ROW_SEL
+ pixel_1975/NB1 pixel_1975/VBIAS pixel_1975/NB2 pixel_1975/AMP_IN pixel_1975/SF_IB
+ pixel_1975/PIX_OUT pixel_1975/CSA_VREF pixel
Xpixel_1964 pixel_1964/gring pixel_1964/VDD pixel_1964/GND pixel_1964/VREF pixel_1964/ROW_SEL
+ pixel_1964/NB1 pixel_1964/VBIAS pixel_1964/NB2 pixel_1964/AMP_IN pixel_1964/SF_IB
+ pixel_1964/PIX_OUT pixel_1964/CSA_VREF pixel
Xpixel_1997 pixel_1997/gring pixel_1997/VDD pixel_1997/GND pixel_1997/VREF pixel_1997/ROW_SEL
+ pixel_1997/NB1 pixel_1997/VBIAS pixel_1997/NB2 pixel_1997/AMP_IN pixel_1997/SF_IB
+ pixel_1997/PIX_OUT pixel_1997/CSA_VREF pixel
Xpixel_5280 pixel_5280/gring pixel_5280/VDD pixel_5280/GND pixel_5280/VREF pixel_5280/ROW_SEL
+ pixel_5280/NB1 pixel_5280/VBIAS pixel_5280/NB2 pixel_5280/AMP_IN pixel_5280/SF_IB
+ pixel_5280/PIX_OUT pixel_5280/CSA_VREF pixel
Xpixel_5291 pixel_5291/gring pixel_5291/VDD pixel_5291/GND pixel_5291/VREF pixel_5291/ROW_SEL
+ pixel_5291/NB1 pixel_5291/VBIAS pixel_5291/NB2 pixel_5291/AMP_IN pixel_5291/SF_IB
+ pixel_5291/PIX_OUT pixel_5291/CSA_VREF pixel
Xpixel_4590 pixel_4590/gring pixel_4590/VDD pixel_4590/GND pixel_4590/VREF pixel_4590/ROW_SEL
+ pixel_4590/NB1 pixel_4590/VBIAS pixel_4590/NB2 pixel_4590/AMP_IN pixel_4590/SF_IB
+ pixel_4590/PIX_OUT pixel_4590/CSA_VREF pixel
Xpixel_6909 pixel_6909/gring pixel_6909/VDD pixel_6909/GND pixel_6909/VREF pixel_6909/ROW_SEL
+ pixel_6909/NB1 pixel_6909/VBIAS pixel_6909/NB2 pixel_6909/AMP_IN pixel_6909/SF_IB
+ pixel_6909/PIX_OUT pixel_6909/CSA_VREF pixel
Xpixel_1205 pixel_1205/gring pixel_1205/VDD pixel_1205/GND pixel_1205/VREF pixel_1205/ROW_SEL
+ pixel_1205/NB1 pixel_1205/VBIAS pixel_1205/NB2 pixel_1205/AMP_IN pixel_1205/SF_IB
+ pixel_1205/PIX_OUT pixel_1205/CSA_VREF pixel
Xpixel_1249 pixel_1249/gring pixel_1249/VDD pixel_1249/GND pixel_1249/VREF pixel_1249/ROW_SEL
+ pixel_1249/NB1 pixel_1249/VBIAS pixel_1249/NB2 pixel_1249/AMP_IN pixel_1249/SF_IB
+ pixel_1249/PIX_OUT pixel_1249/CSA_VREF pixel
Xpixel_1238 pixel_1238/gring pixel_1238/VDD pixel_1238/GND pixel_1238/VREF pixel_1238/ROW_SEL
+ pixel_1238/NB1 pixel_1238/VBIAS pixel_1238/NB2 pixel_1238/AMP_IN pixel_1238/SF_IB
+ pixel_1238/PIX_OUT pixel_1238/CSA_VREF pixel
Xpixel_1227 pixel_1227/gring pixel_1227/VDD pixel_1227/GND pixel_1227/VREF pixel_1227/ROW_SEL
+ pixel_1227/NB1 pixel_1227/VBIAS pixel_1227/NB2 pixel_1227/AMP_IN pixel_1227/SF_IB
+ pixel_1227/PIX_OUT pixel_1227/CSA_VREF pixel
Xpixel_1216 pixel_1216/gring pixel_1216/VDD pixel_1216/GND pixel_1216/VREF pixel_1216/ROW_SEL
+ pixel_1216/NB1 pixel_1216/VBIAS pixel_1216/NB2 pixel_1216/AMP_IN pixel_1216/SF_IB
+ pixel_1216/PIX_OUT pixel_1216/CSA_VREF pixel
Xpixel_9513 pixel_9513/gring pixel_9513/VDD pixel_9513/GND pixel_9513/VREF pixel_9513/ROW_SEL
+ pixel_9513/NB1 pixel_9513/VBIAS pixel_9513/NB2 pixel_9513/AMP_IN pixel_9513/SF_IB
+ pixel_9513/PIX_OUT pixel_9513/CSA_VREF pixel
Xpixel_9502 pixel_9502/gring pixel_9502/VDD pixel_9502/GND pixel_9502/VREF pixel_9502/ROW_SEL
+ pixel_9502/NB1 pixel_9502/VBIAS pixel_9502/NB2 pixel_9502/AMP_IN pixel_9502/SF_IB
+ pixel_9502/PIX_OUT pixel_9502/CSA_VREF pixel
Xpixel_8812 pixel_8812/gring pixel_8812/VDD pixel_8812/GND pixel_8812/VREF pixel_8812/ROW_SEL
+ pixel_8812/NB1 pixel_8812/VBIAS pixel_8812/NB2 pixel_8812/AMP_IN pixel_8812/SF_IB
+ pixel_8812/PIX_OUT pixel_8812/CSA_VREF pixel
Xpixel_8801 pixel_8801/gring pixel_8801/VDD pixel_8801/GND pixel_8801/VREF pixel_8801/ROW_SEL
+ pixel_8801/NB1 pixel_8801/VBIAS pixel_8801/NB2 pixel_8801/AMP_IN pixel_8801/SF_IB
+ pixel_8801/PIX_OUT pixel_8801/CSA_VREF pixel
Xpixel_9557 pixel_9557/gring pixel_9557/VDD pixel_9557/GND pixel_9557/VREF pixel_9557/ROW_SEL
+ pixel_9557/NB1 pixel_9557/VBIAS pixel_9557/NB2 pixel_9557/AMP_IN pixel_9557/SF_IB
+ pixel_9557/PIX_OUT pixel_9557/CSA_VREF pixel
Xpixel_9546 pixel_9546/gring pixel_9546/VDD pixel_9546/GND pixel_9546/VREF pixel_9546/ROW_SEL
+ pixel_9546/NB1 pixel_9546/VBIAS pixel_9546/NB2 pixel_9546/AMP_IN pixel_9546/SF_IB
+ pixel_9546/PIX_OUT pixel_9546/CSA_VREF pixel
Xpixel_9535 pixel_9535/gring pixel_9535/VDD pixel_9535/GND pixel_9535/VREF pixel_9535/ROW_SEL
+ pixel_9535/NB1 pixel_9535/VBIAS pixel_9535/NB2 pixel_9535/AMP_IN pixel_9535/SF_IB
+ pixel_9535/PIX_OUT pixel_9535/CSA_VREF pixel
Xpixel_9524 pixel_9524/gring pixel_9524/VDD pixel_9524/GND pixel_9524/VREF pixel_9524/ROW_SEL
+ pixel_9524/NB1 pixel_9524/VBIAS pixel_9524/NB2 pixel_9524/AMP_IN pixel_9524/SF_IB
+ pixel_9524/PIX_OUT pixel_9524/CSA_VREF pixel
Xpixel_8845 pixel_8845/gring pixel_8845/VDD pixel_8845/GND pixel_8845/VREF pixel_8845/ROW_SEL
+ pixel_8845/NB1 pixel_8845/VBIAS pixel_8845/NB2 pixel_8845/AMP_IN pixel_8845/SF_IB
+ pixel_8845/PIX_OUT pixel_8845/CSA_VREF pixel
Xpixel_8834 pixel_8834/gring pixel_8834/VDD pixel_8834/GND pixel_8834/VREF pixel_8834/ROW_SEL
+ pixel_8834/NB1 pixel_8834/VBIAS pixel_8834/NB2 pixel_8834/AMP_IN pixel_8834/SF_IB
+ pixel_8834/PIX_OUT pixel_8834/CSA_VREF pixel
Xpixel_8823 pixel_8823/gring pixel_8823/VDD pixel_8823/GND pixel_8823/VREF pixel_8823/ROW_SEL
+ pixel_8823/NB1 pixel_8823/VBIAS pixel_8823/NB2 pixel_8823/AMP_IN pixel_8823/SF_IB
+ pixel_8823/PIX_OUT pixel_8823/CSA_VREF pixel
Xpixel_9579 pixel_9579/gring pixel_9579/VDD pixel_9579/GND pixel_9579/VREF pixel_9579/ROW_SEL
+ pixel_9579/NB1 pixel_9579/VBIAS pixel_9579/NB2 pixel_9579/AMP_IN pixel_9579/SF_IB
+ pixel_9579/PIX_OUT pixel_9579/CSA_VREF pixel
Xpixel_9568 pixel_9568/gring pixel_9568/VDD pixel_9568/GND pixel_9568/VREF pixel_9568/ROW_SEL
+ pixel_9568/NB1 pixel_9568/VBIAS pixel_9568/NB2 pixel_9568/AMP_IN pixel_9568/SF_IB
+ pixel_9568/PIX_OUT pixel_9568/CSA_VREF pixel
Xpixel_8878 pixel_8878/gring pixel_8878/VDD pixel_8878/GND pixel_8878/VREF pixel_8878/ROW_SEL
+ pixel_8878/NB1 pixel_8878/VBIAS pixel_8878/NB2 pixel_8878/AMP_IN pixel_8878/SF_IB
+ pixel_8878/PIX_OUT pixel_8878/CSA_VREF pixel
Xpixel_8867 pixel_8867/gring pixel_8867/VDD pixel_8867/GND pixel_8867/VREF pixel_8867/ROW_SEL
+ pixel_8867/NB1 pixel_8867/VBIAS pixel_8867/NB2 pixel_8867/AMP_IN pixel_8867/SF_IB
+ pixel_8867/PIX_OUT pixel_8867/CSA_VREF pixel
Xpixel_8856 pixel_8856/gring pixel_8856/VDD pixel_8856/GND pixel_8856/VREF pixel_8856/ROW_SEL
+ pixel_8856/NB1 pixel_8856/VBIAS pixel_8856/NB2 pixel_8856/AMP_IN pixel_8856/SF_IB
+ pixel_8856/PIX_OUT pixel_8856/CSA_VREF pixel
Xpixel_8889 pixel_8889/gring pixel_8889/VDD pixel_8889/GND pixel_8889/VREF pixel_8889/ROW_SEL
+ pixel_8889/NB1 pixel_8889/VBIAS pixel_8889/NB2 pixel_8889/AMP_IN pixel_8889/SF_IB
+ pixel_8889/PIX_OUT pixel_8889/CSA_VREF pixel
Xpixel_3141 pixel_3141/gring pixel_3141/VDD pixel_3141/GND pixel_3141/VREF pixel_3141/ROW_SEL
+ pixel_3141/NB1 pixel_3141/VBIAS pixel_3141/NB2 pixel_3141/AMP_IN pixel_3141/SF_IB
+ pixel_3141/PIX_OUT pixel_3141/CSA_VREF pixel
Xpixel_3130 pixel_3130/gring pixel_3130/VDD pixel_3130/GND pixel_3130/VREF pixel_3130/ROW_SEL
+ pixel_3130/NB1 pixel_3130/VBIAS pixel_3130/NB2 pixel_3130/AMP_IN pixel_3130/SF_IB
+ pixel_3130/PIX_OUT pixel_3130/CSA_VREF pixel
Xpixel_3174 pixel_3174/gring pixel_3174/VDD pixel_3174/GND pixel_3174/VREF pixel_3174/ROW_SEL
+ pixel_3174/NB1 pixel_3174/VBIAS pixel_3174/NB2 pixel_3174/AMP_IN pixel_3174/SF_IB
+ pixel_3174/PIX_OUT pixel_3174/CSA_VREF pixel
Xpixel_3163 pixel_3163/gring pixel_3163/VDD pixel_3163/GND pixel_3163/VREF pixel_3163/ROW_SEL
+ pixel_3163/NB1 pixel_3163/VBIAS pixel_3163/NB2 pixel_3163/AMP_IN pixel_3163/SF_IB
+ pixel_3163/PIX_OUT pixel_3163/CSA_VREF pixel
Xpixel_3152 pixel_3152/gring pixel_3152/VDD pixel_3152/GND pixel_3152/VREF pixel_3152/ROW_SEL
+ pixel_3152/NB1 pixel_3152/VBIAS pixel_3152/NB2 pixel_3152/AMP_IN pixel_3152/SF_IB
+ pixel_3152/PIX_OUT pixel_3152/CSA_VREF pixel
Xpixel_2473 pixel_2473/gring pixel_2473/VDD pixel_2473/GND pixel_2473/VREF pixel_2473/ROW_SEL
+ pixel_2473/NB1 pixel_2473/VBIAS pixel_2473/NB2 pixel_2473/AMP_IN pixel_2473/SF_IB
+ pixel_2473/PIX_OUT pixel_2473/CSA_VREF pixel
Xpixel_2462 pixel_2462/gring pixel_2462/VDD pixel_2462/GND pixel_2462/VREF pixel_2462/ROW_SEL
+ pixel_2462/NB1 pixel_2462/VBIAS pixel_2462/NB2 pixel_2462/AMP_IN pixel_2462/SF_IB
+ pixel_2462/PIX_OUT pixel_2462/CSA_VREF pixel
Xpixel_2451 pixel_2451/gring pixel_2451/VDD pixel_2451/GND pixel_2451/VREF pixel_2451/ROW_SEL
+ pixel_2451/NB1 pixel_2451/VBIAS pixel_2451/NB2 pixel_2451/AMP_IN pixel_2451/SF_IB
+ pixel_2451/PIX_OUT pixel_2451/CSA_VREF pixel
Xpixel_2440 pixel_2440/gring pixel_2440/VDD pixel_2440/GND pixel_2440/VREF pixel_2440/ROW_SEL
+ pixel_2440/NB1 pixel_2440/VBIAS pixel_2440/NB2 pixel_2440/AMP_IN pixel_2440/SF_IB
+ pixel_2440/PIX_OUT pixel_2440/CSA_VREF pixel
Xpixel_3196 pixel_3196/gring pixel_3196/VDD pixel_3196/GND pixel_3196/VREF pixel_3196/ROW_SEL
+ pixel_3196/NB1 pixel_3196/VBIAS pixel_3196/NB2 pixel_3196/AMP_IN pixel_3196/SF_IB
+ pixel_3196/PIX_OUT pixel_3196/CSA_VREF pixel
Xpixel_3185 pixel_3185/gring pixel_3185/VDD pixel_3185/GND pixel_3185/VREF pixel_3185/ROW_SEL
+ pixel_3185/NB1 pixel_3185/VBIAS pixel_3185/NB2 pixel_3185/AMP_IN pixel_3185/SF_IB
+ pixel_3185/PIX_OUT pixel_3185/CSA_VREF pixel
Xpixel_1761 pixel_1761/gring pixel_1761/VDD pixel_1761/GND pixel_1761/VREF pixel_1761/ROW_SEL
+ pixel_1761/NB1 pixel_1761/VBIAS pixel_1761/NB2 pixel_1761/AMP_IN pixel_1761/SF_IB
+ pixel_1761/PIX_OUT pixel_1761/CSA_VREF pixel
Xpixel_1750 pixel_1750/gring pixel_1750/VDD pixel_1750/GND pixel_1750/VREF pixel_1750/ROW_SEL
+ pixel_1750/NB1 pixel_1750/VBIAS pixel_1750/NB2 pixel_1750/AMP_IN pixel_1750/SF_IB
+ pixel_1750/PIX_OUT pixel_1750/CSA_VREF pixel
Xpixel_2495 pixel_2495/gring pixel_2495/VDD pixel_2495/GND pixel_2495/VREF pixel_2495/ROW_SEL
+ pixel_2495/NB1 pixel_2495/VBIAS pixel_2495/NB2 pixel_2495/AMP_IN pixel_2495/SF_IB
+ pixel_2495/PIX_OUT pixel_2495/CSA_VREF pixel
Xpixel_2484 pixel_2484/gring pixel_2484/VDD pixel_2484/GND pixel_2484/VREF pixel_2484/ROW_SEL
+ pixel_2484/NB1 pixel_2484/VBIAS pixel_2484/NB2 pixel_2484/AMP_IN pixel_2484/SF_IB
+ pixel_2484/PIX_OUT pixel_2484/CSA_VREF pixel
Xpixel_1794 pixel_1794/gring pixel_1794/VDD pixel_1794/GND pixel_1794/VREF pixel_1794/ROW_SEL
+ pixel_1794/NB1 pixel_1794/VBIAS pixel_1794/NB2 pixel_1794/AMP_IN pixel_1794/SF_IB
+ pixel_1794/PIX_OUT pixel_1794/CSA_VREF pixel
Xpixel_1783 pixel_1783/gring pixel_1783/VDD pixel_1783/GND pixel_1783/VREF pixel_1783/ROW_SEL
+ pixel_1783/NB1 pixel_1783/VBIAS pixel_1783/NB2 pixel_1783/AMP_IN pixel_1783/SF_IB
+ pixel_1783/PIX_OUT pixel_1783/CSA_VREF pixel
Xpixel_1772 pixel_1772/gring pixel_1772/VDD pixel_1772/GND pixel_1772/VREF pixel_1772/ROW_SEL
+ pixel_1772/NB1 pixel_1772/VBIAS pixel_1772/NB2 pixel_1772/AMP_IN pixel_1772/SF_IB
+ pixel_1772/PIX_OUT pixel_1772/CSA_VREF pixel
Xpixel_809 pixel_809/gring pixel_809/VDD pixel_809/GND pixel_809/VREF pixel_809/ROW_SEL
+ pixel_809/NB1 pixel_809/VBIAS pixel_809/NB2 pixel_809/AMP_IN pixel_809/SF_IB pixel_809/PIX_OUT
+ pixel_809/CSA_VREF pixel
Xpixel_8108 pixel_8108/gring pixel_8108/VDD pixel_8108/GND pixel_8108/VREF pixel_8108/ROW_SEL
+ pixel_8108/NB1 pixel_8108/VBIAS pixel_8108/NB2 pixel_8108/AMP_IN pixel_8108/SF_IB
+ pixel_8108/PIX_OUT pixel_8108/CSA_VREF pixel
Xpixel_8119 pixel_8119/gring pixel_8119/VDD pixel_8119/GND pixel_8119/VREF pixel_8119/ROW_SEL
+ pixel_8119/NB1 pixel_8119/VBIAS pixel_8119/NB2 pixel_8119/AMP_IN pixel_8119/SF_IB
+ pixel_8119/PIX_OUT pixel_8119/CSA_VREF pixel
Xpixel_7407 pixel_7407/gring pixel_7407/VDD pixel_7407/GND pixel_7407/VREF pixel_7407/ROW_SEL
+ pixel_7407/NB1 pixel_7407/VBIAS pixel_7407/NB2 pixel_7407/AMP_IN pixel_7407/SF_IB
+ pixel_7407/PIX_OUT pixel_7407/CSA_VREF pixel
Xpixel_7418 pixel_7418/gring pixel_7418/VDD pixel_7418/GND pixel_7418/VREF pixel_7418/ROW_SEL
+ pixel_7418/NB1 pixel_7418/VBIAS pixel_7418/NB2 pixel_7418/AMP_IN pixel_7418/SF_IB
+ pixel_7418/PIX_OUT pixel_7418/CSA_VREF pixel
Xpixel_7429 pixel_7429/gring pixel_7429/VDD pixel_7429/GND pixel_7429/VREF pixel_7429/ROW_SEL
+ pixel_7429/NB1 pixel_7429/VBIAS pixel_7429/NB2 pixel_7429/AMP_IN pixel_7429/SF_IB
+ pixel_7429/PIX_OUT pixel_7429/CSA_VREF pixel
Xpixel_6706 pixel_6706/gring pixel_6706/VDD pixel_6706/GND pixel_6706/VREF pixel_6706/ROW_SEL
+ pixel_6706/NB1 pixel_6706/VBIAS pixel_6706/NB2 pixel_6706/AMP_IN pixel_6706/SF_IB
+ pixel_6706/PIX_OUT pixel_6706/CSA_VREF pixel
Xpixel_6717 pixel_6717/gring pixel_6717/VDD pixel_6717/GND pixel_6717/VREF pixel_6717/ROW_SEL
+ pixel_6717/NB1 pixel_6717/VBIAS pixel_6717/NB2 pixel_6717/AMP_IN pixel_6717/SF_IB
+ pixel_6717/PIX_OUT pixel_6717/CSA_VREF pixel
Xpixel_6728 pixel_6728/gring pixel_6728/VDD pixel_6728/GND pixel_6728/VREF pixel_6728/ROW_SEL
+ pixel_6728/NB1 pixel_6728/VBIAS pixel_6728/NB2 pixel_6728/AMP_IN pixel_6728/SF_IB
+ pixel_6728/PIX_OUT pixel_6728/CSA_VREF pixel
Xpixel_6739 pixel_6739/gring pixel_6739/VDD pixel_6739/GND pixel_6739/VREF pixel_6739/ROW_SEL
+ pixel_6739/NB1 pixel_6739/VBIAS pixel_6739/NB2 pixel_6739/AMP_IN pixel_6739/SF_IB
+ pixel_6739/PIX_OUT pixel_6739/CSA_VREF pixel
Xpixel_1024 pixel_1024/gring pixel_1024/VDD pixel_1024/GND pixel_1024/VREF pixel_1024/ROW_SEL
+ pixel_1024/NB1 pixel_1024/VBIAS pixel_1024/NB2 pixel_1024/AMP_IN pixel_1024/SF_IB
+ pixel_1024/PIX_OUT pixel_1024/CSA_VREF pixel
Xpixel_1013 pixel_1013/gring pixel_1013/VDD pixel_1013/GND pixel_1013/VREF pixel_1013/ROW_SEL
+ pixel_1013/NB1 pixel_1013/VBIAS pixel_1013/NB2 pixel_1013/AMP_IN pixel_1013/SF_IB
+ pixel_1013/PIX_OUT pixel_1013/CSA_VREF pixel
Xpixel_1002 pixel_1002/gring pixel_1002/VDD pixel_1002/GND pixel_1002/VREF pixel_1002/ROW_SEL
+ pixel_1002/NB1 pixel_1002/VBIAS pixel_1002/NB2 pixel_1002/AMP_IN pixel_1002/SF_IB
+ pixel_1002/PIX_OUT pixel_1002/CSA_VREF pixel
Xpixel_1057 pixel_1057/gring pixel_1057/VDD pixel_1057/GND pixel_1057/VREF pixel_1057/ROW_SEL
+ pixel_1057/NB1 pixel_1057/VBIAS pixel_1057/NB2 pixel_1057/AMP_IN pixel_1057/SF_IB
+ pixel_1057/PIX_OUT pixel_1057/CSA_VREF pixel
Xpixel_1046 pixel_1046/gring pixel_1046/VDD pixel_1046/GND pixel_1046/VREF pixel_1046/ROW_SEL
+ pixel_1046/NB1 pixel_1046/VBIAS pixel_1046/NB2 pixel_1046/AMP_IN pixel_1046/SF_IB
+ pixel_1046/PIX_OUT pixel_1046/CSA_VREF pixel
Xpixel_1035 pixel_1035/gring pixel_1035/VDD pixel_1035/GND pixel_1035/VREF pixel_1035/ROW_SEL
+ pixel_1035/NB1 pixel_1035/VBIAS pixel_1035/NB2 pixel_1035/AMP_IN pixel_1035/SF_IB
+ pixel_1035/PIX_OUT pixel_1035/CSA_VREF pixel
Xpixel_1079 pixel_1079/gring pixel_1079/VDD pixel_1079/GND pixel_1079/VREF pixel_1079/ROW_SEL
+ pixel_1079/NB1 pixel_1079/VBIAS pixel_1079/NB2 pixel_1079/AMP_IN pixel_1079/SF_IB
+ pixel_1079/PIX_OUT pixel_1079/CSA_VREF pixel
Xpixel_1068 pixel_1068/gring pixel_1068/VDD pixel_1068/GND pixel_1068/VREF pixel_1068/ROW_SEL
+ pixel_1068/NB1 pixel_1068/VBIAS pixel_1068/NB2 pixel_1068/AMP_IN pixel_1068/SF_IB
+ pixel_1068/PIX_OUT pixel_1068/CSA_VREF pixel
Xpixel_9321 pixel_9321/gring pixel_9321/VDD pixel_9321/GND pixel_9321/VREF pixel_9321/ROW_SEL
+ pixel_9321/NB1 pixel_9321/VBIAS pixel_9321/NB2 pixel_9321/AMP_IN pixel_9321/SF_IB
+ pixel_9321/PIX_OUT pixel_9321/CSA_VREF pixel
Xpixel_9310 pixel_9310/gring pixel_9310/VDD pixel_9310/GND pixel_9310/VREF pixel_9310/ROW_SEL
+ pixel_9310/NB1 pixel_9310/VBIAS pixel_9310/NB2 pixel_9310/AMP_IN pixel_9310/SF_IB
+ pixel_9310/PIX_OUT pixel_9310/CSA_VREF pixel
Xpixel_8620 pixel_8620/gring pixel_8620/VDD pixel_8620/GND pixel_8620/VREF pixel_8620/ROW_SEL
+ pixel_8620/NB1 pixel_8620/VBIAS pixel_8620/NB2 pixel_8620/AMP_IN pixel_8620/SF_IB
+ pixel_8620/PIX_OUT pixel_8620/CSA_VREF pixel
Xpixel_9365 pixel_9365/gring pixel_9365/VDD pixel_9365/GND pixel_9365/VREF pixel_9365/ROW_SEL
+ pixel_9365/NB1 pixel_9365/VBIAS pixel_9365/NB2 pixel_9365/AMP_IN pixel_9365/SF_IB
+ pixel_9365/PIX_OUT pixel_9365/CSA_VREF pixel
Xpixel_9354 pixel_9354/gring pixel_9354/VDD pixel_9354/GND pixel_9354/VREF pixel_9354/ROW_SEL
+ pixel_9354/NB1 pixel_9354/VBIAS pixel_9354/NB2 pixel_9354/AMP_IN pixel_9354/SF_IB
+ pixel_9354/PIX_OUT pixel_9354/CSA_VREF pixel
Xpixel_9343 pixel_9343/gring pixel_9343/VDD pixel_9343/GND pixel_9343/VREF pixel_9343/ROW_SEL
+ pixel_9343/NB1 pixel_9343/VBIAS pixel_9343/NB2 pixel_9343/AMP_IN pixel_9343/SF_IB
+ pixel_9343/PIX_OUT pixel_9343/CSA_VREF pixel
Xpixel_9332 pixel_9332/gring pixel_9332/VDD pixel_9332/GND pixel_9332/VREF pixel_9332/ROW_SEL
+ pixel_9332/NB1 pixel_9332/VBIAS pixel_9332/NB2 pixel_9332/AMP_IN pixel_9332/SF_IB
+ pixel_9332/PIX_OUT pixel_9332/CSA_VREF pixel
Xpixel_8653 pixel_8653/gring pixel_8653/VDD pixel_8653/GND pixel_8653/VREF pixel_8653/ROW_SEL
+ pixel_8653/NB1 pixel_8653/VBIAS pixel_8653/NB2 pixel_8653/AMP_IN pixel_8653/SF_IB
+ pixel_8653/PIX_OUT pixel_8653/CSA_VREF pixel
Xpixel_8642 pixel_8642/gring pixel_8642/VDD pixel_8642/GND pixel_8642/VREF pixel_8642/ROW_SEL
+ pixel_8642/NB1 pixel_8642/VBIAS pixel_8642/NB2 pixel_8642/AMP_IN pixel_8642/SF_IB
+ pixel_8642/PIX_OUT pixel_8642/CSA_VREF pixel
Xpixel_8631 pixel_8631/gring pixel_8631/VDD pixel_8631/GND pixel_8631/VREF pixel_8631/ROW_SEL
+ pixel_8631/NB1 pixel_8631/VBIAS pixel_8631/NB2 pixel_8631/AMP_IN pixel_8631/SF_IB
+ pixel_8631/PIX_OUT pixel_8631/CSA_VREF pixel
Xpixel_9398 pixel_9398/gring pixel_9398/VDD pixel_9398/GND pixel_9398/VREF pixel_9398/ROW_SEL
+ pixel_9398/NB1 pixel_9398/VBIAS pixel_9398/NB2 pixel_9398/AMP_IN pixel_9398/SF_IB
+ pixel_9398/PIX_OUT pixel_9398/CSA_VREF pixel
Xpixel_9387 pixel_9387/gring pixel_9387/VDD pixel_9387/GND pixel_9387/VREF pixel_9387/ROW_SEL
+ pixel_9387/NB1 pixel_9387/VBIAS pixel_9387/NB2 pixel_9387/AMP_IN pixel_9387/SF_IB
+ pixel_9387/PIX_OUT pixel_9387/CSA_VREF pixel
Xpixel_9376 pixel_9376/gring pixel_9376/VDD pixel_9376/GND pixel_9376/VREF pixel_9376/ROW_SEL
+ pixel_9376/NB1 pixel_9376/VBIAS pixel_9376/NB2 pixel_9376/AMP_IN pixel_9376/SF_IB
+ pixel_9376/PIX_OUT pixel_9376/CSA_VREF pixel
Xpixel_8697 pixel_8697/gring pixel_8697/VDD pixel_8697/GND pixel_8697/VREF pixel_8697/ROW_SEL
+ pixel_8697/NB1 pixel_8697/VBIAS pixel_8697/NB2 pixel_8697/AMP_IN pixel_8697/SF_IB
+ pixel_8697/PIX_OUT pixel_8697/CSA_VREF pixel
Xpixel_8686 pixel_8686/gring pixel_8686/VDD pixel_8686/GND pixel_8686/VREF pixel_8686/ROW_SEL
+ pixel_8686/NB1 pixel_8686/VBIAS pixel_8686/NB2 pixel_8686/AMP_IN pixel_8686/SF_IB
+ pixel_8686/PIX_OUT pixel_8686/CSA_VREF pixel
Xpixel_8675 pixel_8675/gring pixel_8675/VDD pixel_8675/GND pixel_8675/VREF pixel_8675/ROW_SEL
+ pixel_8675/NB1 pixel_8675/VBIAS pixel_8675/NB2 pixel_8675/AMP_IN pixel_8675/SF_IB
+ pixel_8675/PIX_OUT pixel_8675/CSA_VREF pixel
Xpixel_8664 pixel_8664/gring pixel_8664/VDD pixel_8664/GND pixel_8664/VREF pixel_8664/ROW_SEL
+ pixel_8664/NB1 pixel_8664/VBIAS pixel_8664/NB2 pixel_8664/AMP_IN pixel_8664/SF_IB
+ pixel_8664/PIX_OUT pixel_8664/CSA_VREF pixel
Xpixel_7930 pixel_7930/gring pixel_7930/VDD pixel_7930/GND pixel_7930/VREF pixel_7930/ROW_SEL
+ pixel_7930/NB1 pixel_7930/VBIAS pixel_7930/NB2 pixel_7930/AMP_IN pixel_7930/SF_IB
+ pixel_7930/PIX_OUT pixel_7930/CSA_VREF pixel
Xpixel_7941 pixel_7941/gring pixel_7941/VDD pixel_7941/GND pixel_7941/VREF pixel_7941/ROW_SEL
+ pixel_7941/NB1 pixel_7941/VBIAS pixel_7941/NB2 pixel_7941/AMP_IN pixel_7941/SF_IB
+ pixel_7941/PIX_OUT pixel_7941/CSA_VREF pixel
Xpixel_7952 pixel_7952/gring pixel_7952/VDD pixel_7952/GND pixel_7952/VREF pixel_7952/ROW_SEL
+ pixel_7952/NB1 pixel_7952/VBIAS pixel_7952/NB2 pixel_7952/AMP_IN pixel_7952/SF_IB
+ pixel_7952/PIX_OUT pixel_7952/CSA_VREF pixel
Xpixel_7963 pixel_7963/gring pixel_7963/VDD pixel_7963/GND pixel_7963/VREF pixel_7963/ROW_SEL
+ pixel_7963/NB1 pixel_7963/VBIAS pixel_7963/NB2 pixel_7963/AMP_IN pixel_7963/SF_IB
+ pixel_7963/PIX_OUT pixel_7963/CSA_VREF pixel
Xpixel_7974 pixel_7974/gring pixel_7974/VDD pixel_7974/GND pixel_7974/VREF pixel_7974/ROW_SEL
+ pixel_7974/NB1 pixel_7974/VBIAS pixel_7974/NB2 pixel_7974/AMP_IN pixel_7974/SF_IB
+ pixel_7974/PIX_OUT pixel_7974/CSA_VREF pixel
Xpixel_7985 pixel_7985/gring pixel_7985/VDD pixel_7985/GND pixel_7985/VREF pixel_7985/ROW_SEL
+ pixel_7985/NB1 pixel_7985/VBIAS pixel_7985/NB2 pixel_7985/AMP_IN pixel_7985/SF_IB
+ pixel_7985/PIX_OUT pixel_7985/CSA_VREF pixel
Xpixel_7996 pixel_7996/gring pixel_7996/VDD pixel_7996/GND pixel_7996/VREF pixel_7996/ROW_SEL
+ pixel_7996/NB1 pixel_7996/VBIAS pixel_7996/NB2 pixel_7996/AMP_IN pixel_7996/SF_IB
+ pixel_7996/PIX_OUT pixel_7996/CSA_VREF pixel
Xpixel_2281 pixel_2281/gring pixel_2281/VDD pixel_2281/GND pixel_2281/VREF pixel_2281/ROW_SEL
+ pixel_2281/NB1 pixel_2281/VBIAS pixel_2281/NB2 pixel_2281/AMP_IN pixel_2281/SF_IB
+ pixel_2281/PIX_OUT pixel_2281/CSA_VREF pixel
Xpixel_2270 pixel_2270/gring pixel_2270/VDD pixel_2270/GND pixel_2270/VREF pixel_2270/ROW_SEL
+ pixel_2270/NB1 pixel_2270/VBIAS pixel_2270/NB2 pixel_2270/AMP_IN pixel_2270/SF_IB
+ pixel_2270/PIX_OUT pixel_2270/CSA_VREF pixel
Xpixel_2292 pixel_2292/gring pixel_2292/VDD pixel_2292/GND pixel_2292/VREF pixel_2292/ROW_SEL
+ pixel_2292/NB1 pixel_2292/VBIAS pixel_2292/NB2 pixel_2292/AMP_IN pixel_2292/SF_IB
+ pixel_2292/PIX_OUT pixel_2292/CSA_VREF pixel
Xpixel_1591 pixel_1591/gring pixel_1591/VDD pixel_1591/GND pixel_1591/VREF pixel_1591/ROW_SEL
+ pixel_1591/NB1 pixel_1591/VBIAS pixel_1591/NB2 pixel_1591/AMP_IN pixel_1591/SF_IB
+ pixel_1591/PIX_OUT pixel_1591/CSA_VREF pixel
Xpixel_1580 pixel_1580/gring pixel_1580/VDD pixel_1580/GND pixel_1580/VREF pixel_1580/ROW_SEL
+ pixel_1580/NB1 pixel_1580/VBIAS pixel_1580/NB2 pixel_1580/AMP_IN pixel_1580/SF_IB
+ pixel_1580/PIX_OUT pixel_1580/CSA_VREF pixel
Xpixel_639 pixel_639/gring pixel_639/VDD pixel_639/GND pixel_639/VREF pixel_639/ROW_SEL
+ pixel_639/NB1 pixel_639/VBIAS pixel_639/NB2 pixel_639/AMP_IN pixel_639/SF_IB pixel_639/PIX_OUT
+ pixel_639/CSA_VREF pixel
Xpixel_628 pixel_628/gring pixel_628/VDD pixel_628/GND pixel_628/VREF pixel_628/ROW_SEL
+ pixel_628/NB1 pixel_628/VBIAS pixel_628/NB2 pixel_628/AMP_IN pixel_628/SF_IB pixel_628/PIX_OUT
+ pixel_628/CSA_VREF pixel
Xpixel_617 pixel_617/gring pixel_617/VDD pixel_617/GND pixel_617/VREF pixel_617/ROW_SEL
+ pixel_617/NB1 pixel_617/VBIAS pixel_617/NB2 pixel_617/AMP_IN pixel_617/SF_IB pixel_617/PIX_OUT
+ pixel_617/CSA_VREF pixel
Xpixel_606 pixel_606/gring pixel_606/VDD pixel_606/GND pixel_606/VREF pixel_606/ROW_SEL
+ pixel_606/NB1 pixel_606/VBIAS pixel_606/NB2 pixel_606/AMP_IN pixel_606/SF_IB pixel_606/PIX_OUT
+ pixel_606/CSA_VREF pixel
Xpixel_7204 pixel_7204/gring pixel_7204/VDD pixel_7204/GND pixel_7204/VREF pixel_7204/ROW_SEL
+ pixel_7204/NB1 pixel_7204/VBIAS pixel_7204/NB2 pixel_7204/AMP_IN pixel_7204/SF_IB
+ pixel_7204/PIX_OUT pixel_7204/CSA_VREF pixel
Xpixel_7215 pixel_7215/gring pixel_7215/VDD pixel_7215/GND pixel_7215/VREF pixel_7215/ROW_SEL
+ pixel_7215/NB1 pixel_7215/VBIAS pixel_7215/NB2 pixel_7215/AMP_IN pixel_7215/SF_IB
+ pixel_7215/PIX_OUT pixel_7215/CSA_VREF pixel
Xpixel_7226 pixel_7226/gring pixel_7226/VDD pixel_7226/GND pixel_7226/VREF pixel_7226/ROW_SEL
+ pixel_7226/NB1 pixel_7226/VBIAS pixel_7226/NB2 pixel_7226/AMP_IN pixel_7226/SF_IB
+ pixel_7226/PIX_OUT pixel_7226/CSA_VREF pixel
Xpixel_7237 pixel_7237/gring pixel_7237/VDD pixel_7237/GND pixel_7237/VREF pixel_7237/ROW_SEL
+ pixel_7237/NB1 pixel_7237/VBIAS pixel_7237/NB2 pixel_7237/AMP_IN pixel_7237/SF_IB
+ pixel_7237/PIX_OUT pixel_7237/CSA_VREF pixel
Xpixel_6503 pixel_6503/gring pixel_6503/VDD pixel_6503/GND pixel_6503/VREF pixel_6503/ROW_SEL
+ pixel_6503/NB1 pixel_6503/VBIAS pixel_6503/NB2 pixel_6503/AMP_IN pixel_6503/SF_IB
+ pixel_6503/PIX_OUT pixel_6503/CSA_VREF pixel
Xpixel_7248 pixel_7248/gring pixel_7248/VDD pixel_7248/GND pixel_7248/VREF pixel_7248/ROW_SEL
+ pixel_7248/NB1 pixel_7248/VBIAS pixel_7248/NB2 pixel_7248/AMP_IN pixel_7248/SF_IB
+ pixel_7248/PIX_OUT pixel_7248/CSA_VREF pixel
Xpixel_7259 pixel_7259/gring pixel_7259/VDD pixel_7259/GND pixel_7259/VREF pixel_7259/ROW_SEL
+ pixel_7259/NB1 pixel_7259/VBIAS pixel_7259/NB2 pixel_7259/AMP_IN pixel_7259/SF_IB
+ pixel_7259/PIX_OUT pixel_7259/CSA_VREF pixel
Xpixel_6514 pixel_6514/gring pixel_6514/VDD pixel_6514/GND pixel_6514/VREF pixel_6514/ROW_SEL
+ pixel_6514/NB1 pixel_6514/VBIAS pixel_6514/NB2 pixel_6514/AMP_IN pixel_6514/SF_IB
+ pixel_6514/PIX_OUT pixel_6514/CSA_VREF pixel
Xpixel_6525 pixel_6525/gring pixel_6525/VDD pixel_6525/GND pixel_6525/VREF pixel_6525/ROW_SEL
+ pixel_6525/NB1 pixel_6525/VBIAS pixel_6525/NB2 pixel_6525/AMP_IN pixel_6525/SF_IB
+ pixel_6525/PIX_OUT pixel_6525/CSA_VREF pixel
Xpixel_6536 pixel_6536/gring pixel_6536/VDD pixel_6536/GND pixel_6536/VREF pixel_6536/ROW_SEL
+ pixel_6536/NB1 pixel_6536/VBIAS pixel_6536/NB2 pixel_6536/AMP_IN pixel_6536/SF_IB
+ pixel_6536/PIX_OUT pixel_6536/CSA_VREF pixel
Xpixel_6547 pixel_6547/gring pixel_6547/VDD pixel_6547/GND pixel_6547/VREF pixel_6547/ROW_SEL
+ pixel_6547/NB1 pixel_6547/VBIAS pixel_6547/NB2 pixel_6547/AMP_IN pixel_6547/SF_IB
+ pixel_6547/PIX_OUT pixel_6547/CSA_VREF pixel
Xpixel_6558 pixel_6558/gring pixel_6558/VDD pixel_6558/GND pixel_6558/VREF pixel_6558/ROW_SEL
+ pixel_6558/NB1 pixel_6558/VBIAS pixel_6558/NB2 pixel_6558/AMP_IN pixel_6558/SF_IB
+ pixel_6558/PIX_OUT pixel_6558/CSA_VREF pixel
Xpixel_6569 pixel_6569/gring pixel_6569/VDD pixel_6569/GND pixel_6569/VREF pixel_6569/ROW_SEL
+ pixel_6569/NB1 pixel_6569/VBIAS pixel_6569/NB2 pixel_6569/AMP_IN pixel_6569/SF_IB
+ pixel_6569/PIX_OUT pixel_6569/CSA_VREF pixel
Xpixel_5802 pixel_5802/gring pixel_5802/VDD pixel_5802/GND pixel_5802/VREF pixel_5802/ROW_SEL
+ pixel_5802/NB1 pixel_5802/VBIAS pixel_5802/NB2 pixel_5802/AMP_IN pixel_5802/SF_IB
+ pixel_5802/PIX_OUT pixel_5802/CSA_VREF pixel
Xpixel_5813 pixel_5813/gring pixel_5813/VDD pixel_5813/GND pixel_5813/VREF pixel_5813/ROW_SEL
+ pixel_5813/NB1 pixel_5813/VBIAS pixel_5813/NB2 pixel_5813/AMP_IN pixel_5813/SF_IB
+ pixel_5813/PIX_OUT pixel_5813/CSA_VREF pixel
Xpixel_5824 pixel_5824/gring pixel_5824/VDD pixel_5824/GND pixel_5824/VREF pixel_5824/ROW_SEL
+ pixel_5824/NB1 pixel_5824/VBIAS pixel_5824/NB2 pixel_5824/AMP_IN pixel_5824/SF_IB
+ pixel_5824/PIX_OUT pixel_5824/CSA_VREF pixel
Xpixel_5835 pixel_5835/gring pixel_5835/VDD pixel_5835/GND pixel_5835/VREF pixel_5835/ROW_SEL
+ pixel_5835/NB1 pixel_5835/VBIAS pixel_5835/NB2 pixel_5835/AMP_IN pixel_5835/SF_IB
+ pixel_5835/PIX_OUT pixel_5835/CSA_VREF pixel
Xpixel_5846 pixel_5846/gring pixel_5846/VDD pixel_5846/GND pixel_5846/VREF pixel_5846/ROW_SEL
+ pixel_5846/NB1 pixel_5846/VBIAS pixel_5846/NB2 pixel_5846/AMP_IN pixel_5846/SF_IB
+ pixel_5846/PIX_OUT pixel_5846/CSA_VREF pixel
Xpixel_5857 pixel_5857/gring pixel_5857/VDD pixel_5857/GND pixel_5857/VREF pixel_5857/ROW_SEL
+ pixel_5857/NB1 pixel_5857/VBIAS pixel_5857/NB2 pixel_5857/AMP_IN pixel_5857/SF_IB
+ pixel_5857/PIX_OUT pixel_5857/CSA_VREF pixel
Xpixel_5868 pixel_5868/gring pixel_5868/VDD pixel_5868/GND pixel_5868/VREF pixel_5868/ROW_SEL
+ pixel_5868/NB1 pixel_5868/VBIAS pixel_5868/NB2 pixel_5868/AMP_IN pixel_5868/SF_IB
+ pixel_5868/PIX_OUT pixel_5868/CSA_VREF pixel
Xpixel_5879 pixel_5879/gring pixel_5879/VDD pixel_5879/GND pixel_5879/VREF pixel_5879/ROW_SEL
+ pixel_5879/NB1 pixel_5879/VBIAS pixel_5879/NB2 pixel_5879/AMP_IN pixel_5879/SF_IB
+ pixel_5879/PIX_OUT pixel_5879/CSA_VREF pixel
Xpixel_9140 pixel_9140/gring pixel_9140/VDD pixel_9140/GND pixel_9140/VREF pixel_9140/ROW_SEL
+ pixel_9140/NB1 pixel_9140/VBIAS pixel_9140/NB2 pixel_9140/AMP_IN pixel_9140/SF_IB
+ pixel_9140/PIX_OUT pixel_9140/CSA_VREF pixel
Xpixel_9173 pixel_9173/gring pixel_9173/VDD pixel_9173/GND pixel_9173/VREF pixel_9173/ROW_SEL
+ pixel_9173/NB1 pixel_9173/VBIAS pixel_9173/NB2 pixel_9173/AMP_IN pixel_9173/SF_IB
+ pixel_9173/PIX_OUT pixel_9173/CSA_VREF pixel
Xpixel_9162 pixel_9162/gring pixel_9162/VDD pixel_9162/GND pixel_9162/VREF pixel_9162/ROW_SEL
+ pixel_9162/NB1 pixel_9162/VBIAS pixel_9162/NB2 pixel_9162/AMP_IN pixel_9162/SF_IB
+ pixel_9162/PIX_OUT pixel_9162/CSA_VREF pixel
Xpixel_9151 pixel_9151/gring pixel_9151/VDD pixel_9151/GND pixel_9151/VREF pixel_9151/ROW_SEL
+ pixel_9151/NB1 pixel_9151/VBIAS pixel_9151/NB2 pixel_9151/AMP_IN pixel_9151/SF_IB
+ pixel_9151/PIX_OUT pixel_9151/CSA_VREF pixel
Xpixel_9195 pixel_9195/gring pixel_9195/VDD pixel_9195/GND pixel_9195/VREF pixel_9195/ROW_SEL
+ pixel_9195/NB1 pixel_9195/VBIAS pixel_9195/NB2 pixel_9195/AMP_IN pixel_9195/SF_IB
+ pixel_9195/PIX_OUT pixel_9195/CSA_VREF pixel
Xpixel_9184 pixel_9184/gring pixel_9184/VDD pixel_9184/GND pixel_9184/VREF pixel_9184/ROW_SEL
+ pixel_9184/NB1 pixel_9184/VBIAS pixel_9184/NB2 pixel_9184/AMP_IN pixel_9184/SF_IB
+ pixel_9184/PIX_OUT pixel_9184/CSA_VREF pixel
Xpixel_8450 pixel_8450/gring pixel_8450/VDD pixel_8450/GND pixel_8450/VREF pixel_8450/ROW_SEL
+ pixel_8450/NB1 pixel_8450/VBIAS pixel_8450/NB2 pixel_8450/AMP_IN pixel_8450/SF_IB
+ pixel_8450/PIX_OUT pixel_8450/CSA_VREF pixel
Xpixel_8461 pixel_8461/gring pixel_8461/VDD pixel_8461/GND pixel_8461/VREF pixel_8461/ROW_SEL
+ pixel_8461/NB1 pixel_8461/VBIAS pixel_8461/NB2 pixel_8461/AMP_IN pixel_8461/SF_IB
+ pixel_8461/PIX_OUT pixel_8461/CSA_VREF pixel
Xpixel_8472 pixel_8472/gring pixel_8472/VDD pixel_8472/GND pixel_8472/VREF pixel_8472/ROW_SEL
+ pixel_8472/NB1 pixel_8472/VBIAS pixel_8472/NB2 pixel_8472/AMP_IN pixel_8472/SF_IB
+ pixel_8472/PIX_OUT pixel_8472/CSA_VREF pixel
Xpixel_8483 pixel_8483/gring pixel_8483/VDD pixel_8483/GND pixel_8483/VREF pixel_8483/ROW_SEL
+ pixel_8483/NB1 pixel_8483/VBIAS pixel_8483/NB2 pixel_8483/AMP_IN pixel_8483/SF_IB
+ pixel_8483/PIX_OUT pixel_8483/CSA_VREF pixel
Xpixel_8494 pixel_8494/gring pixel_8494/VDD pixel_8494/GND pixel_8494/VREF pixel_8494/ROW_SEL
+ pixel_8494/NB1 pixel_8494/VBIAS pixel_8494/NB2 pixel_8494/AMP_IN pixel_8494/SF_IB
+ pixel_8494/PIX_OUT pixel_8494/CSA_VREF pixel
Xpixel_7760 pixel_7760/gring pixel_7760/VDD pixel_7760/GND pixel_7760/VREF pixel_7760/ROW_SEL
+ pixel_7760/NB1 pixel_7760/VBIAS pixel_7760/NB2 pixel_7760/AMP_IN pixel_7760/SF_IB
+ pixel_7760/PIX_OUT pixel_7760/CSA_VREF pixel
Xpixel_7771 pixel_7771/gring pixel_7771/VDD pixel_7771/GND pixel_7771/VREF pixel_7771/ROW_SEL
+ pixel_7771/NB1 pixel_7771/VBIAS pixel_7771/NB2 pixel_7771/AMP_IN pixel_7771/SF_IB
+ pixel_7771/PIX_OUT pixel_7771/CSA_VREF pixel
Xpixel_7782 pixel_7782/gring pixel_7782/VDD pixel_7782/GND pixel_7782/VREF pixel_7782/ROW_SEL
+ pixel_7782/NB1 pixel_7782/VBIAS pixel_7782/NB2 pixel_7782/AMP_IN pixel_7782/SF_IB
+ pixel_7782/PIX_OUT pixel_7782/CSA_VREF pixel
Xpixel_7793 pixel_7793/gring pixel_7793/VDD pixel_7793/GND pixel_7793/VREF pixel_7793/ROW_SEL
+ pixel_7793/NB1 pixel_7793/VBIAS pixel_7793/NB2 pixel_7793/AMP_IN pixel_7793/SF_IB
+ pixel_7793/PIX_OUT pixel_7793/CSA_VREF pixel
Xpixel_5109 pixel_5109/gring pixel_5109/VDD pixel_5109/GND pixel_5109/VREF pixel_5109/ROW_SEL
+ pixel_5109/NB1 pixel_5109/VBIAS pixel_5109/NB2 pixel_5109/AMP_IN pixel_5109/SF_IB
+ pixel_5109/PIX_OUT pixel_5109/CSA_VREF pixel
Xpixel_414 pixel_414/gring pixel_414/VDD pixel_414/GND pixel_414/VREF pixel_414/ROW_SEL
+ pixel_414/NB1 pixel_414/VBIAS pixel_414/NB2 pixel_414/AMP_IN pixel_414/SF_IB pixel_414/PIX_OUT
+ pixel_414/CSA_VREF pixel
Xpixel_403 pixel_403/gring pixel_403/VDD pixel_403/GND pixel_403/VREF pixel_403/ROW_SEL
+ pixel_403/NB1 pixel_403/VBIAS pixel_403/NB2 pixel_403/AMP_IN pixel_403/SF_IB pixel_403/PIX_OUT
+ pixel_403/CSA_VREF pixel
Xpixel_4408 pixel_4408/gring pixel_4408/VDD pixel_4408/GND pixel_4408/VREF pixel_4408/ROW_SEL
+ pixel_4408/NB1 pixel_4408/VBIAS pixel_4408/NB2 pixel_4408/AMP_IN pixel_4408/SF_IB
+ pixel_4408/PIX_OUT pixel_4408/CSA_VREF pixel
Xpixel_447 pixel_447/gring pixel_447/VDD pixel_447/GND pixel_447/VREF pixel_447/ROW_SEL
+ pixel_447/NB1 pixel_447/VBIAS pixel_447/NB2 pixel_447/AMP_IN pixel_447/SF_IB pixel_447/PIX_OUT
+ pixel_447/CSA_VREF pixel
Xpixel_436 pixel_436/gring pixel_436/VDD pixel_436/GND pixel_436/VREF pixel_436/ROW_SEL
+ pixel_436/NB1 pixel_436/VBIAS pixel_436/NB2 pixel_436/AMP_IN pixel_436/SF_IB pixel_436/PIX_OUT
+ pixel_436/CSA_VREF pixel
Xpixel_425 pixel_425/gring pixel_425/VDD pixel_425/GND pixel_425/VREF pixel_425/ROW_SEL
+ pixel_425/NB1 pixel_425/VBIAS pixel_425/NB2 pixel_425/AMP_IN pixel_425/SF_IB pixel_425/PIX_OUT
+ pixel_425/CSA_VREF pixel
Xpixel_3707 pixel_3707/gring pixel_3707/VDD pixel_3707/GND pixel_3707/VREF pixel_3707/ROW_SEL
+ pixel_3707/NB1 pixel_3707/VBIAS pixel_3707/NB2 pixel_3707/AMP_IN pixel_3707/SF_IB
+ pixel_3707/PIX_OUT pixel_3707/CSA_VREF pixel
Xpixel_4419 pixel_4419/gring pixel_4419/VDD pixel_4419/GND pixel_4419/VREF pixel_4419/ROW_SEL
+ pixel_4419/NB1 pixel_4419/VBIAS pixel_4419/NB2 pixel_4419/AMP_IN pixel_4419/SF_IB
+ pixel_4419/PIX_OUT pixel_4419/CSA_VREF pixel
Xpixel_469 pixel_469/gring pixel_469/VDD pixel_469/GND pixel_469/VREF pixel_469/ROW_SEL
+ pixel_469/NB1 pixel_469/VBIAS pixel_469/NB2 pixel_469/AMP_IN pixel_469/SF_IB pixel_469/PIX_OUT
+ pixel_469/CSA_VREF pixel
Xpixel_458 pixel_458/gring pixel_458/VDD pixel_458/GND pixel_458/VREF pixel_458/ROW_SEL
+ pixel_458/NB1 pixel_458/VBIAS pixel_458/NB2 pixel_458/AMP_IN pixel_458/SF_IB pixel_458/PIX_OUT
+ pixel_458/CSA_VREF pixel
Xpixel_3729 pixel_3729/gring pixel_3729/VDD pixel_3729/GND pixel_3729/VREF pixel_3729/ROW_SEL
+ pixel_3729/NB1 pixel_3729/VBIAS pixel_3729/NB2 pixel_3729/AMP_IN pixel_3729/SF_IB
+ pixel_3729/PIX_OUT pixel_3729/CSA_VREF pixel
Xpixel_3718 pixel_3718/gring pixel_3718/VDD pixel_3718/GND pixel_3718/VREF pixel_3718/ROW_SEL
+ pixel_3718/NB1 pixel_3718/VBIAS pixel_3718/NB2 pixel_3718/AMP_IN pixel_3718/SF_IB
+ pixel_3718/PIX_OUT pixel_3718/CSA_VREF pixel
Xpixel_7001 pixel_7001/gring pixel_7001/VDD pixel_7001/GND pixel_7001/VREF pixel_7001/ROW_SEL
+ pixel_7001/NB1 pixel_7001/VBIAS pixel_7001/NB2 pixel_7001/AMP_IN pixel_7001/SF_IB
+ pixel_7001/PIX_OUT pixel_7001/CSA_VREF pixel
Xpixel_7012 pixel_7012/gring pixel_7012/VDD pixel_7012/GND pixel_7012/VREF pixel_7012/ROW_SEL
+ pixel_7012/NB1 pixel_7012/VBIAS pixel_7012/NB2 pixel_7012/AMP_IN pixel_7012/SF_IB
+ pixel_7012/PIX_OUT pixel_7012/CSA_VREF pixel
Xpixel_7023 pixel_7023/gring pixel_7023/VDD pixel_7023/GND pixel_7023/VREF pixel_7023/ROW_SEL
+ pixel_7023/NB1 pixel_7023/VBIAS pixel_7023/NB2 pixel_7023/AMP_IN pixel_7023/SF_IB
+ pixel_7023/PIX_OUT pixel_7023/CSA_VREF pixel
Xpixel_7034 pixel_7034/gring pixel_7034/VDD pixel_7034/GND pixel_7034/VREF pixel_7034/ROW_SEL
+ pixel_7034/NB1 pixel_7034/VBIAS pixel_7034/NB2 pixel_7034/AMP_IN pixel_7034/SF_IB
+ pixel_7034/PIX_OUT pixel_7034/CSA_VREF pixel
Xpixel_7045 pixel_7045/gring pixel_7045/VDD pixel_7045/GND pixel_7045/VREF pixel_7045/ROW_SEL
+ pixel_7045/NB1 pixel_7045/VBIAS pixel_7045/NB2 pixel_7045/AMP_IN pixel_7045/SF_IB
+ pixel_7045/PIX_OUT pixel_7045/CSA_VREF pixel
Xpixel_7056 pixel_7056/gring pixel_7056/VDD pixel_7056/GND pixel_7056/VREF pixel_7056/ROW_SEL
+ pixel_7056/NB1 pixel_7056/VBIAS pixel_7056/NB2 pixel_7056/AMP_IN pixel_7056/SF_IB
+ pixel_7056/PIX_OUT pixel_7056/CSA_VREF pixel
Xpixel_6300 pixel_6300/gring pixel_6300/VDD pixel_6300/GND pixel_6300/VREF pixel_6300/ROW_SEL
+ pixel_6300/NB1 pixel_6300/VBIAS pixel_6300/NB2 pixel_6300/AMP_IN pixel_6300/SF_IB
+ pixel_6300/PIX_OUT pixel_6300/CSA_VREF pixel
Xpixel_6311 pixel_6311/gring pixel_6311/VDD pixel_6311/GND pixel_6311/VREF pixel_6311/ROW_SEL
+ pixel_6311/NB1 pixel_6311/VBIAS pixel_6311/NB2 pixel_6311/AMP_IN pixel_6311/SF_IB
+ pixel_6311/PIX_OUT pixel_6311/CSA_VREF pixel
Xpixel_7067 pixel_7067/gring pixel_7067/VDD pixel_7067/GND pixel_7067/VREF pixel_7067/ROW_SEL
+ pixel_7067/NB1 pixel_7067/VBIAS pixel_7067/NB2 pixel_7067/AMP_IN pixel_7067/SF_IB
+ pixel_7067/PIX_OUT pixel_7067/CSA_VREF pixel
Xpixel_7078 pixel_7078/gring pixel_7078/VDD pixel_7078/GND pixel_7078/VREF pixel_7078/ROW_SEL
+ pixel_7078/NB1 pixel_7078/VBIAS pixel_7078/NB2 pixel_7078/AMP_IN pixel_7078/SF_IB
+ pixel_7078/PIX_OUT pixel_7078/CSA_VREF pixel
Xpixel_7089 pixel_7089/gring pixel_7089/VDD pixel_7089/GND pixel_7089/VREF pixel_7089/ROW_SEL
+ pixel_7089/NB1 pixel_7089/VBIAS pixel_7089/NB2 pixel_7089/AMP_IN pixel_7089/SF_IB
+ pixel_7089/PIX_OUT pixel_7089/CSA_VREF pixel
Xpixel_6322 pixel_6322/gring pixel_6322/VDD pixel_6322/GND pixel_6322/VREF pixel_6322/ROW_SEL
+ pixel_6322/NB1 pixel_6322/VBIAS pixel_6322/NB2 pixel_6322/AMP_IN pixel_6322/SF_IB
+ pixel_6322/PIX_OUT pixel_6322/CSA_VREF pixel
Xpixel_6333 pixel_6333/gring pixel_6333/VDD pixel_6333/GND pixel_6333/VREF pixel_6333/ROW_SEL
+ pixel_6333/NB1 pixel_6333/VBIAS pixel_6333/NB2 pixel_6333/AMP_IN pixel_6333/SF_IB
+ pixel_6333/PIX_OUT pixel_6333/CSA_VREF pixel
Xpixel_6344 pixel_6344/gring pixel_6344/VDD pixel_6344/GND pixel_6344/VREF pixel_6344/ROW_SEL
+ pixel_6344/NB1 pixel_6344/VBIAS pixel_6344/NB2 pixel_6344/AMP_IN pixel_6344/SF_IB
+ pixel_6344/PIX_OUT pixel_6344/CSA_VREF pixel
Xpixel_6355 pixel_6355/gring pixel_6355/VDD pixel_6355/GND pixel_6355/VREF pixel_6355/ROW_SEL
+ pixel_6355/NB1 pixel_6355/VBIAS pixel_6355/NB2 pixel_6355/AMP_IN pixel_6355/SF_IB
+ pixel_6355/PIX_OUT pixel_6355/CSA_VREF pixel
Xpixel_6366 pixel_6366/gring pixel_6366/VDD pixel_6366/GND pixel_6366/VREF pixel_6366/ROW_SEL
+ pixel_6366/NB1 pixel_6366/VBIAS pixel_6366/NB2 pixel_6366/AMP_IN pixel_6366/SF_IB
+ pixel_6366/PIX_OUT pixel_6366/CSA_VREF pixel
Xpixel_6377 pixel_6377/gring pixel_6377/VDD pixel_6377/GND pixel_6377/VREF pixel_6377/ROW_SEL
+ pixel_6377/NB1 pixel_6377/VBIAS pixel_6377/NB2 pixel_6377/AMP_IN pixel_6377/SF_IB
+ pixel_6377/PIX_OUT pixel_6377/CSA_VREF pixel
Xpixel_5610 pixel_5610/gring pixel_5610/VDD pixel_5610/GND pixel_5610/VREF pixel_5610/ROW_SEL
+ pixel_5610/NB1 pixel_5610/VBIAS pixel_5610/NB2 pixel_5610/AMP_IN pixel_5610/SF_IB
+ pixel_5610/PIX_OUT pixel_5610/CSA_VREF pixel
Xpixel_5621 pixel_5621/gring pixel_5621/VDD pixel_5621/GND pixel_5621/VREF pixel_5621/ROW_SEL
+ pixel_5621/NB1 pixel_5621/VBIAS pixel_5621/NB2 pixel_5621/AMP_IN pixel_5621/SF_IB
+ pixel_5621/PIX_OUT pixel_5621/CSA_VREF pixel
Xpixel_5632 pixel_5632/gring pixel_5632/VDD pixel_5632/GND pixel_5632/VREF pixel_5632/ROW_SEL
+ pixel_5632/NB1 pixel_5632/VBIAS pixel_5632/NB2 pixel_5632/AMP_IN pixel_5632/SF_IB
+ pixel_5632/PIX_OUT pixel_5632/CSA_VREF pixel
Xpixel_6388 pixel_6388/gring pixel_6388/VDD pixel_6388/GND pixel_6388/VREF pixel_6388/ROW_SEL
+ pixel_6388/NB1 pixel_6388/VBIAS pixel_6388/NB2 pixel_6388/AMP_IN pixel_6388/SF_IB
+ pixel_6388/PIX_OUT pixel_6388/CSA_VREF pixel
Xpixel_6399 pixel_6399/gring pixel_6399/VDD pixel_6399/GND pixel_6399/VREF pixel_6399/ROW_SEL
+ pixel_6399/NB1 pixel_6399/VBIAS pixel_6399/NB2 pixel_6399/AMP_IN pixel_6399/SF_IB
+ pixel_6399/PIX_OUT pixel_6399/CSA_VREF pixel
Xpixel_5643 pixel_5643/gring pixel_5643/VDD pixel_5643/GND pixel_5643/VREF pixel_5643/ROW_SEL
+ pixel_5643/NB1 pixel_5643/VBIAS pixel_5643/NB2 pixel_5643/AMP_IN pixel_5643/SF_IB
+ pixel_5643/PIX_OUT pixel_5643/CSA_VREF pixel
Xpixel_5654 pixel_5654/gring pixel_5654/VDD pixel_5654/GND pixel_5654/VREF pixel_5654/ROW_SEL
+ pixel_5654/NB1 pixel_5654/VBIAS pixel_5654/NB2 pixel_5654/AMP_IN pixel_5654/SF_IB
+ pixel_5654/PIX_OUT pixel_5654/CSA_VREF pixel
Xpixel_5665 pixel_5665/gring pixel_5665/VDD pixel_5665/GND pixel_5665/VREF pixel_5665/ROW_SEL
+ pixel_5665/NB1 pixel_5665/VBIAS pixel_5665/NB2 pixel_5665/AMP_IN pixel_5665/SF_IB
+ pixel_5665/PIX_OUT pixel_5665/CSA_VREF pixel
Xpixel_5676 pixel_5676/gring pixel_5676/VDD pixel_5676/GND pixel_5676/VREF pixel_5676/ROW_SEL
+ pixel_5676/NB1 pixel_5676/VBIAS pixel_5676/NB2 pixel_5676/AMP_IN pixel_5676/SF_IB
+ pixel_5676/PIX_OUT pixel_5676/CSA_VREF pixel
Xpixel_4920 pixel_4920/gring pixel_4920/VDD pixel_4920/GND pixel_4920/VREF pixel_4920/ROW_SEL
+ pixel_4920/NB1 pixel_4920/VBIAS pixel_4920/NB2 pixel_4920/AMP_IN pixel_4920/SF_IB
+ pixel_4920/PIX_OUT pixel_4920/CSA_VREF pixel
Xpixel_4931 pixel_4931/gring pixel_4931/VDD pixel_4931/GND pixel_4931/VREF pixel_4931/ROW_SEL
+ pixel_4931/NB1 pixel_4931/VBIAS pixel_4931/NB2 pixel_4931/AMP_IN pixel_4931/SF_IB
+ pixel_4931/PIX_OUT pixel_4931/CSA_VREF pixel
Xpixel_5687 pixel_5687/gring pixel_5687/VDD pixel_5687/GND pixel_5687/VREF pixel_5687/ROW_SEL
+ pixel_5687/NB1 pixel_5687/VBIAS pixel_5687/NB2 pixel_5687/AMP_IN pixel_5687/SF_IB
+ pixel_5687/PIX_OUT pixel_5687/CSA_VREF pixel
Xpixel_5698 pixel_5698/gring pixel_5698/VDD pixel_5698/GND pixel_5698/VREF pixel_5698/ROW_SEL
+ pixel_5698/NB1 pixel_5698/VBIAS pixel_5698/NB2 pixel_5698/AMP_IN pixel_5698/SF_IB
+ pixel_5698/PIX_OUT pixel_5698/CSA_VREF pixel
Xpixel_4942 pixel_4942/gring pixel_4942/VDD pixel_4942/GND pixel_4942/VREF pixel_4942/ROW_SEL
+ pixel_4942/NB1 pixel_4942/VBIAS pixel_4942/NB2 pixel_4942/AMP_IN pixel_4942/SF_IB
+ pixel_4942/PIX_OUT pixel_4942/CSA_VREF pixel
Xpixel_4953 pixel_4953/gring pixel_4953/VDD pixel_4953/GND pixel_4953/VREF pixel_4953/ROW_SEL
+ pixel_4953/NB1 pixel_4953/VBIAS pixel_4953/NB2 pixel_4953/AMP_IN pixel_4953/SF_IB
+ pixel_4953/PIX_OUT pixel_4953/CSA_VREF pixel
Xpixel_4964 pixel_4964/gring pixel_4964/VDD pixel_4964/GND pixel_4964/VREF pixel_4964/ROW_SEL
+ pixel_4964/NB1 pixel_4964/VBIAS pixel_4964/NB2 pixel_4964/AMP_IN pixel_4964/SF_IB
+ pixel_4964/PIX_OUT pixel_4964/CSA_VREF pixel
Xpixel_992 pixel_992/gring pixel_992/VDD pixel_992/GND pixel_992/VREF pixel_992/ROW_SEL
+ pixel_992/NB1 pixel_992/VBIAS pixel_992/NB2 pixel_992/AMP_IN pixel_992/SF_IB pixel_992/PIX_OUT
+ pixel_992/CSA_VREF pixel
Xpixel_981 pixel_981/gring pixel_981/VDD pixel_981/GND pixel_981/VREF pixel_981/ROW_SEL
+ pixel_981/NB1 pixel_981/VBIAS pixel_981/NB2 pixel_981/AMP_IN pixel_981/SF_IB pixel_981/PIX_OUT
+ pixel_981/CSA_VREF pixel
Xpixel_970 pixel_970/gring pixel_970/VDD pixel_970/GND pixel_970/VREF pixel_970/ROW_SEL
+ pixel_970/NB1 pixel_970/VBIAS pixel_970/NB2 pixel_970/AMP_IN pixel_970/SF_IB pixel_970/PIX_OUT
+ pixel_970/CSA_VREF pixel
Xpixel_4975 pixel_4975/gring pixel_4975/VDD pixel_4975/GND pixel_4975/VREF pixel_4975/ROW_SEL
+ pixel_4975/NB1 pixel_4975/VBIAS pixel_4975/NB2 pixel_4975/AMP_IN pixel_4975/SF_IB
+ pixel_4975/PIX_OUT pixel_4975/CSA_VREF pixel
Xpixel_4986 pixel_4986/gring pixel_4986/VDD pixel_4986/GND pixel_4986/VREF pixel_4986/ROW_SEL
+ pixel_4986/NB1 pixel_4986/VBIAS pixel_4986/NB2 pixel_4986/AMP_IN pixel_4986/SF_IB
+ pixel_4986/PIX_OUT pixel_4986/CSA_VREF pixel
Xpixel_4997 pixel_4997/gring pixel_4997/VDD pixel_4997/GND pixel_4997/VREF pixel_4997/ROW_SEL
+ pixel_4997/NB1 pixel_4997/VBIAS pixel_4997/NB2 pixel_4997/AMP_IN pixel_4997/SF_IB
+ pixel_4997/PIX_OUT pixel_4997/CSA_VREF pixel
Xpixel_8280 pixel_8280/gring pixel_8280/VDD pixel_8280/GND pixel_8280/VREF pixel_8280/ROW_SEL
+ pixel_8280/NB1 pixel_8280/VBIAS pixel_8280/NB2 pixel_8280/AMP_IN pixel_8280/SF_IB
+ pixel_8280/PIX_OUT pixel_8280/CSA_VREF pixel
Xpixel_8291 pixel_8291/gring pixel_8291/VDD pixel_8291/GND pixel_8291/VREF pixel_8291/ROW_SEL
+ pixel_8291/NB1 pixel_8291/VBIAS pixel_8291/NB2 pixel_8291/AMP_IN pixel_8291/SF_IB
+ pixel_8291/PIX_OUT pixel_8291/CSA_VREF pixel
Xpixel_7590 pixel_7590/gring pixel_7590/VDD pixel_7590/GND pixel_7590/VREF pixel_7590/ROW_SEL
+ pixel_7590/NB1 pixel_7590/VBIAS pixel_7590/NB2 pixel_7590/AMP_IN pixel_7590/SF_IB
+ pixel_7590/PIX_OUT pixel_7590/CSA_VREF pixel
Xpixel_9909 pixel_9909/gring pixel_9909/VDD pixel_9909/GND pixel_9909/VREF pixel_9909/ROW_SEL
+ pixel_9909/NB1 pixel_9909/VBIAS pixel_9909/NB2 pixel_9909/AMP_IN pixel_9909/SF_IB
+ pixel_9909/PIX_OUT pixel_9909/CSA_VREF pixel
Xpixel_222 pixel_222/gring pixel_222/VDD pixel_222/GND pixel_222/VREF pixel_222/ROW_SEL
+ pixel_222/NB1 pixel_222/VBIAS pixel_222/NB2 pixel_222/AMP_IN pixel_222/SF_IB pixel_222/PIX_OUT
+ pixel_222/CSA_VREF pixel
Xpixel_211 pixel_211/gring pixel_211/VDD pixel_211/GND pixel_211/VREF pixel_211/ROW_SEL
+ pixel_211/NB1 pixel_211/VBIAS pixel_211/NB2 pixel_211/AMP_IN pixel_211/SF_IB pixel_211/PIX_OUT
+ pixel_211/CSA_VREF pixel
Xpixel_200 pixel_200/gring pixel_200/VDD pixel_200/GND pixel_200/VREF pixel_200/ROW_SEL
+ pixel_200/NB1 pixel_200/VBIAS pixel_200/NB2 pixel_200/AMP_IN pixel_200/SF_IB pixel_200/PIX_OUT
+ pixel_200/CSA_VREF pixel
Xpixel_4205 pixel_4205/gring pixel_4205/VDD pixel_4205/GND pixel_4205/VREF pixel_4205/ROW_SEL
+ pixel_4205/NB1 pixel_4205/VBIAS pixel_4205/NB2 pixel_4205/AMP_IN pixel_4205/SF_IB
+ pixel_4205/PIX_OUT pixel_4205/CSA_VREF pixel
Xpixel_4216 pixel_4216/gring pixel_4216/VDD pixel_4216/GND pixel_4216/VREF pixel_4216/ROW_SEL
+ pixel_4216/NB1 pixel_4216/VBIAS pixel_4216/NB2 pixel_4216/AMP_IN pixel_4216/SF_IB
+ pixel_4216/PIX_OUT pixel_4216/CSA_VREF pixel
Xpixel_4227 pixel_4227/gring pixel_4227/VDD pixel_4227/GND pixel_4227/VREF pixel_4227/ROW_SEL
+ pixel_4227/NB1 pixel_4227/VBIAS pixel_4227/NB2 pixel_4227/AMP_IN pixel_4227/SF_IB
+ pixel_4227/PIX_OUT pixel_4227/CSA_VREF pixel
Xpixel_255 pixel_255/gring pixel_255/VDD pixel_255/GND pixel_255/VREF pixel_255/ROW_SEL
+ pixel_255/NB1 pixel_255/VBIAS pixel_255/NB2 pixel_255/AMP_IN pixel_255/SF_IB pixel_255/PIX_OUT
+ pixel_255/CSA_VREF pixel
Xpixel_244 pixel_244/gring pixel_244/VDD pixel_244/GND pixel_244/VREF pixel_244/ROW_SEL
+ pixel_244/NB1 pixel_244/VBIAS pixel_244/NB2 pixel_244/AMP_IN pixel_244/SF_IB pixel_244/PIX_OUT
+ pixel_244/CSA_VREF pixel
Xpixel_233 pixel_233/gring pixel_233/VDD pixel_233/GND pixel_233/VREF pixel_233/ROW_SEL
+ pixel_233/NB1 pixel_233/VBIAS pixel_233/NB2 pixel_233/AMP_IN pixel_233/SF_IB pixel_233/PIX_OUT
+ pixel_233/CSA_VREF pixel
Xpixel_3515 pixel_3515/gring pixel_3515/VDD pixel_3515/GND pixel_3515/VREF pixel_3515/ROW_SEL
+ pixel_3515/NB1 pixel_3515/VBIAS pixel_3515/NB2 pixel_3515/AMP_IN pixel_3515/SF_IB
+ pixel_3515/PIX_OUT pixel_3515/CSA_VREF pixel
Xpixel_3504 pixel_3504/gring pixel_3504/VDD pixel_3504/GND pixel_3504/VREF pixel_3504/ROW_SEL
+ pixel_3504/NB1 pixel_3504/VBIAS pixel_3504/NB2 pixel_3504/AMP_IN pixel_3504/SF_IB
+ pixel_3504/PIX_OUT pixel_3504/CSA_VREF pixel
Xpixel_4238 pixel_4238/gring pixel_4238/VDD pixel_4238/GND pixel_4238/VREF pixel_4238/ROW_SEL
+ pixel_4238/NB1 pixel_4238/VBIAS pixel_4238/NB2 pixel_4238/AMP_IN pixel_4238/SF_IB
+ pixel_4238/PIX_OUT pixel_4238/CSA_VREF pixel
Xpixel_4249 pixel_4249/gring pixel_4249/VDD pixel_4249/GND pixel_4249/VREF pixel_4249/ROW_SEL
+ pixel_4249/NB1 pixel_4249/VBIAS pixel_4249/NB2 pixel_4249/AMP_IN pixel_4249/SF_IB
+ pixel_4249/PIX_OUT pixel_4249/CSA_VREF pixel
Xpixel_288 pixel_288/gring pixel_288/VDD pixel_288/GND pixel_288/VREF pixel_288/ROW_SEL
+ pixel_288/NB1 pixel_288/VBIAS pixel_288/NB2 pixel_288/AMP_IN pixel_288/SF_IB pixel_288/PIX_OUT
+ pixel_288/CSA_VREF pixel
Xpixel_277 pixel_277/gring pixel_277/VDD pixel_277/GND pixel_277/VREF pixel_277/ROW_SEL
+ pixel_277/NB1 pixel_277/VBIAS pixel_277/NB2 pixel_277/AMP_IN pixel_277/SF_IB pixel_277/PIX_OUT
+ pixel_277/CSA_VREF pixel
Xpixel_266 pixel_266/gring pixel_266/VDD pixel_266/GND pixel_266/VREF pixel_266/ROW_SEL
+ pixel_266/NB1 pixel_266/VBIAS pixel_266/NB2 pixel_266/AMP_IN pixel_266/SF_IB pixel_266/PIX_OUT
+ pixel_266/CSA_VREF pixel
Xpixel_2803 pixel_2803/gring pixel_2803/VDD pixel_2803/GND pixel_2803/VREF pixel_2803/ROW_SEL
+ pixel_2803/NB1 pixel_2803/VBIAS pixel_2803/NB2 pixel_2803/AMP_IN pixel_2803/SF_IB
+ pixel_2803/PIX_OUT pixel_2803/CSA_VREF pixel
Xpixel_3548 pixel_3548/gring pixel_3548/VDD pixel_3548/GND pixel_3548/VREF pixel_3548/ROW_SEL
+ pixel_3548/NB1 pixel_3548/VBIAS pixel_3548/NB2 pixel_3548/AMP_IN pixel_3548/SF_IB
+ pixel_3548/PIX_OUT pixel_3548/CSA_VREF pixel
Xpixel_3537 pixel_3537/gring pixel_3537/VDD pixel_3537/GND pixel_3537/VREF pixel_3537/ROW_SEL
+ pixel_3537/NB1 pixel_3537/VBIAS pixel_3537/NB2 pixel_3537/AMP_IN pixel_3537/SF_IB
+ pixel_3537/PIX_OUT pixel_3537/CSA_VREF pixel
Xpixel_3526 pixel_3526/gring pixel_3526/VDD pixel_3526/GND pixel_3526/VREF pixel_3526/ROW_SEL
+ pixel_3526/NB1 pixel_3526/VBIAS pixel_3526/NB2 pixel_3526/AMP_IN pixel_3526/SF_IB
+ pixel_3526/PIX_OUT pixel_3526/CSA_VREF pixel
Xpixel_299 pixel_299/gring pixel_299/VDD pixel_299/GND pixel_299/VREF pixel_299/ROW_SEL
+ pixel_299/NB1 pixel_299/VBIAS pixel_299/NB2 pixel_299/AMP_IN pixel_299/SF_IB pixel_299/PIX_OUT
+ pixel_299/CSA_VREF pixel
Xpixel_2847 pixel_2847/gring pixel_2847/VDD pixel_2847/GND pixel_2847/VREF pixel_2847/ROW_SEL
+ pixel_2847/NB1 pixel_2847/VBIAS pixel_2847/NB2 pixel_2847/AMP_IN pixel_2847/SF_IB
+ pixel_2847/PIX_OUT pixel_2847/CSA_VREF pixel
Xpixel_2836 pixel_2836/gring pixel_2836/VDD pixel_2836/GND pixel_2836/VREF pixel_2836/ROW_SEL
+ pixel_2836/NB1 pixel_2836/VBIAS pixel_2836/NB2 pixel_2836/AMP_IN pixel_2836/SF_IB
+ pixel_2836/PIX_OUT pixel_2836/CSA_VREF pixel
Xpixel_2825 pixel_2825/gring pixel_2825/VDD pixel_2825/GND pixel_2825/VREF pixel_2825/ROW_SEL
+ pixel_2825/NB1 pixel_2825/VBIAS pixel_2825/NB2 pixel_2825/AMP_IN pixel_2825/SF_IB
+ pixel_2825/PIX_OUT pixel_2825/CSA_VREF pixel
Xpixel_2814 pixel_2814/gring pixel_2814/VDD pixel_2814/GND pixel_2814/VREF pixel_2814/ROW_SEL
+ pixel_2814/NB1 pixel_2814/VBIAS pixel_2814/NB2 pixel_2814/AMP_IN pixel_2814/SF_IB
+ pixel_2814/PIX_OUT pixel_2814/CSA_VREF pixel
Xpixel_3559 pixel_3559/gring pixel_3559/VDD pixel_3559/GND pixel_3559/VREF pixel_3559/ROW_SEL
+ pixel_3559/NB1 pixel_3559/VBIAS pixel_3559/NB2 pixel_3559/AMP_IN pixel_3559/SF_IB
+ pixel_3559/PIX_OUT pixel_3559/CSA_VREF pixel
Xpixel_2869 pixel_2869/gring pixel_2869/VDD pixel_2869/GND pixel_2869/VREF pixel_2869/ROW_SEL
+ pixel_2869/NB1 pixel_2869/VBIAS pixel_2869/NB2 pixel_2869/AMP_IN pixel_2869/SF_IB
+ pixel_2869/PIX_OUT pixel_2869/CSA_VREF pixel
Xpixel_2858 pixel_2858/gring pixel_2858/VDD pixel_2858/GND pixel_2858/VREF pixel_2858/ROW_SEL
+ pixel_2858/NB1 pixel_2858/VBIAS pixel_2858/NB2 pixel_2858/AMP_IN pixel_2858/SF_IB
+ pixel_2858/PIX_OUT pixel_2858/CSA_VREF pixel
Xpixel_6130 pixel_6130/gring pixel_6130/VDD pixel_6130/GND pixel_6130/VREF pixel_6130/ROW_SEL
+ pixel_6130/NB1 pixel_6130/VBIAS pixel_6130/NB2 pixel_6130/AMP_IN pixel_6130/SF_IB
+ pixel_6130/PIX_OUT pixel_6130/CSA_VREF pixel
Xpixel_6141 pixel_6141/gring pixel_6141/VDD pixel_6141/GND pixel_6141/VREF pixel_6141/ROW_SEL
+ pixel_6141/NB1 pixel_6141/VBIAS pixel_6141/NB2 pixel_6141/AMP_IN pixel_6141/SF_IB
+ pixel_6141/PIX_OUT pixel_6141/CSA_VREF pixel
Xpixel_6152 pixel_6152/gring pixel_6152/VDD pixel_6152/GND pixel_6152/VREF pixel_6152/ROW_SEL
+ pixel_6152/NB1 pixel_6152/VBIAS pixel_6152/NB2 pixel_6152/AMP_IN pixel_6152/SF_IB
+ pixel_6152/PIX_OUT pixel_6152/CSA_VREF pixel
Xpixel_6163 pixel_6163/gring pixel_6163/VDD pixel_6163/GND pixel_6163/VREF pixel_6163/ROW_SEL
+ pixel_6163/NB1 pixel_6163/VBIAS pixel_6163/NB2 pixel_6163/AMP_IN pixel_6163/SF_IB
+ pixel_6163/PIX_OUT pixel_6163/CSA_VREF pixel
Xpixel_6174 pixel_6174/gring pixel_6174/VDD pixel_6174/GND pixel_6174/VREF pixel_6174/ROW_SEL
+ pixel_6174/NB1 pixel_6174/VBIAS pixel_6174/NB2 pixel_6174/AMP_IN pixel_6174/SF_IB
+ pixel_6174/PIX_OUT pixel_6174/CSA_VREF pixel
Xpixel_6185 pixel_6185/gring pixel_6185/VDD pixel_6185/GND pixel_6185/VREF pixel_6185/ROW_SEL
+ pixel_6185/NB1 pixel_6185/VBIAS pixel_6185/NB2 pixel_6185/AMP_IN pixel_6185/SF_IB
+ pixel_6185/PIX_OUT pixel_6185/CSA_VREF pixel
Xpixel_6196 pixel_6196/gring pixel_6196/VDD pixel_6196/GND pixel_6196/VREF pixel_6196/ROW_SEL
+ pixel_6196/NB1 pixel_6196/VBIAS pixel_6196/NB2 pixel_6196/AMP_IN pixel_6196/SF_IB
+ pixel_6196/PIX_OUT pixel_6196/CSA_VREF pixel
Xpixel_5440 pixel_5440/gring pixel_5440/VDD pixel_5440/GND pixel_5440/VREF pixel_5440/ROW_SEL
+ pixel_5440/NB1 pixel_5440/VBIAS pixel_5440/NB2 pixel_5440/AMP_IN pixel_5440/SF_IB
+ pixel_5440/PIX_OUT pixel_5440/CSA_VREF pixel
Xpixel_5451 pixel_5451/gring pixel_5451/VDD pixel_5451/GND pixel_5451/VREF pixel_5451/ROW_SEL
+ pixel_5451/NB1 pixel_5451/VBIAS pixel_5451/NB2 pixel_5451/AMP_IN pixel_5451/SF_IB
+ pixel_5451/PIX_OUT pixel_5451/CSA_VREF pixel
Xpixel_5462 pixel_5462/gring pixel_5462/VDD pixel_5462/GND pixel_5462/VREF pixel_5462/ROW_SEL
+ pixel_5462/NB1 pixel_5462/VBIAS pixel_5462/NB2 pixel_5462/AMP_IN pixel_5462/SF_IB
+ pixel_5462/PIX_OUT pixel_5462/CSA_VREF pixel
Xpixel_5473 pixel_5473/gring pixel_5473/VDD pixel_5473/GND pixel_5473/VREF pixel_5473/ROW_SEL
+ pixel_5473/NB1 pixel_5473/VBIAS pixel_5473/NB2 pixel_5473/AMP_IN pixel_5473/SF_IB
+ pixel_5473/PIX_OUT pixel_5473/CSA_VREF pixel
Xpixel_5484 pixel_5484/gring pixel_5484/VDD pixel_5484/GND pixel_5484/VREF pixel_5484/ROW_SEL
+ pixel_5484/NB1 pixel_5484/VBIAS pixel_5484/NB2 pixel_5484/AMP_IN pixel_5484/SF_IB
+ pixel_5484/PIX_OUT pixel_5484/CSA_VREF pixel
Xpixel_5495 pixel_5495/gring pixel_5495/VDD pixel_5495/GND pixel_5495/VREF pixel_5495/ROW_SEL
+ pixel_5495/NB1 pixel_5495/VBIAS pixel_5495/NB2 pixel_5495/AMP_IN pixel_5495/SF_IB
+ pixel_5495/PIX_OUT pixel_5495/CSA_VREF pixel
Xpixel_4750 pixel_4750/gring pixel_4750/VDD pixel_4750/GND pixel_4750/VREF pixel_4750/ROW_SEL
+ pixel_4750/NB1 pixel_4750/VBIAS pixel_4750/NB2 pixel_4750/AMP_IN pixel_4750/SF_IB
+ pixel_4750/PIX_OUT pixel_4750/CSA_VREF pixel
Xpixel_4761 pixel_4761/gring pixel_4761/VDD pixel_4761/GND pixel_4761/VREF pixel_4761/ROW_SEL
+ pixel_4761/NB1 pixel_4761/VBIAS pixel_4761/NB2 pixel_4761/AMP_IN pixel_4761/SF_IB
+ pixel_4761/PIX_OUT pixel_4761/CSA_VREF pixel
Xpixel_4772 pixel_4772/gring pixel_4772/VDD pixel_4772/GND pixel_4772/VREF pixel_4772/ROW_SEL
+ pixel_4772/NB1 pixel_4772/VBIAS pixel_4772/NB2 pixel_4772/AMP_IN pixel_4772/SF_IB
+ pixel_4772/PIX_OUT pixel_4772/CSA_VREF pixel
Xpixel_4783 pixel_4783/gring pixel_4783/VDD pixel_4783/GND pixel_4783/VREF pixel_4783/ROW_SEL
+ pixel_4783/NB1 pixel_4783/VBIAS pixel_4783/NB2 pixel_4783/AMP_IN pixel_4783/SF_IB
+ pixel_4783/PIX_OUT pixel_4783/CSA_VREF pixel
Xpixel_4794 pixel_4794/gring pixel_4794/VDD pixel_4794/GND pixel_4794/VREF pixel_4794/ROW_SEL
+ pixel_4794/NB1 pixel_4794/VBIAS pixel_4794/NB2 pixel_4794/AMP_IN pixel_4794/SF_IB
+ pixel_4794/PIX_OUT pixel_4794/CSA_VREF pixel
Xpixel_1409 pixel_1409/gring pixel_1409/VDD pixel_1409/GND pixel_1409/VREF pixel_1409/ROW_SEL
+ pixel_1409/NB1 pixel_1409/VBIAS pixel_1409/NB2 pixel_1409/AMP_IN pixel_1409/SF_IB
+ pixel_1409/PIX_OUT pixel_1409/CSA_VREF pixel
Xpixel_9706 pixel_9706/gring pixel_9706/VDD pixel_9706/GND pixel_9706/VREF pixel_9706/ROW_SEL
+ pixel_9706/NB1 pixel_9706/VBIAS pixel_9706/NB2 pixel_9706/AMP_IN pixel_9706/SF_IB
+ pixel_9706/PIX_OUT pixel_9706/CSA_VREF pixel
Xpixel_9717 pixel_9717/gring pixel_9717/VDD pixel_9717/GND pixel_9717/VREF pixel_9717/ROW_SEL
+ pixel_9717/NB1 pixel_9717/VBIAS pixel_9717/NB2 pixel_9717/AMP_IN pixel_9717/SF_IB
+ pixel_9717/PIX_OUT pixel_9717/CSA_VREF pixel
Xpixel_9728 pixel_9728/gring pixel_9728/VDD pixel_9728/GND pixel_9728/VREF pixel_9728/ROW_SEL
+ pixel_9728/NB1 pixel_9728/VBIAS pixel_9728/NB2 pixel_9728/AMP_IN pixel_9728/SF_IB
+ pixel_9728/PIX_OUT pixel_9728/CSA_VREF pixel
Xpixel_9739 pixel_9739/gring pixel_9739/VDD pixel_9739/GND pixel_9739/VREF pixel_9739/ROW_SEL
+ pixel_9739/NB1 pixel_9739/VBIAS pixel_9739/NB2 pixel_9739/AMP_IN pixel_9739/SF_IB
+ pixel_9739/PIX_OUT pixel_9739/CSA_VREF pixel
Xpixel_4002 pixel_4002/gring pixel_4002/VDD pixel_4002/GND pixel_4002/VREF pixel_4002/ROW_SEL
+ pixel_4002/NB1 pixel_4002/VBIAS pixel_4002/NB2 pixel_4002/AMP_IN pixel_4002/SF_IB
+ pixel_4002/PIX_OUT pixel_4002/CSA_VREF pixel
Xpixel_4013 pixel_4013/gring pixel_4013/VDD pixel_4013/GND pixel_4013/VREF pixel_4013/ROW_SEL
+ pixel_4013/NB1 pixel_4013/VBIAS pixel_4013/NB2 pixel_4013/AMP_IN pixel_4013/SF_IB
+ pixel_4013/PIX_OUT pixel_4013/CSA_VREF pixel
Xpixel_4024 pixel_4024/gring pixel_4024/VDD pixel_4024/GND pixel_4024/VREF pixel_4024/ROW_SEL
+ pixel_4024/NB1 pixel_4024/VBIAS pixel_4024/NB2 pixel_4024/AMP_IN pixel_4024/SF_IB
+ pixel_4024/PIX_OUT pixel_4024/CSA_VREF pixel
Xpixel_4035 pixel_4035/gring pixel_4035/VDD pixel_4035/GND pixel_4035/VREF pixel_4035/ROW_SEL
+ pixel_4035/NB1 pixel_4035/VBIAS pixel_4035/NB2 pixel_4035/AMP_IN pixel_4035/SF_IB
+ pixel_4035/PIX_OUT pixel_4035/CSA_VREF pixel
Xpixel_3323 pixel_3323/gring pixel_3323/VDD pixel_3323/GND pixel_3323/VREF pixel_3323/ROW_SEL
+ pixel_3323/NB1 pixel_3323/VBIAS pixel_3323/NB2 pixel_3323/AMP_IN pixel_3323/SF_IB
+ pixel_3323/PIX_OUT pixel_3323/CSA_VREF pixel
Xpixel_3312 pixel_3312/gring pixel_3312/VDD pixel_3312/GND pixel_3312/VREF pixel_3312/ROW_SEL
+ pixel_3312/NB1 pixel_3312/VBIAS pixel_3312/NB2 pixel_3312/AMP_IN pixel_3312/SF_IB
+ pixel_3312/PIX_OUT pixel_3312/CSA_VREF pixel
Xpixel_3301 pixel_3301/gring pixel_3301/VDD pixel_3301/GND pixel_3301/VREF pixel_3301/ROW_SEL
+ pixel_3301/NB1 pixel_3301/VBIAS pixel_3301/NB2 pixel_3301/AMP_IN pixel_3301/SF_IB
+ pixel_3301/PIX_OUT pixel_3301/CSA_VREF pixel
Xpixel_4046 pixel_4046/gring pixel_4046/VDD pixel_4046/GND pixel_4046/VREF pixel_4046/ROW_SEL
+ pixel_4046/NB1 pixel_4046/VBIAS pixel_4046/NB2 pixel_4046/AMP_IN pixel_4046/SF_IB
+ pixel_4046/PIX_OUT pixel_4046/CSA_VREF pixel
Xpixel_4057 pixel_4057/gring pixel_4057/VDD pixel_4057/GND pixel_4057/VREF pixel_4057/ROW_SEL
+ pixel_4057/NB1 pixel_4057/VBIAS pixel_4057/NB2 pixel_4057/AMP_IN pixel_4057/SF_IB
+ pixel_4057/PIX_OUT pixel_4057/CSA_VREF pixel
Xpixel_4068 pixel_4068/gring pixel_4068/VDD pixel_4068/GND pixel_4068/VREF pixel_4068/ROW_SEL
+ pixel_4068/NB1 pixel_4068/VBIAS pixel_4068/NB2 pixel_4068/AMP_IN pixel_4068/SF_IB
+ pixel_4068/PIX_OUT pixel_4068/CSA_VREF pixel
Xpixel_2622 pixel_2622/gring pixel_2622/VDD pixel_2622/GND pixel_2622/VREF pixel_2622/ROW_SEL
+ pixel_2622/NB1 pixel_2622/VBIAS pixel_2622/NB2 pixel_2622/AMP_IN pixel_2622/SF_IB
+ pixel_2622/PIX_OUT pixel_2622/CSA_VREF pixel
Xpixel_2611 pixel_2611/gring pixel_2611/VDD pixel_2611/GND pixel_2611/VREF pixel_2611/ROW_SEL
+ pixel_2611/NB1 pixel_2611/VBIAS pixel_2611/NB2 pixel_2611/AMP_IN pixel_2611/SF_IB
+ pixel_2611/PIX_OUT pixel_2611/CSA_VREF pixel
Xpixel_2600 pixel_2600/gring pixel_2600/VDD pixel_2600/GND pixel_2600/VREF pixel_2600/ROW_SEL
+ pixel_2600/NB1 pixel_2600/VBIAS pixel_2600/NB2 pixel_2600/AMP_IN pixel_2600/SF_IB
+ pixel_2600/PIX_OUT pixel_2600/CSA_VREF pixel
Xpixel_3367 pixel_3367/gring pixel_3367/VDD pixel_3367/GND pixel_3367/VREF pixel_3367/ROW_SEL
+ pixel_3367/NB1 pixel_3367/VBIAS pixel_3367/NB2 pixel_3367/AMP_IN pixel_3367/SF_IB
+ pixel_3367/PIX_OUT pixel_3367/CSA_VREF pixel
Xpixel_3356 pixel_3356/gring pixel_3356/VDD pixel_3356/GND pixel_3356/VREF pixel_3356/ROW_SEL
+ pixel_3356/NB1 pixel_3356/VBIAS pixel_3356/NB2 pixel_3356/AMP_IN pixel_3356/SF_IB
+ pixel_3356/PIX_OUT pixel_3356/CSA_VREF pixel
Xpixel_3345 pixel_3345/gring pixel_3345/VDD pixel_3345/GND pixel_3345/VREF pixel_3345/ROW_SEL
+ pixel_3345/NB1 pixel_3345/VBIAS pixel_3345/NB2 pixel_3345/AMP_IN pixel_3345/SF_IB
+ pixel_3345/PIX_OUT pixel_3345/CSA_VREF pixel
Xpixel_3334 pixel_3334/gring pixel_3334/VDD pixel_3334/GND pixel_3334/VREF pixel_3334/ROW_SEL
+ pixel_3334/NB1 pixel_3334/VBIAS pixel_3334/NB2 pixel_3334/AMP_IN pixel_3334/SF_IB
+ pixel_3334/PIX_OUT pixel_3334/CSA_VREF pixel
Xpixel_4079 pixel_4079/gring pixel_4079/VDD pixel_4079/GND pixel_4079/VREF pixel_4079/ROW_SEL
+ pixel_4079/NB1 pixel_4079/VBIAS pixel_4079/NB2 pixel_4079/AMP_IN pixel_4079/SF_IB
+ pixel_4079/PIX_OUT pixel_4079/CSA_VREF pixel
Xpixel_1910 pixel_1910/gring pixel_1910/VDD pixel_1910/GND pixel_1910/VREF pixel_1910/ROW_SEL
+ pixel_1910/NB1 pixel_1910/VBIAS pixel_1910/NB2 pixel_1910/AMP_IN pixel_1910/SF_IB
+ pixel_1910/PIX_OUT pixel_1910/CSA_VREF pixel
Xpixel_2655 pixel_2655/gring pixel_2655/VDD pixel_2655/GND pixel_2655/VREF pixel_2655/ROW_SEL
+ pixel_2655/NB1 pixel_2655/VBIAS pixel_2655/NB2 pixel_2655/AMP_IN pixel_2655/SF_IB
+ pixel_2655/PIX_OUT pixel_2655/CSA_VREF pixel
Xpixel_2644 pixel_2644/gring pixel_2644/VDD pixel_2644/GND pixel_2644/VREF pixel_2644/ROW_SEL
+ pixel_2644/NB1 pixel_2644/VBIAS pixel_2644/NB2 pixel_2644/AMP_IN pixel_2644/SF_IB
+ pixel_2644/PIX_OUT pixel_2644/CSA_VREF pixel
Xpixel_2633 pixel_2633/gring pixel_2633/VDD pixel_2633/GND pixel_2633/VREF pixel_2633/ROW_SEL
+ pixel_2633/NB1 pixel_2633/VBIAS pixel_2633/NB2 pixel_2633/AMP_IN pixel_2633/SF_IB
+ pixel_2633/PIX_OUT pixel_2633/CSA_VREF pixel
Xpixel_3389 pixel_3389/gring pixel_3389/VDD pixel_3389/GND pixel_3389/VREF pixel_3389/ROW_SEL
+ pixel_3389/NB1 pixel_3389/VBIAS pixel_3389/NB2 pixel_3389/AMP_IN pixel_3389/SF_IB
+ pixel_3389/PIX_OUT pixel_3389/CSA_VREF pixel
Xpixel_3378 pixel_3378/gring pixel_3378/VDD pixel_3378/GND pixel_3378/VREF pixel_3378/ROW_SEL
+ pixel_3378/NB1 pixel_3378/VBIAS pixel_3378/NB2 pixel_3378/AMP_IN pixel_3378/SF_IB
+ pixel_3378/PIX_OUT pixel_3378/CSA_VREF pixel
Xpixel_1943 pixel_1943/gring pixel_1943/VDD pixel_1943/GND pixel_1943/VREF pixel_1943/ROW_SEL
+ pixel_1943/NB1 pixel_1943/VBIAS pixel_1943/NB2 pixel_1943/AMP_IN pixel_1943/SF_IB
+ pixel_1943/PIX_OUT pixel_1943/CSA_VREF pixel
Xpixel_1932 pixel_1932/gring pixel_1932/VDD pixel_1932/GND pixel_1932/VREF pixel_1932/ROW_SEL
+ pixel_1932/NB1 pixel_1932/VBIAS pixel_1932/NB2 pixel_1932/AMP_IN pixel_1932/SF_IB
+ pixel_1932/PIX_OUT pixel_1932/CSA_VREF pixel
Xpixel_1921 pixel_1921/gring pixel_1921/VDD pixel_1921/GND pixel_1921/VREF pixel_1921/ROW_SEL
+ pixel_1921/NB1 pixel_1921/VBIAS pixel_1921/NB2 pixel_1921/AMP_IN pixel_1921/SF_IB
+ pixel_1921/PIX_OUT pixel_1921/CSA_VREF pixel
Xpixel_2688 pixel_2688/gring pixel_2688/VDD pixel_2688/GND pixel_2688/VREF pixel_2688/ROW_SEL
+ pixel_2688/NB1 pixel_2688/VBIAS pixel_2688/NB2 pixel_2688/AMP_IN pixel_2688/SF_IB
+ pixel_2688/PIX_OUT pixel_2688/CSA_VREF pixel
Xpixel_2677 pixel_2677/gring pixel_2677/VDD pixel_2677/GND pixel_2677/VREF pixel_2677/ROW_SEL
+ pixel_2677/NB1 pixel_2677/VBIAS pixel_2677/NB2 pixel_2677/AMP_IN pixel_2677/SF_IB
+ pixel_2677/PIX_OUT pixel_2677/CSA_VREF pixel
Xpixel_2666 pixel_2666/gring pixel_2666/VDD pixel_2666/GND pixel_2666/VREF pixel_2666/ROW_SEL
+ pixel_2666/NB1 pixel_2666/VBIAS pixel_2666/NB2 pixel_2666/AMP_IN pixel_2666/SF_IB
+ pixel_2666/PIX_OUT pixel_2666/CSA_VREF pixel
Xpixel_1987 pixel_1987/gring pixel_1987/VDD pixel_1987/GND pixel_1987/VREF pixel_1987/ROW_SEL
+ pixel_1987/NB1 pixel_1987/VBIAS pixel_1987/NB2 pixel_1987/AMP_IN pixel_1987/SF_IB
+ pixel_1987/PIX_OUT pixel_1987/CSA_VREF pixel
Xpixel_1976 pixel_1976/gring pixel_1976/VDD pixel_1976/GND pixel_1976/VREF pixel_1976/ROW_SEL
+ pixel_1976/NB1 pixel_1976/VBIAS pixel_1976/NB2 pixel_1976/AMP_IN pixel_1976/SF_IB
+ pixel_1976/PIX_OUT pixel_1976/CSA_VREF pixel
Xpixel_1965 pixel_1965/gring pixel_1965/VDD pixel_1965/GND pixel_1965/VREF pixel_1965/ROW_SEL
+ pixel_1965/NB1 pixel_1965/VBIAS pixel_1965/NB2 pixel_1965/AMP_IN pixel_1965/SF_IB
+ pixel_1965/PIX_OUT pixel_1965/CSA_VREF pixel
Xpixel_1954 pixel_1954/gring pixel_1954/VDD pixel_1954/GND pixel_1954/VREF pixel_1954/ROW_SEL
+ pixel_1954/NB1 pixel_1954/VBIAS pixel_1954/NB2 pixel_1954/AMP_IN pixel_1954/SF_IB
+ pixel_1954/PIX_OUT pixel_1954/CSA_VREF pixel
Xpixel_2699 pixel_2699/gring pixel_2699/VDD pixel_2699/GND pixel_2699/VREF pixel_2699/ROW_SEL
+ pixel_2699/NB1 pixel_2699/VBIAS pixel_2699/NB2 pixel_2699/AMP_IN pixel_2699/SF_IB
+ pixel_2699/PIX_OUT pixel_2699/CSA_VREF pixel
Xpixel_1998 pixel_1998/gring pixel_1998/VDD pixel_1998/GND pixel_1998/VREF pixel_1998/ROW_SEL
+ pixel_1998/NB1 pixel_1998/VBIAS pixel_1998/NB2 pixel_1998/AMP_IN pixel_1998/SF_IB
+ pixel_1998/PIX_OUT pixel_1998/CSA_VREF pixel
Xpixel_5270 pixel_5270/gring pixel_5270/VDD pixel_5270/GND pixel_5270/VREF pixel_5270/ROW_SEL
+ pixel_5270/NB1 pixel_5270/VBIAS pixel_5270/NB2 pixel_5270/AMP_IN pixel_5270/SF_IB
+ pixel_5270/PIX_OUT pixel_5270/CSA_VREF pixel
Xpixel_5281 pixel_5281/gring pixel_5281/VDD pixel_5281/GND pixel_5281/VREF pixel_5281/ROW_SEL
+ pixel_5281/NB1 pixel_5281/VBIAS pixel_5281/NB2 pixel_5281/AMP_IN pixel_5281/SF_IB
+ pixel_5281/PIX_OUT pixel_5281/CSA_VREF pixel
Xpixel_5292 pixel_5292/gring pixel_5292/VDD pixel_5292/GND pixel_5292/VREF pixel_5292/ROW_SEL
+ pixel_5292/NB1 pixel_5292/VBIAS pixel_5292/NB2 pixel_5292/AMP_IN pixel_5292/SF_IB
+ pixel_5292/PIX_OUT pixel_5292/CSA_VREF pixel
Xpixel_4580 pixel_4580/gring pixel_4580/VDD pixel_4580/GND pixel_4580/VREF pixel_4580/ROW_SEL
+ pixel_4580/NB1 pixel_4580/VBIAS pixel_4580/NB2 pixel_4580/AMP_IN pixel_4580/SF_IB
+ pixel_4580/PIX_OUT pixel_4580/CSA_VREF pixel
Xpixel_4591 pixel_4591/gring pixel_4591/VDD pixel_4591/GND pixel_4591/VREF pixel_4591/ROW_SEL
+ pixel_4591/NB1 pixel_4591/VBIAS pixel_4591/NB2 pixel_4591/AMP_IN pixel_4591/SF_IB
+ pixel_4591/PIX_OUT pixel_4591/CSA_VREF pixel
Xpixel_3890 pixel_3890/gring pixel_3890/VDD pixel_3890/GND pixel_3890/VREF pixel_3890/ROW_SEL
+ pixel_3890/NB1 pixel_3890/VBIAS pixel_3890/NB2 pixel_3890/AMP_IN pixel_3890/SF_IB
+ pixel_3890/PIX_OUT pixel_3890/CSA_VREF pixel
Xpixel_1206 pixel_1206/gring pixel_1206/VDD pixel_1206/GND pixel_1206/VREF pixel_1206/ROW_SEL
+ pixel_1206/NB1 pixel_1206/VBIAS pixel_1206/NB2 pixel_1206/AMP_IN pixel_1206/SF_IB
+ pixel_1206/PIX_OUT pixel_1206/CSA_VREF pixel
Xpixel_1239 pixel_1239/gring pixel_1239/VDD pixel_1239/GND pixel_1239/VREF pixel_1239/ROW_SEL
+ pixel_1239/NB1 pixel_1239/VBIAS pixel_1239/NB2 pixel_1239/AMP_IN pixel_1239/SF_IB
+ pixel_1239/PIX_OUT pixel_1239/CSA_VREF pixel
Xpixel_1228 pixel_1228/gring pixel_1228/VDD pixel_1228/GND pixel_1228/VREF pixel_1228/ROW_SEL
+ pixel_1228/NB1 pixel_1228/VBIAS pixel_1228/NB2 pixel_1228/AMP_IN pixel_1228/SF_IB
+ pixel_1228/PIX_OUT pixel_1228/CSA_VREF pixel
Xpixel_1217 pixel_1217/gring pixel_1217/VDD pixel_1217/GND pixel_1217/VREF pixel_1217/ROW_SEL
+ pixel_1217/NB1 pixel_1217/VBIAS pixel_1217/NB2 pixel_1217/AMP_IN pixel_1217/SF_IB
+ pixel_1217/PIX_OUT pixel_1217/CSA_VREF pixel
Xpixel_9514 pixel_9514/gring pixel_9514/VDD pixel_9514/GND pixel_9514/VREF pixel_9514/ROW_SEL
+ pixel_9514/NB1 pixel_9514/VBIAS pixel_9514/NB2 pixel_9514/AMP_IN pixel_9514/SF_IB
+ pixel_9514/PIX_OUT pixel_9514/CSA_VREF pixel
Xpixel_9503 pixel_9503/gring pixel_9503/VDD pixel_9503/GND pixel_9503/VREF pixel_9503/ROW_SEL
+ pixel_9503/NB1 pixel_9503/VBIAS pixel_9503/NB2 pixel_9503/AMP_IN pixel_9503/SF_IB
+ pixel_9503/PIX_OUT pixel_9503/CSA_VREF pixel
Xpixel_8802 pixel_8802/gring pixel_8802/VDD pixel_8802/GND pixel_8802/VREF pixel_8802/ROW_SEL
+ pixel_8802/NB1 pixel_8802/VBIAS pixel_8802/NB2 pixel_8802/AMP_IN pixel_8802/SF_IB
+ pixel_8802/PIX_OUT pixel_8802/CSA_VREF pixel
Xpixel_9547 pixel_9547/gring pixel_9547/VDD pixel_9547/GND pixel_9547/VREF pixel_9547/ROW_SEL
+ pixel_9547/NB1 pixel_9547/VBIAS pixel_9547/NB2 pixel_9547/AMP_IN pixel_9547/SF_IB
+ pixel_9547/PIX_OUT pixel_9547/CSA_VREF pixel
Xpixel_9536 pixel_9536/gring pixel_9536/VDD pixel_9536/GND pixel_9536/VREF pixel_9536/ROW_SEL
+ pixel_9536/NB1 pixel_9536/VBIAS pixel_9536/NB2 pixel_9536/AMP_IN pixel_9536/SF_IB
+ pixel_9536/PIX_OUT pixel_9536/CSA_VREF pixel
Xpixel_9525 pixel_9525/gring pixel_9525/VDD pixel_9525/GND pixel_9525/VREF pixel_9525/ROW_SEL
+ pixel_9525/NB1 pixel_9525/VBIAS pixel_9525/NB2 pixel_9525/AMP_IN pixel_9525/SF_IB
+ pixel_9525/PIX_OUT pixel_9525/CSA_VREF pixel
Xpixel_8846 pixel_8846/gring pixel_8846/VDD pixel_8846/GND pixel_8846/VREF pixel_8846/ROW_SEL
+ pixel_8846/NB1 pixel_8846/VBIAS pixel_8846/NB2 pixel_8846/AMP_IN pixel_8846/SF_IB
+ pixel_8846/PIX_OUT pixel_8846/CSA_VREF pixel
Xpixel_8835 pixel_8835/gring pixel_8835/VDD pixel_8835/GND pixel_8835/VREF pixel_8835/ROW_SEL
+ pixel_8835/NB1 pixel_8835/VBIAS pixel_8835/NB2 pixel_8835/AMP_IN pixel_8835/SF_IB
+ pixel_8835/PIX_OUT pixel_8835/CSA_VREF pixel
Xpixel_8824 pixel_8824/gring pixel_8824/VDD pixel_8824/GND pixel_8824/VREF pixel_8824/ROW_SEL
+ pixel_8824/NB1 pixel_8824/VBIAS pixel_8824/NB2 pixel_8824/AMP_IN pixel_8824/SF_IB
+ pixel_8824/PIX_OUT pixel_8824/CSA_VREF pixel
Xpixel_8813 pixel_8813/gring pixel_8813/VDD pixel_8813/GND pixel_8813/VREF pixel_8813/ROW_SEL
+ pixel_8813/NB1 pixel_8813/VBIAS pixel_8813/NB2 pixel_8813/AMP_IN pixel_8813/SF_IB
+ pixel_8813/PIX_OUT pixel_8813/CSA_VREF pixel
Xpixel_9569 pixel_9569/gring pixel_9569/VDD pixel_9569/GND pixel_9569/VREF pixel_9569/ROW_SEL
+ pixel_9569/NB1 pixel_9569/VBIAS pixel_9569/NB2 pixel_9569/AMP_IN pixel_9569/SF_IB
+ pixel_9569/PIX_OUT pixel_9569/CSA_VREF pixel
Xpixel_9558 pixel_9558/gring pixel_9558/VDD pixel_9558/GND pixel_9558/VREF pixel_9558/ROW_SEL
+ pixel_9558/NB1 pixel_9558/VBIAS pixel_9558/NB2 pixel_9558/AMP_IN pixel_9558/SF_IB
+ pixel_9558/PIX_OUT pixel_9558/CSA_VREF pixel
Xpixel_8879 pixel_8879/gring pixel_8879/VDD pixel_8879/GND pixel_8879/VREF pixel_8879/ROW_SEL
+ pixel_8879/NB1 pixel_8879/VBIAS pixel_8879/NB2 pixel_8879/AMP_IN pixel_8879/SF_IB
+ pixel_8879/PIX_OUT pixel_8879/CSA_VREF pixel
Xpixel_8868 pixel_8868/gring pixel_8868/VDD pixel_8868/GND pixel_8868/VREF pixel_8868/ROW_SEL
+ pixel_8868/NB1 pixel_8868/VBIAS pixel_8868/NB2 pixel_8868/AMP_IN pixel_8868/SF_IB
+ pixel_8868/PIX_OUT pixel_8868/CSA_VREF pixel
Xpixel_8857 pixel_8857/gring pixel_8857/VDD pixel_8857/GND pixel_8857/VREF pixel_8857/ROW_SEL
+ pixel_8857/NB1 pixel_8857/VBIAS pixel_8857/NB2 pixel_8857/AMP_IN pixel_8857/SF_IB
+ pixel_8857/PIX_OUT pixel_8857/CSA_VREF pixel
Xpixel_3131 pixel_3131/gring pixel_3131/VDD pixel_3131/GND pixel_3131/VREF pixel_3131/ROW_SEL
+ pixel_3131/NB1 pixel_3131/VBIAS pixel_3131/NB2 pixel_3131/AMP_IN pixel_3131/SF_IB
+ pixel_3131/PIX_OUT pixel_3131/CSA_VREF pixel
Xpixel_3120 pixel_3120/gring pixel_3120/VDD pixel_3120/GND pixel_3120/VREF pixel_3120/ROW_SEL
+ pixel_3120/NB1 pixel_3120/VBIAS pixel_3120/NB2 pixel_3120/AMP_IN pixel_3120/SF_IB
+ pixel_3120/PIX_OUT pixel_3120/CSA_VREF pixel
Xpixel_2430 pixel_2430/gring pixel_2430/VDD pixel_2430/GND pixel_2430/VREF pixel_2430/ROW_SEL
+ pixel_2430/NB1 pixel_2430/VBIAS pixel_2430/NB2 pixel_2430/AMP_IN pixel_2430/SF_IB
+ pixel_2430/PIX_OUT pixel_2430/CSA_VREF pixel
Xpixel_3175 pixel_3175/gring pixel_3175/VDD pixel_3175/GND pixel_3175/VREF pixel_3175/ROW_SEL
+ pixel_3175/NB1 pixel_3175/VBIAS pixel_3175/NB2 pixel_3175/AMP_IN pixel_3175/SF_IB
+ pixel_3175/PIX_OUT pixel_3175/CSA_VREF pixel
Xpixel_3164 pixel_3164/gring pixel_3164/VDD pixel_3164/GND pixel_3164/VREF pixel_3164/ROW_SEL
+ pixel_3164/NB1 pixel_3164/VBIAS pixel_3164/NB2 pixel_3164/AMP_IN pixel_3164/SF_IB
+ pixel_3164/PIX_OUT pixel_3164/CSA_VREF pixel
Xpixel_3153 pixel_3153/gring pixel_3153/VDD pixel_3153/GND pixel_3153/VREF pixel_3153/ROW_SEL
+ pixel_3153/NB1 pixel_3153/VBIAS pixel_3153/NB2 pixel_3153/AMP_IN pixel_3153/SF_IB
+ pixel_3153/PIX_OUT pixel_3153/CSA_VREF pixel
Xpixel_3142 pixel_3142/gring pixel_3142/VDD pixel_3142/GND pixel_3142/VREF pixel_3142/ROW_SEL
+ pixel_3142/NB1 pixel_3142/VBIAS pixel_3142/NB2 pixel_3142/AMP_IN pixel_3142/SF_IB
+ pixel_3142/PIX_OUT pixel_3142/CSA_VREF pixel
Xpixel_2463 pixel_2463/gring pixel_2463/VDD pixel_2463/GND pixel_2463/VREF pixel_2463/ROW_SEL
+ pixel_2463/NB1 pixel_2463/VBIAS pixel_2463/NB2 pixel_2463/AMP_IN pixel_2463/SF_IB
+ pixel_2463/PIX_OUT pixel_2463/CSA_VREF pixel
Xpixel_2452 pixel_2452/gring pixel_2452/VDD pixel_2452/GND pixel_2452/VREF pixel_2452/ROW_SEL
+ pixel_2452/NB1 pixel_2452/VBIAS pixel_2452/NB2 pixel_2452/AMP_IN pixel_2452/SF_IB
+ pixel_2452/PIX_OUT pixel_2452/CSA_VREF pixel
Xpixel_2441 pixel_2441/gring pixel_2441/VDD pixel_2441/GND pixel_2441/VREF pixel_2441/ROW_SEL
+ pixel_2441/NB1 pixel_2441/VBIAS pixel_2441/NB2 pixel_2441/AMP_IN pixel_2441/SF_IB
+ pixel_2441/PIX_OUT pixel_2441/CSA_VREF pixel
Xpixel_3197 pixel_3197/gring pixel_3197/VDD pixel_3197/GND pixel_3197/VREF pixel_3197/ROW_SEL
+ pixel_3197/NB1 pixel_3197/VBIAS pixel_3197/NB2 pixel_3197/AMP_IN pixel_3197/SF_IB
+ pixel_3197/PIX_OUT pixel_3197/CSA_VREF pixel
Xpixel_3186 pixel_3186/gring pixel_3186/VDD pixel_3186/GND pixel_3186/VREF pixel_3186/ROW_SEL
+ pixel_3186/NB1 pixel_3186/VBIAS pixel_3186/NB2 pixel_3186/AMP_IN pixel_3186/SF_IB
+ pixel_3186/PIX_OUT pixel_3186/CSA_VREF pixel
Xpixel_1762 pixel_1762/gring pixel_1762/VDD pixel_1762/GND pixel_1762/VREF pixel_1762/ROW_SEL
+ pixel_1762/NB1 pixel_1762/VBIAS pixel_1762/NB2 pixel_1762/AMP_IN pixel_1762/SF_IB
+ pixel_1762/PIX_OUT pixel_1762/CSA_VREF pixel
Xpixel_1751 pixel_1751/gring pixel_1751/VDD pixel_1751/GND pixel_1751/VREF pixel_1751/ROW_SEL
+ pixel_1751/NB1 pixel_1751/VBIAS pixel_1751/NB2 pixel_1751/AMP_IN pixel_1751/SF_IB
+ pixel_1751/PIX_OUT pixel_1751/CSA_VREF pixel
Xpixel_1740 pixel_1740/gring pixel_1740/VDD pixel_1740/GND pixel_1740/VREF pixel_1740/ROW_SEL
+ pixel_1740/NB1 pixel_1740/VBIAS pixel_1740/NB2 pixel_1740/AMP_IN pixel_1740/SF_IB
+ pixel_1740/PIX_OUT pixel_1740/CSA_VREF pixel
Xpixel_2496 pixel_2496/gring pixel_2496/VDD pixel_2496/GND pixel_2496/VREF pixel_2496/ROW_SEL
+ pixel_2496/NB1 pixel_2496/VBIAS pixel_2496/NB2 pixel_2496/AMP_IN pixel_2496/SF_IB
+ pixel_2496/PIX_OUT pixel_2496/CSA_VREF pixel
Xpixel_2485 pixel_2485/gring pixel_2485/VDD pixel_2485/GND pixel_2485/VREF pixel_2485/ROW_SEL
+ pixel_2485/NB1 pixel_2485/VBIAS pixel_2485/NB2 pixel_2485/AMP_IN pixel_2485/SF_IB
+ pixel_2485/PIX_OUT pixel_2485/CSA_VREF pixel
Xpixel_2474 pixel_2474/gring pixel_2474/VDD pixel_2474/GND pixel_2474/VREF pixel_2474/ROW_SEL
+ pixel_2474/NB1 pixel_2474/VBIAS pixel_2474/NB2 pixel_2474/AMP_IN pixel_2474/SF_IB
+ pixel_2474/PIX_OUT pixel_2474/CSA_VREF pixel
Xpixel_1795 pixel_1795/gring pixel_1795/VDD pixel_1795/GND pixel_1795/VREF pixel_1795/ROW_SEL
+ pixel_1795/NB1 pixel_1795/VBIAS pixel_1795/NB2 pixel_1795/AMP_IN pixel_1795/SF_IB
+ pixel_1795/PIX_OUT pixel_1795/CSA_VREF pixel
Xpixel_1784 pixel_1784/gring pixel_1784/VDD pixel_1784/GND pixel_1784/VREF pixel_1784/ROW_SEL
+ pixel_1784/NB1 pixel_1784/VBIAS pixel_1784/NB2 pixel_1784/AMP_IN pixel_1784/SF_IB
+ pixel_1784/PIX_OUT pixel_1784/CSA_VREF pixel
Xpixel_1773 pixel_1773/gring pixel_1773/VDD pixel_1773/GND pixel_1773/VREF pixel_1773/ROW_SEL
+ pixel_1773/NB1 pixel_1773/VBIAS pixel_1773/NB2 pixel_1773/AMP_IN pixel_1773/SF_IB
+ pixel_1773/PIX_OUT pixel_1773/CSA_VREF pixel
Xpixel_8109 pixel_8109/gring pixel_8109/VDD pixel_8109/GND pixel_8109/VREF pixel_8109/ROW_SEL
+ pixel_8109/NB1 pixel_8109/VBIAS pixel_8109/NB2 pixel_8109/AMP_IN pixel_8109/SF_IB
+ pixel_8109/PIX_OUT pixel_8109/CSA_VREF pixel
Xpixel_7408 pixel_7408/gring pixel_7408/VDD pixel_7408/GND pixel_7408/VREF pixel_7408/ROW_SEL
+ pixel_7408/NB1 pixel_7408/VBIAS pixel_7408/NB2 pixel_7408/AMP_IN pixel_7408/SF_IB
+ pixel_7408/PIX_OUT pixel_7408/CSA_VREF pixel
Xpixel_7419 pixel_7419/gring pixel_7419/VDD pixel_7419/GND pixel_7419/VREF pixel_7419/ROW_SEL
+ pixel_7419/NB1 pixel_7419/VBIAS pixel_7419/NB2 pixel_7419/AMP_IN pixel_7419/SF_IB
+ pixel_7419/PIX_OUT pixel_7419/CSA_VREF pixel
Xpixel_6707 pixel_6707/gring pixel_6707/VDD pixel_6707/GND pixel_6707/VREF pixel_6707/ROW_SEL
+ pixel_6707/NB1 pixel_6707/VBIAS pixel_6707/NB2 pixel_6707/AMP_IN pixel_6707/SF_IB
+ pixel_6707/PIX_OUT pixel_6707/CSA_VREF pixel
Xpixel_6718 pixel_6718/gring pixel_6718/VDD pixel_6718/GND pixel_6718/VREF pixel_6718/ROW_SEL
+ pixel_6718/NB1 pixel_6718/VBIAS pixel_6718/NB2 pixel_6718/AMP_IN pixel_6718/SF_IB
+ pixel_6718/PIX_OUT pixel_6718/CSA_VREF pixel
Xpixel_6729 pixel_6729/gring pixel_6729/VDD pixel_6729/GND pixel_6729/VREF pixel_6729/ROW_SEL
+ pixel_6729/NB1 pixel_6729/VBIAS pixel_6729/NB2 pixel_6729/AMP_IN pixel_6729/SF_IB
+ pixel_6729/PIX_OUT pixel_6729/CSA_VREF pixel
Xpixel_1014 pixel_1014/gring pixel_1014/VDD pixel_1014/GND pixel_1014/VREF pixel_1014/ROW_SEL
+ pixel_1014/NB1 pixel_1014/VBIAS pixel_1014/NB2 pixel_1014/AMP_IN pixel_1014/SF_IB
+ pixel_1014/PIX_OUT pixel_1014/CSA_VREF pixel
Xpixel_1003 pixel_1003/gring pixel_1003/VDD pixel_1003/GND pixel_1003/VREF pixel_1003/ROW_SEL
+ pixel_1003/NB1 pixel_1003/VBIAS pixel_1003/NB2 pixel_1003/AMP_IN pixel_1003/SF_IB
+ pixel_1003/PIX_OUT pixel_1003/CSA_VREF pixel
Xpixel_1047 pixel_1047/gring pixel_1047/VDD pixel_1047/GND pixel_1047/VREF pixel_1047/ROW_SEL
+ pixel_1047/NB1 pixel_1047/VBIAS pixel_1047/NB2 pixel_1047/AMP_IN pixel_1047/SF_IB
+ pixel_1047/PIX_OUT pixel_1047/CSA_VREF pixel
Xpixel_1036 pixel_1036/gring pixel_1036/VDD pixel_1036/GND pixel_1036/VREF pixel_1036/ROW_SEL
+ pixel_1036/NB1 pixel_1036/VBIAS pixel_1036/NB2 pixel_1036/AMP_IN pixel_1036/SF_IB
+ pixel_1036/PIX_OUT pixel_1036/CSA_VREF pixel
Xpixel_1025 pixel_1025/gring pixel_1025/VDD pixel_1025/GND pixel_1025/VREF pixel_1025/ROW_SEL
+ pixel_1025/NB1 pixel_1025/VBIAS pixel_1025/NB2 pixel_1025/AMP_IN pixel_1025/SF_IB
+ pixel_1025/PIX_OUT pixel_1025/CSA_VREF pixel
Xpixel_1069 pixel_1069/gring pixel_1069/VDD pixel_1069/GND pixel_1069/VREF pixel_1069/ROW_SEL
+ pixel_1069/NB1 pixel_1069/VBIAS pixel_1069/NB2 pixel_1069/AMP_IN pixel_1069/SF_IB
+ pixel_1069/PIX_OUT pixel_1069/CSA_VREF pixel
Xpixel_1058 pixel_1058/gring pixel_1058/VDD pixel_1058/GND pixel_1058/VREF pixel_1058/ROW_SEL
+ pixel_1058/NB1 pixel_1058/VBIAS pixel_1058/NB2 pixel_1058/AMP_IN pixel_1058/SF_IB
+ pixel_1058/PIX_OUT pixel_1058/CSA_VREF pixel
Xpixel_9322 pixel_9322/gring pixel_9322/VDD pixel_9322/GND pixel_9322/VREF pixel_9322/ROW_SEL
+ pixel_9322/NB1 pixel_9322/VBIAS pixel_9322/NB2 pixel_9322/AMP_IN pixel_9322/SF_IB
+ pixel_9322/PIX_OUT pixel_9322/CSA_VREF pixel
Xpixel_9311 pixel_9311/gring pixel_9311/VDD pixel_9311/GND pixel_9311/VREF pixel_9311/ROW_SEL
+ pixel_9311/NB1 pixel_9311/VBIAS pixel_9311/NB2 pixel_9311/AMP_IN pixel_9311/SF_IB
+ pixel_9311/PIX_OUT pixel_9311/CSA_VREF pixel
Xpixel_9300 pixel_9300/gring pixel_9300/VDD pixel_9300/GND pixel_9300/VREF pixel_9300/ROW_SEL
+ pixel_9300/NB1 pixel_9300/VBIAS pixel_9300/NB2 pixel_9300/AMP_IN pixel_9300/SF_IB
+ pixel_9300/PIX_OUT pixel_9300/CSA_VREF pixel
Xpixel_8610 pixel_8610/gring pixel_8610/VDD pixel_8610/GND pixel_8610/VREF pixel_8610/ROW_SEL
+ pixel_8610/NB1 pixel_8610/VBIAS pixel_8610/NB2 pixel_8610/AMP_IN pixel_8610/SF_IB
+ pixel_8610/PIX_OUT pixel_8610/CSA_VREF pixel
Xpixel_9355 pixel_9355/gring pixel_9355/VDD pixel_9355/GND pixel_9355/VREF pixel_9355/ROW_SEL
+ pixel_9355/NB1 pixel_9355/VBIAS pixel_9355/NB2 pixel_9355/AMP_IN pixel_9355/SF_IB
+ pixel_9355/PIX_OUT pixel_9355/CSA_VREF pixel
Xpixel_9344 pixel_9344/gring pixel_9344/VDD pixel_9344/GND pixel_9344/VREF pixel_9344/ROW_SEL
+ pixel_9344/NB1 pixel_9344/VBIAS pixel_9344/NB2 pixel_9344/AMP_IN pixel_9344/SF_IB
+ pixel_9344/PIX_OUT pixel_9344/CSA_VREF pixel
Xpixel_9333 pixel_9333/gring pixel_9333/VDD pixel_9333/GND pixel_9333/VREF pixel_9333/ROW_SEL
+ pixel_9333/NB1 pixel_9333/VBIAS pixel_9333/NB2 pixel_9333/AMP_IN pixel_9333/SF_IB
+ pixel_9333/PIX_OUT pixel_9333/CSA_VREF pixel
Xpixel_8654 pixel_8654/gring pixel_8654/VDD pixel_8654/GND pixel_8654/VREF pixel_8654/ROW_SEL
+ pixel_8654/NB1 pixel_8654/VBIAS pixel_8654/NB2 pixel_8654/AMP_IN pixel_8654/SF_IB
+ pixel_8654/PIX_OUT pixel_8654/CSA_VREF pixel
Xpixel_8643 pixel_8643/gring pixel_8643/VDD pixel_8643/GND pixel_8643/VREF pixel_8643/ROW_SEL
+ pixel_8643/NB1 pixel_8643/VBIAS pixel_8643/NB2 pixel_8643/AMP_IN pixel_8643/SF_IB
+ pixel_8643/PIX_OUT pixel_8643/CSA_VREF pixel
Xpixel_8632 pixel_8632/gring pixel_8632/VDD pixel_8632/GND pixel_8632/VREF pixel_8632/ROW_SEL
+ pixel_8632/NB1 pixel_8632/VBIAS pixel_8632/NB2 pixel_8632/AMP_IN pixel_8632/SF_IB
+ pixel_8632/PIX_OUT pixel_8632/CSA_VREF pixel
Xpixel_8621 pixel_8621/gring pixel_8621/VDD pixel_8621/GND pixel_8621/VREF pixel_8621/ROW_SEL
+ pixel_8621/NB1 pixel_8621/VBIAS pixel_8621/NB2 pixel_8621/AMP_IN pixel_8621/SF_IB
+ pixel_8621/PIX_OUT pixel_8621/CSA_VREF pixel
Xpixel_9399 pixel_9399/gring pixel_9399/VDD pixel_9399/GND pixel_9399/VREF pixel_9399/ROW_SEL
+ pixel_9399/NB1 pixel_9399/VBIAS pixel_9399/NB2 pixel_9399/AMP_IN pixel_9399/SF_IB
+ pixel_9399/PIX_OUT pixel_9399/CSA_VREF pixel
Xpixel_9388 pixel_9388/gring pixel_9388/VDD pixel_9388/GND pixel_9388/VREF pixel_9388/ROW_SEL
+ pixel_9388/NB1 pixel_9388/VBIAS pixel_9388/NB2 pixel_9388/AMP_IN pixel_9388/SF_IB
+ pixel_9388/PIX_OUT pixel_9388/CSA_VREF pixel
Xpixel_9377 pixel_9377/gring pixel_9377/VDD pixel_9377/GND pixel_9377/VREF pixel_9377/ROW_SEL
+ pixel_9377/NB1 pixel_9377/VBIAS pixel_9377/NB2 pixel_9377/AMP_IN pixel_9377/SF_IB
+ pixel_9377/PIX_OUT pixel_9377/CSA_VREF pixel
Xpixel_9366 pixel_9366/gring pixel_9366/VDD pixel_9366/GND pixel_9366/VREF pixel_9366/ROW_SEL
+ pixel_9366/NB1 pixel_9366/VBIAS pixel_9366/NB2 pixel_9366/AMP_IN pixel_9366/SF_IB
+ pixel_9366/PIX_OUT pixel_9366/CSA_VREF pixel
Xpixel_8687 pixel_8687/gring pixel_8687/VDD pixel_8687/GND pixel_8687/VREF pixel_8687/ROW_SEL
+ pixel_8687/NB1 pixel_8687/VBIAS pixel_8687/NB2 pixel_8687/AMP_IN pixel_8687/SF_IB
+ pixel_8687/PIX_OUT pixel_8687/CSA_VREF pixel
Xpixel_8676 pixel_8676/gring pixel_8676/VDD pixel_8676/GND pixel_8676/VREF pixel_8676/ROW_SEL
+ pixel_8676/NB1 pixel_8676/VBIAS pixel_8676/NB2 pixel_8676/AMP_IN pixel_8676/SF_IB
+ pixel_8676/PIX_OUT pixel_8676/CSA_VREF pixel
Xpixel_8665 pixel_8665/gring pixel_8665/VDD pixel_8665/GND pixel_8665/VREF pixel_8665/ROW_SEL
+ pixel_8665/NB1 pixel_8665/VBIAS pixel_8665/NB2 pixel_8665/AMP_IN pixel_8665/SF_IB
+ pixel_8665/PIX_OUT pixel_8665/CSA_VREF pixel
Xpixel_7920 pixel_7920/gring pixel_7920/VDD pixel_7920/GND pixel_7920/VREF pixel_7920/ROW_SEL
+ pixel_7920/NB1 pixel_7920/VBIAS pixel_7920/NB2 pixel_7920/AMP_IN pixel_7920/SF_IB
+ pixel_7920/PIX_OUT pixel_7920/CSA_VREF pixel
Xpixel_7931 pixel_7931/gring pixel_7931/VDD pixel_7931/GND pixel_7931/VREF pixel_7931/ROW_SEL
+ pixel_7931/NB1 pixel_7931/VBIAS pixel_7931/NB2 pixel_7931/AMP_IN pixel_7931/SF_IB
+ pixel_7931/PIX_OUT pixel_7931/CSA_VREF pixel
Xpixel_7942 pixel_7942/gring pixel_7942/VDD pixel_7942/GND pixel_7942/VREF pixel_7942/ROW_SEL
+ pixel_7942/NB1 pixel_7942/VBIAS pixel_7942/NB2 pixel_7942/AMP_IN pixel_7942/SF_IB
+ pixel_7942/PIX_OUT pixel_7942/CSA_VREF pixel
Xpixel_8698 pixel_8698/gring pixel_8698/VDD pixel_8698/GND pixel_8698/VREF pixel_8698/ROW_SEL
+ pixel_8698/NB1 pixel_8698/VBIAS pixel_8698/NB2 pixel_8698/AMP_IN pixel_8698/SF_IB
+ pixel_8698/PIX_OUT pixel_8698/CSA_VREF pixel
Xpixel_7953 pixel_7953/gring pixel_7953/VDD pixel_7953/GND pixel_7953/VREF pixel_7953/ROW_SEL
+ pixel_7953/NB1 pixel_7953/VBIAS pixel_7953/NB2 pixel_7953/AMP_IN pixel_7953/SF_IB
+ pixel_7953/PIX_OUT pixel_7953/CSA_VREF pixel
Xpixel_7964 pixel_7964/gring pixel_7964/VDD pixel_7964/GND pixel_7964/VREF pixel_7964/ROW_SEL
+ pixel_7964/NB1 pixel_7964/VBIAS pixel_7964/NB2 pixel_7964/AMP_IN pixel_7964/SF_IB
+ pixel_7964/PIX_OUT pixel_7964/CSA_VREF pixel
Xpixel_7975 pixel_7975/gring pixel_7975/VDD pixel_7975/GND pixel_7975/VREF pixel_7975/ROW_SEL
+ pixel_7975/NB1 pixel_7975/VBIAS pixel_7975/NB2 pixel_7975/AMP_IN pixel_7975/SF_IB
+ pixel_7975/PIX_OUT pixel_7975/CSA_VREF pixel
Xpixel_7986 pixel_7986/gring pixel_7986/VDD pixel_7986/GND pixel_7986/VREF pixel_7986/ROW_SEL
+ pixel_7986/NB1 pixel_7986/VBIAS pixel_7986/NB2 pixel_7986/AMP_IN pixel_7986/SF_IB
+ pixel_7986/PIX_OUT pixel_7986/CSA_VREF pixel
Xpixel_7997 pixel_7997/gring pixel_7997/VDD pixel_7997/GND pixel_7997/VREF pixel_7997/ROW_SEL
+ pixel_7997/NB1 pixel_7997/VBIAS pixel_7997/NB2 pixel_7997/AMP_IN pixel_7997/SF_IB
+ pixel_7997/PIX_OUT pixel_7997/CSA_VREF pixel
Xpixel_2271 pixel_2271/gring pixel_2271/VDD pixel_2271/GND pixel_2271/VREF pixel_2271/ROW_SEL
+ pixel_2271/NB1 pixel_2271/VBIAS pixel_2271/NB2 pixel_2271/AMP_IN pixel_2271/SF_IB
+ pixel_2271/PIX_OUT pixel_2271/CSA_VREF pixel
Xpixel_2260 pixel_2260/gring pixel_2260/VDD pixel_2260/GND pixel_2260/VREF pixel_2260/ROW_SEL
+ pixel_2260/NB1 pixel_2260/VBIAS pixel_2260/NB2 pixel_2260/AMP_IN pixel_2260/SF_IB
+ pixel_2260/PIX_OUT pixel_2260/CSA_VREF pixel
Xpixel_1570 pixel_1570/gring pixel_1570/VDD pixel_1570/GND pixel_1570/VREF pixel_1570/ROW_SEL
+ pixel_1570/NB1 pixel_1570/VBIAS pixel_1570/NB2 pixel_1570/AMP_IN pixel_1570/SF_IB
+ pixel_1570/PIX_OUT pixel_1570/CSA_VREF pixel
Xpixel_2293 pixel_2293/gring pixel_2293/VDD pixel_2293/GND pixel_2293/VREF pixel_2293/ROW_SEL
+ pixel_2293/NB1 pixel_2293/VBIAS pixel_2293/NB2 pixel_2293/AMP_IN pixel_2293/SF_IB
+ pixel_2293/PIX_OUT pixel_2293/CSA_VREF pixel
Xpixel_2282 pixel_2282/gring pixel_2282/VDD pixel_2282/GND pixel_2282/VREF pixel_2282/ROW_SEL
+ pixel_2282/NB1 pixel_2282/VBIAS pixel_2282/NB2 pixel_2282/AMP_IN pixel_2282/SF_IB
+ pixel_2282/PIX_OUT pixel_2282/CSA_VREF pixel
Xpixel_1592 pixel_1592/gring pixel_1592/VDD pixel_1592/GND pixel_1592/VREF pixel_1592/ROW_SEL
+ pixel_1592/NB1 pixel_1592/VBIAS pixel_1592/NB2 pixel_1592/AMP_IN pixel_1592/SF_IB
+ pixel_1592/PIX_OUT pixel_1592/CSA_VREF pixel
Xpixel_1581 pixel_1581/gring pixel_1581/VDD pixel_1581/GND pixel_1581/VREF pixel_1581/ROW_SEL
+ pixel_1581/NB1 pixel_1581/VBIAS pixel_1581/NB2 pixel_1581/AMP_IN pixel_1581/SF_IB
+ pixel_1581/PIX_OUT pixel_1581/CSA_VREF pixel
Xpixel_629 pixel_629/gring pixel_629/VDD pixel_629/GND pixel_629/VREF pixel_629/ROW_SEL
+ pixel_629/NB1 pixel_629/VBIAS pixel_629/NB2 pixel_629/AMP_IN pixel_629/SF_IB pixel_629/PIX_OUT
+ pixel_629/CSA_VREF pixel
Xpixel_618 pixel_618/gring pixel_618/VDD pixel_618/GND pixel_618/VREF pixel_618/ROW_SEL
+ pixel_618/NB1 pixel_618/VBIAS pixel_618/NB2 pixel_618/AMP_IN pixel_618/SF_IB pixel_618/PIX_OUT
+ pixel_618/CSA_VREF pixel
Xpixel_607 pixel_607/gring pixel_607/VDD pixel_607/GND pixel_607/VREF pixel_607/ROW_SEL
+ pixel_607/NB1 pixel_607/VBIAS pixel_607/NB2 pixel_607/AMP_IN pixel_607/SF_IB pixel_607/PIX_OUT
+ pixel_607/CSA_VREF pixel
Xpixel_7205 pixel_7205/gring pixel_7205/VDD pixel_7205/GND pixel_7205/VREF pixel_7205/ROW_SEL
+ pixel_7205/NB1 pixel_7205/VBIAS pixel_7205/NB2 pixel_7205/AMP_IN pixel_7205/SF_IB
+ pixel_7205/PIX_OUT pixel_7205/CSA_VREF pixel
Xpixel_7216 pixel_7216/gring pixel_7216/VDD pixel_7216/GND pixel_7216/VREF pixel_7216/ROW_SEL
+ pixel_7216/NB1 pixel_7216/VBIAS pixel_7216/NB2 pixel_7216/AMP_IN pixel_7216/SF_IB
+ pixel_7216/PIX_OUT pixel_7216/CSA_VREF pixel
Xpixel_7227 pixel_7227/gring pixel_7227/VDD pixel_7227/GND pixel_7227/VREF pixel_7227/ROW_SEL
+ pixel_7227/NB1 pixel_7227/VBIAS pixel_7227/NB2 pixel_7227/AMP_IN pixel_7227/SF_IB
+ pixel_7227/PIX_OUT pixel_7227/CSA_VREF pixel
Xpixel_7238 pixel_7238/gring pixel_7238/VDD pixel_7238/GND pixel_7238/VREF pixel_7238/ROW_SEL
+ pixel_7238/NB1 pixel_7238/VBIAS pixel_7238/NB2 pixel_7238/AMP_IN pixel_7238/SF_IB
+ pixel_7238/PIX_OUT pixel_7238/CSA_VREF pixel
Xpixel_7249 pixel_7249/gring pixel_7249/VDD pixel_7249/GND pixel_7249/VREF pixel_7249/ROW_SEL
+ pixel_7249/NB1 pixel_7249/VBIAS pixel_7249/NB2 pixel_7249/AMP_IN pixel_7249/SF_IB
+ pixel_7249/PIX_OUT pixel_7249/CSA_VREF pixel
Xpixel_6504 pixel_6504/gring pixel_6504/VDD pixel_6504/GND pixel_6504/VREF pixel_6504/ROW_SEL
+ pixel_6504/NB1 pixel_6504/VBIAS pixel_6504/NB2 pixel_6504/AMP_IN pixel_6504/SF_IB
+ pixel_6504/PIX_OUT pixel_6504/CSA_VREF pixel
Xpixel_6515 pixel_6515/gring pixel_6515/VDD pixel_6515/GND pixel_6515/VREF pixel_6515/ROW_SEL
+ pixel_6515/NB1 pixel_6515/VBIAS pixel_6515/NB2 pixel_6515/AMP_IN pixel_6515/SF_IB
+ pixel_6515/PIX_OUT pixel_6515/CSA_VREF pixel
Xpixel_6526 pixel_6526/gring pixel_6526/VDD pixel_6526/GND pixel_6526/VREF pixel_6526/ROW_SEL
+ pixel_6526/NB1 pixel_6526/VBIAS pixel_6526/NB2 pixel_6526/AMP_IN pixel_6526/SF_IB
+ pixel_6526/PIX_OUT pixel_6526/CSA_VREF pixel
Xpixel_6537 pixel_6537/gring pixel_6537/VDD pixel_6537/GND pixel_6537/VREF pixel_6537/ROW_SEL
+ pixel_6537/NB1 pixel_6537/VBIAS pixel_6537/NB2 pixel_6537/AMP_IN pixel_6537/SF_IB
+ pixel_6537/PIX_OUT pixel_6537/CSA_VREF pixel
Xpixel_6548 pixel_6548/gring pixel_6548/VDD pixel_6548/GND pixel_6548/VREF pixel_6548/ROW_SEL
+ pixel_6548/NB1 pixel_6548/VBIAS pixel_6548/NB2 pixel_6548/AMP_IN pixel_6548/SF_IB
+ pixel_6548/PIX_OUT pixel_6548/CSA_VREF pixel
Xpixel_6559 pixel_6559/gring pixel_6559/VDD pixel_6559/GND pixel_6559/VREF pixel_6559/ROW_SEL
+ pixel_6559/NB1 pixel_6559/VBIAS pixel_6559/NB2 pixel_6559/AMP_IN pixel_6559/SF_IB
+ pixel_6559/PIX_OUT pixel_6559/CSA_VREF pixel
Xpixel_5803 pixel_5803/gring pixel_5803/VDD pixel_5803/GND pixel_5803/VREF pixel_5803/ROW_SEL
+ pixel_5803/NB1 pixel_5803/VBIAS pixel_5803/NB2 pixel_5803/AMP_IN pixel_5803/SF_IB
+ pixel_5803/PIX_OUT pixel_5803/CSA_VREF pixel
Xpixel_5814 pixel_5814/gring pixel_5814/VDD pixel_5814/GND pixel_5814/VREF pixel_5814/ROW_SEL
+ pixel_5814/NB1 pixel_5814/VBIAS pixel_5814/NB2 pixel_5814/AMP_IN pixel_5814/SF_IB
+ pixel_5814/PIX_OUT pixel_5814/CSA_VREF pixel
Xpixel_5825 pixel_5825/gring pixel_5825/VDD pixel_5825/GND pixel_5825/VREF pixel_5825/ROW_SEL
+ pixel_5825/NB1 pixel_5825/VBIAS pixel_5825/NB2 pixel_5825/AMP_IN pixel_5825/SF_IB
+ pixel_5825/PIX_OUT pixel_5825/CSA_VREF pixel
Xpixel_5836 pixel_5836/gring pixel_5836/VDD pixel_5836/GND pixel_5836/VREF pixel_5836/ROW_SEL
+ pixel_5836/NB1 pixel_5836/VBIAS pixel_5836/NB2 pixel_5836/AMP_IN pixel_5836/SF_IB
+ pixel_5836/PIX_OUT pixel_5836/CSA_VREF pixel
Xpixel_5847 pixel_5847/gring pixel_5847/VDD pixel_5847/GND pixel_5847/VREF pixel_5847/ROW_SEL
+ pixel_5847/NB1 pixel_5847/VBIAS pixel_5847/NB2 pixel_5847/AMP_IN pixel_5847/SF_IB
+ pixel_5847/PIX_OUT pixel_5847/CSA_VREF pixel
Xpixel_5858 pixel_5858/gring pixel_5858/VDD pixel_5858/GND pixel_5858/VREF pixel_5858/ROW_SEL
+ pixel_5858/NB1 pixel_5858/VBIAS pixel_5858/NB2 pixel_5858/AMP_IN pixel_5858/SF_IB
+ pixel_5858/PIX_OUT pixel_5858/CSA_VREF pixel
Xpixel_5869 pixel_5869/gring pixel_5869/VDD pixel_5869/GND pixel_5869/VREF pixel_5869/ROW_SEL
+ pixel_5869/NB1 pixel_5869/VBIAS pixel_5869/NB2 pixel_5869/AMP_IN pixel_5869/SF_IB
+ pixel_5869/PIX_OUT pixel_5869/CSA_VREF pixel
Xpixel_9130 pixel_9130/gring pixel_9130/VDD pixel_9130/GND pixel_9130/VREF pixel_9130/ROW_SEL
+ pixel_9130/NB1 pixel_9130/VBIAS pixel_9130/NB2 pixel_9130/AMP_IN pixel_9130/SF_IB
+ pixel_9130/PIX_OUT pixel_9130/CSA_VREF pixel
Xpixel_9163 pixel_9163/gring pixel_9163/VDD pixel_9163/GND pixel_9163/VREF pixel_9163/ROW_SEL
+ pixel_9163/NB1 pixel_9163/VBIAS pixel_9163/NB2 pixel_9163/AMP_IN pixel_9163/SF_IB
+ pixel_9163/PIX_OUT pixel_9163/CSA_VREF pixel
Xpixel_9152 pixel_9152/gring pixel_9152/VDD pixel_9152/GND pixel_9152/VREF pixel_9152/ROW_SEL
+ pixel_9152/NB1 pixel_9152/VBIAS pixel_9152/NB2 pixel_9152/AMP_IN pixel_9152/SF_IB
+ pixel_9152/PIX_OUT pixel_9152/CSA_VREF pixel
Xpixel_9141 pixel_9141/gring pixel_9141/VDD pixel_9141/GND pixel_9141/VREF pixel_9141/ROW_SEL
+ pixel_9141/NB1 pixel_9141/VBIAS pixel_9141/NB2 pixel_9141/AMP_IN pixel_9141/SF_IB
+ pixel_9141/PIX_OUT pixel_9141/CSA_VREF pixel
Xpixel_9196 pixel_9196/gring pixel_9196/VDD pixel_9196/GND pixel_9196/VREF pixel_9196/ROW_SEL
+ pixel_9196/NB1 pixel_9196/VBIAS pixel_9196/NB2 pixel_9196/AMP_IN pixel_9196/SF_IB
+ pixel_9196/PIX_OUT pixel_9196/CSA_VREF pixel
Xpixel_9185 pixel_9185/gring pixel_9185/VDD pixel_9185/GND pixel_9185/VREF pixel_9185/ROW_SEL
+ pixel_9185/NB1 pixel_9185/VBIAS pixel_9185/NB2 pixel_9185/AMP_IN pixel_9185/SF_IB
+ pixel_9185/PIX_OUT pixel_9185/CSA_VREF pixel
Xpixel_9174 pixel_9174/gring pixel_9174/VDD pixel_9174/GND pixel_9174/VREF pixel_9174/ROW_SEL
+ pixel_9174/NB1 pixel_9174/VBIAS pixel_9174/NB2 pixel_9174/AMP_IN pixel_9174/SF_IB
+ pixel_9174/PIX_OUT pixel_9174/CSA_VREF pixel
Xpixel_8440 pixel_8440/gring pixel_8440/VDD pixel_8440/GND pixel_8440/VREF pixel_8440/ROW_SEL
+ pixel_8440/NB1 pixel_8440/VBIAS pixel_8440/NB2 pixel_8440/AMP_IN pixel_8440/SF_IB
+ pixel_8440/PIX_OUT pixel_8440/CSA_VREF pixel
Xpixel_8451 pixel_8451/gring pixel_8451/VDD pixel_8451/GND pixel_8451/VREF pixel_8451/ROW_SEL
+ pixel_8451/NB1 pixel_8451/VBIAS pixel_8451/NB2 pixel_8451/AMP_IN pixel_8451/SF_IB
+ pixel_8451/PIX_OUT pixel_8451/CSA_VREF pixel
Xpixel_8462 pixel_8462/gring pixel_8462/VDD pixel_8462/GND pixel_8462/VREF pixel_8462/ROW_SEL
+ pixel_8462/NB1 pixel_8462/VBIAS pixel_8462/NB2 pixel_8462/AMP_IN pixel_8462/SF_IB
+ pixel_8462/PIX_OUT pixel_8462/CSA_VREF pixel
Xpixel_8473 pixel_8473/gring pixel_8473/VDD pixel_8473/GND pixel_8473/VREF pixel_8473/ROW_SEL
+ pixel_8473/NB1 pixel_8473/VBIAS pixel_8473/NB2 pixel_8473/AMP_IN pixel_8473/SF_IB
+ pixel_8473/PIX_OUT pixel_8473/CSA_VREF pixel
Xpixel_8484 pixel_8484/gring pixel_8484/VDD pixel_8484/GND pixel_8484/VREF pixel_8484/ROW_SEL
+ pixel_8484/NB1 pixel_8484/VBIAS pixel_8484/NB2 pixel_8484/AMP_IN pixel_8484/SF_IB
+ pixel_8484/PIX_OUT pixel_8484/CSA_VREF pixel
Xpixel_8495 pixel_8495/gring pixel_8495/VDD pixel_8495/GND pixel_8495/VREF pixel_8495/ROW_SEL
+ pixel_8495/NB1 pixel_8495/VBIAS pixel_8495/NB2 pixel_8495/AMP_IN pixel_8495/SF_IB
+ pixel_8495/PIX_OUT pixel_8495/CSA_VREF pixel
Xpixel_7750 pixel_7750/gring pixel_7750/VDD pixel_7750/GND pixel_7750/VREF pixel_7750/ROW_SEL
+ pixel_7750/NB1 pixel_7750/VBIAS pixel_7750/NB2 pixel_7750/AMP_IN pixel_7750/SF_IB
+ pixel_7750/PIX_OUT pixel_7750/CSA_VREF pixel
Xpixel_7761 pixel_7761/gring pixel_7761/VDD pixel_7761/GND pixel_7761/VREF pixel_7761/ROW_SEL
+ pixel_7761/NB1 pixel_7761/VBIAS pixel_7761/NB2 pixel_7761/AMP_IN pixel_7761/SF_IB
+ pixel_7761/PIX_OUT pixel_7761/CSA_VREF pixel
Xpixel_7772 pixel_7772/gring pixel_7772/VDD pixel_7772/GND pixel_7772/VREF pixel_7772/ROW_SEL
+ pixel_7772/NB1 pixel_7772/VBIAS pixel_7772/NB2 pixel_7772/AMP_IN pixel_7772/SF_IB
+ pixel_7772/PIX_OUT pixel_7772/CSA_VREF pixel
Xpixel_7783 pixel_7783/gring pixel_7783/VDD pixel_7783/GND pixel_7783/VREF pixel_7783/ROW_SEL
+ pixel_7783/NB1 pixel_7783/VBIAS pixel_7783/NB2 pixel_7783/AMP_IN pixel_7783/SF_IB
+ pixel_7783/PIX_OUT pixel_7783/CSA_VREF pixel
Xpixel_7794 pixel_7794/gring pixel_7794/VDD pixel_7794/GND pixel_7794/VREF pixel_7794/ROW_SEL
+ pixel_7794/NB1 pixel_7794/VBIAS pixel_7794/NB2 pixel_7794/AMP_IN pixel_7794/SF_IB
+ pixel_7794/PIX_OUT pixel_7794/CSA_VREF pixel
Xpixel_2090 pixel_2090/gring pixel_2090/VDD pixel_2090/GND pixel_2090/VREF pixel_2090/ROW_SEL
+ pixel_2090/NB1 pixel_2090/VBIAS pixel_2090/NB2 pixel_2090/AMP_IN pixel_2090/SF_IB
+ pixel_2090/PIX_OUT pixel_2090/CSA_VREF pixel
Xpixel_404 pixel_404/gring pixel_404/VDD pixel_404/GND pixel_404/VREF pixel_404/ROW_SEL
+ pixel_404/NB1 pixel_404/VBIAS pixel_404/NB2 pixel_404/AMP_IN pixel_404/SF_IB pixel_404/PIX_OUT
+ pixel_404/CSA_VREF pixel
Xpixel_4409 pixel_4409/gring pixel_4409/VDD pixel_4409/GND pixel_4409/VREF pixel_4409/ROW_SEL
+ pixel_4409/NB1 pixel_4409/VBIAS pixel_4409/NB2 pixel_4409/AMP_IN pixel_4409/SF_IB
+ pixel_4409/PIX_OUT pixel_4409/CSA_VREF pixel
Xpixel_437 pixel_437/gring pixel_437/VDD pixel_437/GND pixel_437/VREF pixel_437/ROW_SEL
+ pixel_437/NB1 pixel_437/VBIAS pixel_437/NB2 pixel_437/AMP_IN pixel_437/SF_IB pixel_437/PIX_OUT
+ pixel_437/CSA_VREF pixel
Xpixel_426 pixel_426/gring pixel_426/VDD pixel_426/GND pixel_426/VREF pixel_426/ROW_SEL
+ pixel_426/NB1 pixel_426/VBIAS pixel_426/NB2 pixel_426/AMP_IN pixel_426/SF_IB pixel_426/PIX_OUT
+ pixel_426/CSA_VREF pixel
Xpixel_415 pixel_415/gring pixel_415/VDD pixel_415/GND pixel_415/VREF pixel_415/ROW_SEL
+ pixel_415/NB1 pixel_415/VBIAS pixel_415/NB2 pixel_415/AMP_IN pixel_415/SF_IB pixel_415/PIX_OUT
+ pixel_415/CSA_VREF pixel
Xpixel_459 pixel_459/gring pixel_459/VDD pixel_459/GND pixel_459/VREF pixel_459/ROW_SEL
+ pixel_459/NB1 pixel_459/VBIAS pixel_459/NB2 pixel_459/AMP_IN pixel_459/SF_IB pixel_459/PIX_OUT
+ pixel_459/CSA_VREF pixel
Xpixel_448 pixel_448/gring pixel_448/VDD pixel_448/GND pixel_448/VREF pixel_448/ROW_SEL
+ pixel_448/NB1 pixel_448/VBIAS pixel_448/NB2 pixel_448/AMP_IN pixel_448/SF_IB pixel_448/PIX_OUT
+ pixel_448/CSA_VREF pixel
Xpixel_3719 pixel_3719/gring pixel_3719/VDD pixel_3719/GND pixel_3719/VREF pixel_3719/ROW_SEL
+ pixel_3719/NB1 pixel_3719/VBIAS pixel_3719/NB2 pixel_3719/AMP_IN pixel_3719/SF_IB
+ pixel_3719/PIX_OUT pixel_3719/CSA_VREF pixel
Xpixel_3708 pixel_3708/gring pixel_3708/VDD pixel_3708/GND pixel_3708/VREF pixel_3708/ROW_SEL
+ pixel_3708/NB1 pixel_3708/VBIAS pixel_3708/NB2 pixel_3708/AMP_IN pixel_3708/SF_IB
+ pixel_3708/PIX_OUT pixel_3708/CSA_VREF pixel
Xpixel_7002 pixel_7002/gring pixel_7002/VDD pixel_7002/GND pixel_7002/VREF pixel_7002/ROW_SEL
+ pixel_7002/NB1 pixel_7002/VBIAS pixel_7002/NB2 pixel_7002/AMP_IN pixel_7002/SF_IB
+ pixel_7002/PIX_OUT pixel_7002/CSA_VREF pixel
Xpixel_7013 pixel_7013/gring pixel_7013/VDD pixel_7013/GND pixel_7013/VREF pixel_7013/ROW_SEL
+ pixel_7013/NB1 pixel_7013/VBIAS pixel_7013/NB2 pixel_7013/AMP_IN pixel_7013/SF_IB
+ pixel_7013/PIX_OUT pixel_7013/CSA_VREF pixel
Xpixel_7024 pixel_7024/gring pixel_7024/VDD pixel_7024/GND pixel_7024/VREF pixel_7024/ROW_SEL
+ pixel_7024/NB1 pixel_7024/VBIAS pixel_7024/NB2 pixel_7024/AMP_IN pixel_7024/SF_IB
+ pixel_7024/PIX_OUT pixel_7024/CSA_VREF pixel
Xpixel_7035 pixel_7035/gring pixel_7035/VDD pixel_7035/GND pixel_7035/VREF pixel_7035/ROW_SEL
+ pixel_7035/NB1 pixel_7035/VBIAS pixel_7035/NB2 pixel_7035/AMP_IN pixel_7035/SF_IB
+ pixel_7035/PIX_OUT pixel_7035/CSA_VREF pixel
Xpixel_7046 pixel_7046/gring pixel_7046/VDD pixel_7046/GND pixel_7046/VREF pixel_7046/ROW_SEL
+ pixel_7046/NB1 pixel_7046/VBIAS pixel_7046/NB2 pixel_7046/AMP_IN pixel_7046/SF_IB
+ pixel_7046/PIX_OUT pixel_7046/CSA_VREF pixel
Xpixel_6301 pixel_6301/gring pixel_6301/VDD pixel_6301/GND pixel_6301/VREF pixel_6301/ROW_SEL
+ pixel_6301/NB1 pixel_6301/VBIAS pixel_6301/NB2 pixel_6301/AMP_IN pixel_6301/SF_IB
+ pixel_6301/PIX_OUT pixel_6301/CSA_VREF pixel
Xpixel_7057 pixel_7057/gring pixel_7057/VDD pixel_7057/GND pixel_7057/VREF pixel_7057/ROW_SEL
+ pixel_7057/NB1 pixel_7057/VBIAS pixel_7057/NB2 pixel_7057/AMP_IN pixel_7057/SF_IB
+ pixel_7057/PIX_OUT pixel_7057/CSA_VREF pixel
Xpixel_7068 pixel_7068/gring pixel_7068/VDD pixel_7068/GND pixel_7068/VREF pixel_7068/ROW_SEL
+ pixel_7068/NB1 pixel_7068/VBIAS pixel_7068/NB2 pixel_7068/AMP_IN pixel_7068/SF_IB
+ pixel_7068/PIX_OUT pixel_7068/CSA_VREF pixel
Xpixel_7079 pixel_7079/gring pixel_7079/VDD pixel_7079/GND pixel_7079/VREF pixel_7079/ROW_SEL
+ pixel_7079/NB1 pixel_7079/VBIAS pixel_7079/NB2 pixel_7079/AMP_IN pixel_7079/SF_IB
+ pixel_7079/PIX_OUT pixel_7079/CSA_VREF pixel
Xpixel_6312 pixel_6312/gring pixel_6312/VDD pixel_6312/GND pixel_6312/VREF pixel_6312/ROW_SEL
+ pixel_6312/NB1 pixel_6312/VBIAS pixel_6312/NB2 pixel_6312/AMP_IN pixel_6312/SF_IB
+ pixel_6312/PIX_OUT pixel_6312/CSA_VREF pixel
Xpixel_6323 pixel_6323/gring pixel_6323/VDD pixel_6323/GND pixel_6323/VREF pixel_6323/ROW_SEL
+ pixel_6323/NB1 pixel_6323/VBIAS pixel_6323/NB2 pixel_6323/AMP_IN pixel_6323/SF_IB
+ pixel_6323/PIX_OUT pixel_6323/CSA_VREF pixel
Xpixel_6334 pixel_6334/gring pixel_6334/VDD pixel_6334/GND pixel_6334/VREF pixel_6334/ROW_SEL
+ pixel_6334/NB1 pixel_6334/VBIAS pixel_6334/NB2 pixel_6334/AMP_IN pixel_6334/SF_IB
+ pixel_6334/PIX_OUT pixel_6334/CSA_VREF pixel
Xpixel_6345 pixel_6345/gring pixel_6345/VDD pixel_6345/GND pixel_6345/VREF pixel_6345/ROW_SEL
+ pixel_6345/NB1 pixel_6345/VBIAS pixel_6345/NB2 pixel_6345/AMP_IN pixel_6345/SF_IB
+ pixel_6345/PIX_OUT pixel_6345/CSA_VREF pixel
Xpixel_5600 pixel_5600/gring pixel_5600/VDD pixel_5600/GND pixel_5600/VREF pixel_5600/ROW_SEL
+ pixel_5600/NB1 pixel_5600/VBIAS pixel_5600/NB2 pixel_5600/AMP_IN pixel_5600/SF_IB
+ pixel_5600/PIX_OUT pixel_5600/CSA_VREF pixel
Xpixel_6356 pixel_6356/gring pixel_6356/VDD pixel_6356/GND pixel_6356/VREF pixel_6356/ROW_SEL
+ pixel_6356/NB1 pixel_6356/VBIAS pixel_6356/NB2 pixel_6356/AMP_IN pixel_6356/SF_IB
+ pixel_6356/PIX_OUT pixel_6356/CSA_VREF pixel
Xpixel_6367 pixel_6367/gring pixel_6367/VDD pixel_6367/GND pixel_6367/VREF pixel_6367/ROW_SEL
+ pixel_6367/NB1 pixel_6367/VBIAS pixel_6367/NB2 pixel_6367/AMP_IN pixel_6367/SF_IB
+ pixel_6367/PIX_OUT pixel_6367/CSA_VREF pixel
Xpixel_6378 pixel_6378/gring pixel_6378/VDD pixel_6378/GND pixel_6378/VREF pixel_6378/ROW_SEL
+ pixel_6378/NB1 pixel_6378/VBIAS pixel_6378/NB2 pixel_6378/AMP_IN pixel_6378/SF_IB
+ pixel_6378/PIX_OUT pixel_6378/CSA_VREF pixel
Xpixel_5611 pixel_5611/gring pixel_5611/VDD pixel_5611/GND pixel_5611/VREF pixel_5611/ROW_SEL
+ pixel_5611/NB1 pixel_5611/VBIAS pixel_5611/NB2 pixel_5611/AMP_IN pixel_5611/SF_IB
+ pixel_5611/PIX_OUT pixel_5611/CSA_VREF pixel
Xpixel_5622 pixel_5622/gring pixel_5622/VDD pixel_5622/GND pixel_5622/VREF pixel_5622/ROW_SEL
+ pixel_5622/NB1 pixel_5622/VBIAS pixel_5622/NB2 pixel_5622/AMP_IN pixel_5622/SF_IB
+ pixel_5622/PIX_OUT pixel_5622/CSA_VREF pixel
Xpixel_5633 pixel_5633/gring pixel_5633/VDD pixel_5633/GND pixel_5633/VREF pixel_5633/ROW_SEL
+ pixel_5633/NB1 pixel_5633/VBIAS pixel_5633/NB2 pixel_5633/AMP_IN pixel_5633/SF_IB
+ pixel_5633/PIX_OUT pixel_5633/CSA_VREF pixel
Xpixel_6389 pixel_6389/gring pixel_6389/VDD pixel_6389/GND pixel_6389/VREF pixel_6389/ROW_SEL
+ pixel_6389/NB1 pixel_6389/VBIAS pixel_6389/NB2 pixel_6389/AMP_IN pixel_6389/SF_IB
+ pixel_6389/PIX_OUT pixel_6389/CSA_VREF pixel
Xpixel_5644 pixel_5644/gring pixel_5644/VDD pixel_5644/GND pixel_5644/VREF pixel_5644/ROW_SEL
+ pixel_5644/NB1 pixel_5644/VBIAS pixel_5644/NB2 pixel_5644/AMP_IN pixel_5644/SF_IB
+ pixel_5644/PIX_OUT pixel_5644/CSA_VREF pixel
Xpixel_5655 pixel_5655/gring pixel_5655/VDD pixel_5655/GND pixel_5655/VREF pixel_5655/ROW_SEL
+ pixel_5655/NB1 pixel_5655/VBIAS pixel_5655/NB2 pixel_5655/AMP_IN pixel_5655/SF_IB
+ pixel_5655/PIX_OUT pixel_5655/CSA_VREF pixel
Xpixel_5666 pixel_5666/gring pixel_5666/VDD pixel_5666/GND pixel_5666/VREF pixel_5666/ROW_SEL
+ pixel_5666/NB1 pixel_5666/VBIAS pixel_5666/NB2 pixel_5666/AMP_IN pixel_5666/SF_IB
+ pixel_5666/PIX_OUT pixel_5666/CSA_VREF pixel
Xpixel_4910 pixel_4910/gring pixel_4910/VDD pixel_4910/GND pixel_4910/VREF pixel_4910/ROW_SEL
+ pixel_4910/NB1 pixel_4910/VBIAS pixel_4910/NB2 pixel_4910/AMP_IN pixel_4910/SF_IB
+ pixel_4910/PIX_OUT pixel_4910/CSA_VREF pixel
Xpixel_4921 pixel_4921/gring pixel_4921/VDD pixel_4921/GND pixel_4921/VREF pixel_4921/ROW_SEL
+ pixel_4921/NB1 pixel_4921/VBIAS pixel_4921/NB2 pixel_4921/AMP_IN pixel_4921/SF_IB
+ pixel_4921/PIX_OUT pixel_4921/CSA_VREF pixel
Xpixel_960 pixel_960/gring pixel_960/VDD pixel_960/GND pixel_960/VREF pixel_960/ROW_SEL
+ pixel_960/NB1 pixel_960/VBIAS pixel_960/NB2 pixel_960/AMP_IN pixel_960/SF_IB pixel_960/PIX_OUT
+ pixel_960/CSA_VREF pixel
Xpixel_5677 pixel_5677/gring pixel_5677/VDD pixel_5677/GND pixel_5677/VREF pixel_5677/ROW_SEL
+ pixel_5677/NB1 pixel_5677/VBIAS pixel_5677/NB2 pixel_5677/AMP_IN pixel_5677/SF_IB
+ pixel_5677/PIX_OUT pixel_5677/CSA_VREF pixel
Xpixel_5688 pixel_5688/gring pixel_5688/VDD pixel_5688/GND pixel_5688/VREF pixel_5688/ROW_SEL
+ pixel_5688/NB1 pixel_5688/VBIAS pixel_5688/NB2 pixel_5688/AMP_IN pixel_5688/SF_IB
+ pixel_5688/PIX_OUT pixel_5688/CSA_VREF pixel
Xpixel_5699 pixel_5699/gring pixel_5699/VDD pixel_5699/GND pixel_5699/VREF pixel_5699/ROW_SEL
+ pixel_5699/NB1 pixel_5699/VBIAS pixel_5699/NB2 pixel_5699/AMP_IN pixel_5699/SF_IB
+ pixel_5699/PIX_OUT pixel_5699/CSA_VREF pixel
Xpixel_4932 pixel_4932/gring pixel_4932/VDD pixel_4932/GND pixel_4932/VREF pixel_4932/ROW_SEL
+ pixel_4932/NB1 pixel_4932/VBIAS pixel_4932/NB2 pixel_4932/AMP_IN pixel_4932/SF_IB
+ pixel_4932/PIX_OUT pixel_4932/CSA_VREF pixel
Xpixel_4943 pixel_4943/gring pixel_4943/VDD pixel_4943/GND pixel_4943/VREF pixel_4943/ROW_SEL
+ pixel_4943/NB1 pixel_4943/VBIAS pixel_4943/NB2 pixel_4943/AMP_IN pixel_4943/SF_IB
+ pixel_4943/PIX_OUT pixel_4943/CSA_VREF pixel
Xpixel_4954 pixel_4954/gring pixel_4954/VDD pixel_4954/GND pixel_4954/VREF pixel_4954/ROW_SEL
+ pixel_4954/NB1 pixel_4954/VBIAS pixel_4954/NB2 pixel_4954/AMP_IN pixel_4954/SF_IB
+ pixel_4954/PIX_OUT pixel_4954/CSA_VREF pixel
Xpixel_4965 pixel_4965/gring pixel_4965/VDD pixel_4965/GND pixel_4965/VREF pixel_4965/ROW_SEL
+ pixel_4965/NB1 pixel_4965/VBIAS pixel_4965/NB2 pixel_4965/AMP_IN pixel_4965/SF_IB
+ pixel_4965/PIX_OUT pixel_4965/CSA_VREF pixel
Xpixel_993 pixel_993/gring pixel_993/VDD pixel_993/GND pixel_993/VREF pixel_993/ROW_SEL
+ pixel_993/NB1 pixel_993/VBIAS pixel_993/NB2 pixel_993/AMP_IN pixel_993/SF_IB pixel_993/PIX_OUT
+ pixel_993/CSA_VREF pixel
Xpixel_982 pixel_982/gring pixel_982/VDD pixel_982/GND pixel_982/VREF pixel_982/ROW_SEL
+ pixel_982/NB1 pixel_982/VBIAS pixel_982/NB2 pixel_982/AMP_IN pixel_982/SF_IB pixel_982/PIX_OUT
+ pixel_982/CSA_VREF pixel
Xpixel_971 pixel_971/gring pixel_971/VDD pixel_971/GND pixel_971/VREF pixel_971/ROW_SEL
+ pixel_971/NB1 pixel_971/VBIAS pixel_971/NB2 pixel_971/AMP_IN pixel_971/SF_IB pixel_971/PIX_OUT
+ pixel_971/CSA_VREF pixel
Xpixel_4976 pixel_4976/gring pixel_4976/VDD pixel_4976/GND pixel_4976/VREF pixel_4976/ROW_SEL
+ pixel_4976/NB1 pixel_4976/VBIAS pixel_4976/NB2 pixel_4976/AMP_IN pixel_4976/SF_IB
+ pixel_4976/PIX_OUT pixel_4976/CSA_VREF pixel
Xpixel_4987 pixel_4987/gring pixel_4987/VDD pixel_4987/GND pixel_4987/VREF pixel_4987/ROW_SEL
+ pixel_4987/NB1 pixel_4987/VBIAS pixel_4987/NB2 pixel_4987/AMP_IN pixel_4987/SF_IB
+ pixel_4987/PIX_OUT pixel_4987/CSA_VREF pixel
Xpixel_4998 pixel_4998/gring pixel_4998/VDD pixel_4998/GND pixel_4998/VREF pixel_4998/ROW_SEL
+ pixel_4998/NB1 pixel_4998/VBIAS pixel_4998/NB2 pixel_4998/AMP_IN pixel_4998/SF_IB
+ pixel_4998/PIX_OUT pixel_4998/CSA_VREF pixel
Xpixel_8270 pixel_8270/gring pixel_8270/VDD pixel_8270/GND pixel_8270/VREF pixel_8270/ROW_SEL
+ pixel_8270/NB1 pixel_8270/VBIAS pixel_8270/NB2 pixel_8270/AMP_IN pixel_8270/SF_IB
+ pixel_8270/PIX_OUT pixel_8270/CSA_VREF pixel
Xpixel_8281 pixel_8281/gring pixel_8281/VDD pixel_8281/GND pixel_8281/VREF pixel_8281/ROW_SEL
+ pixel_8281/NB1 pixel_8281/VBIAS pixel_8281/NB2 pixel_8281/AMP_IN pixel_8281/SF_IB
+ pixel_8281/PIX_OUT pixel_8281/CSA_VREF pixel
Xpixel_8292 pixel_8292/gring pixel_8292/VDD pixel_8292/GND pixel_8292/VREF pixel_8292/ROW_SEL
+ pixel_8292/NB1 pixel_8292/VBIAS pixel_8292/NB2 pixel_8292/AMP_IN pixel_8292/SF_IB
+ pixel_8292/PIX_OUT pixel_8292/CSA_VREF pixel
Xpixel_7580 pixel_7580/gring pixel_7580/VDD pixel_7580/GND pixel_7580/VREF pixel_7580/ROW_SEL
+ pixel_7580/NB1 pixel_7580/VBIAS pixel_7580/NB2 pixel_7580/AMP_IN pixel_7580/SF_IB
+ pixel_7580/PIX_OUT pixel_7580/CSA_VREF pixel
Xpixel_7591 pixel_7591/gring pixel_7591/VDD pixel_7591/GND pixel_7591/VREF pixel_7591/ROW_SEL
+ pixel_7591/NB1 pixel_7591/VBIAS pixel_7591/NB2 pixel_7591/AMP_IN pixel_7591/SF_IB
+ pixel_7591/PIX_OUT pixel_7591/CSA_VREF pixel
Xpixel_6890 pixel_6890/gring pixel_6890/VDD pixel_6890/GND pixel_6890/VREF pixel_6890/ROW_SEL
+ pixel_6890/NB1 pixel_6890/VBIAS pixel_6890/NB2 pixel_6890/AMP_IN pixel_6890/SF_IB
+ pixel_6890/PIX_OUT pixel_6890/CSA_VREF pixel
Xpixel_212 pixel_212/gring pixel_212/VDD pixel_212/GND pixel_212/VREF pixel_212/ROW_SEL
+ pixel_212/NB1 pixel_212/VBIAS pixel_212/NB2 pixel_212/AMP_IN pixel_212/SF_IB pixel_212/PIX_OUT
+ pixel_212/CSA_VREF pixel
Xpixel_201 pixel_201/gring pixel_201/VDD pixel_201/GND pixel_201/VREF pixel_201/ROW_SEL
+ pixel_201/NB1 pixel_201/VBIAS pixel_201/NB2 pixel_201/AMP_IN pixel_201/SF_IB pixel_201/PIX_OUT
+ pixel_201/CSA_VREF pixel
Xpixel_4206 pixel_4206/gring pixel_4206/VDD pixel_4206/GND pixel_4206/VREF pixel_4206/ROW_SEL
+ pixel_4206/NB1 pixel_4206/VBIAS pixel_4206/NB2 pixel_4206/AMP_IN pixel_4206/SF_IB
+ pixel_4206/PIX_OUT pixel_4206/CSA_VREF pixel
Xpixel_4217 pixel_4217/gring pixel_4217/VDD pixel_4217/GND pixel_4217/VREF pixel_4217/ROW_SEL
+ pixel_4217/NB1 pixel_4217/VBIAS pixel_4217/NB2 pixel_4217/AMP_IN pixel_4217/SF_IB
+ pixel_4217/PIX_OUT pixel_4217/CSA_VREF pixel
Xpixel_256 pixel_256/gring pixel_256/VDD pixel_256/GND pixel_256/VREF pixel_256/ROW_SEL
+ pixel_256/NB1 pixel_256/VBIAS pixel_256/NB2 pixel_256/AMP_IN pixel_256/SF_IB pixel_256/PIX_OUT
+ pixel_256/CSA_VREF pixel
Xpixel_245 pixel_245/gring pixel_245/VDD pixel_245/GND pixel_245/VREF pixel_245/ROW_SEL
+ pixel_245/NB1 pixel_245/VBIAS pixel_245/NB2 pixel_245/AMP_IN pixel_245/SF_IB pixel_245/PIX_OUT
+ pixel_245/CSA_VREF pixel
Xpixel_234 pixel_234/gring pixel_234/VDD pixel_234/GND pixel_234/VREF pixel_234/ROW_SEL
+ pixel_234/NB1 pixel_234/VBIAS pixel_234/NB2 pixel_234/AMP_IN pixel_234/SF_IB pixel_234/PIX_OUT
+ pixel_234/CSA_VREF pixel
Xpixel_223 pixel_223/gring pixel_223/VDD pixel_223/GND pixel_223/VREF pixel_223/ROW_SEL
+ pixel_223/NB1 pixel_223/VBIAS pixel_223/NB2 pixel_223/AMP_IN pixel_223/SF_IB pixel_223/PIX_OUT
+ pixel_223/CSA_VREF pixel
Xpixel_3516 pixel_3516/gring pixel_3516/VDD pixel_3516/GND pixel_3516/VREF pixel_3516/ROW_SEL
+ pixel_3516/NB1 pixel_3516/VBIAS pixel_3516/NB2 pixel_3516/AMP_IN pixel_3516/SF_IB
+ pixel_3516/PIX_OUT pixel_3516/CSA_VREF pixel
Xpixel_3505 pixel_3505/gring pixel_3505/VDD pixel_3505/GND pixel_3505/VREF pixel_3505/ROW_SEL
+ pixel_3505/NB1 pixel_3505/VBIAS pixel_3505/NB2 pixel_3505/AMP_IN pixel_3505/SF_IB
+ pixel_3505/PIX_OUT pixel_3505/CSA_VREF pixel
Xpixel_4228 pixel_4228/gring pixel_4228/VDD pixel_4228/GND pixel_4228/VREF pixel_4228/ROW_SEL
+ pixel_4228/NB1 pixel_4228/VBIAS pixel_4228/NB2 pixel_4228/AMP_IN pixel_4228/SF_IB
+ pixel_4228/PIX_OUT pixel_4228/CSA_VREF pixel
Xpixel_4239 pixel_4239/gring pixel_4239/VDD pixel_4239/GND pixel_4239/VREF pixel_4239/ROW_SEL
+ pixel_4239/NB1 pixel_4239/VBIAS pixel_4239/NB2 pixel_4239/AMP_IN pixel_4239/SF_IB
+ pixel_4239/PIX_OUT pixel_4239/CSA_VREF pixel
Xpixel_289 pixel_289/gring pixel_289/VDD pixel_289/GND pixel_289/VREF pixel_289/ROW_SEL
+ pixel_289/NB1 pixel_289/VBIAS pixel_289/NB2 pixel_289/AMP_IN pixel_289/SF_IB pixel_289/PIX_OUT
+ pixel_289/CSA_VREF pixel
Xpixel_278 pixel_278/gring pixel_278/VDD pixel_278/GND pixel_278/VREF pixel_278/ROW_SEL
+ pixel_278/NB1 pixel_278/VBIAS pixel_278/NB2 pixel_278/AMP_IN pixel_278/SF_IB pixel_278/PIX_OUT
+ pixel_278/CSA_VREF pixel
Xpixel_267 pixel_267/gring pixel_267/VDD pixel_267/GND pixel_267/VREF pixel_267/ROW_SEL
+ pixel_267/NB1 pixel_267/VBIAS pixel_267/NB2 pixel_267/AMP_IN pixel_267/SF_IB pixel_267/PIX_OUT
+ pixel_267/CSA_VREF pixel
Xpixel_2804 pixel_2804/gring pixel_2804/VDD pixel_2804/GND pixel_2804/VREF pixel_2804/ROW_SEL
+ pixel_2804/NB1 pixel_2804/VBIAS pixel_2804/NB2 pixel_2804/AMP_IN pixel_2804/SF_IB
+ pixel_2804/PIX_OUT pixel_2804/CSA_VREF pixel
Xpixel_3549 pixel_3549/gring pixel_3549/VDD pixel_3549/GND pixel_3549/VREF pixel_3549/ROW_SEL
+ pixel_3549/NB1 pixel_3549/VBIAS pixel_3549/NB2 pixel_3549/AMP_IN pixel_3549/SF_IB
+ pixel_3549/PIX_OUT pixel_3549/CSA_VREF pixel
Xpixel_3538 pixel_3538/gring pixel_3538/VDD pixel_3538/GND pixel_3538/VREF pixel_3538/ROW_SEL
+ pixel_3538/NB1 pixel_3538/VBIAS pixel_3538/NB2 pixel_3538/AMP_IN pixel_3538/SF_IB
+ pixel_3538/PIX_OUT pixel_3538/CSA_VREF pixel
Xpixel_3527 pixel_3527/gring pixel_3527/VDD pixel_3527/GND pixel_3527/VREF pixel_3527/ROW_SEL
+ pixel_3527/NB1 pixel_3527/VBIAS pixel_3527/NB2 pixel_3527/AMP_IN pixel_3527/SF_IB
+ pixel_3527/PIX_OUT pixel_3527/CSA_VREF pixel
Xpixel_2837 pixel_2837/gring pixel_2837/VDD pixel_2837/GND pixel_2837/VREF pixel_2837/ROW_SEL
+ pixel_2837/NB1 pixel_2837/VBIAS pixel_2837/NB2 pixel_2837/AMP_IN pixel_2837/SF_IB
+ pixel_2837/PIX_OUT pixel_2837/CSA_VREF pixel
Xpixel_2826 pixel_2826/gring pixel_2826/VDD pixel_2826/GND pixel_2826/VREF pixel_2826/ROW_SEL
+ pixel_2826/NB1 pixel_2826/VBIAS pixel_2826/NB2 pixel_2826/AMP_IN pixel_2826/SF_IB
+ pixel_2826/PIX_OUT pixel_2826/CSA_VREF pixel
Xpixel_2815 pixel_2815/gring pixel_2815/VDD pixel_2815/GND pixel_2815/VREF pixel_2815/ROW_SEL
+ pixel_2815/NB1 pixel_2815/VBIAS pixel_2815/NB2 pixel_2815/AMP_IN pixel_2815/SF_IB
+ pixel_2815/PIX_OUT pixel_2815/CSA_VREF pixel
Xpixel_2859 pixel_2859/gring pixel_2859/VDD pixel_2859/GND pixel_2859/VREF pixel_2859/ROW_SEL
+ pixel_2859/NB1 pixel_2859/VBIAS pixel_2859/NB2 pixel_2859/AMP_IN pixel_2859/SF_IB
+ pixel_2859/PIX_OUT pixel_2859/CSA_VREF pixel
Xpixel_2848 pixel_2848/gring pixel_2848/VDD pixel_2848/GND pixel_2848/VREF pixel_2848/ROW_SEL
+ pixel_2848/NB1 pixel_2848/VBIAS pixel_2848/NB2 pixel_2848/AMP_IN pixel_2848/SF_IB
+ pixel_2848/PIX_OUT pixel_2848/CSA_VREF pixel
Xpixel_6120 pixel_6120/gring pixel_6120/VDD pixel_6120/GND pixel_6120/VREF pixel_6120/ROW_SEL
+ pixel_6120/NB1 pixel_6120/VBIAS pixel_6120/NB2 pixel_6120/AMP_IN pixel_6120/SF_IB
+ pixel_6120/PIX_OUT pixel_6120/CSA_VREF pixel
Xpixel_6131 pixel_6131/gring pixel_6131/VDD pixel_6131/GND pixel_6131/VREF pixel_6131/ROW_SEL
+ pixel_6131/NB1 pixel_6131/VBIAS pixel_6131/NB2 pixel_6131/AMP_IN pixel_6131/SF_IB
+ pixel_6131/PIX_OUT pixel_6131/CSA_VREF pixel
Xpixel_6142 pixel_6142/gring pixel_6142/VDD pixel_6142/GND pixel_6142/VREF pixel_6142/ROW_SEL
+ pixel_6142/NB1 pixel_6142/VBIAS pixel_6142/NB2 pixel_6142/AMP_IN pixel_6142/SF_IB
+ pixel_6142/PIX_OUT pixel_6142/CSA_VREF pixel
Xpixel_6153 pixel_6153/gring pixel_6153/VDD pixel_6153/GND pixel_6153/VREF pixel_6153/ROW_SEL
+ pixel_6153/NB1 pixel_6153/VBIAS pixel_6153/NB2 pixel_6153/AMP_IN pixel_6153/SF_IB
+ pixel_6153/PIX_OUT pixel_6153/CSA_VREF pixel
Xpixel_6164 pixel_6164/gring pixel_6164/VDD pixel_6164/GND pixel_6164/VREF pixel_6164/ROW_SEL
+ pixel_6164/NB1 pixel_6164/VBIAS pixel_6164/NB2 pixel_6164/AMP_IN pixel_6164/SF_IB
+ pixel_6164/PIX_OUT pixel_6164/CSA_VREF pixel
Xpixel_6175 pixel_6175/gring pixel_6175/VDD pixel_6175/GND pixel_6175/VREF pixel_6175/ROW_SEL
+ pixel_6175/NB1 pixel_6175/VBIAS pixel_6175/NB2 pixel_6175/AMP_IN pixel_6175/SF_IB
+ pixel_6175/PIX_OUT pixel_6175/CSA_VREF pixel
Xpixel_6186 pixel_6186/gring pixel_6186/VDD pixel_6186/GND pixel_6186/VREF pixel_6186/ROW_SEL
+ pixel_6186/NB1 pixel_6186/VBIAS pixel_6186/NB2 pixel_6186/AMP_IN pixel_6186/SF_IB
+ pixel_6186/PIX_OUT pixel_6186/CSA_VREF pixel
Xpixel_5430 pixel_5430/gring pixel_5430/VDD pixel_5430/GND pixel_5430/VREF pixel_5430/ROW_SEL
+ pixel_5430/NB1 pixel_5430/VBIAS pixel_5430/NB2 pixel_5430/AMP_IN pixel_5430/SF_IB
+ pixel_5430/PIX_OUT pixel_5430/CSA_VREF pixel
Xpixel_5441 pixel_5441/gring pixel_5441/VDD pixel_5441/GND pixel_5441/VREF pixel_5441/ROW_SEL
+ pixel_5441/NB1 pixel_5441/VBIAS pixel_5441/NB2 pixel_5441/AMP_IN pixel_5441/SF_IB
+ pixel_5441/PIX_OUT pixel_5441/CSA_VREF pixel
Xpixel_6197 pixel_6197/gring pixel_6197/VDD pixel_6197/GND pixel_6197/VREF pixel_6197/ROW_SEL
+ pixel_6197/NB1 pixel_6197/VBIAS pixel_6197/NB2 pixel_6197/AMP_IN pixel_6197/SF_IB
+ pixel_6197/PIX_OUT pixel_6197/CSA_VREF pixel
Xpixel_5452 pixel_5452/gring pixel_5452/VDD pixel_5452/GND pixel_5452/VREF pixel_5452/ROW_SEL
+ pixel_5452/NB1 pixel_5452/VBIAS pixel_5452/NB2 pixel_5452/AMP_IN pixel_5452/SF_IB
+ pixel_5452/PIX_OUT pixel_5452/CSA_VREF pixel
Xpixel_5463 pixel_5463/gring pixel_5463/VDD pixel_5463/GND pixel_5463/VREF pixel_5463/ROW_SEL
+ pixel_5463/NB1 pixel_5463/VBIAS pixel_5463/NB2 pixel_5463/AMP_IN pixel_5463/SF_IB
+ pixel_5463/PIX_OUT pixel_5463/CSA_VREF pixel
Xpixel_5474 pixel_5474/gring pixel_5474/VDD pixel_5474/GND pixel_5474/VREF pixel_5474/ROW_SEL
+ pixel_5474/NB1 pixel_5474/VBIAS pixel_5474/NB2 pixel_5474/AMP_IN pixel_5474/SF_IB
+ pixel_5474/PIX_OUT pixel_5474/CSA_VREF pixel
Xpixel_4740 pixel_4740/gring pixel_4740/VDD pixel_4740/GND pixel_4740/VREF pixel_4740/ROW_SEL
+ pixel_4740/NB1 pixel_4740/VBIAS pixel_4740/NB2 pixel_4740/AMP_IN pixel_4740/SF_IB
+ pixel_4740/PIX_OUT pixel_4740/CSA_VREF pixel
Xpixel_5485 pixel_5485/gring pixel_5485/VDD pixel_5485/GND pixel_5485/VREF pixel_5485/ROW_SEL
+ pixel_5485/NB1 pixel_5485/VBIAS pixel_5485/NB2 pixel_5485/AMP_IN pixel_5485/SF_IB
+ pixel_5485/PIX_OUT pixel_5485/CSA_VREF pixel
Xpixel_5496 pixel_5496/gring pixel_5496/VDD pixel_5496/GND pixel_5496/VREF pixel_5496/ROW_SEL
+ pixel_5496/NB1 pixel_5496/VBIAS pixel_5496/NB2 pixel_5496/AMP_IN pixel_5496/SF_IB
+ pixel_5496/PIX_OUT pixel_5496/CSA_VREF pixel
Xpixel_4751 pixel_4751/gring pixel_4751/VDD pixel_4751/GND pixel_4751/VREF pixel_4751/ROW_SEL
+ pixel_4751/NB1 pixel_4751/VBIAS pixel_4751/NB2 pixel_4751/AMP_IN pixel_4751/SF_IB
+ pixel_4751/PIX_OUT pixel_4751/CSA_VREF pixel
Xpixel_4762 pixel_4762/gring pixel_4762/VDD pixel_4762/GND pixel_4762/VREF pixel_4762/ROW_SEL
+ pixel_4762/NB1 pixel_4762/VBIAS pixel_4762/NB2 pixel_4762/AMP_IN pixel_4762/SF_IB
+ pixel_4762/PIX_OUT pixel_4762/CSA_VREF pixel
Xpixel_4773 pixel_4773/gring pixel_4773/VDD pixel_4773/GND pixel_4773/VREF pixel_4773/ROW_SEL
+ pixel_4773/NB1 pixel_4773/VBIAS pixel_4773/NB2 pixel_4773/AMP_IN pixel_4773/SF_IB
+ pixel_4773/PIX_OUT pixel_4773/CSA_VREF pixel
Xpixel_790 pixel_790/gring pixel_790/VDD pixel_790/GND pixel_790/VREF pixel_790/ROW_SEL
+ pixel_790/NB1 pixel_790/VBIAS pixel_790/NB2 pixel_790/AMP_IN pixel_790/SF_IB pixel_790/PIX_OUT
+ pixel_790/CSA_VREF pixel
Xpixel_4784 pixel_4784/gring pixel_4784/VDD pixel_4784/GND pixel_4784/VREF pixel_4784/ROW_SEL
+ pixel_4784/NB1 pixel_4784/VBIAS pixel_4784/NB2 pixel_4784/AMP_IN pixel_4784/SF_IB
+ pixel_4784/PIX_OUT pixel_4784/CSA_VREF pixel
Xpixel_4795 pixel_4795/gring pixel_4795/VDD pixel_4795/GND pixel_4795/VREF pixel_4795/ROW_SEL
+ pixel_4795/NB1 pixel_4795/VBIAS pixel_4795/NB2 pixel_4795/AMP_IN pixel_4795/SF_IB
+ pixel_4795/PIX_OUT pixel_4795/CSA_VREF pixel
Xpixel_9707 pixel_9707/gring pixel_9707/VDD pixel_9707/GND pixel_9707/VREF pixel_9707/ROW_SEL
+ pixel_9707/NB1 pixel_9707/VBIAS pixel_9707/NB2 pixel_9707/AMP_IN pixel_9707/SF_IB
+ pixel_9707/PIX_OUT pixel_9707/CSA_VREF pixel
Xpixel_9718 pixel_9718/gring pixel_9718/VDD pixel_9718/GND pixel_9718/VREF pixel_9718/ROW_SEL
+ pixel_9718/NB1 pixel_9718/VBIAS pixel_9718/NB2 pixel_9718/AMP_IN pixel_9718/SF_IB
+ pixel_9718/PIX_OUT pixel_9718/CSA_VREF pixel
Xpixel_9729 pixel_9729/gring pixel_9729/VDD pixel_9729/GND pixel_9729/VREF pixel_9729/ROW_SEL
+ pixel_9729/NB1 pixel_9729/VBIAS pixel_9729/NB2 pixel_9729/AMP_IN pixel_9729/SF_IB
+ pixel_9729/PIX_OUT pixel_9729/CSA_VREF pixel
Xpixel_4003 pixel_4003/gring pixel_4003/VDD pixel_4003/GND pixel_4003/VREF pixel_4003/ROW_SEL
+ pixel_4003/NB1 pixel_4003/VBIAS pixel_4003/NB2 pixel_4003/AMP_IN pixel_4003/SF_IB
+ pixel_4003/PIX_OUT pixel_4003/CSA_VREF pixel
Xpixel_4014 pixel_4014/gring pixel_4014/VDD pixel_4014/GND pixel_4014/VREF pixel_4014/ROW_SEL
+ pixel_4014/NB1 pixel_4014/VBIAS pixel_4014/NB2 pixel_4014/AMP_IN pixel_4014/SF_IB
+ pixel_4014/PIX_OUT pixel_4014/CSA_VREF pixel
Xpixel_4025 pixel_4025/gring pixel_4025/VDD pixel_4025/GND pixel_4025/VREF pixel_4025/ROW_SEL
+ pixel_4025/NB1 pixel_4025/VBIAS pixel_4025/NB2 pixel_4025/AMP_IN pixel_4025/SF_IB
+ pixel_4025/PIX_OUT pixel_4025/CSA_VREF pixel
Xpixel_3324 pixel_3324/gring pixel_3324/VDD pixel_3324/GND pixel_3324/VREF pixel_3324/ROW_SEL
+ pixel_3324/NB1 pixel_3324/VBIAS pixel_3324/NB2 pixel_3324/AMP_IN pixel_3324/SF_IB
+ pixel_3324/PIX_OUT pixel_3324/CSA_VREF pixel
Xpixel_3313 pixel_3313/gring pixel_3313/VDD pixel_3313/GND pixel_3313/VREF pixel_3313/ROW_SEL
+ pixel_3313/NB1 pixel_3313/VBIAS pixel_3313/NB2 pixel_3313/AMP_IN pixel_3313/SF_IB
+ pixel_3313/PIX_OUT pixel_3313/CSA_VREF pixel
Xpixel_3302 pixel_3302/gring pixel_3302/VDD pixel_3302/GND pixel_3302/VREF pixel_3302/ROW_SEL
+ pixel_3302/NB1 pixel_3302/VBIAS pixel_3302/NB2 pixel_3302/AMP_IN pixel_3302/SF_IB
+ pixel_3302/PIX_OUT pixel_3302/CSA_VREF pixel
Xpixel_4036 pixel_4036/gring pixel_4036/VDD pixel_4036/GND pixel_4036/VREF pixel_4036/ROW_SEL
+ pixel_4036/NB1 pixel_4036/VBIAS pixel_4036/NB2 pixel_4036/AMP_IN pixel_4036/SF_IB
+ pixel_4036/PIX_OUT pixel_4036/CSA_VREF pixel
Xpixel_4047 pixel_4047/gring pixel_4047/VDD pixel_4047/GND pixel_4047/VREF pixel_4047/ROW_SEL
+ pixel_4047/NB1 pixel_4047/VBIAS pixel_4047/NB2 pixel_4047/AMP_IN pixel_4047/SF_IB
+ pixel_4047/PIX_OUT pixel_4047/CSA_VREF pixel
Xpixel_4058 pixel_4058/gring pixel_4058/VDD pixel_4058/GND pixel_4058/VREF pixel_4058/ROW_SEL
+ pixel_4058/NB1 pixel_4058/VBIAS pixel_4058/NB2 pixel_4058/AMP_IN pixel_4058/SF_IB
+ pixel_4058/PIX_OUT pixel_4058/CSA_VREF pixel
Xpixel_4069 pixel_4069/gring pixel_4069/VDD pixel_4069/GND pixel_4069/VREF pixel_4069/ROW_SEL
+ pixel_4069/NB1 pixel_4069/VBIAS pixel_4069/NB2 pixel_4069/AMP_IN pixel_4069/SF_IB
+ pixel_4069/PIX_OUT pixel_4069/CSA_VREF pixel
Xpixel_2612 pixel_2612/gring pixel_2612/VDD pixel_2612/GND pixel_2612/VREF pixel_2612/ROW_SEL
+ pixel_2612/NB1 pixel_2612/VBIAS pixel_2612/NB2 pixel_2612/AMP_IN pixel_2612/SF_IB
+ pixel_2612/PIX_OUT pixel_2612/CSA_VREF pixel
Xpixel_2601 pixel_2601/gring pixel_2601/VDD pixel_2601/GND pixel_2601/VREF pixel_2601/ROW_SEL
+ pixel_2601/NB1 pixel_2601/VBIAS pixel_2601/NB2 pixel_2601/AMP_IN pixel_2601/SF_IB
+ pixel_2601/PIX_OUT pixel_2601/CSA_VREF pixel
Xpixel_3357 pixel_3357/gring pixel_3357/VDD pixel_3357/GND pixel_3357/VREF pixel_3357/ROW_SEL
+ pixel_3357/NB1 pixel_3357/VBIAS pixel_3357/NB2 pixel_3357/AMP_IN pixel_3357/SF_IB
+ pixel_3357/PIX_OUT pixel_3357/CSA_VREF pixel
Xpixel_3346 pixel_3346/gring pixel_3346/VDD pixel_3346/GND pixel_3346/VREF pixel_3346/ROW_SEL
+ pixel_3346/NB1 pixel_3346/VBIAS pixel_3346/NB2 pixel_3346/AMP_IN pixel_3346/SF_IB
+ pixel_3346/PIX_OUT pixel_3346/CSA_VREF pixel
Xpixel_3335 pixel_3335/gring pixel_3335/VDD pixel_3335/GND pixel_3335/VREF pixel_3335/ROW_SEL
+ pixel_3335/NB1 pixel_3335/VBIAS pixel_3335/NB2 pixel_3335/AMP_IN pixel_3335/SF_IB
+ pixel_3335/PIX_OUT pixel_3335/CSA_VREF pixel
Xpixel_1911 pixel_1911/gring pixel_1911/VDD pixel_1911/GND pixel_1911/VREF pixel_1911/ROW_SEL
+ pixel_1911/NB1 pixel_1911/VBIAS pixel_1911/NB2 pixel_1911/AMP_IN pixel_1911/SF_IB
+ pixel_1911/PIX_OUT pixel_1911/CSA_VREF pixel
Xpixel_1900 pixel_1900/gring pixel_1900/VDD pixel_1900/GND pixel_1900/VREF pixel_1900/ROW_SEL
+ pixel_1900/NB1 pixel_1900/VBIAS pixel_1900/NB2 pixel_1900/AMP_IN pixel_1900/SF_IB
+ pixel_1900/PIX_OUT pixel_1900/CSA_VREF pixel
Xpixel_2645 pixel_2645/gring pixel_2645/VDD pixel_2645/GND pixel_2645/VREF pixel_2645/ROW_SEL
+ pixel_2645/NB1 pixel_2645/VBIAS pixel_2645/NB2 pixel_2645/AMP_IN pixel_2645/SF_IB
+ pixel_2645/PIX_OUT pixel_2645/CSA_VREF pixel
Xpixel_2634 pixel_2634/gring pixel_2634/VDD pixel_2634/GND pixel_2634/VREF pixel_2634/ROW_SEL
+ pixel_2634/NB1 pixel_2634/VBIAS pixel_2634/NB2 pixel_2634/AMP_IN pixel_2634/SF_IB
+ pixel_2634/PIX_OUT pixel_2634/CSA_VREF pixel
Xpixel_2623 pixel_2623/gring pixel_2623/VDD pixel_2623/GND pixel_2623/VREF pixel_2623/ROW_SEL
+ pixel_2623/NB1 pixel_2623/VBIAS pixel_2623/NB2 pixel_2623/AMP_IN pixel_2623/SF_IB
+ pixel_2623/PIX_OUT pixel_2623/CSA_VREF pixel
Xpixel_3379 pixel_3379/gring pixel_3379/VDD pixel_3379/GND pixel_3379/VREF pixel_3379/ROW_SEL
+ pixel_3379/NB1 pixel_3379/VBIAS pixel_3379/NB2 pixel_3379/AMP_IN pixel_3379/SF_IB
+ pixel_3379/PIX_OUT pixel_3379/CSA_VREF pixel
Xpixel_3368 pixel_3368/gring pixel_3368/VDD pixel_3368/GND pixel_3368/VREF pixel_3368/ROW_SEL
+ pixel_3368/NB1 pixel_3368/VBIAS pixel_3368/NB2 pixel_3368/AMP_IN pixel_3368/SF_IB
+ pixel_3368/PIX_OUT pixel_3368/CSA_VREF pixel
Xpixel_1944 pixel_1944/gring pixel_1944/VDD pixel_1944/GND pixel_1944/VREF pixel_1944/ROW_SEL
+ pixel_1944/NB1 pixel_1944/VBIAS pixel_1944/NB2 pixel_1944/AMP_IN pixel_1944/SF_IB
+ pixel_1944/PIX_OUT pixel_1944/CSA_VREF pixel
Xpixel_1933 pixel_1933/gring pixel_1933/VDD pixel_1933/GND pixel_1933/VREF pixel_1933/ROW_SEL
+ pixel_1933/NB1 pixel_1933/VBIAS pixel_1933/NB2 pixel_1933/AMP_IN pixel_1933/SF_IB
+ pixel_1933/PIX_OUT pixel_1933/CSA_VREF pixel
Xpixel_1922 pixel_1922/gring pixel_1922/VDD pixel_1922/GND pixel_1922/VREF pixel_1922/ROW_SEL
+ pixel_1922/NB1 pixel_1922/VBIAS pixel_1922/NB2 pixel_1922/AMP_IN pixel_1922/SF_IB
+ pixel_1922/PIX_OUT pixel_1922/CSA_VREF pixel
Xpixel_2689 pixel_2689/gring pixel_2689/VDD pixel_2689/GND pixel_2689/VREF pixel_2689/ROW_SEL
+ pixel_2689/NB1 pixel_2689/VBIAS pixel_2689/NB2 pixel_2689/AMP_IN pixel_2689/SF_IB
+ pixel_2689/PIX_OUT pixel_2689/CSA_VREF pixel
Xpixel_2678 pixel_2678/gring pixel_2678/VDD pixel_2678/GND pixel_2678/VREF pixel_2678/ROW_SEL
+ pixel_2678/NB1 pixel_2678/VBIAS pixel_2678/NB2 pixel_2678/AMP_IN pixel_2678/SF_IB
+ pixel_2678/PIX_OUT pixel_2678/CSA_VREF pixel
Xpixel_2667 pixel_2667/gring pixel_2667/VDD pixel_2667/GND pixel_2667/VREF pixel_2667/ROW_SEL
+ pixel_2667/NB1 pixel_2667/VBIAS pixel_2667/NB2 pixel_2667/AMP_IN pixel_2667/SF_IB
+ pixel_2667/PIX_OUT pixel_2667/CSA_VREF pixel
Xpixel_2656 pixel_2656/gring pixel_2656/VDD pixel_2656/GND pixel_2656/VREF pixel_2656/ROW_SEL
+ pixel_2656/NB1 pixel_2656/VBIAS pixel_2656/NB2 pixel_2656/AMP_IN pixel_2656/SF_IB
+ pixel_2656/PIX_OUT pixel_2656/CSA_VREF pixel
Xpixel_1977 pixel_1977/gring pixel_1977/VDD pixel_1977/GND pixel_1977/VREF pixel_1977/ROW_SEL
+ pixel_1977/NB1 pixel_1977/VBIAS pixel_1977/NB2 pixel_1977/AMP_IN pixel_1977/SF_IB
+ pixel_1977/PIX_OUT pixel_1977/CSA_VREF pixel
Xpixel_1966 pixel_1966/gring pixel_1966/VDD pixel_1966/GND pixel_1966/VREF pixel_1966/ROW_SEL
+ pixel_1966/NB1 pixel_1966/VBIAS pixel_1966/NB2 pixel_1966/AMP_IN pixel_1966/SF_IB
+ pixel_1966/PIX_OUT pixel_1966/CSA_VREF pixel
Xpixel_1955 pixel_1955/gring pixel_1955/VDD pixel_1955/GND pixel_1955/VREF pixel_1955/ROW_SEL
+ pixel_1955/NB1 pixel_1955/VBIAS pixel_1955/NB2 pixel_1955/AMP_IN pixel_1955/SF_IB
+ pixel_1955/PIX_OUT pixel_1955/CSA_VREF pixel
Xpixel_1999 pixel_1999/gring pixel_1999/VDD pixel_1999/GND pixel_1999/VREF pixel_1999/ROW_SEL
+ pixel_1999/NB1 pixel_1999/VBIAS pixel_1999/NB2 pixel_1999/AMP_IN pixel_1999/SF_IB
+ pixel_1999/PIX_OUT pixel_1999/CSA_VREF pixel
Xpixel_1988 pixel_1988/gring pixel_1988/VDD pixel_1988/GND pixel_1988/VREF pixel_1988/ROW_SEL
+ pixel_1988/NB1 pixel_1988/VBIAS pixel_1988/NB2 pixel_1988/AMP_IN pixel_1988/SF_IB
+ pixel_1988/PIX_OUT pixel_1988/CSA_VREF pixel
Xpixel_5260 pixel_5260/gring pixel_5260/VDD pixel_5260/GND pixel_5260/VREF pixel_5260/ROW_SEL
+ pixel_5260/NB1 pixel_5260/VBIAS pixel_5260/NB2 pixel_5260/AMP_IN pixel_5260/SF_IB
+ pixel_5260/PIX_OUT pixel_5260/CSA_VREF pixel
Xpixel_5271 pixel_5271/gring pixel_5271/VDD pixel_5271/GND pixel_5271/VREF pixel_5271/ROW_SEL
+ pixel_5271/NB1 pixel_5271/VBIAS pixel_5271/NB2 pixel_5271/AMP_IN pixel_5271/SF_IB
+ pixel_5271/PIX_OUT pixel_5271/CSA_VREF pixel
Xpixel_5282 pixel_5282/gring pixel_5282/VDD pixel_5282/GND pixel_5282/VREF pixel_5282/ROW_SEL
+ pixel_5282/NB1 pixel_5282/VBIAS pixel_5282/NB2 pixel_5282/AMP_IN pixel_5282/SF_IB
+ pixel_5282/PIX_OUT pixel_5282/CSA_VREF pixel
Xpixel_5293 pixel_5293/gring pixel_5293/VDD pixel_5293/GND pixel_5293/VREF pixel_5293/ROW_SEL
+ pixel_5293/NB1 pixel_5293/VBIAS pixel_5293/NB2 pixel_5293/AMP_IN pixel_5293/SF_IB
+ pixel_5293/PIX_OUT pixel_5293/CSA_VREF pixel
Xpixel_4570 pixel_4570/gring pixel_4570/VDD pixel_4570/GND pixel_4570/VREF pixel_4570/ROW_SEL
+ pixel_4570/NB1 pixel_4570/VBIAS pixel_4570/NB2 pixel_4570/AMP_IN pixel_4570/SF_IB
+ pixel_4570/PIX_OUT pixel_4570/CSA_VREF pixel
Xpixel_4581 pixel_4581/gring pixel_4581/VDD pixel_4581/GND pixel_4581/VREF pixel_4581/ROW_SEL
+ pixel_4581/NB1 pixel_4581/VBIAS pixel_4581/NB2 pixel_4581/AMP_IN pixel_4581/SF_IB
+ pixel_4581/PIX_OUT pixel_4581/CSA_VREF pixel
Xpixel_3880 pixel_3880/gring pixel_3880/VDD pixel_3880/GND pixel_3880/VREF pixel_3880/ROW_SEL
+ pixel_3880/NB1 pixel_3880/VBIAS pixel_3880/NB2 pixel_3880/AMP_IN pixel_3880/SF_IB
+ pixel_3880/PIX_OUT pixel_3880/CSA_VREF pixel
Xpixel_4592 pixel_4592/gring pixel_4592/VDD pixel_4592/GND pixel_4592/VREF pixel_4592/ROW_SEL
+ pixel_4592/NB1 pixel_4592/VBIAS pixel_4592/NB2 pixel_4592/AMP_IN pixel_4592/SF_IB
+ pixel_4592/PIX_OUT pixel_4592/CSA_VREF pixel
Xpixel_3891 pixel_3891/gring pixel_3891/VDD pixel_3891/GND pixel_3891/VREF pixel_3891/ROW_SEL
+ pixel_3891/NB1 pixel_3891/VBIAS pixel_3891/NB2 pixel_3891/AMP_IN pixel_3891/SF_IB
+ pixel_3891/PIX_OUT pixel_3891/CSA_VREF pixel
Xpixel_1229 pixel_1229/gring pixel_1229/VDD pixel_1229/GND pixel_1229/VREF pixel_1229/ROW_SEL
+ pixel_1229/NB1 pixel_1229/VBIAS pixel_1229/NB2 pixel_1229/AMP_IN pixel_1229/SF_IB
+ pixel_1229/PIX_OUT pixel_1229/CSA_VREF pixel
Xpixel_1218 pixel_1218/gring pixel_1218/VDD pixel_1218/GND pixel_1218/VREF pixel_1218/ROW_SEL
+ pixel_1218/NB1 pixel_1218/VBIAS pixel_1218/NB2 pixel_1218/AMP_IN pixel_1218/SF_IB
+ pixel_1218/PIX_OUT pixel_1218/CSA_VREF pixel
Xpixel_1207 pixel_1207/gring pixel_1207/VDD pixel_1207/GND pixel_1207/VREF pixel_1207/ROW_SEL
+ pixel_1207/NB1 pixel_1207/VBIAS pixel_1207/NB2 pixel_1207/AMP_IN pixel_1207/SF_IB
+ pixel_1207/PIX_OUT pixel_1207/CSA_VREF pixel
Xpixel_9504 pixel_9504/gring pixel_9504/VDD pixel_9504/GND pixel_9504/VREF pixel_9504/ROW_SEL
+ pixel_9504/NB1 pixel_9504/VBIAS pixel_9504/NB2 pixel_9504/AMP_IN pixel_9504/SF_IB
+ pixel_9504/PIX_OUT pixel_9504/CSA_VREF pixel
Xpixel_8803 pixel_8803/gring pixel_8803/VDD pixel_8803/GND pixel_8803/VREF pixel_8803/ROW_SEL
+ pixel_8803/NB1 pixel_8803/VBIAS pixel_8803/NB2 pixel_8803/AMP_IN pixel_8803/SF_IB
+ pixel_8803/PIX_OUT pixel_8803/CSA_VREF pixel
Xpixel_9548 pixel_9548/gring pixel_9548/VDD pixel_9548/GND pixel_9548/VREF pixel_9548/ROW_SEL
+ pixel_9548/NB1 pixel_9548/VBIAS pixel_9548/NB2 pixel_9548/AMP_IN pixel_9548/SF_IB
+ pixel_9548/PIX_OUT pixel_9548/CSA_VREF pixel
Xpixel_9537 pixel_9537/gring pixel_9537/VDD pixel_9537/GND pixel_9537/VREF pixel_9537/ROW_SEL
+ pixel_9537/NB1 pixel_9537/VBIAS pixel_9537/NB2 pixel_9537/AMP_IN pixel_9537/SF_IB
+ pixel_9537/PIX_OUT pixel_9537/CSA_VREF pixel
Xpixel_9526 pixel_9526/gring pixel_9526/VDD pixel_9526/GND pixel_9526/VREF pixel_9526/ROW_SEL
+ pixel_9526/NB1 pixel_9526/VBIAS pixel_9526/NB2 pixel_9526/AMP_IN pixel_9526/SF_IB
+ pixel_9526/PIX_OUT pixel_9526/CSA_VREF pixel
Xpixel_9515 pixel_9515/gring pixel_9515/VDD pixel_9515/GND pixel_9515/VREF pixel_9515/ROW_SEL
+ pixel_9515/NB1 pixel_9515/VBIAS pixel_9515/NB2 pixel_9515/AMP_IN pixel_9515/SF_IB
+ pixel_9515/PIX_OUT pixel_9515/CSA_VREF pixel
Xpixel_8836 pixel_8836/gring pixel_8836/VDD pixel_8836/GND pixel_8836/VREF pixel_8836/ROW_SEL
+ pixel_8836/NB1 pixel_8836/VBIAS pixel_8836/NB2 pixel_8836/AMP_IN pixel_8836/SF_IB
+ pixel_8836/PIX_OUT pixel_8836/CSA_VREF pixel
Xpixel_8825 pixel_8825/gring pixel_8825/VDD pixel_8825/GND pixel_8825/VREF pixel_8825/ROW_SEL
+ pixel_8825/NB1 pixel_8825/VBIAS pixel_8825/NB2 pixel_8825/AMP_IN pixel_8825/SF_IB
+ pixel_8825/PIX_OUT pixel_8825/CSA_VREF pixel
Xpixel_8814 pixel_8814/gring pixel_8814/VDD pixel_8814/GND pixel_8814/VREF pixel_8814/ROW_SEL
+ pixel_8814/NB1 pixel_8814/VBIAS pixel_8814/NB2 pixel_8814/AMP_IN pixel_8814/SF_IB
+ pixel_8814/PIX_OUT pixel_8814/CSA_VREF pixel
Xpixel_9559 pixel_9559/gring pixel_9559/VDD pixel_9559/GND pixel_9559/VREF pixel_9559/ROW_SEL
+ pixel_9559/NB1 pixel_9559/VBIAS pixel_9559/NB2 pixel_9559/AMP_IN pixel_9559/SF_IB
+ pixel_9559/PIX_OUT pixel_9559/CSA_VREF pixel
Xpixel_8869 pixel_8869/gring pixel_8869/VDD pixel_8869/GND pixel_8869/VREF pixel_8869/ROW_SEL
+ pixel_8869/NB1 pixel_8869/VBIAS pixel_8869/NB2 pixel_8869/AMP_IN pixel_8869/SF_IB
+ pixel_8869/PIX_OUT pixel_8869/CSA_VREF pixel
Xpixel_8858 pixel_8858/gring pixel_8858/VDD pixel_8858/GND pixel_8858/VREF pixel_8858/ROW_SEL
+ pixel_8858/NB1 pixel_8858/VBIAS pixel_8858/NB2 pixel_8858/AMP_IN pixel_8858/SF_IB
+ pixel_8858/PIX_OUT pixel_8858/CSA_VREF pixel
Xpixel_8847 pixel_8847/gring pixel_8847/VDD pixel_8847/GND pixel_8847/VREF pixel_8847/ROW_SEL
+ pixel_8847/NB1 pixel_8847/VBIAS pixel_8847/NB2 pixel_8847/AMP_IN pixel_8847/SF_IB
+ pixel_8847/PIX_OUT pixel_8847/CSA_VREF pixel
Xpixel_3132 pixel_3132/gring pixel_3132/VDD pixel_3132/GND pixel_3132/VREF pixel_3132/ROW_SEL
+ pixel_3132/NB1 pixel_3132/VBIAS pixel_3132/NB2 pixel_3132/AMP_IN pixel_3132/SF_IB
+ pixel_3132/PIX_OUT pixel_3132/CSA_VREF pixel
Xpixel_3121 pixel_3121/gring pixel_3121/VDD pixel_3121/GND pixel_3121/VREF pixel_3121/ROW_SEL
+ pixel_3121/NB1 pixel_3121/VBIAS pixel_3121/NB2 pixel_3121/AMP_IN pixel_3121/SF_IB
+ pixel_3121/PIX_OUT pixel_3121/CSA_VREF pixel
Xpixel_3110 pixel_3110/gring pixel_3110/VDD pixel_3110/GND pixel_3110/VREF pixel_3110/ROW_SEL
+ pixel_3110/NB1 pixel_3110/VBIAS pixel_3110/NB2 pixel_3110/AMP_IN pixel_3110/SF_IB
+ pixel_3110/PIX_OUT pixel_3110/CSA_VREF pixel
Xpixel_2420 pixel_2420/gring pixel_2420/VDD pixel_2420/GND pixel_2420/VREF pixel_2420/ROW_SEL
+ pixel_2420/NB1 pixel_2420/VBIAS pixel_2420/NB2 pixel_2420/AMP_IN pixel_2420/SF_IB
+ pixel_2420/PIX_OUT pixel_2420/CSA_VREF pixel
Xpixel_3165 pixel_3165/gring pixel_3165/VDD pixel_3165/GND pixel_3165/VREF pixel_3165/ROW_SEL
+ pixel_3165/NB1 pixel_3165/VBIAS pixel_3165/NB2 pixel_3165/AMP_IN pixel_3165/SF_IB
+ pixel_3165/PIX_OUT pixel_3165/CSA_VREF pixel
Xpixel_3154 pixel_3154/gring pixel_3154/VDD pixel_3154/GND pixel_3154/VREF pixel_3154/ROW_SEL
+ pixel_3154/NB1 pixel_3154/VBIAS pixel_3154/NB2 pixel_3154/AMP_IN pixel_3154/SF_IB
+ pixel_3154/PIX_OUT pixel_3154/CSA_VREF pixel
Xpixel_3143 pixel_3143/gring pixel_3143/VDD pixel_3143/GND pixel_3143/VREF pixel_3143/ROW_SEL
+ pixel_3143/NB1 pixel_3143/VBIAS pixel_3143/NB2 pixel_3143/AMP_IN pixel_3143/SF_IB
+ pixel_3143/PIX_OUT pixel_3143/CSA_VREF pixel
Xpixel_2464 pixel_2464/gring pixel_2464/VDD pixel_2464/GND pixel_2464/VREF pixel_2464/ROW_SEL
+ pixel_2464/NB1 pixel_2464/VBIAS pixel_2464/NB2 pixel_2464/AMP_IN pixel_2464/SF_IB
+ pixel_2464/PIX_OUT pixel_2464/CSA_VREF pixel
Xpixel_2453 pixel_2453/gring pixel_2453/VDD pixel_2453/GND pixel_2453/VREF pixel_2453/ROW_SEL
+ pixel_2453/NB1 pixel_2453/VBIAS pixel_2453/NB2 pixel_2453/AMP_IN pixel_2453/SF_IB
+ pixel_2453/PIX_OUT pixel_2453/CSA_VREF pixel
Xpixel_2442 pixel_2442/gring pixel_2442/VDD pixel_2442/GND pixel_2442/VREF pixel_2442/ROW_SEL
+ pixel_2442/NB1 pixel_2442/VBIAS pixel_2442/NB2 pixel_2442/AMP_IN pixel_2442/SF_IB
+ pixel_2442/PIX_OUT pixel_2442/CSA_VREF pixel
Xpixel_2431 pixel_2431/gring pixel_2431/VDD pixel_2431/GND pixel_2431/VREF pixel_2431/ROW_SEL
+ pixel_2431/NB1 pixel_2431/VBIAS pixel_2431/NB2 pixel_2431/AMP_IN pixel_2431/SF_IB
+ pixel_2431/PIX_OUT pixel_2431/CSA_VREF pixel
Xpixel_3198 pixel_3198/gring pixel_3198/VDD pixel_3198/GND pixel_3198/VREF pixel_3198/ROW_SEL
+ pixel_3198/NB1 pixel_3198/VBIAS pixel_3198/NB2 pixel_3198/AMP_IN pixel_3198/SF_IB
+ pixel_3198/PIX_OUT pixel_3198/CSA_VREF pixel
Xpixel_3187 pixel_3187/gring pixel_3187/VDD pixel_3187/GND pixel_3187/VREF pixel_3187/ROW_SEL
+ pixel_3187/NB1 pixel_3187/VBIAS pixel_3187/NB2 pixel_3187/AMP_IN pixel_3187/SF_IB
+ pixel_3187/PIX_OUT pixel_3187/CSA_VREF pixel
Xpixel_3176 pixel_3176/gring pixel_3176/VDD pixel_3176/GND pixel_3176/VREF pixel_3176/ROW_SEL
+ pixel_3176/NB1 pixel_3176/VBIAS pixel_3176/NB2 pixel_3176/AMP_IN pixel_3176/SF_IB
+ pixel_3176/PIX_OUT pixel_3176/CSA_VREF pixel
Xpixel_1752 pixel_1752/gring pixel_1752/VDD pixel_1752/GND pixel_1752/VREF pixel_1752/ROW_SEL
+ pixel_1752/NB1 pixel_1752/VBIAS pixel_1752/NB2 pixel_1752/AMP_IN pixel_1752/SF_IB
+ pixel_1752/PIX_OUT pixel_1752/CSA_VREF pixel
Xpixel_1741 pixel_1741/gring pixel_1741/VDD pixel_1741/GND pixel_1741/VREF pixel_1741/ROW_SEL
+ pixel_1741/NB1 pixel_1741/VBIAS pixel_1741/NB2 pixel_1741/AMP_IN pixel_1741/SF_IB
+ pixel_1741/PIX_OUT pixel_1741/CSA_VREF pixel
Xpixel_1730 pixel_1730/gring pixel_1730/VDD pixel_1730/GND pixel_1730/VREF pixel_1730/ROW_SEL
+ pixel_1730/NB1 pixel_1730/VBIAS pixel_1730/NB2 pixel_1730/AMP_IN pixel_1730/SF_IB
+ pixel_1730/PIX_OUT pixel_1730/CSA_VREF pixel
Xpixel_2497 pixel_2497/gring pixel_2497/VDD pixel_2497/GND pixel_2497/VREF pixel_2497/ROW_SEL
+ pixel_2497/NB1 pixel_2497/VBIAS pixel_2497/NB2 pixel_2497/AMP_IN pixel_2497/SF_IB
+ pixel_2497/PIX_OUT pixel_2497/CSA_VREF pixel
Xpixel_2486 pixel_2486/gring pixel_2486/VDD pixel_2486/GND pixel_2486/VREF pixel_2486/ROW_SEL
+ pixel_2486/NB1 pixel_2486/VBIAS pixel_2486/NB2 pixel_2486/AMP_IN pixel_2486/SF_IB
+ pixel_2486/PIX_OUT pixel_2486/CSA_VREF pixel
Xpixel_2475 pixel_2475/gring pixel_2475/VDD pixel_2475/GND pixel_2475/VREF pixel_2475/ROW_SEL
+ pixel_2475/NB1 pixel_2475/VBIAS pixel_2475/NB2 pixel_2475/AMP_IN pixel_2475/SF_IB
+ pixel_2475/PIX_OUT pixel_2475/CSA_VREF pixel
Xpixel_1785 pixel_1785/gring pixel_1785/VDD pixel_1785/GND pixel_1785/VREF pixel_1785/ROW_SEL
+ pixel_1785/NB1 pixel_1785/VBIAS pixel_1785/NB2 pixel_1785/AMP_IN pixel_1785/SF_IB
+ pixel_1785/PIX_OUT pixel_1785/CSA_VREF pixel
Xpixel_1774 pixel_1774/gring pixel_1774/VDD pixel_1774/GND pixel_1774/VREF pixel_1774/ROW_SEL
+ pixel_1774/NB1 pixel_1774/VBIAS pixel_1774/NB2 pixel_1774/AMP_IN pixel_1774/SF_IB
+ pixel_1774/PIX_OUT pixel_1774/CSA_VREF pixel
Xpixel_1763 pixel_1763/gring pixel_1763/VDD pixel_1763/GND pixel_1763/VREF pixel_1763/ROW_SEL
+ pixel_1763/NB1 pixel_1763/VBIAS pixel_1763/NB2 pixel_1763/AMP_IN pixel_1763/SF_IB
+ pixel_1763/PIX_OUT pixel_1763/CSA_VREF pixel
Xpixel_1796 pixel_1796/gring pixel_1796/VDD pixel_1796/GND pixel_1796/VREF pixel_1796/ROW_SEL
+ pixel_1796/NB1 pixel_1796/VBIAS pixel_1796/NB2 pixel_1796/AMP_IN pixel_1796/SF_IB
+ pixel_1796/PIX_OUT pixel_1796/CSA_VREF pixel
Xpixel_5090 pixel_5090/gring pixel_5090/VDD pixel_5090/GND pixel_5090/VREF pixel_5090/ROW_SEL
+ pixel_5090/NB1 pixel_5090/VBIAS pixel_5090/NB2 pixel_5090/AMP_IN pixel_5090/SF_IB
+ pixel_5090/PIX_OUT pixel_5090/CSA_VREF pixel
Xpixel_7409 pixel_7409/gring pixel_7409/VDD pixel_7409/GND pixel_7409/VREF pixel_7409/ROW_SEL
+ pixel_7409/NB1 pixel_7409/VBIAS pixel_7409/NB2 pixel_7409/AMP_IN pixel_7409/SF_IB
+ pixel_7409/PIX_OUT pixel_7409/CSA_VREF pixel
Xpixel_6708 pixel_6708/gring pixel_6708/VDD pixel_6708/GND pixel_6708/VREF pixel_6708/ROW_SEL
+ pixel_6708/NB1 pixel_6708/VBIAS pixel_6708/NB2 pixel_6708/AMP_IN pixel_6708/SF_IB
+ pixel_6708/PIX_OUT pixel_6708/CSA_VREF pixel
Xpixel_6719 pixel_6719/gring pixel_6719/VDD pixel_6719/GND pixel_6719/VREF pixel_6719/ROW_SEL
+ pixel_6719/NB1 pixel_6719/VBIAS pixel_6719/NB2 pixel_6719/AMP_IN pixel_6719/SF_IB
+ pixel_6719/PIX_OUT pixel_6719/CSA_VREF pixel
Xpixel_1004 pixel_1004/gring pixel_1004/VDD pixel_1004/GND pixel_1004/VREF pixel_1004/ROW_SEL
+ pixel_1004/NB1 pixel_1004/VBIAS pixel_1004/NB2 pixel_1004/AMP_IN pixel_1004/SF_IB
+ pixel_1004/PIX_OUT pixel_1004/CSA_VREF pixel
Xpixel_1048 pixel_1048/gring pixel_1048/VDD pixel_1048/GND pixel_1048/VREF pixel_1048/ROW_SEL
+ pixel_1048/NB1 pixel_1048/VBIAS pixel_1048/NB2 pixel_1048/AMP_IN pixel_1048/SF_IB
+ pixel_1048/PIX_OUT pixel_1048/CSA_VREF pixel
Xpixel_1037 pixel_1037/gring pixel_1037/VDD pixel_1037/GND pixel_1037/VREF pixel_1037/ROW_SEL
+ pixel_1037/NB1 pixel_1037/VBIAS pixel_1037/NB2 pixel_1037/AMP_IN pixel_1037/SF_IB
+ pixel_1037/PIX_OUT pixel_1037/CSA_VREF pixel
Xpixel_1026 pixel_1026/gring pixel_1026/VDD pixel_1026/GND pixel_1026/VREF pixel_1026/ROW_SEL
+ pixel_1026/NB1 pixel_1026/VBIAS pixel_1026/NB2 pixel_1026/AMP_IN pixel_1026/SF_IB
+ pixel_1026/PIX_OUT pixel_1026/CSA_VREF pixel
Xpixel_1015 pixel_1015/gring pixel_1015/VDD pixel_1015/GND pixel_1015/VREF pixel_1015/ROW_SEL
+ pixel_1015/NB1 pixel_1015/VBIAS pixel_1015/NB2 pixel_1015/AMP_IN pixel_1015/SF_IB
+ pixel_1015/PIX_OUT pixel_1015/CSA_VREF pixel
Xpixel_1059 pixel_1059/gring pixel_1059/VDD pixel_1059/GND pixel_1059/VREF pixel_1059/ROW_SEL
+ pixel_1059/NB1 pixel_1059/VBIAS pixel_1059/NB2 pixel_1059/AMP_IN pixel_1059/SF_IB
+ pixel_1059/PIX_OUT pixel_1059/CSA_VREF pixel
Xpixel_9312 pixel_9312/gring pixel_9312/VDD pixel_9312/GND pixel_9312/VREF pixel_9312/ROW_SEL
+ pixel_9312/NB1 pixel_9312/VBIAS pixel_9312/NB2 pixel_9312/AMP_IN pixel_9312/SF_IB
+ pixel_9312/PIX_OUT pixel_9312/CSA_VREF pixel
Xpixel_9301 pixel_9301/gring pixel_9301/VDD pixel_9301/GND pixel_9301/VREF pixel_9301/ROW_SEL
+ pixel_9301/NB1 pixel_9301/VBIAS pixel_9301/NB2 pixel_9301/AMP_IN pixel_9301/SF_IB
+ pixel_9301/PIX_OUT pixel_9301/CSA_VREF pixel
Xpixel_8611 pixel_8611/gring pixel_8611/VDD pixel_8611/GND pixel_8611/VREF pixel_8611/ROW_SEL
+ pixel_8611/NB1 pixel_8611/VBIAS pixel_8611/NB2 pixel_8611/AMP_IN pixel_8611/SF_IB
+ pixel_8611/PIX_OUT pixel_8611/CSA_VREF pixel
Xpixel_8600 pixel_8600/gring pixel_8600/VDD pixel_8600/GND pixel_8600/VREF pixel_8600/ROW_SEL
+ pixel_8600/NB1 pixel_8600/VBIAS pixel_8600/NB2 pixel_8600/AMP_IN pixel_8600/SF_IB
+ pixel_8600/PIX_OUT pixel_8600/CSA_VREF pixel
Xpixel_9356 pixel_9356/gring pixel_9356/VDD pixel_9356/GND pixel_9356/VREF pixel_9356/ROW_SEL
+ pixel_9356/NB1 pixel_9356/VBIAS pixel_9356/NB2 pixel_9356/AMP_IN pixel_9356/SF_IB
+ pixel_9356/PIX_OUT pixel_9356/CSA_VREF pixel
Xpixel_9345 pixel_9345/gring pixel_9345/VDD pixel_9345/GND pixel_9345/VREF pixel_9345/ROW_SEL
+ pixel_9345/NB1 pixel_9345/VBIAS pixel_9345/NB2 pixel_9345/AMP_IN pixel_9345/SF_IB
+ pixel_9345/PIX_OUT pixel_9345/CSA_VREF pixel
Xpixel_9334 pixel_9334/gring pixel_9334/VDD pixel_9334/GND pixel_9334/VREF pixel_9334/ROW_SEL
+ pixel_9334/NB1 pixel_9334/VBIAS pixel_9334/NB2 pixel_9334/AMP_IN pixel_9334/SF_IB
+ pixel_9334/PIX_OUT pixel_9334/CSA_VREF pixel
Xpixel_9323 pixel_9323/gring pixel_9323/VDD pixel_9323/GND pixel_9323/VREF pixel_9323/ROW_SEL
+ pixel_9323/NB1 pixel_9323/VBIAS pixel_9323/NB2 pixel_9323/AMP_IN pixel_9323/SF_IB
+ pixel_9323/PIX_OUT pixel_9323/CSA_VREF pixel
Xpixel_8644 pixel_8644/gring pixel_8644/VDD pixel_8644/GND pixel_8644/VREF pixel_8644/ROW_SEL
+ pixel_8644/NB1 pixel_8644/VBIAS pixel_8644/NB2 pixel_8644/AMP_IN pixel_8644/SF_IB
+ pixel_8644/PIX_OUT pixel_8644/CSA_VREF pixel
Xpixel_8633 pixel_8633/gring pixel_8633/VDD pixel_8633/GND pixel_8633/VREF pixel_8633/ROW_SEL
+ pixel_8633/NB1 pixel_8633/VBIAS pixel_8633/NB2 pixel_8633/AMP_IN pixel_8633/SF_IB
+ pixel_8633/PIX_OUT pixel_8633/CSA_VREF pixel
Xpixel_8622 pixel_8622/gring pixel_8622/VDD pixel_8622/GND pixel_8622/VREF pixel_8622/ROW_SEL
+ pixel_8622/NB1 pixel_8622/VBIAS pixel_8622/NB2 pixel_8622/AMP_IN pixel_8622/SF_IB
+ pixel_8622/PIX_OUT pixel_8622/CSA_VREF pixel
Xpixel_9389 pixel_9389/gring pixel_9389/VDD pixel_9389/GND pixel_9389/VREF pixel_9389/ROW_SEL
+ pixel_9389/NB1 pixel_9389/VBIAS pixel_9389/NB2 pixel_9389/AMP_IN pixel_9389/SF_IB
+ pixel_9389/PIX_OUT pixel_9389/CSA_VREF pixel
Xpixel_9378 pixel_9378/gring pixel_9378/VDD pixel_9378/GND pixel_9378/VREF pixel_9378/ROW_SEL
+ pixel_9378/NB1 pixel_9378/VBIAS pixel_9378/NB2 pixel_9378/AMP_IN pixel_9378/SF_IB
+ pixel_9378/PIX_OUT pixel_9378/CSA_VREF pixel
Xpixel_9367 pixel_9367/gring pixel_9367/VDD pixel_9367/GND pixel_9367/VREF pixel_9367/ROW_SEL
+ pixel_9367/NB1 pixel_9367/VBIAS pixel_9367/NB2 pixel_9367/AMP_IN pixel_9367/SF_IB
+ pixel_9367/PIX_OUT pixel_9367/CSA_VREF pixel
Xpixel_8688 pixel_8688/gring pixel_8688/VDD pixel_8688/GND pixel_8688/VREF pixel_8688/ROW_SEL
+ pixel_8688/NB1 pixel_8688/VBIAS pixel_8688/NB2 pixel_8688/AMP_IN pixel_8688/SF_IB
+ pixel_8688/PIX_OUT pixel_8688/CSA_VREF pixel
Xpixel_8677 pixel_8677/gring pixel_8677/VDD pixel_8677/GND pixel_8677/VREF pixel_8677/ROW_SEL
+ pixel_8677/NB1 pixel_8677/VBIAS pixel_8677/NB2 pixel_8677/AMP_IN pixel_8677/SF_IB
+ pixel_8677/PIX_OUT pixel_8677/CSA_VREF pixel
Xpixel_8666 pixel_8666/gring pixel_8666/VDD pixel_8666/GND pixel_8666/VREF pixel_8666/ROW_SEL
+ pixel_8666/NB1 pixel_8666/VBIAS pixel_8666/NB2 pixel_8666/AMP_IN pixel_8666/SF_IB
+ pixel_8666/PIX_OUT pixel_8666/CSA_VREF pixel
Xpixel_8655 pixel_8655/gring pixel_8655/VDD pixel_8655/GND pixel_8655/VREF pixel_8655/ROW_SEL
+ pixel_8655/NB1 pixel_8655/VBIAS pixel_8655/NB2 pixel_8655/AMP_IN pixel_8655/SF_IB
+ pixel_8655/PIX_OUT pixel_8655/CSA_VREF pixel
Xpixel_7910 pixel_7910/gring pixel_7910/VDD pixel_7910/GND pixel_7910/VREF pixel_7910/ROW_SEL
+ pixel_7910/NB1 pixel_7910/VBIAS pixel_7910/NB2 pixel_7910/AMP_IN pixel_7910/SF_IB
+ pixel_7910/PIX_OUT pixel_7910/CSA_VREF pixel
Xpixel_7921 pixel_7921/gring pixel_7921/VDD pixel_7921/GND pixel_7921/VREF pixel_7921/ROW_SEL
+ pixel_7921/NB1 pixel_7921/VBIAS pixel_7921/NB2 pixel_7921/AMP_IN pixel_7921/SF_IB
+ pixel_7921/PIX_OUT pixel_7921/CSA_VREF pixel
Xpixel_7932 pixel_7932/gring pixel_7932/VDD pixel_7932/GND pixel_7932/VREF pixel_7932/ROW_SEL
+ pixel_7932/NB1 pixel_7932/VBIAS pixel_7932/NB2 pixel_7932/AMP_IN pixel_7932/SF_IB
+ pixel_7932/PIX_OUT pixel_7932/CSA_VREF pixel
Xpixel_7943 pixel_7943/gring pixel_7943/VDD pixel_7943/GND pixel_7943/VREF pixel_7943/ROW_SEL
+ pixel_7943/NB1 pixel_7943/VBIAS pixel_7943/NB2 pixel_7943/AMP_IN pixel_7943/SF_IB
+ pixel_7943/PIX_OUT pixel_7943/CSA_VREF pixel
Xpixel_8699 pixel_8699/gring pixel_8699/VDD pixel_8699/GND pixel_8699/VREF pixel_8699/ROW_SEL
+ pixel_8699/NB1 pixel_8699/VBIAS pixel_8699/NB2 pixel_8699/AMP_IN pixel_8699/SF_IB
+ pixel_8699/PIX_OUT pixel_8699/CSA_VREF pixel
Xpixel_7954 pixel_7954/gring pixel_7954/VDD pixel_7954/GND pixel_7954/VREF pixel_7954/ROW_SEL
+ pixel_7954/NB1 pixel_7954/VBIAS pixel_7954/NB2 pixel_7954/AMP_IN pixel_7954/SF_IB
+ pixel_7954/PIX_OUT pixel_7954/CSA_VREF pixel
Xpixel_7965 pixel_7965/gring pixel_7965/VDD pixel_7965/GND pixel_7965/VREF pixel_7965/ROW_SEL
+ pixel_7965/NB1 pixel_7965/VBIAS pixel_7965/NB2 pixel_7965/AMP_IN pixel_7965/SF_IB
+ pixel_7965/PIX_OUT pixel_7965/CSA_VREF pixel
Xpixel_7976 pixel_7976/gring pixel_7976/VDD pixel_7976/GND pixel_7976/VREF pixel_7976/ROW_SEL
+ pixel_7976/NB1 pixel_7976/VBIAS pixel_7976/NB2 pixel_7976/AMP_IN pixel_7976/SF_IB
+ pixel_7976/PIX_OUT pixel_7976/CSA_VREF pixel
Xpixel_7987 pixel_7987/gring pixel_7987/VDD pixel_7987/GND pixel_7987/VREF pixel_7987/ROW_SEL
+ pixel_7987/NB1 pixel_7987/VBIAS pixel_7987/NB2 pixel_7987/AMP_IN pixel_7987/SF_IB
+ pixel_7987/PIX_OUT pixel_7987/CSA_VREF pixel
Xpixel_7998 pixel_7998/gring pixel_7998/VDD pixel_7998/GND pixel_7998/VREF pixel_7998/ROW_SEL
+ pixel_7998/NB1 pixel_7998/VBIAS pixel_7998/NB2 pixel_7998/AMP_IN pixel_7998/SF_IB
+ pixel_7998/PIX_OUT pixel_7998/CSA_VREF pixel
Xpixel_2272 pixel_2272/gring pixel_2272/VDD pixel_2272/GND pixel_2272/VREF pixel_2272/ROW_SEL
+ pixel_2272/NB1 pixel_2272/VBIAS pixel_2272/NB2 pixel_2272/AMP_IN pixel_2272/SF_IB
+ pixel_2272/PIX_OUT pixel_2272/CSA_VREF pixel
Xpixel_2261 pixel_2261/gring pixel_2261/VDD pixel_2261/GND pixel_2261/VREF pixel_2261/ROW_SEL
+ pixel_2261/NB1 pixel_2261/VBIAS pixel_2261/NB2 pixel_2261/AMP_IN pixel_2261/SF_IB
+ pixel_2261/PIX_OUT pixel_2261/CSA_VREF pixel
Xpixel_2250 pixel_2250/gring pixel_2250/VDD pixel_2250/GND pixel_2250/VREF pixel_2250/ROW_SEL
+ pixel_2250/NB1 pixel_2250/VBIAS pixel_2250/NB2 pixel_2250/AMP_IN pixel_2250/SF_IB
+ pixel_2250/PIX_OUT pixel_2250/CSA_VREF pixel
Xpixel_1560 pixel_1560/gring pixel_1560/VDD pixel_1560/GND pixel_1560/VREF pixel_1560/ROW_SEL
+ pixel_1560/NB1 pixel_1560/VBIAS pixel_1560/NB2 pixel_1560/AMP_IN pixel_1560/SF_IB
+ pixel_1560/PIX_OUT pixel_1560/CSA_VREF pixel
Xpixel_2294 pixel_2294/gring pixel_2294/VDD pixel_2294/GND pixel_2294/VREF pixel_2294/ROW_SEL
+ pixel_2294/NB1 pixel_2294/VBIAS pixel_2294/NB2 pixel_2294/AMP_IN pixel_2294/SF_IB
+ pixel_2294/PIX_OUT pixel_2294/CSA_VREF pixel
Xpixel_2283 pixel_2283/gring pixel_2283/VDD pixel_2283/GND pixel_2283/VREF pixel_2283/ROW_SEL
+ pixel_2283/NB1 pixel_2283/VBIAS pixel_2283/NB2 pixel_2283/AMP_IN pixel_2283/SF_IB
+ pixel_2283/PIX_OUT pixel_2283/CSA_VREF pixel
Xpixel_1593 pixel_1593/gring pixel_1593/VDD pixel_1593/GND pixel_1593/VREF pixel_1593/ROW_SEL
+ pixel_1593/NB1 pixel_1593/VBIAS pixel_1593/NB2 pixel_1593/AMP_IN pixel_1593/SF_IB
+ pixel_1593/PIX_OUT pixel_1593/CSA_VREF pixel
Xpixel_1582 pixel_1582/gring pixel_1582/VDD pixel_1582/GND pixel_1582/VREF pixel_1582/ROW_SEL
+ pixel_1582/NB1 pixel_1582/VBIAS pixel_1582/NB2 pixel_1582/AMP_IN pixel_1582/SF_IB
+ pixel_1582/PIX_OUT pixel_1582/CSA_VREF pixel
Xpixel_1571 pixel_1571/gring pixel_1571/VDD pixel_1571/GND pixel_1571/VREF pixel_1571/ROW_SEL
+ pixel_1571/NB1 pixel_1571/VBIAS pixel_1571/NB2 pixel_1571/AMP_IN pixel_1571/SF_IB
+ pixel_1571/PIX_OUT pixel_1571/CSA_VREF pixel
Xpixel_9890 pixel_9890/gring pixel_9890/VDD pixel_9890/GND pixel_9890/VREF pixel_9890/ROW_SEL
+ pixel_9890/NB1 pixel_9890/VBIAS pixel_9890/NB2 pixel_9890/AMP_IN pixel_9890/SF_IB
+ pixel_9890/PIX_OUT pixel_9890/CSA_VREF pixel
Xpixel_619 pixel_619/gring pixel_619/VDD pixel_619/GND pixel_619/VREF pixel_619/ROW_SEL
+ pixel_619/NB1 pixel_619/VBIAS pixel_619/NB2 pixel_619/AMP_IN pixel_619/SF_IB pixel_619/PIX_OUT
+ pixel_619/CSA_VREF pixel
Xpixel_608 pixel_608/gring pixel_608/VDD pixel_608/GND pixel_608/VREF pixel_608/ROW_SEL
+ pixel_608/NB1 pixel_608/VBIAS pixel_608/NB2 pixel_608/AMP_IN pixel_608/SF_IB pixel_608/PIX_OUT
+ pixel_608/CSA_VREF pixel
Xpixel_7206 pixel_7206/gring pixel_7206/VDD pixel_7206/GND pixel_7206/VREF pixel_7206/ROW_SEL
+ pixel_7206/NB1 pixel_7206/VBIAS pixel_7206/NB2 pixel_7206/AMP_IN pixel_7206/SF_IB
+ pixel_7206/PIX_OUT pixel_7206/CSA_VREF pixel
Xpixel_7217 pixel_7217/gring pixel_7217/VDD pixel_7217/GND pixel_7217/VREF pixel_7217/ROW_SEL
+ pixel_7217/NB1 pixel_7217/VBIAS pixel_7217/NB2 pixel_7217/AMP_IN pixel_7217/SF_IB
+ pixel_7217/PIX_OUT pixel_7217/CSA_VREF pixel
Xpixel_7228 pixel_7228/gring pixel_7228/VDD pixel_7228/GND pixel_7228/VREF pixel_7228/ROW_SEL
+ pixel_7228/NB1 pixel_7228/VBIAS pixel_7228/NB2 pixel_7228/AMP_IN pixel_7228/SF_IB
+ pixel_7228/PIX_OUT pixel_7228/CSA_VREF pixel
Xpixel_7239 pixel_7239/gring pixel_7239/VDD pixel_7239/GND pixel_7239/VREF pixel_7239/ROW_SEL
+ pixel_7239/NB1 pixel_7239/VBIAS pixel_7239/NB2 pixel_7239/AMP_IN pixel_7239/SF_IB
+ pixel_7239/PIX_OUT pixel_7239/CSA_VREF pixel
Xpixel_6505 pixel_6505/gring pixel_6505/VDD pixel_6505/GND pixel_6505/VREF pixel_6505/ROW_SEL
+ pixel_6505/NB1 pixel_6505/VBIAS pixel_6505/NB2 pixel_6505/AMP_IN pixel_6505/SF_IB
+ pixel_6505/PIX_OUT pixel_6505/CSA_VREF pixel
Xpixel_6516 pixel_6516/gring pixel_6516/VDD pixel_6516/GND pixel_6516/VREF pixel_6516/ROW_SEL
+ pixel_6516/NB1 pixel_6516/VBIAS pixel_6516/NB2 pixel_6516/AMP_IN pixel_6516/SF_IB
+ pixel_6516/PIX_OUT pixel_6516/CSA_VREF pixel
Xpixel_6527 pixel_6527/gring pixel_6527/VDD pixel_6527/GND pixel_6527/VREF pixel_6527/ROW_SEL
+ pixel_6527/NB1 pixel_6527/VBIAS pixel_6527/NB2 pixel_6527/AMP_IN pixel_6527/SF_IB
+ pixel_6527/PIX_OUT pixel_6527/CSA_VREF pixel
Xpixel_6538 pixel_6538/gring pixel_6538/VDD pixel_6538/GND pixel_6538/VREF pixel_6538/ROW_SEL
+ pixel_6538/NB1 pixel_6538/VBIAS pixel_6538/NB2 pixel_6538/AMP_IN pixel_6538/SF_IB
+ pixel_6538/PIX_OUT pixel_6538/CSA_VREF pixel
Xpixel_6549 pixel_6549/gring pixel_6549/VDD pixel_6549/GND pixel_6549/VREF pixel_6549/ROW_SEL
+ pixel_6549/NB1 pixel_6549/VBIAS pixel_6549/NB2 pixel_6549/AMP_IN pixel_6549/SF_IB
+ pixel_6549/PIX_OUT pixel_6549/CSA_VREF pixel
Xpixel_5804 pixel_5804/gring pixel_5804/VDD pixel_5804/GND pixel_5804/VREF pixel_5804/ROW_SEL
+ pixel_5804/NB1 pixel_5804/VBIAS pixel_5804/NB2 pixel_5804/AMP_IN pixel_5804/SF_IB
+ pixel_5804/PIX_OUT pixel_5804/CSA_VREF pixel
Xpixel_5815 pixel_5815/gring pixel_5815/VDD pixel_5815/GND pixel_5815/VREF pixel_5815/ROW_SEL
+ pixel_5815/NB1 pixel_5815/VBIAS pixel_5815/NB2 pixel_5815/AMP_IN pixel_5815/SF_IB
+ pixel_5815/PIX_OUT pixel_5815/CSA_VREF pixel
Xpixel_5826 pixel_5826/gring pixel_5826/VDD pixel_5826/GND pixel_5826/VREF pixel_5826/ROW_SEL
+ pixel_5826/NB1 pixel_5826/VBIAS pixel_5826/NB2 pixel_5826/AMP_IN pixel_5826/SF_IB
+ pixel_5826/PIX_OUT pixel_5826/CSA_VREF pixel
Xpixel_5837 pixel_5837/gring pixel_5837/VDD pixel_5837/GND pixel_5837/VREF pixel_5837/ROW_SEL
+ pixel_5837/NB1 pixel_5837/VBIAS pixel_5837/NB2 pixel_5837/AMP_IN pixel_5837/SF_IB
+ pixel_5837/PIX_OUT pixel_5837/CSA_VREF pixel
Xpixel_5848 pixel_5848/gring pixel_5848/VDD pixel_5848/GND pixel_5848/VREF pixel_5848/ROW_SEL
+ pixel_5848/NB1 pixel_5848/VBIAS pixel_5848/NB2 pixel_5848/AMP_IN pixel_5848/SF_IB
+ pixel_5848/PIX_OUT pixel_5848/CSA_VREF pixel
Xpixel_5859 pixel_5859/gring pixel_5859/VDD pixel_5859/GND pixel_5859/VREF pixel_5859/ROW_SEL
+ pixel_5859/NB1 pixel_5859/VBIAS pixel_5859/NB2 pixel_5859/AMP_IN pixel_5859/SF_IB
+ pixel_5859/PIX_OUT pixel_5859/CSA_VREF pixel
Xpixel_9131 pixel_9131/gring pixel_9131/VDD pixel_9131/GND pixel_9131/VREF pixel_9131/ROW_SEL
+ pixel_9131/NB1 pixel_9131/VBIAS pixel_9131/NB2 pixel_9131/AMP_IN pixel_9131/SF_IB
+ pixel_9131/PIX_OUT pixel_9131/CSA_VREF pixel
Xpixel_9120 pixel_9120/gring pixel_9120/VDD pixel_9120/GND pixel_9120/VREF pixel_9120/ROW_SEL
+ pixel_9120/NB1 pixel_9120/VBIAS pixel_9120/NB2 pixel_9120/AMP_IN pixel_9120/SF_IB
+ pixel_9120/PIX_OUT pixel_9120/CSA_VREF pixel
Xpixel_9164 pixel_9164/gring pixel_9164/VDD pixel_9164/GND pixel_9164/VREF pixel_9164/ROW_SEL
+ pixel_9164/NB1 pixel_9164/VBIAS pixel_9164/NB2 pixel_9164/AMP_IN pixel_9164/SF_IB
+ pixel_9164/PIX_OUT pixel_9164/CSA_VREF pixel
Xpixel_9153 pixel_9153/gring pixel_9153/VDD pixel_9153/GND pixel_9153/VREF pixel_9153/ROW_SEL
+ pixel_9153/NB1 pixel_9153/VBIAS pixel_9153/NB2 pixel_9153/AMP_IN pixel_9153/SF_IB
+ pixel_9153/PIX_OUT pixel_9153/CSA_VREF pixel
Xpixel_9142 pixel_9142/gring pixel_9142/VDD pixel_9142/GND pixel_9142/VREF pixel_9142/ROW_SEL
+ pixel_9142/NB1 pixel_9142/VBIAS pixel_9142/NB2 pixel_9142/AMP_IN pixel_9142/SF_IB
+ pixel_9142/PIX_OUT pixel_9142/CSA_VREF pixel
Xpixel_8430 pixel_8430/gring pixel_8430/VDD pixel_8430/GND pixel_8430/VREF pixel_8430/ROW_SEL
+ pixel_8430/NB1 pixel_8430/VBIAS pixel_8430/NB2 pixel_8430/AMP_IN pixel_8430/SF_IB
+ pixel_8430/PIX_OUT pixel_8430/CSA_VREF pixel
Xpixel_9197 pixel_9197/gring pixel_9197/VDD pixel_9197/GND pixel_9197/VREF pixel_9197/ROW_SEL
+ pixel_9197/NB1 pixel_9197/VBIAS pixel_9197/NB2 pixel_9197/AMP_IN pixel_9197/SF_IB
+ pixel_9197/PIX_OUT pixel_9197/CSA_VREF pixel
Xpixel_9186 pixel_9186/gring pixel_9186/VDD pixel_9186/GND pixel_9186/VREF pixel_9186/ROW_SEL
+ pixel_9186/NB1 pixel_9186/VBIAS pixel_9186/NB2 pixel_9186/AMP_IN pixel_9186/SF_IB
+ pixel_9186/PIX_OUT pixel_9186/CSA_VREF pixel
Xpixel_9175 pixel_9175/gring pixel_9175/VDD pixel_9175/GND pixel_9175/VREF pixel_9175/ROW_SEL
+ pixel_9175/NB1 pixel_9175/VBIAS pixel_9175/NB2 pixel_9175/AMP_IN pixel_9175/SF_IB
+ pixel_9175/PIX_OUT pixel_9175/CSA_VREF pixel
Xpixel_8441 pixel_8441/gring pixel_8441/VDD pixel_8441/GND pixel_8441/VREF pixel_8441/ROW_SEL
+ pixel_8441/NB1 pixel_8441/VBIAS pixel_8441/NB2 pixel_8441/AMP_IN pixel_8441/SF_IB
+ pixel_8441/PIX_OUT pixel_8441/CSA_VREF pixel
Xpixel_8452 pixel_8452/gring pixel_8452/VDD pixel_8452/GND pixel_8452/VREF pixel_8452/ROW_SEL
+ pixel_8452/NB1 pixel_8452/VBIAS pixel_8452/NB2 pixel_8452/AMP_IN pixel_8452/SF_IB
+ pixel_8452/PIX_OUT pixel_8452/CSA_VREF pixel
Xpixel_8463 pixel_8463/gring pixel_8463/VDD pixel_8463/GND pixel_8463/VREF pixel_8463/ROW_SEL
+ pixel_8463/NB1 pixel_8463/VBIAS pixel_8463/NB2 pixel_8463/AMP_IN pixel_8463/SF_IB
+ pixel_8463/PIX_OUT pixel_8463/CSA_VREF pixel
Xpixel_8474 pixel_8474/gring pixel_8474/VDD pixel_8474/GND pixel_8474/VREF pixel_8474/ROW_SEL
+ pixel_8474/NB1 pixel_8474/VBIAS pixel_8474/NB2 pixel_8474/AMP_IN pixel_8474/SF_IB
+ pixel_8474/PIX_OUT pixel_8474/CSA_VREF pixel
Xpixel_8485 pixel_8485/gring pixel_8485/VDD pixel_8485/GND pixel_8485/VREF pixel_8485/ROW_SEL
+ pixel_8485/NB1 pixel_8485/VBIAS pixel_8485/NB2 pixel_8485/AMP_IN pixel_8485/SF_IB
+ pixel_8485/PIX_OUT pixel_8485/CSA_VREF pixel
Xpixel_8496 pixel_8496/gring pixel_8496/VDD pixel_8496/GND pixel_8496/VREF pixel_8496/ROW_SEL
+ pixel_8496/NB1 pixel_8496/VBIAS pixel_8496/NB2 pixel_8496/AMP_IN pixel_8496/SF_IB
+ pixel_8496/PIX_OUT pixel_8496/CSA_VREF pixel
Xpixel_7740 pixel_7740/gring pixel_7740/VDD pixel_7740/GND pixel_7740/VREF pixel_7740/ROW_SEL
+ pixel_7740/NB1 pixel_7740/VBIAS pixel_7740/NB2 pixel_7740/AMP_IN pixel_7740/SF_IB
+ pixel_7740/PIX_OUT pixel_7740/CSA_VREF pixel
Xpixel_7751 pixel_7751/gring pixel_7751/VDD pixel_7751/GND pixel_7751/VREF pixel_7751/ROW_SEL
+ pixel_7751/NB1 pixel_7751/VBIAS pixel_7751/NB2 pixel_7751/AMP_IN pixel_7751/SF_IB
+ pixel_7751/PIX_OUT pixel_7751/CSA_VREF pixel
Xpixel_7762 pixel_7762/gring pixel_7762/VDD pixel_7762/GND pixel_7762/VREF pixel_7762/ROW_SEL
+ pixel_7762/NB1 pixel_7762/VBIAS pixel_7762/NB2 pixel_7762/AMP_IN pixel_7762/SF_IB
+ pixel_7762/PIX_OUT pixel_7762/CSA_VREF pixel
Xpixel_7773 pixel_7773/gring pixel_7773/VDD pixel_7773/GND pixel_7773/VREF pixel_7773/ROW_SEL
+ pixel_7773/NB1 pixel_7773/VBIAS pixel_7773/NB2 pixel_7773/AMP_IN pixel_7773/SF_IB
+ pixel_7773/PIX_OUT pixel_7773/CSA_VREF pixel
Xpixel_7784 pixel_7784/gring pixel_7784/VDD pixel_7784/GND pixel_7784/VREF pixel_7784/ROW_SEL
+ pixel_7784/NB1 pixel_7784/VBIAS pixel_7784/NB2 pixel_7784/AMP_IN pixel_7784/SF_IB
+ pixel_7784/PIX_OUT pixel_7784/CSA_VREF pixel
Xpixel_7795 pixel_7795/gring pixel_7795/VDD pixel_7795/GND pixel_7795/VREF pixel_7795/ROW_SEL
+ pixel_7795/NB1 pixel_7795/VBIAS pixel_7795/NB2 pixel_7795/AMP_IN pixel_7795/SF_IB
+ pixel_7795/PIX_OUT pixel_7795/CSA_VREF pixel
Xpixel_2080 pixel_2080/gring pixel_2080/VDD pixel_2080/GND pixel_2080/VREF pixel_2080/ROW_SEL
+ pixel_2080/NB1 pixel_2080/VBIAS pixel_2080/NB2 pixel_2080/AMP_IN pixel_2080/SF_IB
+ pixel_2080/PIX_OUT pixel_2080/CSA_VREF pixel
Xpixel_2091 pixel_2091/gring pixel_2091/VDD pixel_2091/GND pixel_2091/VREF pixel_2091/ROW_SEL
+ pixel_2091/NB1 pixel_2091/VBIAS pixel_2091/NB2 pixel_2091/AMP_IN pixel_2091/SF_IB
+ pixel_2091/PIX_OUT pixel_2091/CSA_VREF pixel
Xpixel_1390 pixel_1390/gring pixel_1390/VDD pixel_1390/GND pixel_1390/VREF pixel_1390/ROW_SEL
+ pixel_1390/NB1 pixel_1390/VBIAS pixel_1390/NB2 pixel_1390/AMP_IN pixel_1390/SF_IB
+ pixel_1390/PIX_OUT pixel_1390/CSA_VREF pixel
Xpixel_405 pixel_405/gring pixel_405/VDD pixel_405/GND pixel_405/VREF pixel_405/ROW_SEL
+ pixel_405/NB1 pixel_405/VBIAS pixel_405/NB2 pixel_405/AMP_IN pixel_405/SF_IB pixel_405/PIX_OUT
+ pixel_405/CSA_VREF pixel
Xpixel_438 pixel_438/gring pixel_438/VDD pixel_438/GND pixel_438/VREF pixel_438/ROW_SEL
+ pixel_438/NB1 pixel_438/VBIAS pixel_438/NB2 pixel_438/AMP_IN pixel_438/SF_IB pixel_438/PIX_OUT
+ pixel_438/CSA_VREF pixel
Xpixel_427 pixel_427/gring pixel_427/VDD pixel_427/GND pixel_427/VREF pixel_427/ROW_SEL
+ pixel_427/NB1 pixel_427/VBIAS pixel_427/NB2 pixel_427/AMP_IN pixel_427/SF_IB pixel_427/PIX_OUT
+ pixel_427/CSA_VREF pixel
Xpixel_416 pixel_416/gring pixel_416/VDD pixel_416/GND pixel_416/VREF pixel_416/ROW_SEL
+ pixel_416/NB1 pixel_416/VBIAS pixel_416/NB2 pixel_416/AMP_IN pixel_416/SF_IB pixel_416/PIX_OUT
+ pixel_416/CSA_VREF pixel
Xpixel_449 pixel_449/gring pixel_449/VDD pixel_449/GND pixel_449/VREF pixel_449/ROW_SEL
+ pixel_449/NB1 pixel_449/VBIAS pixel_449/NB2 pixel_449/AMP_IN pixel_449/SF_IB pixel_449/PIX_OUT
+ pixel_449/CSA_VREF pixel
Xpixel_3709 pixel_3709/gring pixel_3709/VDD pixel_3709/GND pixel_3709/VREF pixel_3709/ROW_SEL
+ pixel_3709/NB1 pixel_3709/VBIAS pixel_3709/NB2 pixel_3709/AMP_IN pixel_3709/SF_IB
+ pixel_3709/PIX_OUT pixel_3709/CSA_VREF pixel
Xpixel_7003 pixel_7003/gring pixel_7003/VDD pixel_7003/GND pixel_7003/VREF pixel_7003/ROW_SEL
+ pixel_7003/NB1 pixel_7003/VBIAS pixel_7003/NB2 pixel_7003/AMP_IN pixel_7003/SF_IB
+ pixel_7003/PIX_OUT pixel_7003/CSA_VREF pixel
Xpixel_7014 pixel_7014/gring pixel_7014/VDD pixel_7014/GND pixel_7014/VREF pixel_7014/ROW_SEL
+ pixel_7014/NB1 pixel_7014/VBIAS pixel_7014/NB2 pixel_7014/AMP_IN pixel_7014/SF_IB
+ pixel_7014/PIX_OUT pixel_7014/CSA_VREF pixel
Xpixel_7025 pixel_7025/gring pixel_7025/VDD pixel_7025/GND pixel_7025/VREF pixel_7025/ROW_SEL
+ pixel_7025/NB1 pixel_7025/VBIAS pixel_7025/NB2 pixel_7025/AMP_IN pixel_7025/SF_IB
+ pixel_7025/PIX_OUT pixel_7025/CSA_VREF pixel
Xpixel_7036 pixel_7036/gring pixel_7036/VDD pixel_7036/GND pixel_7036/VREF pixel_7036/ROW_SEL
+ pixel_7036/NB1 pixel_7036/VBIAS pixel_7036/NB2 pixel_7036/AMP_IN pixel_7036/SF_IB
+ pixel_7036/PIX_OUT pixel_7036/CSA_VREF pixel
Xpixel_7047 pixel_7047/gring pixel_7047/VDD pixel_7047/GND pixel_7047/VREF pixel_7047/ROW_SEL
+ pixel_7047/NB1 pixel_7047/VBIAS pixel_7047/NB2 pixel_7047/AMP_IN pixel_7047/SF_IB
+ pixel_7047/PIX_OUT pixel_7047/CSA_VREF pixel
Xpixel_6302 pixel_6302/gring pixel_6302/VDD pixel_6302/GND pixel_6302/VREF pixel_6302/ROW_SEL
+ pixel_6302/NB1 pixel_6302/VBIAS pixel_6302/NB2 pixel_6302/AMP_IN pixel_6302/SF_IB
+ pixel_6302/PIX_OUT pixel_6302/CSA_VREF pixel
Xpixel_7058 pixel_7058/gring pixel_7058/VDD pixel_7058/GND pixel_7058/VREF pixel_7058/ROW_SEL
+ pixel_7058/NB1 pixel_7058/VBIAS pixel_7058/NB2 pixel_7058/AMP_IN pixel_7058/SF_IB
+ pixel_7058/PIX_OUT pixel_7058/CSA_VREF pixel
Xpixel_7069 pixel_7069/gring pixel_7069/VDD pixel_7069/GND pixel_7069/VREF pixel_7069/ROW_SEL
+ pixel_7069/NB1 pixel_7069/VBIAS pixel_7069/NB2 pixel_7069/AMP_IN pixel_7069/SF_IB
+ pixel_7069/PIX_OUT pixel_7069/CSA_VREF pixel
Xpixel_6313 pixel_6313/gring pixel_6313/VDD pixel_6313/GND pixel_6313/VREF pixel_6313/ROW_SEL
+ pixel_6313/NB1 pixel_6313/VBIAS pixel_6313/NB2 pixel_6313/AMP_IN pixel_6313/SF_IB
+ pixel_6313/PIX_OUT pixel_6313/CSA_VREF pixel
Xpixel_6324 pixel_6324/gring pixel_6324/VDD pixel_6324/GND pixel_6324/VREF pixel_6324/ROW_SEL
+ pixel_6324/NB1 pixel_6324/VBIAS pixel_6324/NB2 pixel_6324/AMP_IN pixel_6324/SF_IB
+ pixel_6324/PIX_OUT pixel_6324/CSA_VREF pixel
Xpixel_6335 pixel_6335/gring pixel_6335/VDD pixel_6335/GND pixel_6335/VREF pixel_6335/ROW_SEL
+ pixel_6335/NB1 pixel_6335/VBIAS pixel_6335/NB2 pixel_6335/AMP_IN pixel_6335/SF_IB
+ pixel_6335/PIX_OUT pixel_6335/CSA_VREF pixel
Xpixel_6346 pixel_6346/gring pixel_6346/VDD pixel_6346/GND pixel_6346/VREF pixel_6346/ROW_SEL
+ pixel_6346/NB1 pixel_6346/VBIAS pixel_6346/NB2 pixel_6346/AMP_IN pixel_6346/SF_IB
+ pixel_6346/PIX_OUT pixel_6346/CSA_VREF pixel
Xpixel_6357 pixel_6357/gring pixel_6357/VDD pixel_6357/GND pixel_6357/VREF pixel_6357/ROW_SEL
+ pixel_6357/NB1 pixel_6357/VBIAS pixel_6357/NB2 pixel_6357/AMP_IN pixel_6357/SF_IB
+ pixel_6357/PIX_OUT pixel_6357/CSA_VREF pixel
Xpixel_6368 pixel_6368/gring pixel_6368/VDD pixel_6368/GND pixel_6368/VREF pixel_6368/ROW_SEL
+ pixel_6368/NB1 pixel_6368/VBIAS pixel_6368/NB2 pixel_6368/AMP_IN pixel_6368/SF_IB
+ pixel_6368/PIX_OUT pixel_6368/CSA_VREF pixel
Xpixel_5601 pixel_5601/gring pixel_5601/VDD pixel_5601/GND pixel_5601/VREF pixel_5601/ROW_SEL
+ pixel_5601/NB1 pixel_5601/VBIAS pixel_5601/NB2 pixel_5601/AMP_IN pixel_5601/SF_IB
+ pixel_5601/PIX_OUT pixel_5601/CSA_VREF pixel
Xpixel_5612 pixel_5612/gring pixel_5612/VDD pixel_5612/GND pixel_5612/VREF pixel_5612/ROW_SEL
+ pixel_5612/NB1 pixel_5612/VBIAS pixel_5612/NB2 pixel_5612/AMP_IN pixel_5612/SF_IB
+ pixel_5612/PIX_OUT pixel_5612/CSA_VREF pixel
Xpixel_5623 pixel_5623/gring pixel_5623/VDD pixel_5623/GND pixel_5623/VREF pixel_5623/ROW_SEL
+ pixel_5623/NB1 pixel_5623/VBIAS pixel_5623/NB2 pixel_5623/AMP_IN pixel_5623/SF_IB
+ pixel_5623/PIX_OUT pixel_5623/CSA_VREF pixel
Xpixel_6379 pixel_6379/gring pixel_6379/VDD pixel_6379/GND pixel_6379/VREF pixel_6379/ROW_SEL
+ pixel_6379/NB1 pixel_6379/VBIAS pixel_6379/NB2 pixel_6379/AMP_IN pixel_6379/SF_IB
+ pixel_6379/PIX_OUT pixel_6379/CSA_VREF pixel
Xpixel_5634 pixel_5634/gring pixel_5634/VDD pixel_5634/GND pixel_5634/VREF pixel_5634/ROW_SEL
+ pixel_5634/NB1 pixel_5634/VBIAS pixel_5634/NB2 pixel_5634/AMP_IN pixel_5634/SF_IB
+ pixel_5634/PIX_OUT pixel_5634/CSA_VREF pixel
Xpixel_5645 pixel_5645/gring pixel_5645/VDD pixel_5645/GND pixel_5645/VREF pixel_5645/ROW_SEL
+ pixel_5645/NB1 pixel_5645/VBIAS pixel_5645/NB2 pixel_5645/AMP_IN pixel_5645/SF_IB
+ pixel_5645/PIX_OUT pixel_5645/CSA_VREF pixel
Xpixel_5656 pixel_5656/gring pixel_5656/VDD pixel_5656/GND pixel_5656/VREF pixel_5656/ROW_SEL
+ pixel_5656/NB1 pixel_5656/VBIAS pixel_5656/NB2 pixel_5656/AMP_IN pixel_5656/SF_IB
+ pixel_5656/PIX_OUT pixel_5656/CSA_VREF pixel
Xpixel_5667 pixel_5667/gring pixel_5667/VDD pixel_5667/GND pixel_5667/VREF pixel_5667/ROW_SEL
+ pixel_5667/NB1 pixel_5667/VBIAS pixel_5667/NB2 pixel_5667/AMP_IN pixel_5667/SF_IB
+ pixel_5667/PIX_OUT pixel_5667/CSA_VREF pixel
Xpixel_4900 pixel_4900/gring pixel_4900/VDD pixel_4900/GND pixel_4900/VREF pixel_4900/ROW_SEL
+ pixel_4900/NB1 pixel_4900/VBIAS pixel_4900/NB2 pixel_4900/AMP_IN pixel_4900/SF_IB
+ pixel_4900/PIX_OUT pixel_4900/CSA_VREF pixel
Xpixel_4911 pixel_4911/gring pixel_4911/VDD pixel_4911/GND pixel_4911/VREF pixel_4911/ROW_SEL
+ pixel_4911/NB1 pixel_4911/VBIAS pixel_4911/NB2 pixel_4911/AMP_IN pixel_4911/SF_IB
+ pixel_4911/PIX_OUT pixel_4911/CSA_VREF pixel
Xpixel_4922 pixel_4922/gring pixel_4922/VDD pixel_4922/GND pixel_4922/VREF pixel_4922/ROW_SEL
+ pixel_4922/NB1 pixel_4922/VBIAS pixel_4922/NB2 pixel_4922/AMP_IN pixel_4922/SF_IB
+ pixel_4922/PIX_OUT pixel_4922/CSA_VREF pixel
Xpixel_950 pixel_950/gring pixel_950/VDD pixel_950/GND pixel_950/VREF pixel_950/ROW_SEL
+ pixel_950/NB1 pixel_950/VBIAS pixel_950/NB2 pixel_950/AMP_IN pixel_950/SF_IB pixel_950/PIX_OUT
+ pixel_950/CSA_VREF pixel
Xpixel_5678 pixel_5678/gring pixel_5678/VDD pixel_5678/GND pixel_5678/VREF pixel_5678/ROW_SEL
+ pixel_5678/NB1 pixel_5678/VBIAS pixel_5678/NB2 pixel_5678/AMP_IN pixel_5678/SF_IB
+ pixel_5678/PIX_OUT pixel_5678/CSA_VREF pixel
Xpixel_5689 pixel_5689/gring pixel_5689/VDD pixel_5689/GND pixel_5689/VREF pixel_5689/ROW_SEL
+ pixel_5689/NB1 pixel_5689/VBIAS pixel_5689/NB2 pixel_5689/AMP_IN pixel_5689/SF_IB
+ pixel_5689/PIX_OUT pixel_5689/CSA_VREF pixel
Xpixel_4933 pixel_4933/gring pixel_4933/VDD pixel_4933/GND pixel_4933/VREF pixel_4933/ROW_SEL
+ pixel_4933/NB1 pixel_4933/VBIAS pixel_4933/NB2 pixel_4933/AMP_IN pixel_4933/SF_IB
+ pixel_4933/PIX_OUT pixel_4933/CSA_VREF pixel
Xpixel_4944 pixel_4944/gring pixel_4944/VDD pixel_4944/GND pixel_4944/VREF pixel_4944/ROW_SEL
+ pixel_4944/NB1 pixel_4944/VBIAS pixel_4944/NB2 pixel_4944/AMP_IN pixel_4944/SF_IB
+ pixel_4944/PIX_OUT pixel_4944/CSA_VREF pixel
Xpixel_4955 pixel_4955/gring pixel_4955/VDD pixel_4955/GND pixel_4955/VREF pixel_4955/ROW_SEL
+ pixel_4955/NB1 pixel_4955/VBIAS pixel_4955/NB2 pixel_4955/AMP_IN pixel_4955/SF_IB
+ pixel_4955/PIX_OUT pixel_4955/CSA_VREF pixel
Xpixel_994 pixel_994/gring pixel_994/VDD pixel_994/GND pixel_994/VREF pixel_994/ROW_SEL
+ pixel_994/NB1 pixel_994/VBIAS pixel_994/NB2 pixel_994/AMP_IN pixel_994/SF_IB pixel_994/PIX_OUT
+ pixel_994/CSA_VREF pixel
Xpixel_983 pixel_983/gring pixel_983/VDD pixel_983/GND pixel_983/VREF pixel_983/ROW_SEL
+ pixel_983/NB1 pixel_983/VBIAS pixel_983/NB2 pixel_983/AMP_IN pixel_983/SF_IB pixel_983/PIX_OUT
+ pixel_983/CSA_VREF pixel
Xpixel_972 pixel_972/gring pixel_972/VDD pixel_972/GND pixel_972/VREF pixel_972/ROW_SEL
+ pixel_972/NB1 pixel_972/VBIAS pixel_972/NB2 pixel_972/AMP_IN pixel_972/SF_IB pixel_972/PIX_OUT
+ pixel_972/CSA_VREF pixel
Xpixel_961 pixel_961/gring pixel_961/VDD pixel_961/GND pixel_961/VREF pixel_961/ROW_SEL
+ pixel_961/NB1 pixel_961/VBIAS pixel_961/NB2 pixel_961/AMP_IN pixel_961/SF_IB pixel_961/PIX_OUT
+ pixel_961/CSA_VREF pixel
Xpixel_4966 pixel_4966/gring pixel_4966/VDD pixel_4966/GND pixel_4966/VREF pixel_4966/ROW_SEL
+ pixel_4966/NB1 pixel_4966/VBIAS pixel_4966/NB2 pixel_4966/AMP_IN pixel_4966/SF_IB
+ pixel_4966/PIX_OUT pixel_4966/CSA_VREF pixel
Xpixel_4977 pixel_4977/gring pixel_4977/VDD pixel_4977/GND pixel_4977/VREF pixel_4977/ROW_SEL
+ pixel_4977/NB1 pixel_4977/VBIAS pixel_4977/NB2 pixel_4977/AMP_IN pixel_4977/SF_IB
+ pixel_4977/PIX_OUT pixel_4977/CSA_VREF pixel
Xpixel_4988 pixel_4988/gring pixel_4988/VDD pixel_4988/GND pixel_4988/VREF pixel_4988/ROW_SEL
+ pixel_4988/NB1 pixel_4988/VBIAS pixel_4988/NB2 pixel_4988/AMP_IN pixel_4988/SF_IB
+ pixel_4988/PIX_OUT pixel_4988/CSA_VREF pixel
Xpixel_4999 pixel_4999/gring pixel_4999/VDD pixel_4999/GND pixel_4999/VREF pixel_4999/ROW_SEL
+ pixel_4999/NB1 pixel_4999/VBIAS pixel_4999/NB2 pixel_4999/AMP_IN pixel_4999/SF_IB
+ pixel_4999/PIX_OUT pixel_4999/CSA_VREF pixel
Xpixel_8260 pixel_8260/gring pixel_8260/VDD pixel_8260/GND pixel_8260/VREF pixel_8260/ROW_SEL
+ pixel_8260/NB1 pixel_8260/VBIAS pixel_8260/NB2 pixel_8260/AMP_IN pixel_8260/SF_IB
+ pixel_8260/PIX_OUT pixel_8260/CSA_VREF pixel
Xpixel_8271 pixel_8271/gring pixel_8271/VDD pixel_8271/GND pixel_8271/VREF pixel_8271/ROW_SEL
+ pixel_8271/NB1 pixel_8271/VBIAS pixel_8271/NB2 pixel_8271/AMP_IN pixel_8271/SF_IB
+ pixel_8271/PIX_OUT pixel_8271/CSA_VREF pixel
Xpixel_8282 pixel_8282/gring pixel_8282/VDD pixel_8282/GND pixel_8282/VREF pixel_8282/ROW_SEL
+ pixel_8282/NB1 pixel_8282/VBIAS pixel_8282/NB2 pixel_8282/AMP_IN pixel_8282/SF_IB
+ pixel_8282/PIX_OUT pixel_8282/CSA_VREF pixel
Xpixel_8293 pixel_8293/gring pixel_8293/VDD pixel_8293/GND pixel_8293/VREF pixel_8293/ROW_SEL
+ pixel_8293/NB1 pixel_8293/VBIAS pixel_8293/NB2 pixel_8293/AMP_IN pixel_8293/SF_IB
+ pixel_8293/PIX_OUT pixel_8293/CSA_VREF pixel
Xpixel_7570 pixel_7570/gring pixel_7570/VDD pixel_7570/GND pixel_7570/VREF pixel_7570/ROW_SEL
+ pixel_7570/NB1 pixel_7570/VBIAS pixel_7570/NB2 pixel_7570/AMP_IN pixel_7570/SF_IB
+ pixel_7570/PIX_OUT pixel_7570/CSA_VREF pixel
Xpixel_7581 pixel_7581/gring pixel_7581/VDD pixel_7581/GND pixel_7581/VREF pixel_7581/ROW_SEL
+ pixel_7581/NB1 pixel_7581/VBIAS pixel_7581/NB2 pixel_7581/AMP_IN pixel_7581/SF_IB
+ pixel_7581/PIX_OUT pixel_7581/CSA_VREF pixel
Xpixel_7592 pixel_7592/gring pixel_7592/VDD pixel_7592/GND pixel_7592/VREF pixel_7592/ROW_SEL
+ pixel_7592/NB1 pixel_7592/VBIAS pixel_7592/NB2 pixel_7592/AMP_IN pixel_7592/SF_IB
+ pixel_7592/PIX_OUT pixel_7592/CSA_VREF pixel
Xpixel_6880 pixel_6880/gring pixel_6880/VDD pixel_6880/GND pixel_6880/VREF pixel_6880/ROW_SEL
+ pixel_6880/NB1 pixel_6880/VBIAS pixel_6880/NB2 pixel_6880/AMP_IN pixel_6880/SF_IB
+ pixel_6880/PIX_OUT pixel_6880/CSA_VREF pixel
Xpixel_6891 pixel_6891/gring pixel_6891/VDD pixel_6891/GND pixel_6891/VREF pixel_6891/ROW_SEL
+ pixel_6891/NB1 pixel_6891/VBIAS pixel_6891/NB2 pixel_6891/AMP_IN pixel_6891/SF_IB
+ pixel_6891/PIX_OUT pixel_6891/CSA_VREF pixel
Xpixel_213 pixel_213/gring pixel_213/VDD pixel_213/GND pixel_213/VREF pixel_213/ROW_SEL
+ pixel_213/NB1 pixel_213/VBIAS pixel_213/NB2 pixel_213/AMP_IN pixel_213/SF_IB pixel_213/PIX_OUT
+ pixel_213/CSA_VREF pixel
Xpixel_202 pixel_202/gring pixel_202/VDD pixel_202/GND pixel_202/VREF pixel_202/ROW_SEL
+ pixel_202/NB1 pixel_202/VBIAS pixel_202/NB2 pixel_202/AMP_IN pixel_202/SF_IB pixel_202/PIX_OUT
+ pixel_202/CSA_VREF pixel
Xpixel_4207 pixel_4207/gring pixel_4207/VDD pixel_4207/GND pixel_4207/VREF pixel_4207/ROW_SEL
+ pixel_4207/NB1 pixel_4207/VBIAS pixel_4207/NB2 pixel_4207/AMP_IN pixel_4207/SF_IB
+ pixel_4207/PIX_OUT pixel_4207/CSA_VREF pixel
Xpixel_4218 pixel_4218/gring pixel_4218/VDD pixel_4218/GND pixel_4218/VREF pixel_4218/ROW_SEL
+ pixel_4218/NB1 pixel_4218/VBIAS pixel_4218/NB2 pixel_4218/AMP_IN pixel_4218/SF_IB
+ pixel_4218/PIX_OUT pixel_4218/CSA_VREF pixel
Xpixel_246 pixel_246/gring pixel_246/VDD pixel_246/GND pixel_246/VREF pixel_246/ROW_SEL
+ pixel_246/NB1 pixel_246/VBIAS pixel_246/NB2 pixel_246/AMP_IN pixel_246/SF_IB pixel_246/PIX_OUT
+ pixel_246/CSA_VREF pixel
Xpixel_235 pixel_235/gring pixel_235/VDD pixel_235/GND pixel_235/VREF pixel_235/ROW_SEL
+ pixel_235/NB1 pixel_235/VBIAS pixel_235/NB2 pixel_235/AMP_IN pixel_235/SF_IB pixel_235/PIX_OUT
+ pixel_235/CSA_VREF pixel
Xpixel_224 pixel_224/gring pixel_224/VDD pixel_224/GND pixel_224/VREF pixel_224/ROW_SEL
+ pixel_224/NB1 pixel_224/VBIAS pixel_224/NB2 pixel_224/AMP_IN pixel_224/SF_IB pixel_224/PIX_OUT
+ pixel_224/CSA_VREF pixel
Xpixel_3506 pixel_3506/gring pixel_3506/VDD pixel_3506/GND pixel_3506/VREF pixel_3506/ROW_SEL
+ pixel_3506/NB1 pixel_3506/VBIAS pixel_3506/NB2 pixel_3506/AMP_IN pixel_3506/SF_IB
+ pixel_3506/PIX_OUT pixel_3506/CSA_VREF pixel
Xpixel_4229 pixel_4229/gring pixel_4229/VDD pixel_4229/GND pixel_4229/VREF pixel_4229/ROW_SEL
+ pixel_4229/NB1 pixel_4229/VBIAS pixel_4229/NB2 pixel_4229/AMP_IN pixel_4229/SF_IB
+ pixel_4229/PIX_OUT pixel_4229/CSA_VREF pixel
Xpixel_279 pixel_279/gring pixel_279/VDD pixel_279/GND pixel_279/VREF pixel_279/ROW_SEL
+ pixel_279/NB1 pixel_279/VBIAS pixel_279/NB2 pixel_279/AMP_IN pixel_279/SF_IB pixel_279/PIX_OUT
+ pixel_279/CSA_VREF pixel
Xpixel_268 pixel_268/gring pixel_268/VDD pixel_268/GND pixel_268/VREF pixel_268/ROW_SEL
+ pixel_268/NB1 pixel_268/VBIAS pixel_268/NB2 pixel_268/AMP_IN pixel_268/SF_IB pixel_268/PIX_OUT
+ pixel_268/CSA_VREF pixel
Xpixel_257 pixel_257/gring pixel_257/VDD pixel_257/GND pixel_257/VREF pixel_257/ROW_SEL
+ pixel_257/NB1 pixel_257/VBIAS pixel_257/NB2 pixel_257/AMP_IN pixel_257/SF_IB pixel_257/PIX_OUT
+ pixel_257/CSA_VREF pixel
Xpixel_3539 pixel_3539/gring pixel_3539/VDD pixel_3539/GND pixel_3539/VREF pixel_3539/ROW_SEL
+ pixel_3539/NB1 pixel_3539/VBIAS pixel_3539/NB2 pixel_3539/AMP_IN pixel_3539/SF_IB
+ pixel_3539/PIX_OUT pixel_3539/CSA_VREF pixel
Xpixel_3528 pixel_3528/gring pixel_3528/VDD pixel_3528/GND pixel_3528/VREF pixel_3528/ROW_SEL
+ pixel_3528/NB1 pixel_3528/VBIAS pixel_3528/NB2 pixel_3528/AMP_IN pixel_3528/SF_IB
+ pixel_3528/PIX_OUT pixel_3528/CSA_VREF pixel
Xpixel_3517 pixel_3517/gring pixel_3517/VDD pixel_3517/GND pixel_3517/VREF pixel_3517/ROW_SEL
+ pixel_3517/NB1 pixel_3517/VBIAS pixel_3517/NB2 pixel_3517/AMP_IN pixel_3517/SF_IB
+ pixel_3517/PIX_OUT pixel_3517/CSA_VREF pixel
Xpixel_2838 pixel_2838/gring pixel_2838/VDD pixel_2838/GND pixel_2838/VREF pixel_2838/ROW_SEL
+ pixel_2838/NB1 pixel_2838/VBIAS pixel_2838/NB2 pixel_2838/AMP_IN pixel_2838/SF_IB
+ pixel_2838/PIX_OUT pixel_2838/CSA_VREF pixel
Xpixel_2827 pixel_2827/gring pixel_2827/VDD pixel_2827/GND pixel_2827/VREF pixel_2827/ROW_SEL
+ pixel_2827/NB1 pixel_2827/VBIAS pixel_2827/NB2 pixel_2827/AMP_IN pixel_2827/SF_IB
+ pixel_2827/PIX_OUT pixel_2827/CSA_VREF pixel
Xpixel_2816 pixel_2816/gring pixel_2816/VDD pixel_2816/GND pixel_2816/VREF pixel_2816/ROW_SEL
+ pixel_2816/NB1 pixel_2816/VBIAS pixel_2816/NB2 pixel_2816/AMP_IN pixel_2816/SF_IB
+ pixel_2816/PIX_OUT pixel_2816/CSA_VREF pixel
Xpixel_2805 pixel_2805/gring pixel_2805/VDD pixel_2805/GND pixel_2805/VREF pixel_2805/ROW_SEL
+ pixel_2805/NB1 pixel_2805/VBIAS pixel_2805/NB2 pixel_2805/AMP_IN pixel_2805/SF_IB
+ pixel_2805/PIX_OUT pixel_2805/CSA_VREF pixel
Xpixel_2849 pixel_2849/gring pixel_2849/VDD pixel_2849/GND pixel_2849/VREF pixel_2849/ROW_SEL
+ pixel_2849/NB1 pixel_2849/VBIAS pixel_2849/NB2 pixel_2849/AMP_IN pixel_2849/SF_IB
+ pixel_2849/PIX_OUT pixel_2849/CSA_VREF pixel
Xpixel_6110 pixel_6110/gring pixel_6110/VDD pixel_6110/GND pixel_6110/VREF pixel_6110/ROW_SEL
+ pixel_6110/NB1 pixel_6110/VBIAS pixel_6110/NB2 pixel_6110/AMP_IN pixel_6110/SF_IB
+ pixel_6110/PIX_OUT pixel_6110/CSA_VREF pixel
Xpixel_6121 pixel_6121/gring pixel_6121/VDD pixel_6121/GND pixel_6121/VREF pixel_6121/ROW_SEL
+ pixel_6121/NB1 pixel_6121/VBIAS pixel_6121/NB2 pixel_6121/AMP_IN pixel_6121/SF_IB
+ pixel_6121/PIX_OUT pixel_6121/CSA_VREF pixel
Xpixel_6132 pixel_6132/gring pixel_6132/VDD pixel_6132/GND pixel_6132/VREF pixel_6132/ROW_SEL
+ pixel_6132/NB1 pixel_6132/VBIAS pixel_6132/NB2 pixel_6132/AMP_IN pixel_6132/SF_IB
+ pixel_6132/PIX_OUT pixel_6132/CSA_VREF pixel
Xpixel_6143 pixel_6143/gring pixel_6143/VDD pixel_6143/GND pixel_6143/VREF pixel_6143/ROW_SEL
+ pixel_6143/NB1 pixel_6143/VBIAS pixel_6143/NB2 pixel_6143/AMP_IN pixel_6143/SF_IB
+ pixel_6143/PIX_OUT pixel_6143/CSA_VREF pixel
Xpixel_6154 pixel_6154/gring pixel_6154/VDD pixel_6154/GND pixel_6154/VREF pixel_6154/ROW_SEL
+ pixel_6154/NB1 pixel_6154/VBIAS pixel_6154/NB2 pixel_6154/AMP_IN pixel_6154/SF_IB
+ pixel_6154/PIX_OUT pixel_6154/CSA_VREF pixel
Xpixel_6165 pixel_6165/gring pixel_6165/VDD pixel_6165/GND pixel_6165/VREF pixel_6165/ROW_SEL
+ pixel_6165/NB1 pixel_6165/VBIAS pixel_6165/NB2 pixel_6165/AMP_IN pixel_6165/SF_IB
+ pixel_6165/PIX_OUT pixel_6165/CSA_VREF pixel
Xpixel_6176 pixel_6176/gring pixel_6176/VDD pixel_6176/GND pixel_6176/VREF pixel_6176/ROW_SEL
+ pixel_6176/NB1 pixel_6176/VBIAS pixel_6176/NB2 pixel_6176/AMP_IN pixel_6176/SF_IB
+ pixel_6176/PIX_OUT pixel_6176/CSA_VREF pixel
Xpixel_6187 pixel_6187/gring pixel_6187/VDD pixel_6187/GND pixel_6187/VREF pixel_6187/ROW_SEL
+ pixel_6187/NB1 pixel_6187/VBIAS pixel_6187/NB2 pixel_6187/AMP_IN pixel_6187/SF_IB
+ pixel_6187/PIX_OUT pixel_6187/CSA_VREF pixel
Xpixel_5420 pixel_5420/gring pixel_5420/VDD pixel_5420/GND pixel_5420/VREF pixel_5420/ROW_SEL
+ pixel_5420/NB1 pixel_5420/VBIAS pixel_5420/NB2 pixel_5420/AMP_IN pixel_5420/SF_IB
+ pixel_5420/PIX_OUT pixel_5420/CSA_VREF pixel
Xpixel_5431 pixel_5431/gring pixel_5431/VDD pixel_5431/GND pixel_5431/VREF pixel_5431/ROW_SEL
+ pixel_5431/NB1 pixel_5431/VBIAS pixel_5431/NB2 pixel_5431/AMP_IN pixel_5431/SF_IB
+ pixel_5431/PIX_OUT pixel_5431/CSA_VREF pixel
Xpixel_5442 pixel_5442/gring pixel_5442/VDD pixel_5442/GND pixel_5442/VREF pixel_5442/ROW_SEL
+ pixel_5442/NB1 pixel_5442/VBIAS pixel_5442/NB2 pixel_5442/AMP_IN pixel_5442/SF_IB
+ pixel_5442/PIX_OUT pixel_5442/CSA_VREF pixel
Xpixel_6198 pixel_6198/gring pixel_6198/VDD pixel_6198/GND pixel_6198/VREF pixel_6198/ROW_SEL
+ pixel_6198/NB1 pixel_6198/VBIAS pixel_6198/NB2 pixel_6198/AMP_IN pixel_6198/SF_IB
+ pixel_6198/PIX_OUT pixel_6198/CSA_VREF pixel
Xpixel_5453 pixel_5453/gring pixel_5453/VDD pixel_5453/GND pixel_5453/VREF pixel_5453/ROW_SEL
+ pixel_5453/NB1 pixel_5453/VBIAS pixel_5453/NB2 pixel_5453/AMP_IN pixel_5453/SF_IB
+ pixel_5453/PIX_OUT pixel_5453/CSA_VREF pixel
Xpixel_5464 pixel_5464/gring pixel_5464/VDD pixel_5464/GND pixel_5464/VREF pixel_5464/ROW_SEL
+ pixel_5464/NB1 pixel_5464/VBIAS pixel_5464/NB2 pixel_5464/AMP_IN pixel_5464/SF_IB
+ pixel_5464/PIX_OUT pixel_5464/CSA_VREF pixel
Xpixel_5475 pixel_5475/gring pixel_5475/VDD pixel_5475/GND pixel_5475/VREF pixel_5475/ROW_SEL
+ pixel_5475/NB1 pixel_5475/VBIAS pixel_5475/NB2 pixel_5475/AMP_IN pixel_5475/SF_IB
+ pixel_5475/PIX_OUT pixel_5475/CSA_VREF pixel
Xpixel_4730 pixel_4730/gring pixel_4730/VDD pixel_4730/GND pixel_4730/VREF pixel_4730/ROW_SEL
+ pixel_4730/NB1 pixel_4730/VBIAS pixel_4730/NB2 pixel_4730/AMP_IN pixel_4730/SF_IB
+ pixel_4730/PIX_OUT pixel_4730/CSA_VREF pixel
Xpixel_5486 pixel_5486/gring pixel_5486/VDD pixel_5486/GND pixel_5486/VREF pixel_5486/ROW_SEL
+ pixel_5486/NB1 pixel_5486/VBIAS pixel_5486/NB2 pixel_5486/AMP_IN pixel_5486/SF_IB
+ pixel_5486/PIX_OUT pixel_5486/CSA_VREF pixel
Xpixel_5497 pixel_5497/gring pixel_5497/VDD pixel_5497/GND pixel_5497/VREF pixel_5497/ROW_SEL
+ pixel_5497/NB1 pixel_5497/VBIAS pixel_5497/NB2 pixel_5497/AMP_IN pixel_5497/SF_IB
+ pixel_5497/PIX_OUT pixel_5497/CSA_VREF pixel
Xpixel_4741 pixel_4741/gring pixel_4741/VDD pixel_4741/GND pixel_4741/VREF pixel_4741/ROW_SEL
+ pixel_4741/NB1 pixel_4741/VBIAS pixel_4741/NB2 pixel_4741/AMP_IN pixel_4741/SF_IB
+ pixel_4741/PIX_OUT pixel_4741/CSA_VREF pixel
Xpixel_4752 pixel_4752/gring pixel_4752/VDD pixel_4752/GND pixel_4752/VREF pixel_4752/ROW_SEL
+ pixel_4752/NB1 pixel_4752/VBIAS pixel_4752/NB2 pixel_4752/AMP_IN pixel_4752/SF_IB
+ pixel_4752/PIX_OUT pixel_4752/CSA_VREF pixel
Xpixel_4763 pixel_4763/gring pixel_4763/VDD pixel_4763/GND pixel_4763/VREF pixel_4763/ROW_SEL
+ pixel_4763/NB1 pixel_4763/VBIAS pixel_4763/NB2 pixel_4763/AMP_IN pixel_4763/SF_IB
+ pixel_4763/PIX_OUT pixel_4763/CSA_VREF pixel
Xpixel_791 pixel_791/gring pixel_791/VDD pixel_791/GND pixel_791/VREF pixel_791/ROW_SEL
+ pixel_791/NB1 pixel_791/VBIAS pixel_791/NB2 pixel_791/AMP_IN pixel_791/SF_IB pixel_791/PIX_OUT
+ pixel_791/CSA_VREF pixel
Xpixel_780 pixel_780/gring pixel_780/VDD pixel_780/GND pixel_780/VREF pixel_780/ROW_SEL
+ pixel_780/NB1 pixel_780/VBIAS pixel_780/NB2 pixel_780/AMP_IN pixel_780/SF_IB pixel_780/PIX_OUT
+ pixel_780/CSA_VREF pixel
Xpixel_4774 pixel_4774/gring pixel_4774/VDD pixel_4774/GND pixel_4774/VREF pixel_4774/ROW_SEL
+ pixel_4774/NB1 pixel_4774/VBIAS pixel_4774/NB2 pixel_4774/AMP_IN pixel_4774/SF_IB
+ pixel_4774/PIX_OUT pixel_4774/CSA_VREF pixel
Xpixel_4785 pixel_4785/gring pixel_4785/VDD pixel_4785/GND pixel_4785/VREF pixel_4785/ROW_SEL
+ pixel_4785/NB1 pixel_4785/VBIAS pixel_4785/NB2 pixel_4785/AMP_IN pixel_4785/SF_IB
+ pixel_4785/PIX_OUT pixel_4785/CSA_VREF pixel
Xpixel_4796 pixel_4796/gring pixel_4796/VDD pixel_4796/GND pixel_4796/VREF pixel_4796/ROW_SEL
+ pixel_4796/NB1 pixel_4796/VBIAS pixel_4796/NB2 pixel_4796/AMP_IN pixel_4796/SF_IB
+ pixel_4796/PIX_OUT pixel_4796/CSA_VREF pixel
Xpixel_8090 pixel_8090/gring pixel_8090/VDD pixel_8090/GND pixel_8090/VREF pixel_8090/ROW_SEL
+ pixel_8090/NB1 pixel_8090/VBIAS pixel_8090/NB2 pixel_8090/AMP_IN pixel_8090/SF_IB
+ pixel_8090/PIX_OUT pixel_8090/CSA_VREF pixel
Xpixel_9708 pixel_9708/gring pixel_9708/VDD pixel_9708/GND pixel_9708/VREF pixel_9708/ROW_SEL
+ pixel_9708/NB1 pixel_9708/VBIAS pixel_9708/NB2 pixel_9708/AMP_IN pixel_9708/SF_IB
+ pixel_9708/PIX_OUT pixel_9708/CSA_VREF pixel
Xpixel_9719 pixel_9719/gring pixel_9719/VDD pixel_9719/GND pixel_9719/VREF pixel_9719/ROW_SEL
+ pixel_9719/NB1 pixel_9719/VBIAS pixel_9719/NB2 pixel_9719/AMP_IN pixel_9719/SF_IB
+ pixel_9719/PIX_OUT pixel_9719/CSA_VREF pixel
Xpixel_4004 pixel_4004/gring pixel_4004/VDD pixel_4004/GND pixel_4004/VREF pixel_4004/ROW_SEL
+ pixel_4004/NB1 pixel_4004/VBIAS pixel_4004/NB2 pixel_4004/AMP_IN pixel_4004/SF_IB
+ pixel_4004/PIX_OUT pixel_4004/CSA_VREF pixel
Xpixel_4015 pixel_4015/gring pixel_4015/VDD pixel_4015/GND pixel_4015/VREF pixel_4015/ROW_SEL
+ pixel_4015/NB1 pixel_4015/VBIAS pixel_4015/NB2 pixel_4015/AMP_IN pixel_4015/SF_IB
+ pixel_4015/PIX_OUT pixel_4015/CSA_VREF pixel
Xpixel_4026 pixel_4026/gring pixel_4026/VDD pixel_4026/GND pixel_4026/VREF pixel_4026/ROW_SEL
+ pixel_4026/NB1 pixel_4026/VBIAS pixel_4026/NB2 pixel_4026/AMP_IN pixel_4026/SF_IB
+ pixel_4026/PIX_OUT pixel_4026/CSA_VREF pixel
Xpixel_3314 pixel_3314/gring pixel_3314/VDD pixel_3314/GND pixel_3314/VREF pixel_3314/ROW_SEL
+ pixel_3314/NB1 pixel_3314/VBIAS pixel_3314/NB2 pixel_3314/AMP_IN pixel_3314/SF_IB
+ pixel_3314/PIX_OUT pixel_3314/CSA_VREF pixel
Xpixel_3303 pixel_3303/gring pixel_3303/VDD pixel_3303/GND pixel_3303/VREF pixel_3303/ROW_SEL
+ pixel_3303/NB1 pixel_3303/VBIAS pixel_3303/NB2 pixel_3303/AMP_IN pixel_3303/SF_IB
+ pixel_3303/PIX_OUT pixel_3303/CSA_VREF pixel
Xpixel_4037 pixel_4037/gring pixel_4037/VDD pixel_4037/GND pixel_4037/VREF pixel_4037/ROW_SEL
+ pixel_4037/NB1 pixel_4037/VBIAS pixel_4037/NB2 pixel_4037/AMP_IN pixel_4037/SF_IB
+ pixel_4037/PIX_OUT pixel_4037/CSA_VREF pixel
Xpixel_4048 pixel_4048/gring pixel_4048/VDD pixel_4048/GND pixel_4048/VREF pixel_4048/ROW_SEL
+ pixel_4048/NB1 pixel_4048/VBIAS pixel_4048/NB2 pixel_4048/AMP_IN pixel_4048/SF_IB
+ pixel_4048/PIX_OUT pixel_4048/CSA_VREF pixel
Xpixel_4059 pixel_4059/gring pixel_4059/VDD pixel_4059/GND pixel_4059/VREF pixel_4059/ROW_SEL
+ pixel_4059/NB1 pixel_4059/VBIAS pixel_4059/NB2 pixel_4059/AMP_IN pixel_4059/SF_IB
+ pixel_4059/PIX_OUT pixel_4059/CSA_VREF pixel
Xpixel_2613 pixel_2613/gring pixel_2613/VDD pixel_2613/GND pixel_2613/VREF pixel_2613/ROW_SEL
+ pixel_2613/NB1 pixel_2613/VBIAS pixel_2613/NB2 pixel_2613/AMP_IN pixel_2613/SF_IB
+ pixel_2613/PIX_OUT pixel_2613/CSA_VREF pixel
Xpixel_2602 pixel_2602/gring pixel_2602/VDD pixel_2602/GND pixel_2602/VREF pixel_2602/ROW_SEL
+ pixel_2602/NB1 pixel_2602/VBIAS pixel_2602/NB2 pixel_2602/AMP_IN pixel_2602/SF_IB
+ pixel_2602/PIX_OUT pixel_2602/CSA_VREF pixel
Xpixel_3358 pixel_3358/gring pixel_3358/VDD pixel_3358/GND pixel_3358/VREF pixel_3358/ROW_SEL
+ pixel_3358/NB1 pixel_3358/VBIAS pixel_3358/NB2 pixel_3358/AMP_IN pixel_3358/SF_IB
+ pixel_3358/PIX_OUT pixel_3358/CSA_VREF pixel
Xpixel_3347 pixel_3347/gring pixel_3347/VDD pixel_3347/GND pixel_3347/VREF pixel_3347/ROW_SEL
+ pixel_3347/NB1 pixel_3347/VBIAS pixel_3347/NB2 pixel_3347/AMP_IN pixel_3347/SF_IB
+ pixel_3347/PIX_OUT pixel_3347/CSA_VREF pixel
Xpixel_3336 pixel_3336/gring pixel_3336/VDD pixel_3336/GND pixel_3336/VREF pixel_3336/ROW_SEL
+ pixel_3336/NB1 pixel_3336/VBIAS pixel_3336/NB2 pixel_3336/AMP_IN pixel_3336/SF_IB
+ pixel_3336/PIX_OUT pixel_3336/CSA_VREF pixel
Xpixel_3325 pixel_3325/gring pixel_3325/VDD pixel_3325/GND pixel_3325/VREF pixel_3325/ROW_SEL
+ pixel_3325/NB1 pixel_3325/VBIAS pixel_3325/NB2 pixel_3325/AMP_IN pixel_3325/SF_IB
+ pixel_3325/PIX_OUT pixel_3325/CSA_VREF pixel
Xpixel_1901 pixel_1901/gring pixel_1901/VDD pixel_1901/GND pixel_1901/VREF pixel_1901/ROW_SEL
+ pixel_1901/NB1 pixel_1901/VBIAS pixel_1901/NB2 pixel_1901/AMP_IN pixel_1901/SF_IB
+ pixel_1901/PIX_OUT pixel_1901/CSA_VREF pixel
Xpixel_2646 pixel_2646/gring pixel_2646/VDD pixel_2646/GND pixel_2646/VREF pixel_2646/ROW_SEL
+ pixel_2646/NB1 pixel_2646/VBIAS pixel_2646/NB2 pixel_2646/AMP_IN pixel_2646/SF_IB
+ pixel_2646/PIX_OUT pixel_2646/CSA_VREF pixel
Xpixel_2635 pixel_2635/gring pixel_2635/VDD pixel_2635/GND pixel_2635/VREF pixel_2635/ROW_SEL
+ pixel_2635/NB1 pixel_2635/VBIAS pixel_2635/NB2 pixel_2635/AMP_IN pixel_2635/SF_IB
+ pixel_2635/PIX_OUT pixel_2635/CSA_VREF pixel
Xpixel_2624 pixel_2624/gring pixel_2624/VDD pixel_2624/GND pixel_2624/VREF pixel_2624/ROW_SEL
+ pixel_2624/NB1 pixel_2624/VBIAS pixel_2624/NB2 pixel_2624/AMP_IN pixel_2624/SF_IB
+ pixel_2624/PIX_OUT pixel_2624/CSA_VREF pixel
Xpixel_3369 pixel_3369/gring pixel_3369/VDD pixel_3369/GND pixel_3369/VREF pixel_3369/ROW_SEL
+ pixel_3369/NB1 pixel_3369/VBIAS pixel_3369/NB2 pixel_3369/AMP_IN pixel_3369/SF_IB
+ pixel_3369/PIX_OUT pixel_3369/CSA_VREF pixel
Xpixel_1934 pixel_1934/gring pixel_1934/VDD pixel_1934/GND pixel_1934/VREF pixel_1934/ROW_SEL
+ pixel_1934/NB1 pixel_1934/VBIAS pixel_1934/NB2 pixel_1934/AMP_IN pixel_1934/SF_IB
+ pixel_1934/PIX_OUT pixel_1934/CSA_VREF pixel
Xpixel_1923 pixel_1923/gring pixel_1923/VDD pixel_1923/GND pixel_1923/VREF pixel_1923/ROW_SEL
+ pixel_1923/NB1 pixel_1923/VBIAS pixel_1923/NB2 pixel_1923/AMP_IN pixel_1923/SF_IB
+ pixel_1923/PIX_OUT pixel_1923/CSA_VREF pixel
Xpixel_1912 pixel_1912/gring pixel_1912/VDD pixel_1912/GND pixel_1912/VREF pixel_1912/ROW_SEL
+ pixel_1912/NB1 pixel_1912/VBIAS pixel_1912/NB2 pixel_1912/AMP_IN pixel_1912/SF_IB
+ pixel_1912/PIX_OUT pixel_1912/CSA_VREF pixel
Xpixel_2679 pixel_2679/gring pixel_2679/VDD pixel_2679/GND pixel_2679/VREF pixel_2679/ROW_SEL
+ pixel_2679/NB1 pixel_2679/VBIAS pixel_2679/NB2 pixel_2679/AMP_IN pixel_2679/SF_IB
+ pixel_2679/PIX_OUT pixel_2679/CSA_VREF pixel
Xpixel_2668 pixel_2668/gring pixel_2668/VDD pixel_2668/GND pixel_2668/VREF pixel_2668/ROW_SEL
+ pixel_2668/NB1 pixel_2668/VBIAS pixel_2668/NB2 pixel_2668/AMP_IN pixel_2668/SF_IB
+ pixel_2668/PIX_OUT pixel_2668/CSA_VREF pixel
Xpixel_2657 pixel_2657/gring pixel_2657/VDD pixel_2657/GND pixel_2657/VREF pixel_2657/ROW_SEL
+ pixel_2657/NB1 pixel_2657/VBIAS pixel_2657/NB2 pixel_2657/AMP_IN pixel_2657/SF_IB
+ pixel_2657/PIX_OUT pixel_2657/CSA_VREF pixel
Xpixel_1978 pixel_1978/gring pixel_1978/VDD pixel_1978/GND pixel_1978/VREF pixel_1978/ROW_SEL
+ pixel_1978/NB1 pixel_1978/VBIAS pixel_1978/NB2 pixel_1978/AMP_IN pixel_1978/SF_IB
+ pixel_1978/PIX_OUT pixel_1978/CSA_VREF pixel
Xpixel_1967 pixel_1967/gring pixel_1967/VDD pixel_1967/GND pixel_1967/VREF pixel_1967/ROW_SEL
+ pixel_1967/NB1 pixel_1967/VBIAS pixel_1967/NB2 pixel_1967/AMP_IN pixel_1967/SF_IB
+ pixel_1967/PIX_OUT pixel_1967/CSA_VREF pixel
Xpixel_1956 pixel_1956/gring pixel_1956/VDD pixel_1956/GND pixel_1956/VREF pixel_1956/ROW_SEL
+ pixel_1956/NB1 pixel_1956/VBIAS pixel_1956/NB2 pixel_1956/AMP_IN pixel_1956/SF_IB
+ pixel_1956/PIX_OUT pixel_1956/CSA_VREF pixel
Xpixel_1945 pixel_1945/gring pixel_1945/VDD pixel_1945/GND pixel_1945/VREF pixel_1945/ROW_SEL
+ pixel_1945/NB1 pixel_1945/VBIAS pixel_1945/NB2 pixel_1945/AMP_IN pixel_1945/SF_IB
+ pixel_1945/PIX_OUT pixel_1945/CSA_VREF pixel
Xpixel_1989 pixel_1989/gring pixel_1989/VDD pixel_1989/GND pixel_1989/VREF pixel_1989/ROW_SEL
+ pixel_1989/NB1 pixel_1989/VBIAS pixel_1989/NB2 pixel_1989/AMP_IN pixel_1989/SF_IB
+ pixel_1989/PIX_OUT pixel_1989/CSA_VREF pixel
Xpixel_5250 pixel_5250/gring pixel_5250/VDD pixel_5250/GND pixel_5250/VREF pixel_5250/ROW_SEL
+ pixel_5250/NB1 pixel_5250/VBIAS pixel_5250/NB2 pixel_5250/AMP_IN pixel_5250/SF_IB
+ pixel_5250/PIX_OUT pixel_5250/CSA_VREF pixel
Xpixel_5261 pixel_5261/gring pixel_5261/VDD pixel_5261/GND pixel_5261/VREF pixel_5261/ROW_SEL
+ pixel_5261/NB1 pixel_5261/VBIAS pixel_5261/NB2 pixel_5261/AMP_IN pixel_5261/SF_IB
+ pixel_5261/PIX_OUT pixel_5261/CSA_VREF pixel
Xpixel_5272 pixel_5272/gring pixel_5272/VDD pixel_5272/GND pixel_5272/VREF pixel_5272/ROW_SEL
+ pixel_5272/NB1 pixel_5272/VBIAS pixel_5272/NB2 pixel_5272/AMP_IN pixel_5272/SF_IB
+ pixel_5272/PIX_OUT pixel_5272/CSA_VREF pixel
Xpixel_5283 pixel_5283/gring pixel_5283/VDD pixel_5283/GND pixel_5283/VREF pixel_5283/ROW_SEL
+ pixel_5283/NB1 pixel_5283/VBIAS pixel_5283/NB2 pixel_5283/AMP_IN pixel_5283/SF_IB
+ pixel_5283/PIX_OUT pixel_5283/CSA_VREF pixel
Xpixel_5294 pixel_5294/gring pixel_5294/VDD pixel_5294/GND pixel_5294/VREF pixel_5294/ROW_SEL
+ pixel_5294/NB1 pixel_5294/VBIAS pixel_5294/NB2 pixel_5294/AMP_IN pixel_5294/SF_IB
+ pixel_5294/PIX_OUT pixel_5294/CSA_VREF pixel
Xpixel_4560 pixel_4560/gring pixel_4560/VDD pixel_4560/GND pixel_4560/VREF pixel_4560/ROW_SEL
+ pixel_4560/NB1 pixel_4560/VBIAS pixel_4560/NB2 pixel_4560/AMP_IN pixel_4560/SF_IB
+ pixel_4560/PIX_OUT pixel_4560/CSA_VREF pixel
Xpixel_4571 pixel_4571/gring pixel_4571/VDD pixel_4571/GND pixel_4571/VREF pixel_4571/ROW_SEL
+ pixel_4571/NB1 pixel_4571/VBIAS pixel_4571/NB2 pixel_4571/AMP_IN pixel_4571/SF_IB
+ pixel_4571/PIX_OUT pixel_4571/CSA_VREF pixel
Xpixel_4582 pixel_4582/gring pixel_4582/VDD pixel_4582/GND pixel_4582/VREF pixel_4582/ROW_SEL
+ pixel_4582/NB1 pixel_4582/VBIAS pixel_4582/NB2 pixel_4582/AMP_IN pixel_4582/SF_IB
+ pixel_4582/PIX_OUT pixel_4582/CSA_VREF pixel
Xpixel_3870 pixel_3870/gring pixel_3870/VDD pixel_3870/GND pixel_3870/VREF pixel_3870/ROW_SEL
+ pixel_3870/NB1 pixel_3870/VBIAS pixel_3870/NB2 pixel_3870/AMP_IN pixel_3870/SF_IB
+ pixel_3870/PIX_OUT pixel_3870/CSA_VREF pixel
Xpixel_4593 pixel_4593/gring pixel_4593/VDD pixel_4593/GND pixel_4593/VREF pixel_4593/ROW_SEL
+ pixel_4593/NB1 pixel_4593/VBIAS pixel_4593/NB2 pixel_4593/AMP_IN pixel_4593/SF_IB
+ pixel_4593/PIX_OUT pixel_4593/CSA_VREF pixel
Xpixel_3892 pixel_3892/gring pixel_3892/VDD pixel_3892/GND pixel_3892/VREF pixel_3892/ROW_SEL
+ pixel_3892/NB1 pixel_3892/VBIAS pixel_3892/NB2 pixel_3892/AMP_IN pixel_3892/SF_IB
+ pixel_3892/PIX_OUT pixel_3892/CSA_VREF pixel
Xpixel_3881 pixel_3881/gring pixel_3881/VDD pixel_3881/GND pixel_3881/VREF pixel_3881/ROW_SEL
+ pixel_3881/NB1 pixel_3881/VBIAS pixel_3881/NB2 pixel_3881/AMP_IN pixel_3881/SF_IB
+ pixel_3881/PIX_OUT pixel_3881/CSA_VREF pixel
Xpixel_1219 pixel_1219/gring pixel_1219/VDD pixel_1219/GND pixel_1219/VREF pixel_1219/ROW_SEL
+ pixel_1219/NB1 pixel_1219/VBIAS pixel_1219/NB2 pixel_1219/AMP_IN pixel_1219/SF_IB
+ pixel_1219/PIX_OUT pixel_1219/CSA_VREF pixel
Xpixel_1208 pixel_1208/gring pixel_1208/VDD pixel_1208/GND pixel_1208/VREF pixel_1208/ROW_SEL
+ pixel_1208/NB1 pixel_1208/VBIAS pixel_1208/NB2 pixel_1208/AMP_IN pixel_1208/SF_IB
+ pixel_1208/PIX_OUT pixel_1208/CSA_VREF pixel
Xpixel_9505 pixel_9505/gring pixel_9505/VDD pixel_9505/GND pixel_9505/VREF pixel_9505/ROW_SEL
+ pixel_9505/NB1 pixel_9505/VBIAS pixel_9505/NB2 pixel_9505/AMP_IN pixel_9505/SF_IB
+ pixel_9505/PIX_OUT pixel_9505/CSA_VREF pixel
Xpixel_9538 pixel_9538/gring pixel_9538/VDD pixel_9538/GND pixel_9538/VREF pixel_9538/ROW_SEL
+ pixel_9538/NB1 pixel_9538/VBIAS pixel_9538/NB2 pixel_9538/AMP_IN pixel_9538/SF_IB
+ pixel_9538/PIX_OUT pixel_9538/CSA_VREF pixel
Xpixel_9527 pixel_9527/gring pixel_9527/VDD pixel_9527/GND pixel_9527/VREF pixel_9527/ROW_SEL
+ pixel_9527/NB1 pixel_9527/VBIAS pixel_9527/NB2 pixel_9527/AMP_IN pixel_9527/SF_IB
+ pixel_9527/PIX_OUT pixel_9527/CSA_VREF pixel
Xpixel_9516 pixel_9516/gring pixel_9516/VDD pixel_9516/GND pixel_9516/VREF pixel_9516/ROW_SEL
+ pixel_9516/NB1 pixel_9516/VBIAS pixel_9516/NB2 pixel_9516/AMP_IN pixel_9516/SF_IB
+ pixel_9516/PIX_OUT pixel_9516/CSA_VREF pixel
Xpixel_8837 pixel_8837/gring pixel_8837/VDD pixel_8837/GND pixel_8837/VREF pixel_8837/ROW_SEL
+ pixel_8837/NB1 pixel_8837/VBIAS pixel_8837/NB2 pixel_8837/AMP_IN pixel_8837/SF_IB
+ pixel_8837/PIX_OUT pixel_8837/CSA_VREF pixel
Xpixel_8826 pixel_8826/gring pixel_8826/VDD pixel_8826/GND pixel_8826/VREF pixel_8826/ROW_SEL
+ pixel_8826/NB1 pixel_8826/VBIAS pixel_8826/NB2 pixel_8826/AMP_IN pixel_8826/SF_IB
+ pixel_8826/PIX_OUT pixel_8826/CSA_VREF pixel
Xpixel_8815 pixel_8815/gring pixel_8815/VDD pixel_8815/GND pixel_8815/VREF pixel_8815/ROW_SEL
+ pixel_8815/NB1 pixel_8815/VBIAS pixel_8815/NB2 pixel_8815/AMP_IN pixel_8815/SF_IB
+ pixel_8815/PIX_OUT pixel_8815/CSA_VREF pixel
Xpixel_8804 pixel_8804/gring pixel_8804/VDD pixel_8804/GND pixel_8804/VREF pixel_8804/ROW_SEL
+ pixel_8804/NB1 pixel_8804/VBIAS pixel_8804/NB2 pixel_8804/AMP_IN pixel_8804/SF_IB
+ pixel_8804/PIX_OUT pixel_8804/CSA_VREF pixel
Xpixel_9549 pixel_9549/gring pixel_9549/VDD pixel_9549/GND pixel_9549/VREF pixel_9549/ROW_SEL
+ pixel_9549/NB1 pixel_9549/VBIAS pixel_9549/NB2 pixel_9549/AMP_IN pixel_9549/SF_IB
+ pixel_9549/PIX_OUT pixel_9549/CSA_VREF pixel
Xpixel_8859 pixel_8859/gring pixel_8859/VDD pixel_8859/GND pixel_8859/VREF pixel_8859/ROW_SEL
+ pixel_8859/NB1 pixel_8859/VBIAS pixel_8859/NB2 pixel_8859/AMP_IN pixel_8859/SF_IB
+ pixel_8859/PIX_OUT pixel_8859/CSA_VREF pixel
Xpixel_8848 pixel_8848/gring pixel_8848/VDD pixel_8848/GND pixel_8848/VREF pixel_8848/ROW_SEL
+ pixel_8848/NB1 pixel_8848/VBIAS pixel_8848/NB2 pixel_8848/AMP_IN pixel_8848/SF_IB
+ pixel_8848/PIX_OUT pixel_8848/CSA_VREF pixel
Xpixel_3122 pixel_3122/gring pixel_3122/VDD pixel_3122/GND pixel_3122/VREF pixel_3122/ROW_SEL
+ pixel_3122/NB1 pixel_3122/VBIAS pixel_3122/NB2 pixel_3122/AMP_IN pixel_3122/SF_IB
+ pixel_3122/PIX_OUT pixel_3122/CSA_VREF pixel
Xpixel_3111 pixel_3111/gring pixel_3111/VDD pixel_3111/GND pixel_3111/VREF pixel_3111/ROW_SEL
+ pixel_3111/NB1 pixel_3111/VBIAS pixel_3111/NB2 pixel_3111/AMP_IN pixel_3111/SF_IB
+ pixel_3111/PIX_OUT pixel_3111/CSA_VREF pixel
Xpixel_3100 pixel_3100/gring pixel_3100/VDD pixel_3100/GND pixel_3100/VREF pixel_3100/ROW_SEL
+ pixel_3100/NB1 pixel_3100/VBIAS pixel_3100/NB2 pixel_3100/AMP_IN pixel_3100/SF_IB
+ pixel_3100/PIX_OUT pixel_3100/CSA_VREF pixel
Xpixel_2421 pixel_2421/gring pixel_2421/VDD pixel_2421/GND pixel_2421/VREF pixel_2421/ROW_SEL
+ pixel_2421/NB1 pixel_2421/VBIAS pixel_2421/NB2 pixel_2421/AMP_IN pixel_2421/SF_IB
+ pixel_2421/PIX_OUT pixel_2421/CSA_VREF pixel
Xpixel_2410 pixel_2410/gring pixel_2410/VDD pixel_2410/GND pixel_2410/VREF pixel_2410/ROW_SEL
+ pixel_2410/NB1 pixel_2410/VBIAS pixel_2410/NB2 pixel_2410/AMP_IN pixel_2410/SF_IB
+ pixel_2410/PIX_OUT pixel_2410/CSA_VREF pixel
Xpixel_3166 pixel_3166/gring pixel_3166/VDD pixel_3166/GND pixel_3166/VREF pixel_3166/ROW_SEL
+ pixel_3166/NB1 pixel_3166/VBIAS pixel_3166/NB2 pixel_3166/AMP_IN pixel_3166/SF_IB
+ pixel_3166/PIX_OUT pixel_3166/CSA_VREF pixel
Xpixel_3155 pixel_3155/gring pixel_3155/VDD pixel_3155/GND pixel_3155/VREF pixel_3155/ROW_SEL
+ pixel_3155/NB1 pixel_3155/VBIAS pixel_3155/NB2 pixel_3155/AMP_IN pixel_3155/SF_IB
+ pixel_3155/PIX_OUT pixel_3155/CSA_VREF pixel
Xpixel_3144 pixel_3144/gring pixel_3144/VDD pixel_3144/GND pixel_3144/VREF pixel_3144/ROW_SEL
+ pixel_3144/NB1 pixel_3144/VBIAS pixel_3144/NB2 pixel_3144/AMP_IN pixel_3144/SF_IB
+ pixel_3144/PIX_OUT pixel_3144/CSA_VREF pixel
Xpixel_3133 pixel_3133/gring pixel_3133/VDD pixel_3133/GND pixel_3133/VREF pixel_3133/ROW_SEL
+ pixel_3133/NB1 pixel_3133/VBIAS pixel_3133/NB2 pixel_3133/AMP_IN pixel_3133/SF_IB
+ pixel_3133/PIX_OUT pixel_3133/CSA_VREF pixel
Xpixel_2454 pixel_2454/gring pixel_2454/VDD pixel_2454/GND pixel_2454/VREF pixel_2454/ROW_SEL
+ pixel_2454/NB1 pixel_2454/VBIAS pixel_2454/NB2 pixel_2454/AMP_IN pixel_2454/SF_IB
+ pixel_2454/PIX_OUT pixel_2454/CSA_VREF pixel
Xpixel_2443 pixel_2443/gring pixel_2443/VDD pixel_2443/GND pixel_2443/VREF pixel_2443/ROW_SEL
+ pixel_2443/NB1 pixel_2443/VBIAS pixel_2443/NB2 pixel_2443/AMP_IN pixel_2443/SF_IB
+ pixel_2443/PIX_OUT pixel_2443/CSA_VREF pixel
Xpixel_2432 pixel_2432/gring pixel_2432/VDD pixel_2432/GND pixel_2432/VREF pixel_2432/ROW_SEL
+ pixel_2432/NB1 pixel_2432/VBIAS pixel_2432/NB2 pixel_2432/AMP_IN pixel_2432/SF_IB
+ pixel_2432/PIX_OUT pixel_2432/CSA_VREF pixel
Xpixel_3199 pixel_3199/gring pixel_3199/VDD pixel_3199/GND pixel_3199/VREF pixel_3199/ROW_SEL
+ pixel_3199/NB1 pixel_3199/VBIAS pixel_3199/NB2 pixel_3199/AMP_IN pixel_3199/SF_IB
+ pixel_3199/PIX_OUT pixel_3199/CSA_VREF pixel
Xpixel_3188 pixel_3188/gring pixel_3188/VDD pixel_3188/GND pixel_3188/VREF pixel_3188/ROW_SEL
+ pixel_3188/NB1 pixel_3188/VBIAS pixel_3188/NB2 pixel_3188/AMP_IN pixel_3188/SF_IB
+ pixel_3188/PIX_OUT pixel_3188/CSA_VREF pixel
Xpixel_3177 pixel_3177/gring pixel_3177/VDD pixel_3177/GND pixel_3177/VREF pixel_3177/ROW_SEL
+ pixel_3177/NB1 pixel_3177/VBIAS pixel_3177/NB2 pixel_3177/AMP_IN pixel_3177/SF_IB
+ pixel_3177/PIX_OUT pixel_3177/CSA_VREF pixel
Xpixel_1753 pixel_1753/gring pixel_1753/VDD pixel_1753/GND pixel_1753/VREF pixel_1753/ROW_SEL
+ pixel_1753/NB1 pixel_1753/VBIAS pixel_1753/NB2 pixel_1753/AMP_IN pixel_1753/SF_IB
+ pixel_1753/PIX_OUT pixel_1753/CSA_VREF pixel
Xpixel_1742 pixel_1742/gring pixel_1742/VDD pixel_1742/GND pixel_1742/VREF pixel_1742/ROW_SEL
+ pixel_1742/NB1 pixel_1742/VBIAS pixel_1742/NB2 pixel_1742/AMP_IN pixel_1742/SF_IB
+ pixel_1742/PIX_OUT pixel_1742/CSA_VREF pixel
Xpixel_1731 pixel_1731/gring pixel_1731/VDD pixel_1731/GND pixel_1731/VREF pixel_1731/ROW_SEL
+ pixel_1731/NB1 pixel_1731/VBIAS pixel_1731/NB2 pixel_1731/AMP_IN pixel_1731/SF_IB
+ pixel_1731/PIX_OUT pixel_1731/CSA_VREF pixel
Xpixel_1720 pixel_1720/gring pixel_1720/VDD pixel_1720/GND pixel_1720/VREF pixel_1720/ROW_SEL
+ pixel_1720/NB1 pixel_1720/VBIAS pixel_1720/NB2 pixel_1720/AMP_IN pixel_1720/SF_IB
+ pixel_1720/PIX_OUT pixel_1720/CSA_VREF pixel
Xpixel_2487 pixel_2487/gring pixel_2487/VDD pixel_2487/GND pixel_2487/VREF pixel_2487/ROW_SEL
+ pixel_2487/NB1 pixel_2487/VBIAS pixel_2487/NB2 pixel_2487/AMP_IN pixel_2487/SF_IB
+ pixel_2487/PIX_OUT pixel_2487/CSA_VREF pixel
Xpixel_2476 pixel_2476/gring pixel_2476/VDD pixel_2476/GND pixel_2476/VREF pixel_2476/ROW_SEL
+ pixel_2476/NB1 pixel_2476/VBIAS pixel_2476/NB2 pixel_2476/AMP_IN pixel_2476/SF_IB
+ pixel_2476/PIX_OUT pixel_2476/CSA_VREF pixel
Xpixel_2465 pixel_2465/gring pixel_2465/VDD pixel_2465/GND pixel_2465/VREF pixel_2465/ROW_SEL
+ pixel_2465/NB1 pixel_2465/VBIAS pixel_2465/NB2 pixel_2465/AMP_IN pixel_2465/SF_IB
+ pixel_2465/PIX_OUT pixel_2465/CSA_VREF pixel
Xpixel_1786 pixel_1786/gring pixel_1786/VDD pixel_1786/GND pixel_1786/VREF pixel_1786/ROW_SEL
+ pixel_1786/NB1 pixel_1786/VBIAS pixel_1786/NB2 pixel_1786/AMP_IN pixel_1786/SF_IB
+ pixel_1786/PIX_OUT pixel_1786/CSA_VREF pixel
Xpixel_1775 pixel_1775/gring pixel_1775/VDD pixel_1775/GND pixel_1775/VREF pixel_1775/ROW_SEL
+ pixel_1775/NB1 pixel_1775/VBIAS pixel_1775/NB2 pixel_1775/AMP_IN pixel_1775/SF_IB
+ pixel_1775/PIX_OUT pixel_1775/CSA_VREF pixel
Xpixel_1764 pixel_1764/gring pixel_1764/VDD pixel_1764/GND pixel_1764/VREF pixel_1764/ROW_SEL
+ pixel_1764/NB1 pixel_1764/VBIAS pixel_1764/NB2 pixel_1764/AMP_IN pixel_1764/SF_IB
+ pixel_1764/PIX_OUT pixel_1764/CSA_VREF pixel
Xpixel_2498 pixel_2498/gring pixel_2498/VDD pixel_2498/GND pixel_2498/VREF pixel_2498/ROW_SEL
+ pixel_2498/NB1 pixel_2498/VBIAS pixel_2498/NB2 pixel_2498/AMP_IN pixel_2498/SF_IB
+ pixel_2498/PIX_OUT pixel_2498/CSA_VREF pixel
Xpixel_1797 pixel_1797/gring pixel_1797/VDD pixel_1797/GND pixel_1797/VREF pixel_1797/ROW_SEL
+ pixel_1797/NB1 pixel_1797/VBIAS pixel_1797/NB2 pixel_1797/AMP_IN pixel_1797/SF_IB
+ pixel_1797/PIX_OUT pixel_1797/CSA_VREF pixel
Xpixel_5080 pixel_5080/gring pixel_5080/VDD pixel_5080/GND pixel_5080/VREF pixel_5080/ROW_SEL
+ pixel_5080/NB1 pixel_5080/VBIAS pixel_5080/NB2 pixel_5080/AMP_IN pixel_5080/SF_IB
+ pixel_5080/PIX_OUT pixel_5080/CSA_VREF pixel
Xpixel_5091 pixel_5091/gring pixel_5091/VDD pixel_5091/GND pixel_5091/VREF pixel_5091/ROW_SEL
+ pixel_5091/NB1 pixel_5091/VBIAS pixel_5091/NB2 pixel_5091/AMP_IN pixel_5091/SF_IB
+ pixel_5091/PIX_OUT pixel_5091/CSA_VREF pixel
Xpixel_4390 pixel_4390/gring pixel_4390/VDD pixel_4390/GND pixel_4390/VREF pixel_4390/ROW_SEL
+ pixel_4390/NB1 pixel_4390/VBIAS pixel_4390/NB2 pixel_4390/AMP_IN pixel_4390/SF_IB
+ pixel_4390/PIX_OUT pixel_4390/CSA_VREF pixel
Xpixel_6709 pixel_6709/gring pixel_6709/VDD pixel_6709/GND pixel_6709/VREF pixel_6709/ROW_SEL
+ pixel_6709/NB1 pixel_6709/VBIAS pixel_6709/NB2 pixel_6709/AMP_IN pixel_6709/SF_IB
+ pixel_6709/PIX_OUT pixel_6709/CSA_VREF pixel
Xpixel_1005 pixel_1005/gring pixel_1005/VDD pixel_1005/GND pixel_1005/VREF pixel_1005/ROW_SEL
+ pixel_1005/NB1 pixel_1005/VBIAS pixel_1005/NB2 pixel_1005/AMP_IN pixel_1005/SF_IB
+ pixel_1005/PIX_OUT pixel_1005/CSA_VREF pixel
Xpixel_1038 pixel_1038/gring pixel_1038/VDD pixel_1038/GND pixel_1038/VREF pixel_1038/ROW_SEL
+ pixel_1038/NB1 pixel_1038/VBIAS pixel_1038/NB2 pixel_1038/AMP_IN pixel_1038/SF_IB
+ pixel_1038/PIX_OUT pixel_1038/CSA_VREF pixel
Xpixel_1027 pixel_1027/gring pixel_1027/VDD pixel_1027/GND pixel_1027/VREF pixel_1027/ROW_SEL
+ pixel_1027/NB1 pixel_1027/VBIAS pixel_1027/NB2 pixel_1027/AMP_IN pixel_1027/SF_IB
+ pixel_1027/PIX_OUT pixel_1027/CSA_VREF pixel
Xpixel_1016 pixel_1016/gring pixel_1016/VDD pixel_1016/GND pixel_1016/VREF pixel_1016/ROW_SEL
+ pixel_1016/NB1 pixel_1016/VBIAS pixel_1016/NB2 pixel_1016/AMP_IN pixel_1016/SF_IB
+ pixel_1016/PIX_OUT pixel_1016/CSA_VREF pixel
Xpixel_1049 pixel_1049/gring pixel_1049/VDD pixel_1049/GND pixel_1049/VREF pixel_1049/ROW_SEL
+ pixel_1049/NB1 pixel_1049/VBIAS pixel_1049/NB2 pixel_1049/AMP_IN pixel_1049/SF_IB
+ pixel_1049/PIX_OUT pixel_1049/CSA_VREF pixel
Xpixel_9313 pixel_9313/gring pixel_9313/VDD pixel_9313/GND pixel_9313/VREF pixel_9313/ROW_SEL
+ pixel_9313/NB1 pixel_9313/VBIAS pixel_9313/NB2 pixel_9313/AMP_IN pixel_9313/SF_IB
+ pixel_9313/PIX_OUT pixel_9313/CSA_VREF pixel
Xpixel_9302 pixel_9302/gring pixel_9302/VDD pixel_9302/GND pixel_9302/VREF pixel_9302/ROW_SEL
+ pixel_9302/NB1 pixel_9302/VBIAS pixel_9302/NB2 pixel_9302/AMP_IN pixel_9302/SF_IB
+ pixel_9302/PIX_OUT pixel_9302/CSA_VREF pixel
Xpixel_8601 pixel_8601/gring pixel_8601/VDD pixel_8601/GND pixel_8601/VREF pixel_8601/ROW_SEL
+ pixel_8601/NB1 pixel_8601/VBIAS pixel_8601/NB2 pixel_8601/AMP_IN pixel_8601/SF_IB
+ pixel_8601/PIX_OUT pixel_8601/CSA_VREF pixel
Xpixel_9346 pixel_9346/gring pixel_9346/VDD pixel_9346/GND pixel_9346/VREF pixel_9346/ROW_SEL
+ pixel_9346/NB1 pixel_9346/VBIAS pixel_9346/NB2 pixel_9346/AMP_IN pixel_9346/SF_IB
+ pixel_9346/PIX_OUT pixel_9346/CSA_VREF pixel
Xpixel_9335 pixel_9335/gring pixel_9335/VDD pixel_9335/GND pixel_9335/VREF pixel_9335/ROW_SEL
+ pixel_9335/NB1 pixel_9335/VBIAS pixel_9335/NB2 pixel_9335/AMP_IN pixel_9335/SF_IB
+ pixel_9335/PIX_OUT pixel_9335/CSA_VREF pixel
Xpixel_9324 pixel_9324/gring pixel_9324/VDD pixel_9324/GND pixel_9324/VREF pixel_9324/ROW_SEL
+ pixel_9324/NB1 pixel_9324/VBIAS pixel_9324/NB2 pixel_9324/AMP_IN pixel_9324/SF_IB
+ pixel_9324/PIX_OUT pixel_9324/CSA_VREF pixel
Xpixel_8645 pixel_8645/gring pixel_8645/VDD pixel_8645/GND pixel_8645/VREF pixel_8645/ROW_SEL
+ pixel_8645/NB1 pixel_8645/VBIAS pixel_8645/NB2 pixel_8645/AMP_IN pixel_8645/SF_IB
+ pixel_8645/PIX_OUT pixel_8645/CSA_VREF pixel
Xpixel_8634 pixel_8634/gring pixel_8634/VDD pixel_8634/GND pixel_8634/VREF pixel_8634/ROW_SEL
+ pixel_8634/NB1 pixel_8634/VBIAS pixel_8634/NB2 pixel_8634/AMP_IN pixel_8634/SF_IB
+ pixel_8634/PIX_OUT pixel_8634/CSA_VREF pixel
Xpixel_8623 pixel_8623/gring pixel_8623/VDD pixel_8623/GND pixel_8623/VREF pixel_8623/ROW_SEL
+ pixel_8623/NB1 pixel_8623/VBIAS pixel_8623/NB2 pixel_8623/AMP_IN pixel_8623/SF_IB
+ pixel_8623/PIX_OUT pixel_8623/CSA_VREF pixel
Xpixel_8612 pixel_8612/gring pixel_8612/VDD pixel_8612/GND pixel_8612/VREF pixel_8612/ROW_SEL
+ pixel_8612/NB1 pixel_8612/VBIAS pixel_8612/NB2 pixel_8612/AMP_IN pixel_8612/SF_IB
+ pixel_8612/PIX_OUT pixel_8612/CSA_VREF pixel
Xpixel_9379 pixel_9379/gring pixel_9379/VDD pixel_9379/GND pixel_9379/VREF pixel_9379/ROW_SEL
+ pixel_9379/NB1 pixel_9379/VBIAS pixel_9379/NB2 pixel_9379/AMP_IN pixel_9379/SF_IB
+ pixel_9379/PIX_OUT pixel_9379/CSA_VREF pixel
Xpixel_9368 pixel_9368/gring pixel_9368/VDD pixel_9368/GND pixel_9368/VREF pixel_9368/ROW_SEL
+ pixel_9368/NB1 pixel_9368/VBIAS pixel_9368/NB2 pixel_9368/AMP_IN pixel_9368/SF_IB
+ pixel_9368/PIX_OUT pixel_9368/CSA_VREF pixel
Xpixel_9357 pixel_9357/gring pixel_9357/VDD pixel_9357/GND pixel_9357/VREF pixel_9357/ROW_SEL
+ pixel_9357/NB1 pixel_9357/VBIAS pixel_9357/NB2 pixel_9357/AMP_IN pixel_9357/SF_IB
+ pixel_9357/PIX_OUT pixel_9357/CSA_VREF pixel
Xpixel_7900 pixel_7900/gring pixel_7900/VDD pixel_7900/GND pixel_7900/VREF pixel_7900/ROW_SEL
+ pixel_7900/NB1 pixel_7900/VBIAS pixel_7900/NB2 pixel_7900/AMP_IN pixel_7900/SF_IB
+ pixel_7900/PIX_OUT pixel_7900/CSA_VREF pixel
Xpixel_8678 pixel_8678/gring pixel_8678/VDD pixel_8678/GND pixel_8678/VREF pixel_8678/ROW_SEL
+ pixel_8678/NB1 pixel_8678/VBIAS pixel_8678/NB2 pixel_8678/AMP_IN pixel_8678/SF_IB
+ pixel_8678/PIX_OUT pixel_8678/CSA_VREF pixel
Xpixel_8667 pixel_8667/gring pixel_8667/VDD pixel_8667/GND pixel_8667/VREF pixel_8667/ROW_SEL
+ pixel_8667/NB1 pixel_8667/VBIAS pixel_8667/NB2 pixel_8667/AMP_IN pixel_8667/SF_IB
+ pixel_8667/PIX_OUT pixel_8667/CSA_VREF pixel
Xpixel_8656 pixel_8656/gring pixel_8656/VDD pixel_8656/GND pixel_8656/VREF pixel_8656/ROW_SEL
+ pixel_8656/NB1 pixel_8656/VBIAS pixel_8656/NB2 pixel_8656/AMP_IN pixel_8656/SF_IB
+ pixel_8656/PIX_OUT pixel_8656/CSA_VREF pixel
Xpixel_7911 pixel_7911/gring pixel_7911/VDD pixel_7911/GND pixel_7911/VREF pixel_7911/ROW_SEL
+ pixel_7911/NB1 pixel_7911/VBIAS pixel_7911/NB2 pixel_7911/AMP_IN pixel_7911/SF_IB
+ pixel_7911/PIX_OUT pixel_7911/CSA_VREF pixel
Xpixel_7922 pixel_7922/gring pixel_7922/VDD pixel_7922/GND pixel_7922/VREF pixel_7922/ROW_SEL
+ pixel_7922/NB1 pixel_7922/VBIAS pixel_7922/NB2 pixel_7922/AMP_IN pixel_7922/SF_IB
+ pixel_7922/PIX_OUT pixel_7922/CSA_VREF pixel
Xpixel_7933 pixel_7933/gring pixel_7933/VDD pixel_7933/GND pixel_7933/VREF pixel_7933/ROW_SEL
+ pixel_7933/NB1 pixel_7933/VBIAS pixel_7933/NB2 pixel_7933/AMP_IN pixel_7933/SF_IB
+ pixel_7933/PIX_OUT pixel_7933/CSA_VREF pixel
Xpixel_8689 pixel_8689/gring pixel_8689/VDD pixel_8689/GND pixel_8689/VREF pixel_8689/ROW_SEL
+ pixel_8689/NB1 pixel_8689/VBIAS pixel_8689/NB2 pixel_8689/AMP_IN pixel_8689/SF_IB
+ pixel_8689/PIX_OUT pixel_8689/CSA_VREF pixel
Xpixel_7944 pixel_7944/gring pixel_7944/VDD pixel_7944/GND pixel_7944/VREF pixel_7944/ROW_SEL
+ pixel_7944/NB1 pixel_7944/VBIAS pixel_7944/NB2 pixel_7944/AMP_IN pixel_7944/SF_IB
+ pixel_7944/PIX_OUT pixel_7944/CSA_VREF pixel
Xpixel_7955 pixel_7955/gring pixel_7955/VDD pixel_7955/GND pixel_7955/VREF pixel_7955/ROW_SEL
+ pixel_7955/NB1 pixel_7955/VBIAS pixel_7955/NB2 pixel_7955/AMP_IN pixel_7955/SF_IB
+ pixel_7955/PIX_OUT pixel_7955/CSA_VREF pixel
Xpixel_7966 pixel_7966/gring pixel_7966/VDD pixel_7966/GND pixel_7966/VREF pixel_7966/ROW_SEL
+ pixel_7966/NB1 pixel_7966/VBIAS pixel_7966/NB2 pixel_7966/AMP_IN pixel_7966/SF_IB
+ pixel_7966/PIX_OUT pixel_7966/CSA_VREF pixel
Xpixel_7977 pixel_7977/gring pixel_7977/VDD pixel_7977/GND pixel_7977/VREF pixel_7977/ROW_SEL
+ pixel_7977/NB1 pixel_7977/VBIAS pixel_7977/NB2 pixel_7977/AMP_IN pixel_7977/SF_IB
+ pixel_7977/PIX_OUT pixel_7977/CSA_VREF pixel
Xpixel_7988 pixel_7988/gring pixel_7988/VDD pixel_7988/GND pixel_7988/VREF pixel_7988/ROW_SEL
+ pixel_7988/NB1 pixel_7988/VBIAS pixel_7988/NB2 pixel_7988/AMP_IN pixel_7988/SF_IB
+ pixel_7988/PIX_OUT pixel_7988/CSA_VREF pixel
Xpixel_7999 pixel_7999/gring pixel_7999/VDD pixel_7999/GND pixel_7999/VREF pixel_7999/ROW_SEL
+ pixel_7999/NB1 pixel_7999/VBIAS pixel_7999/NB2 pixel_7999/AMP_IN pixel_7999/SF_IB
+ pixel_7999/PIX_OUT pixel_7999/CSA_VREF pixel
Xpixel_2262 pixel_2262/gring pixel_2262/VDD pixel_2262/GND pixel_2262/VREF pixel_2262/ROW_SEL
+ pixel_2262/NB1 pixel_2262/VBIAS pixel_2262/NB2 pixel_2262/AMP_IN pixel_2262/SF_IB
+ pixel_2262/PIX_OUT pixel_2262/CSA_VREF pixel
Xpixel_2251 pixel_2251/gring pixel_2251/VDD pixel_2251/GND pixel_2251/VREF pixel_2251/ROW_SEL
+ pixel_2251/NB1 pixel_2251/VBIAS pixel_2251/NB2 pixel_2251/AMP_IN pixel_2251/SF_IB
+ pixel_2251/PIX_OUT pixel_2251/CSA_VREF pixel
Xpixel_2240 pixel_2240/gring pixel_2240/VDD pixel_2240/GND pixel_2240/VREF pixel_2240/ROW_SEL
+ pixel_2240/NB1 pixel_2240/VBIAS pixel_2240/NB2 pixel_2240/AMP_IN pixel_2240/SF_IB
+ pixel_2240/PIX_OUT pixel_2240/CSA_VREF pixel
Xpixel_1561 pixel_1561/gring pixel_1561/VDD pixel_1561/GND pixel_1561/VREF pixel_1561/ROW_SEL
+ pixel_1561/NB1 pixel_1561/VBIAS pixel_1561/NB2 pixel_1561/AMP_IN pixel_1561/SF_IB
+ pixel_1561/PIX_OUT pixel_1561/CSA_VREF pixel
Xpixel_1550 pixel_1550/gring pixel_1550/VDD pixel_1550/GND pixel_1550/VREF pixel_1550/ROW_SEL
+ pixel_1550/NB1 pixel_1550/VBIAS pixel_1550/NB2 pixel_1550/AMP_IN pixel_1550/SF_IB
+ pixel_1550/PIX_OUT pixel_1550/CSA_VREF pixel
Xpixel_2295 pixel_2295/gring pixel_2295/VDD pixel_2295/GND pixel_2295/VREF pixel_2295/ROW_SEL
+ pixel_2295/NB1 pixel_2295/VBIAS pixel_2295/NB2 pixel_2295/AMP_IN pixel_2295/SF_IB
+ pixel_2295/PIX_OUT pixel_2295/CSA_VREF pixel
Xpixel_2284 pixel_2284/gring pixel_2284/VDD pixel_2284/GND pixel_2284/VREF pixel_2284/ROW_SEL
+ pixel_2284/NB1 pixel_2284/VBIAS pixel_2284/NB2 pixel_2284/AMP_IN pixel_2284/SF_IB
+ pixel_2284/PIX_OUT pixel_2284/CSA_VREF pixel
Xpixel_2273 pixel_2273/gring pixel_2273/VDD pixel_2273/GND pixel_2273/VREF pixel_2273/ROW_SEL
+ pixel_2273/NB1 pixel_2273/VBIAS pixel_2273/NB2 pixel_2273/AMP_IN pixel_2273/SF_IB
+ pixel_2273/PIX_OUT pixel_2273/CSA_VREF pixel
Xpixel_1594 pixel_1594/gring pixel_1594/VDD pixel_1594/GND pixel_1594/VREF pixel_1594/ROW_SEL
+ pixel_1594/NB1 pixel_1594/VBIAS pixel_1594/NB2 pixel_1594/AMP_IN pixel_1594/SF_IB
+ pixel_1594/PIX_OUT pixel_1594/CSA_VREF pixel
Xpixel_1583 pixel_1583/gring pixel_1583/VDD pixel_1583/GND pixel_1583/VREF pixel_1583/ROW_SEL
+ pixel_1583/NB1 pixel_1583/VBIAS pixel_1583/NB2 pixel_1583/AMP_IN pixel_1583/SF_IB
+ pixel_1583/PIX_OUT pixel_1583/CSA_VREF pixel
Xpixel_1572 pixel_1572/gring pixel_1572/VDD pixel_1572/GND pixel_1572/VREF pixel_1572/ROW_SEL
+ pixel_1572/NB1 pixel_1572/VBIAS pixel_1572/NB2 pixel_1572/AMP_IN pixel_1572/SF_IB
+ pixel_1572/PIX_OUT pixel_1572/CSA_VREF pixel
Xpixel_9880 pixel_9880/gring pixel_9880/VDD pixel_9880/GND pixel_9880/VREF pixel_9880/ROW_SEL
+ pixel_9880/NB1 pixel_9880/VBIAS pixel_9880/NB2 pixel_9880/AMP_IN pixel_9880/SF_IB
+ pixel_9880/PIX_OUT pixel_9880/CSA_VREF pixel
Xpixel_9891 pixel_9891/gring pixel_9891/VDD pixel_9891/GND pixel_9891/VREF pixel_9891/ROW_SEL
+ pixel_9891/NB1 pixel_9891/VBIAS pixel_9891/NB2 pixel_9891/AMP_IN pixel_9891/SF_IB
+ pixel_9891/PIX_OUT pixel_9891/CSA_VREF pixel
Xpixel_609 pixel_609/gring pixel_609/VDD pixel_609/GND pixel_609/VREF pixel_609/ROW_SEL
+ pixel_609/NB1 pixel_609/VBIAS pixel_609/NB2 pixel_609/AMP_IN pixel_609/SF_IB pixel_609/PIX_OUT
+ pixel_609/CSA_VREF pixel
Xpixel_7207 pixel_7207/gring pixel_7207/VDD pixel_7207/GND pixel_7207/VREF pixel_7207/ROW_SEL
+ pixel_7207/NB1 pixel_7207/VBIAS pixel_7207/NB2 pixel_7207/AMP_IN pixel_7207/SF_IB
+ pixel_7207/PIX_OUT pixel_7207/CSA_VREF pixel
Xpixel_7218 pixel_7218/gring pixel_7218/VDD pixel_7218/GND pixel_7218/VREF pixel_7218/ROW_SEL
+ pixel_7218/NB1 pixel_7218/VBIAS pixel_7218/NB2 pixel_7218/AMP_IN pixel_7218/SF_IB
+ pixel_7218/PIX_OUT pixel_7218/CSA_VREF pixel
Xpixel_7229 pixel_7229/gring pixel_7229/VDD pixel_7229/GND pixel_7229/VREF pixel_7229/ROW_SEL
+ pixel_7229/NB1 pixel_7229/VBIAS pixel_7229/NB2 pixel_7229/AMP_IN pixel_7229/SF_IB
+ pixel_7229/PIX_OUT pixel_7229/CSA_VREF pixel
Xpixel_6506 pixel_6506/gring pixel_6506/VDD pixel_6506/GND pixel_6506/VREF pixel_6506/ROW_SEL
+ pixel_6506/NB1 pixel_6506/VBIAS pixel_6506/NB2 pixel_6506/AMP_IN pixel_6506/SF_IB
+ pixel_6506/PIX_OUT pixel_6506/CSA_VREF pixel
Xpixel_6517 pixel_6517/gring pixel_6517/VDD pixel_6517/GND pixel_6517/VREF pixel_6517/ROW_SEL
+ pixel_6517/NB1 pixel_6517/VBIAS pixel_6517/NB2 pixel_6517/AMP_IN pixel_6517/SF_IB
+ pixel_6517/PIX_OUT pixel_6517/CSA_VREF pixel
Xpixel_6528 pixel_6528/gring pixel_6528/VDD pixel_6528/GND pixel_6528/VREF pixel_6528/ROW_SEL
+ pixel_6528/NB1 pixel_6528/VBIAS pixel_6528/NB2 pixel_6528/AMP_IN pixel_6528/SF_IB
+ pixel_6528/PIX_OUT pixel_6528/CSA_VREF pixel
Xpixel_6539 pixel_6539/gring pixel_6539/VDD pixel_6539/GND pixel_6539/VREF pixel_6539/ROW_SEL
+ pixel_6539/NB1 pixel_6539/VBIAS pixel_6539/NB2 pixel_6539/AMP_IN pixel_6539/SF_IB
+ pixel_6539/PIX_OUT pixel_6539/CSA_VREF pixel
Xpixel_5805 pixel_5805/gring pixel_5805/VDD pixel_5805/GND pixel_5805/VREF pixel_5805/ROW_SEL
+ pixel_5805/NB1 pixel_5805/VBIAS pixel_5805/NB2 pixel_5805/AMP_IN pixel_5805/SF_IB
+ pixel_5805/PIX_OUT pixel_5805/CSA_VREF pixel
Xpixel_5816 pixel_5816/gring pixel_5816/VDD pixel_5816/GND pixel_5816/VREF pixel_5816/ROW_SEL
+ pixel_5816/NB1 pixel_5816/VBIAS pixel_5816/NB2 pixel_5816/AMP_IN pixel_5816/SF_IB
+ pixel_5816/PIX_OUT pixel_5816/CSA_VREF pixel
Xpixel_5827 pixel_5827/gring pixel_5827/VDD pixel_5827/GND pixel_5827/VREF pixel_5827/ROW_SEL
+ pixel_5827/NB1 pixel_5827/VBIAS pixel_5827/NB2 pixel_5827/AMP_IN pixel_5827/SF_IB
+ pixel_5827/PIX_OUT pixel_5827/CSA_VREF pixel
Xpixel_5838 pixel_5838/gring pixel_5838/VDD pixel_5838/GND pixel_5838/VREF pixel_5838/ROW_SEL
+ pixel_5838/NB1 pixel_5838/VBIAS pixel_5838/NB2 pixel_5838/AMP_IN pixel_5838/SF_IB
+ pixel_5838/PIX_OUT pixel_5838/CSA_VREF pixel
Xpixel_5849 pixel_5849/gring pixel_5849/VDD pixel_5849/GND pixel_5849/VREF pixel_5849/ROW_SEL
+ pixel_5849/NB1 pixel_5849/VBIAS pixel_5849/NB2 pixel_5849/AMP_IN pixel_5849/SF_IB
+ pixel_5849/PIX_OUT pixel_5849/CSA_VREF pixel
Xpixel_9121 pixel_9121/gring pixel_9121/VDD pixel_9121/GND pixel_9121/VREF pixel_9121/ROW_SEL
+ pixel_9121/NB1 pixel_9121/VBIAS pixel_9121/NB2 pixel_9121/AMP_IN pixel_9121/SF_IB
+ pixel_9121/PIX_OUT pixel_9121/CSA_VREF pixel
Xpixel_9110 pixel_9110/gring pixel_9110/VDD pixel_9110/GND pixel_9110/VREF pixel_9110/ROW_SEL
+ pixel_9110/NB1 pixel_9110/VBIAS pixel_9110/NB2 pixel_9110/AMP_IN pixel_9110/SF_IB
+ pixel_9110/PIX_OUT pixel_9110/CSA_VREF pixel
Xpixel_8420 pixel_8420/gring pixel_8420/VDD pixel_8420/GND pixel_8420/VREF pixel_8420/ROW_SEL
+ pixel_8420/NB1 pixel_8420/VBIAS pixel_8420/NB2 pixel_8420/AMP_IN pixel_8420/SF_IB
+ pixel_8420/PIX_OUT pixel_8420/CSA_VREF pixel
Xpixel_9154 pixel_9154/gring pixel_9154/VDD pixel_9154/GND pixel_9154/VREF pixel_9154/ROW_SEL
+ pixel_9154/NB1 pixel_9154/VBIAS pixel_9154/NB2 pixel_9154/AMP_IN pixel_9154/SF_IB
+ pixel_9154/PIX_OUT pixel_9154/CSA_VREF pixel
Xpixel_9143 pixel_9143/gring pixel_9143/VDD pixel_9143/GND pixel_9143/VREF pixel_9143/ROW_SEL
+ pixel_9143/NB1 pixel_9143/VBIAS pixel_9143/NB2 pixel_9143/AMP_IN pixel_9143/SF_IB
+ pixel_9143/PIX_OUT pixel_9143/CSA_VREF pixel
Xpixel_9132 pixel_9132/gring pixel_9132/VDD pixel_9132/GND pixel_9132/VREF pixel_9132/ROW_SEL
+ pixel_9132/NB1 pixel_9132/VBIAS pixel_9132/NB2 pixel_9132/AMP_IN pixel_9132/SF_IB
+ pixel_9132/PIX_OUT pixel_9132/CSA_VREF pixel
Xpixel_8431 pixel_8431/gring pixel_8431/VDD pixel_8431/GND pixel_8431/VREF pixel_8431/ROW_SEL
+ pixel_8431/NB1 pixel_8431/VBIAS pixel_8431/NB2 pixel_8431/AMP_IN pixel_8431/SF_IB
+ pixel_8431/PIX_OUT pixel_8431/CSA_VREF pixel
Xpixel_9198 pixel_9198/gring pixel_9198/VDD pixel_9198/GND pixel_9198/VREF pixel_9198/ROW_SEL
+ pixel_9198/NB1 pixel_9198/VBIAS pixel_9198/NB2 pixel_9198/AMP_IN pixel_9198/SF_IB
+ pixel_9198/PIX_OUT pixel_9198/CSA_VREF pixel
Xpixel_9187 pixel_9187/gring pixel_9187/VDD pixel_9187/GND pixel_9187/VREF pixel_9187/ROW_SEL
+ pixel_9187/NB1 pixel_9187/VBIAS pixel_9187/NB2 pixel_9187/AMP_IN pixel_9187/SF_IB
+ pixel_9187/PIX_OUT pixel_9187/CSA_VREF pixel
Xpixel_9176 pixel_9176/gring pixel_9176/VDD pixel_9176/GND pixel_9176/VREF pixel_9176/ROW_SEL
+ pixel_9176/NB1 pixel_9176/VBIAS pixel_9176/NB2 pixel_9176/AMP_IN pixel_9176/SF_IB
+ pixel_9176/PIX_OUT pixel_9176/CSA_VREF pixel
Xpixel_9165 pixel_9165/gring pixel_9165/VDD pixel_9165/GND pixel_9165/VREF pixel_9165/ROW_SEL
+ pixel_9165/NB1 pixel_9165/VBIAS pixel_9165/NB2 pixel_9165/AMP_IN pixel_9165/SF_IB
+ pixel_9165/PIX_OUT pixel_9165/CSA_VREF pixel
Xpixel_8442 pixel_8442/gring pixel_8442/VDD pixel_8442/GND pixel_8442/VREF pixel_8442/ROW_SEL
+ pixel_8442/NB1 pixel_8442/VBIAS pixel_8442/NB2 pixel_8442/AMP_IN pixel_8442/SF_IB
+ pixel_8442/PIX_OUT pixel_8442/CSA_VREF pixel
Xpixel_8453 pixel_8453/gring pixel_8453/VDD pixel_8453/GND pixel_8453/VREF pixel_8453/ROW_SEL
+ pixel_8453/NB1 pixel_8453/VBIAS pixel_8453/NB2 pixel_8453/AMP_IN pixel_8453/SF_IB
+ pixel_8453/PIX_OUT pixel_8453/CSA_VREF pixel
Xpixel_8464 pixel_8464/gring pixel_8464/VDD pixel_8464/GND pixel_8464/VREF pixel_8464/ROW_SEL
+ pixel_8464/NB1 pixel_8464/VBIAS pixel_8464/NB2 pixel_8464/AMP_IN pixel_8464/SF_IB
+ pixel_8464/PIX_OUT pixel_8464/CSA_VREF pixel
Xpixel_8475 pixel_8475/gring pixel_8475/VDD pixel_8475/GND pixel_8475/VREF pixel_8475/ROW_SEL
+ pixel_8475/NB1 pixel_8475/VBIAS pixel_8475/NB2 pixel_8475/AMP_IN pixel_8475/SF_IB
+ pixel_8475/PIX_OUT pixel_8475/CSA_VREF pixel
Xpixel_8486 pixel_8486/gring pixel_8486/VDD pixel_8486/GND pixel_8486/VREF pixel_8486/ROW_SEL
+ pixel_8486/NB1 pixel_8486/VBIAS pixel_8486/NB2 pixel_8486/AMP_IN pixel_8486/SF_IB
+ pixel_8486/PIX_OUT pixel_8486/CSA_VREF pixel
Xpixel_7730 pixel_7730/gring pixel_7730/VDD pixel_7730/GND pixel_7730/VREF pixel_7730/ROW_SEL
+ pixel_7730/NB1 pixel_7730/VBIAS pixel_7730/NB2 pixel_7730/AMP_IN pixel_7730/SF_IB
+ pixel_7730/PIX_OUT pixel_7730/CSA_VREF pixel
Xpixel_7741 pixel_7741/gring pixel_7741/VDD pixel_7741/GND pixel_7741/VREF pixel_7741/ROW_SEL
+ pixel_7741/NB1 pixel_7741/VBIAS pixel_7741/NB2 pixel_7741/AMP_IN pixel_7741/SF_IB
+ pixel_7741/PIX_OUT pixel_7741/CSA_VREF pixel
Xpixel_8497 pixel_8497/gring pixel_8497/VDD pixel_8497/GND pixel_8497/VREF pixel_8497/ROW_SEL
+ pixel_8497/NB1 pixel_8497/VBIAS pixel_8497/NB2 pixel_8497/AMP_IN pixel_8497/SF_IB
+ pixel_8497/PIX_OUT pixel_8497/CSA_VREF pixel
Xpixel_7752 pixel_7752/gring pixel_7752/VDD pixel_7752/GND pixel_7752/VREF pixel_7752/ROW_SEL
+ pixel_7752/NB1 pixel_7752/VBIAS pixel_7752/NB2 pixel_7752/AMP_IN pixel_7752/SF_IB
+ pixel_7752/PIX_OUT pixel_7752/CSA_VREF pixel
Xpixel_7763 pixel_7763/gring pixel_7763/VDD pixel_7763/GND pixel_7763/VREF pixel_7763/ROW_SEL
+ pixel_7763/NB1 pixel_7763/VBIAS pixel_7763/NB2 pixel_7763/AMP_IN pixel_7763/SF_IB
+ pixel_7763/PIX_OUT pixel_7763/CSA_VREF pixel
Xpixel_7774 pixel_7774/gring pixel_7774/VDD pixel_7774/GND pixel_7774/VREF pixel_7774/ROW_SEL
+ pixel_7774/NB1 pixel_7774/VBIAS pixel_7774/NB2 pixel_7774/AMP_IN pixel_7774/SF_IB
+ pixel_7774/PIX_OUT pixel_7774/CSA_VREF pixel
Xpixel_7785 pixel_7785/gring pixel_7785/VDD pixel_7785/GND pixel_7785/VREF pixel_7785/ROW_SEL
+ pixel_7785/NB1 pixel_7785/VBIAS pixel_7785/NB2 pixel_7785/AMP_IN pixel_7785/SF_IB
+ pixel_7785/PIX_OUT pixel_7785/CSA_VREF pixel
Xpixel_7796 pixel_7796/gring pixel_7796/VDD pixel_7796/GND pixel_7796/VREF pixel_7796/ROW_SEL
+ pixel_7796/NB1 pixel_7796/VBIAS pixel_7796/NB2 pixel_7796/AMP_IN pixel_7796/SF_IB
+ pixel_7796/PIX_OUT pixel_7796/CSA_VREF pixel
Xpixel_2081 pixel_2081/gring pixel_2081/VDD pixel_2081/GND pixel_2081/VREF pixel_2081/ROW_SEL
+ pixel_2081/NB1 pixel_2081/VBIAS pixel_2081/NB2 pixel_2081/AMP_IN pixel_2081/SF_IB
+ pixel_2081/PIX_OUT pixel_2081/CSA_VREF pixel
Xpixel_2070 pixel_2070/gring pixel_2070/VDD pixel_2070/GND pixel_2070/VREF pixel_2070/ROW_SEL
+ pixel_2070/NB1 pixel_2070/VBIAS pixel_2070/NB2 pixel_2070/AMP_IN pixel_2070/SF_IB
+ pixel_2070/PIX_OUT pixel_2070/CSA_VREF pixel
Xpixel_2092 pixel_2092/gring pixel_2092/VDD pixel_2092/GND pixel_2092/VREF pixel_2092/ROW_SEL
+ pixel_2092/NB1 pixel_2092/VBIAS pixel_2092/NB2 pixel_2092/AMP_IN pixel_2092/SF_IB
+ pixel_2092/PIX_OUT pixel_2092/CSA_VREF pixel
Xpixel_1391 pixel_1391/gring pixel_1391/VDD pixel_1391/GND pixel_1391/VREF pixel_1391/ROW_SEL
+ pixel_1391/NB1 pixel_1391/VBIAS pixel_1391/NB2 pixel_1391/AMP_IN pixel_1391/SF_IB
+ pixel_1391/PIX_OUT pixel_1391/CSA_VREF pixel
Xpixel_1380 pixel_1380/gring pixel_1380/VDD pixel_1380/GND pixel_1380/VREF pixel_1380/ROW_SEL
+ pixel_1380/NB1 pixel_1380/VBIAS pixel_1380/NB2 pixel_1380/AMP_IN pixel_1380/SF_IB
+ pixel_1380/PIX_OUT pixel_1380/CSA_VREF pixel
Xpixel_428 pixel_428/gring pixel_428/VDD pixel_428/GND pixel_428/VREF pixel_428/ROW_SEL
+ pixel_428/NB1 pixel_428/VBIAS pixel_428/NB2 pixel_428/AMP_IN pixel_428/SF_IB pixel_428/PIX_OUT
+ pixel_428/CSA_VREF pixel
Xpixel_417 pixel_417/gring pixel_417/VDD pixel_417/GND pixel_417/VREF pixel_417/ROW_SEL
+ pixel_417/NB1 pixel_417/VBIAS pixel_417/NB2 pixel_417/AMP_IN pixel_417/SF_IB pixel_417/PIX_OUT
+ pixel_417/CSA_VREF pixel
Xpixel_406 pixel_406/gring pixel_406/VDD pixel_406/GND pixel_406/VREF pixel_406/ROW_SEL
+ pixel_406/NB1 pixel_406/VBIAS pixel_406/NB2 pixel_406/AMP_IN pixel_406/SF_IB pixel_406/PIX_OUT
+ pixel_406/CSA_VREF pixel
Xpixel_439 pixel_439/gring pixel_439/VDD pixel_439/GND pixel_439/VREF pixel_439/ROW_SEL
+ pixel_439/NB1 pixel_439/VBIAS pixel_439/NB2 pixel_439/AMP_IN pixel_439/SF_IB pixel_439/PIX_OUT
+ pixel_439/CSA_VREF pixel
Xpixel_7004 pixel_7004/gring pixel_7004/VDD pixel_7004/GND pixel_7004/VREF pixel_7004/ROW_SEL
+ pixel_7004/NB1 pixel_7004/VBIAS pixel_7004/NB2 pixel_7004/AMP_IN pixel_7004/SF_IB
+ pixel_7004/PIX_OUT pixel_7004/CSA_VREF pixel
Xpixel_7015 pixel_7015/gring pixel_7015/VDD pixel_7015/GND pixel_7015/VREF pixel_7015/ROW_SEL
+ pixel_7015/NB1 pixel_7015/VBIAS pixel_7015/NB2 pixel_7015/AMP_IN pixel_7015/SF_IB
+ pixel_7015/PIX_OUT pixel_7015/CSA_VREF pixel
Xpixel_7026 pixel_7026/gring pixel_7026/VDD pixel_7026/GND pixel_7026/VREF pixel_7026/ROW_SEL
+ pixel_7026/NB1 pixel_7026/VBIAS pixel_7026/NB2 pixel_7026/AMP_IN pixel_7026/SF_IB
+ pixel_7026/PIX_OUT pixel_7026/CSA_VREF pixel
Xpixel_7037 pixel_7037/gring pixel_7037/VDD pixel_7037/GND pixel_7037/VREF pixel_7037/ROW_SEL
+ pixel_7037/NB1 pixel_7037/VBIAS pixel_7037/NB2 pixel_7037/AMP_IN pixel_7037/SF_IB
+ pixel_7037/PIX_OUT pixel_7037/CSA_VREF pixel
Xpixel_7048 pixel_7048/gring pixel_7048/VDD pixel_7048/GND pixel_7048/VREF pixel_7048/ROW_SEL
+ pixel_7048/NB1 pixel_7048/VBIAS pixel_7048/NB2 pixel_7048/AMP_IN pixel_7048/SF_IB
+ pixel_7048/PIX_OUT pixel_7048/CSA_VREF pixel
Xpixel_7059 pixel_7059/gring pixel_7059/VDD pixel_7059/GND pixel_7059/VREF pixel_7059/ROW_SEL
+ pixel_7059/NB1 pixel_7059/VBIAS pixel_7059/NB2 pixel_7059/AMP_IN pixel_7059/SF_IB
+ pixel_7059/PIX_OUT pixel_7059/CSA_VREF pixel
Xpixel_6303 pixel_6303/gring pixel_6303/VDD pixel_6303/GND pixel_6303/VREF pixel_6303/ROW_SEL
+ pixel_6303/NB1 pixel_6303/VBIAS pixel_6303/NB2 pixel_6303/AMP_IN pixel_6303/SF_IB
+ pixel_6303/PIX_OUT pixel_6303/CSA_VREF pixel
Xpixel_6314 pixel_6314/gring pixel_6314/VDD pixel_6314/GND pixel_6314/VREF pixel_6314/ROW_SEL
+ pixel_6314/NB1 pixel_6314/VBIAS pixel_6314/NB2 pixel_6314/AMP_IN pixel_6314/SF_IB
+ pixel_6314/PIX_OUT pixel_6314/CSA_VREF pixel
Xpixel_6325 pixel_6325/gring pixel_6325/VDD pixel_6325/GND pixel_6325/VREF pixel_6325/ROW_SEL
+ pixel_6325/NB1 pixel_6325/VBIAS pixel_6325/NB2 pixel_6325/AMP_IN pixel_6325/SF_IB
+ pixel_6325/PIX_OUT pixel_6325/CSA_VREF pixel
Xpixel_6336 pixel_6336/gring pixel_6336/VDD pixel_6336/GND pixel_6336/VREF pixel_6336/ROW_SEL
+ pixel_6336/NB1 pixel_6336/VBIAS pixel_6336/NB2 pixel_6336/AMP_IN pixel_6336/SF_IB
+ pixel_6336/PIX_OUT pixel_6336/CSA_VREF pixel
Xpixel_6347 pixel_6347/gring pixel_6347/VDD pixel_6347/GND pixel_6347/VREF pixel_6347/ROW_SEL
+ pixel_6347/NB1 pixel_6347/VBIAS pixel_6347/NB2 pixel_6347/AMP_IN pixel_6347/SF_IB
+ pixel_6347/PIX_OUT pixel_6347/CSA_VREF pixel
Xpixel_6358 pixel_6358/gring pixel_6358/VDD pixel_6358/GND pixel_6358/VREF pixel_6358/ROW_SEL
+ pixel_6358/NB1 pixel_6358/VBIAS pixel_6358/NB2 pixel_6358/AMP_IN pixel_6358/SF_IB
+ pixel_6358/PIX_OUT pixel_6358/CSA_VREF pixel
Xpixel_6369 pixel_6369/gring pixel_6369/VDD pixel_6369/GND pixel_6369/VREF pixel_6369/ROW_SEL
+ pixel_6369/NB1 pixel_6369/VBIAS pixel_6369/NB2 pixel_6369/AMP_IN pixel_6369/SF_IB
+ pixel_6369/PIX_OUT pixel_6369/CSA_VREF pixel
Xpixel_5602 pixel_5602/gring pixel_5602/VDD pixel_5602/GND pixel_5602/VREF pixel_5602/ROW_SEL
+ pixel_5602/NB1 pixel_5602/VBIAS pixel_5602/NB2 pixel_5602/AMP_IN pixel_5602/SF_IB
+ pixel_5602/PIX_OUT pixel_5602/CSA_VREF pixel
Xpixel_5613 pixel_5613/gring pixel_5613/VDD pixel_5613/GND pixel_5613/VREF pixel_5613/ROW_SEL
+ pixel_5613/NB1 pixel_5613/VBIAS pixel_5613/NB2 pixel_5613/AMP_IN pixel_5613/SF_IB
+ pixel_5613/PIX_OUT pixel_5613/CSA_VREF pixel
Xpixel_5624 pixel_5624/gring pixel_5624/VDD pixel_5624/GND pixel_5624/VREF pixel_5624/ROW_SEL
+ pixel_5624/NB1 pixel_5624/VBIAS pixel_5624/NB2 pixel_5624/AMP_IN pixel_5624/SF_IB
+ pixel_5624/PIX_OUT pixel_5624/CSA_VREF pixel
Xpixel_5635 pixel_5635/gring pixel_5635/VDD pixel_5635/GND pixel_5635/VREF pixel_5635/ROW_SEL
+ pixel_5635/NB1 pixel_5635/VBIAS pixel_5635/NB2 pixel_5635/AMP_IN pixel_5635/SF_IB
+ pixel_5635/PIX_OUT pixel_5635/CSA_VREF pixel
Xpixel_5646 pixel_5646/gring pixel_5646/VDD pixel_5646/GND pixel_5646/VREF pixel_5646/ROW_SEL
+ pixel_5646/NB1 pixel_5646/VBIAS pixel_5646/NB2 pixel_5646/AMP_IN pixel_5646/SF_IB
+ pixel_5646/PIX_OUT pixel_5646/CSA_VREF pixel
Xpixel_5657 pixel_5657/gring pixel_5657/VDD pixel_5657/GND pixel_5657/VREF pixel_5657/ROW_SEL
+ pixel_5657/NB1 pixel_5657/VBIAS pixel_5657/NB2 pixel_5657/AMP_IN pixel_5657/SF_IB
+ pixel_5657/PIX_OUT pixel_5657/CSA_VREF pixel
Xpixel_4901 pixel_4901/gring pixel_4901/VDD pixel_4901/GND pixel_4901/VREF pixel_4901/ROW_SEL
+ pixel_4901/NB1 pixel_4901/VBIAS pixel_4901/NB2 pixel_4901/AMP_IN pixel_4901/SF_IB
+ pixel_4901/PIX_OUT pixel_4901/CSA_VREF pixel
Xpixel_4912 pixel_4912/gring pixel_4912/VDD pixel_4912/GND pixel_4912/VREF pixel_4912/ROW_SEL
+ pixel_4912/NB1 pixel_4912/VBIAS pixel_4912/NB2 pixel_4912/AMP_IN pixel_4912/SF_IB
+ pixel_4912/PIX_OUT pixel_4912/CSA_VREF pixel
Xpixel_951 pixel_951/gring pixel_951/VDD pixel_951/GND pixel_951/VREF pixel_951/ROW_SEL
+ pixel_951/NB1 pixel_951/VBIAS pixel_951/NB2 pixel_951/AMP_IN pixel_951/SF_IB pixel_951/PIX_OUT
+ pixel_951/CSA_VREF pixel
Xpixel_940 pixel_940/gring pixel_940/VDD pixel_940/GND pixel_940/VREF pixel_940/ROW_SEL
+ pixel_940/NB1 pixel_940/VBIAS pixel_940/NB2 pixel_940/AMP_IN pixel_940/SF_IB pixel_940/PIX_OUT
+ pixel_940/CSA_VREF pixel
Xpixel_5668 pixel_5668/gring pixel_5668/VDD pixel_5668/GND pixel_5668/VREF pixel_5668/ROW_SEL
+ pixel_5668/NB1 pixel_5668/VBIAS pixel_5668/NB2 pixel_5668/AMP_IN pixel_5668/SF_IB
+ pixel_5668/PIX_OUT pixel_5668/CSA_VREF pixel
Xpixel_5679 pixel_5679/gring pixel_5679/VDD pixel_5679/GND pixel_5679/VREF pixel_5679/ROW_SEL
+ pixel_5679/NB1 pixel_5679/VBIAS pixel_5679/NB2 pixel_5679/AMP_IN pixel_5679/SF_IB
+ pixel_5679/PIX_OUT pixel_5679/CSA_VREF pixel
Xpixel_4923 pixel_4923/gring pixel_4923/VDD pixel_4923/GND pixel_4923/VREF pixel_4923/ROW_SEL
+ pixel_4923/NB1 pixel_4923/VBIAS pixel_4923/NB2 pixel_4923/AMP_IN pixel_4923/SF_IB
+ pixel_4923/PIX_OUT pixel_4923/CSA_VREF pixel
Xpixel_4934 pixel_4934/gring pixel_4934/VDD pixel_4934/GND pixel_4934/VREF pixel_4934/ROW_SEL
+ pixel_4934/NB1 pixel_4934/VBIAS pixel_4934/NB2 pixel_4934/AMP_IN pixel_4934/SF_IB
+ pixel_4934/PIX_OUT pixel_4934/CSA_VREF pixel
Xpixel_4945 pixel_4945/gring pixel_4945/VDD pixel_4945/GND pixel_4945/VREF pixel_4945/ROW_SEL
+ pixel_4945/NB1 pixel_4945/VBIAS pixel_4945/NB2 pixel_4945/AMP_IN pixel_4945/SF_IB
+ pixel_4945/PIX_OUT pixel_4945/CSA_VREF pixel
Xpixel_4956 pixel_4956/gring pixel_4956/VDD pixel_4956/GND pixel_4956/VREF pixel_4956/ROW_SEL
+ pixel_4956/NB1 pixel_4956/VBIAS pixel_4956/NB2 pixel_4956/AMP_IN pixel_4956/SF_IB
+ pixel_4956/PIX_OUT pixel_4956/CSA_VREF pixel
Xpixel_984 pixel_984/gring pixel_984/VDD pixel_984/GND pixel_984/VREF pixel_984/ROW_SEL
+ pixel_984/NB1 pixel_984/VBIAS pixel_984/NB2 pixel_984/AMP_IN pixel_984/SF_IB pixel_984/PIX_OUT
+ pixel_984/CSA_VREF pixel
Xpixel_973 pixel_973/gring pixel_973/VDD pixel_973/GND pixel_973/VREF pixel_973/ROW_SEL
+ pixel_973/NB1 pixel_973/VBIAS pixel_973/NB2 pixel_973/AMP_IN pixel_973/SF_IB pixel_973/PIX_OUT
+ pixel_973/CSA_VREF pixel
Xpixel_962 pixel_962/gring pixel_962/VDD pixel_962/GND pixel_962/VREF pixel_962/ROW_SEL
+ pixel_962/NB1 pixel_962/VBIAS pixel_962/NB2 pixel_962/AMP_IN pixel_962/SF_IB pixel_962/PIX_OUT
+ pixel_962/CSA_VREF pixel
Xpixel_4967 pixel_4967/gring pixel_4967/VDD pixel_4967/GND pixel_4967/VREF pixel_4967/ROW_SEL
+ pixel_4967/NB1 pixel_4967/VBIAS pixel_4967/NB2 pixel_4967/AMP_IN pixel_4967/SF_IB
+ pixel_4967/PIX_OUT pixel_4967/CSA_VREF pixel
Xpixel_4978 pixel_4978/gring pixel_4978/VDD pixel_4978/GND pixel_4978/VREF pixel_4978/ROW_SEL
+ pixel_4978/NB1 pixel_4978/VBIAS pixel_4978/NB2 pixel_4978/AMP_IN pixel_4978/SF_IB
+ pixel_4978/PIX_OUT pixel_4978/CSA_VREF pixel
Xpixel_4989 pixel_4989/gring pixel_4989/VDD pixel_4989/GND pixel_4989/VREF pixel_4989/ROW_SEL
+ pixel_4989/NB1 pixel_4989/VBIAS pixel_4989/NB2 pixel_4989/AMP_IN pixel_4989/SF_IB
+ pixel_4989/PIX_OUT pixel_4989/CSA_VREF pixel
Xpixel_995 pixel_995/gring pixel_995/VDD pixel_995/GND pixel_995/VREF pixel_995/ROW_SEL
+ pixel_995/NB1 pixel_995/VBIAS pixel_995/NB2 pixel_995/AMP_IN pixel_995/SF_IB pixel_995/PIX_OUT
+ pixel_995/CSA_VREF pixel
Xpixel_8250 pixel_8250/gring pixel_8250/VDD pixel_8250/GND pixel_8250/VREF pixel_8250/ROW_SEL
+ pixel_8250/NB1 pixel_8250/VBIAS pixel_8250/NB2 pixel_8250/AMP_IN pixel_8250/SF_IB
+ pixel_8250/PIX_OUT pixel_8250/CSA_VREF pixel
Xpixel_8261 pixel_8261/gring pixel_8261/VDD pixel_8261/GND pixel_8261/VREF pixel_8261/ROW_SEL
+ pixel_8261/NB1 pixel_8261/VBIAS pixel_8261/NB2 pixel_8261/AMP_IN pixel_8261/SF_IB
+ pixel_8261/PIX_OUT pixel_8261/CSA_VREF pixel
Xpixel_8272 pixel_8272/gring pixel_8272/VDD pixel_8272/GND pixel_8272/VREF pixel_8272/ROW_SEL
+ pixel_8272/NB1 pixel_8272/VBIAS pixel_8272/NB2 pixel_8272/AMP_IN pixel_8272/SF_IB
+ pixel_8272/PIX_OUT pixel_8272/CSA_VREF pixel
Xpixel_8283 pixel_8283/gring pixel_8283/VDD pixel_8283/GND pixel_8283/VREF pixel_8283/ROW_SEL
+ pixel_8283/NB1 pixel_8283/VBIAS pixel_8283/NB2 pixel_8283/AMP_IN pixel_8283/SF_IB
+ pixel_8283/PIX_OUT pixel_8283/CSA_VREF pixel
Xpixel_8294 pixel_8294/gring pixel_8294/VDD pixel_8294/GND pixel_8294/VREF pixel_8294/ROW_SEL
+ pixel_8294/NB1 pixel_8294/VBIAS pixel_8294/NB2 pixel_8294/AMP_IN pixel_8294/SF_IB
+ pixel_8294/PIX_OUT pixel_8294/CSA_VREF pixel
Xpixel_7560 pixel_7560/gring pixel_7560/VDD pixel_7560/GND pixel_7560/VREF pixel_7560/ROW_SEL
+ pixel_7560/NB1 pixel_7560/VBIAS pixel_7560/NB2 pixel_7560/AMP_IN pixel_7560/SF_IB
+ pixel_7560/PIX_OUT pixel_7560/CSA_VREF pixel
Xpixel_7571 pixel_7571/gring pixel_7571/VDD pixel_7571/GND pixel_7571/VREF pixel_7571/ROW_SEL
+ pixel_7571/NB1 pixel_7571/VBIAS pixel_7571/NB2 pixel_7571/AMP_IN pixel_7571/SF_IB
+ pixel_7571/PIX_OUT pixel_7571/CSA_VREF pixel
Xpixel_7582 pixel_7582/gring pixel_7582/VDD pixel_7582/GND pixel_7582/VREF pixel_7582/ROW_SEL
+ pixel_7582/NB1 pixel_7582/VBIAS pixel_7582/NB2 pixel_7582/AMP_IN pixel_7582/SF_IB
+ pixel_7582/PIX_OUT pixel_7582/CSA_VREF pixel
Xpixel_7593 pixel_7593/gring pixel_7593/VDD pixel_7593/GND pixel_7593/VREF pixel_7593/ROW_SEL
+ pixel_7593/NB1 pixel_7593/VBIAS pixel_7593/NB2 pixel_7593/AMP_IN pixel_7593/SF_IB
+ pixel_7593/PIX_OUT pixel_7593/CSA_VREF pixel
Xpixel_6870 pixel_6870/gring pixel_6870/VDD pixel_6870/GND pixel_6870/VREF pixel_6870/ROW_SEL
+ pixel_6870/NB1 pixel_6870/VBIAS pixel_6870/NB2 pixel_6870/AMP_IN pixel_6870/SF_IB
+ pixel_6870/PIX_OUT pixel_6870/CSA_VREF pixel
Xpixel_6881 pixel_6881/gring pixel_6881/VDD pixel_6881/GND pixel_6881/VREF pixel_6881/ROW_SEL
+ pixel_6881/NB1 pixel_6881/VBIAS pixel_6881/NB2 pixel_6881/AMP_IN pixel_6881/SF_IB
+ pixel_6881/PIX_OUT pixel_6881/CSA_VREF pixel
Xpixel_6892 pixel_6892/gring pixel_6892/VDD pixel_6892/GND pixel_6892/VREF pixel_6892/ROW_SEL
+ pixel_6892/NB1 pixel_6892/VBIAS pixel_6892/NB2 pixel_6892/AMP_IN pixel_6892/SF_IB
+ pixel_6892/PIX_OUT pixel_6892/CSA_VREF pixel
Xpixel_203 pixel_203/gring pixel_203/VDD pixel_203/GND pixel_203/VREF pixel_203/ROW_SEL
+ pixel_203/NB1 pixel_203/VBIAS pixel_203/NB2 pixel_203/AMP_IN pixel_203/SF_IB pixel_203/PIX_OUT
+ pixel_203/CSA_VREF pixel
Xpixel_4208 pixel_4208/gring pixel_4208/VDD pixel_4208/GND pixel_4208/VREF pixel_4208/ROW_SEL
+ pixel_4208/NB1 pixel_4208/VBIAS pixel_4208/NB2 pixel_4208/AMP_IN pixel_4208/SF_IB
+ pixel_4208/PIX_OUT pixel_4208/CSA_VREF pixel
Xpixel_247 pixel_247/gring pixel_247/VDD pixel_247/GND pixel_247/VREF pixel_247/ROW_SEL
+ pixel_247/NB1 pixel_247/VBIAS pixel_247/NB2 pixel_247/AMP_IN pixel_247/SF_IB pixel_247/PIX_OUT
+ pixel_247/CSA_VREF pixel
Xpixel_236 pixel_236/gring pixel_236/VDD pixel_236/GND pixel_236/VREF pixel_236/ROW_SEL
+ pixel_236/NB1 pixel_236/VBIAS pixel_236/NB2 pixel_236/AMP_IN pixel_236/SF_IB pixel_236/PIX_OUT
+ pixel_236/CSA_VREF pixel
Xpixel_225 pixel_225/gring pixel_225/VDD pixel_225/GND pixel_225/VREF pixel_225/ROW_SEL
+ pixel_225/NB1 pixel_225/VBIAS pixel_225/NB2 pixel_225/AMP_IN pixel_225/SF_IB pixel_225/PIX_OUT
+ pixel_225/CSA_VREF pixel
Xpixel_214 pixel_214/gring pixel_214/VDD pixel_214/GND pixel_214/VREF pixel_214/ROW_SEL
+ pixel_214/NB1 pixel_214/VBIAS pixel_214/NB2 pixel_214/AMP_IN pixel_214/SF_IB pixel_214/PIX_OUT
+ pixel_214/CSA_VREF pixel
Xpixel_3507 pixel_3507/gring pixel_3507/VDD pixel_3507/GND pixel_3507/VREF pixel_3507/ROW_SEL
+ pixel_3507/NB1 pixel_3507/VBIAS pixel_3507/NB2 pixel_3507/AMP_IN pixel_3507/SF_IB
+ pixel_3507/PIX_OUT pixel_3507/CSA_VREF pixel
Xpixel_4219 pixel_4219/gring pixel_4219/VDD pixel_4219/GND pixel_4219/VREF pixel_4219/ROW_SEL
+ pixel_4219/NB1 pixel_4219/VBIAS pixel_4219/NB2 pixel_4219/AMP_IN pixel_4219/SF_IB
+ pixel_4219/PIX_OUT pixel_4219/CSA_VREF pixel
Xpixel_269 pixel_269/gring pixel_269/VDD pixel_269/GND pixel_269/VREF pixel_269/ROW_SEL
+ pixel_269/NB1 pixel_269/VBIAS pixel_269/NB2 pixel_269/AMP_IN pixel_269/SF_IB pixel_269/PIX_OUT
+ pixel_269/CSA_VREF pixel
Xpixel_258 pixel_258/gring pixel_258/VDD pixel_258/GND pixel_258/VREF pixel_258/ROW_SEL
+ pixel_258/NB1 pixel_258/VBIAS pixel_258/NB2 pixel_258/AMP_IN pixel_258/SF_IB pixel_258/PIX_OUT
+ pixel_258/CSA_VREF pixel
Xpixel_3529 pixel_3529/gring pixel_3529/VDD pixel_3529/GND pixel_3529/VREF pixel_3529/ROW_SEL
+ pixel_3529/NB1 pixel_3529/VBIAS pixel_3529/NB2 pixel_3529/AMP_IN pixel_3529/SF_IB
+ pixel_3529/PIX_OUT pixel_3529/CSA_VREF pixel
Xpixel_3518 pixel_3518/gring pixel_3518/VDD pixel_3518/GND pixel_3518/VREF pixel_3518/ROW_SEL
+ pixel_3518/NB1 pixel_3518/VBIAS pixel_3518/NB2 pixel_3518/AMP_IN pixel_3518/SF_IB
+ pixel_3518/PIX_OUT pixel_3518/CSA_VREF pixel
Xpixel_2828 pixel_2828/gring pixel_2828/VDD pixel_2828/GND pixel_2828/VREF pixel_2828/ROW_SEL
+ pixel_2828/NB1 pixel_2828/VBIAS pixel_2828/NB2 pixel_2828/AMP_IN pixel_2828/SF_IB
+ pixel_2828/PIX_OUT pixel_2828/CSA_VREF pixel
Xpixel_2817 pixel_2817/gring pixel_2817/VDD pixel_2817/GND pixel_2817/VREF pixel_2817/ROW_SEL
+ pixel_2817/NB1 pixel_2817/VBIAS pixel_2817/NB2 pixel_2817/AMP_IN pixel_2817/SF_IB
+ pixel_2817/PIX_OUT pixel_2817/CSA_VREF pixel
Xpixel_2806 pixel_2806/gring pixel_2806/VDD pixel_2806/GND pixel_2806/VREF pixel_2806/ROW_SEL
+ pixel_2806/NB1 pixel_2806/VBIAS pixel_2806/NB2 pixel_2806/AMP_IN pixel_2806/SF_IB
+ pixel_2806/PIX_OUT pixel_2806/CSA_VREF pixel
Xpixel_2839 pixel_2839/gring pixel_2839/VDD pixel_2839/GND pixel_2839/VREF pixel_2839/ROW_SEL
+ pixel_2839/NB1 pixel_2839/VBIAS pixel_2839/NB2 pixel_2839/AMP_IN pixel_2839/SF_IB
+ pixel_2839/PIX_OUT pixel_2839/CSA_VREF pixel
Xpixel_6100 pixel_6100/gring pixel_6100/VDD pixel_6100/GND pixel_6100/VREF pixel_6100/ROW_SEL
+ pixel_6100/NB1 pixel_6100/VBIAS pixel_6100/NB2 pixel_6100/AMP_IN pixel_6100/SF_IB
+ pixel_6100/PIX_OUT pixel_6100/CSA_VREF pixel
Xpixel_6111 pixel_6111/gring pixel_6111/VDD pixel_6111/GND pixel_6111/VREF pixel_6111/ROW_SEL
+ pixel_6111/NB1 pixel_6111/VBIAS pixel_6111/NB2 pixel_6111/AMP_IN pixel_6111/SF_IB
+ pixel_6111/PIX_OUT pixel_6111/CSA_VREF pixel
Xpixel_6122 pixel_6122/gring pixel_6122/VDD pixel_6122/GND pixel_6122/VREF pixel_6122/ROW_SEL
+ pixel_6122/NB1 pixel_6122/VBIAS pixel_6122/NB2 pixel_6122/AMP_IN pixel_6122/SF_IB
+ pixel_6122/PIX_OUT pixel_6122/CSA_VREF pixel
Xpixel_6133 pixel_6133/gring pixel_6133/VDD pixel_6133/GND pixel_6133/VREF pixel_6133/ROW_SEL
+ pixel_6133/NB1 pixel_6133/VBIAS pixel_6133/NB2 pixel_6133/AMP_IN pixel_6133/SF_IB
+ pixel_6133/PIX_OUT pixel_6133/CSA_VREF pixel
Xpixel_6144 pixel_6144/gring pixel_6144/VDD pixel_6144/GND pixel_6144/VREF pixel_6144/ROW_SEL
+ pixel_6144/NB1 pixel_6144/VBIAS pixel_6144/NB2 pixel_6144/AMP_IN pixel_6144/SF_IB
+ pixel_6144/PIX_OUT pixel_6144/CSA_VREF pixel
Xpixel_6155 pixel_6155/gring pixel_6155/VDD pixel_6155/GND pixel_6155/VREF pixel_6155/ROW_SEL
+ pixel_6155/NB1 pixel_6155/VBIAS pixel_6155/NB2 pixel_6155/AMP_IN pixel_6155/SF_IB
+ pixel_6155/PIX_OUT pixel_6155/CSA_VREF pixel
Xpixel_6166 pixel_6166/gring pixel_6166/VDD pixel_6166/GND pixel_6166/VREF pixel_6166/ROW_SEL
+ pixel_6166/NB1 pixel_6166/VBIAS pixel_6166/NB2 pixel_6166/AMP_IN pixel_6166/SF_IB
+ pixel_6166/PIX_OUT pixel_6166/CSA_VREF pixel
Xpixel_6177 pixel_6177/gring pixel_6177/VDD pixel_6177/GND pixel_6177/VREF pixel_6177/ROW_SEL
+ pixel_6177/NB1 pixel_6177/VBIAS pixel_6177/NB2 pixel_6177/AMP_IN pixel_6177/SF_IB
+ pixel_6177/PIX_OUT pixel_6177/CSA_VREF pixel
Xpixel_5410 pixel_5410/gring pixel_5410/VDD pixel_5410/GND pixel_5410/VREF pixel_5410/ROW_SEL
+ pixel_5410/NB1 pixel_5410/VBIAS pixel_5410/NB2 pixel_5410/AMP_IN pixel_5410/SF_IB
+ pixel_5410/PIX_OUT pixel_5410/CSA_VREF pixel
Xpixel_5421 pixel_5421/gring pixel_5421/VDD pixel_5421/GND pixel_5421/VREF pixel_5421/ROW_SEL
+ pixel_5421/NB1 pixel_5421/VBIAS pixel_5421/NB2 pixel_5421/AMP_IN pixel_5421/SF_IB
+ pixel_5421/PIX_OUT pixel_5421/CSA_VREF pixel
Xpixel_5432 pixel_5432/gring pixel_5432/VDD pixel_5432/GND pixel_5432/VREF pixel_5432/ROW_SEL
+ pixel_5432/NB1 pixel_5432/VBIAS pixel_5432/NB2 pixel_5432/AMP_IN pixel_5432/SF_IB
+ pixel_5432/PIX_OUT pixel_5432/CSA_VREF pixel
Xpixel_6188 pixel_6188/gring pixel_6188/VDD pixel_6188/GND pixel_6188/VREF pixel_6188/ROW_SEL
+ pixel_6188/NB1 pixel_6188/VBIAS pixel_6188/NB2 pixel_6188/AMP_IN pixel_6188/SF_IB
+ pixel_6188/PIX_OUT pixel_6188/CSA_VREF pixel
Xpixel_6199 pixel_6199/gring pixel_6199/VDD pixel_6199/GND pixel_6199/VREF pixel_6199/ROW_SEL
+ pixel_6199/NB1 pixel_6199/VBIAS pixel_6199/NB2 pixel_6199/AMP_IN pixel_6199/SF_IB
+ pixel_6199/PIX_OUT pixel_6199/CSA_VREF pixel
Xpixel_5443 pixel_5443/gring pixel_5443/VDD pixel_5443/GND pixel_5443/VREF pixel_5443/ROW_SEL
+ pixel_5443/NB1 pixel_5443/VBIAS pixel_5443/NB2 pixel_5443/AMP_IN pixel_5443/SF_IB
+ pixel_5443/PIX_OUT pixel_5443/CSA_VREF pixel
Xpixel_5454 pixel_5454/gring pixel_5454/VDD pixel_5454/GND pixel_5454/VREF pixel_5454/ROW_SEL
+ pixel_5454/NB1 pixel_5454/VBIAS pixel_5454/NB2 pixel_5454/AMP_IN pixel_5454/SF_IB
+ pixel_5454/PIX_OUT pixel_5454/CSA_VREF pixel
Xpixel_5465 pixel_5465/gring pixel_5465/VDD pixel_5465/GND pixel_5465/VREF pixel_5465/ROW_SEL
+ pixel_5465/NB1 pixel_5465/VBIAS pixel_5465/NB2 pixel_5465/AMP_IN pixel_5465/SF_IB
+ pixel_5465/PIX_OUT pixel_5465/CSA_VREF pixel
Xpixel_4720 pixel_4720/gring pixel_4720/VDD pixel_4720/GND pixel_4720/VREF pixel_4720/ROW_SEL
+ pixel_4720/NB1 pixel_4720/VBIAS pixel_4720/NB2 pixel_4720/AMP_IN pixel_4720/SF_IB
+ pixel_4720/PIX_OUT pixel_4720/CSA_VREF pixel
Xpixel_4731 pixel_4731/gring pixel_4731/VDD pixel_4731/GND pixel_4731/VREF pixel_4731/ROW_SEL
+ pixel_4731/NB1 pixel_4731/VBIAS pixel_4731/NB2 pixel_4731/AMP_IN pixel_4731/SF_IB
+ pixel_4731/PIX_OUT pixel_4731/CSA_VREF pixel
Xpixel_5476 pixel_5476/gring pixel_5476/VDD pixel_5476/GND pixel_5476/VREF pixel_5476/ROW_SEL
+ pixel_5476/NB1 pixel_5476/VBIAS pixel_5476/NB2 pixel_5476/AMP_IN pixel_5476/SF_IB
+ pixel_5476/PIX_OUT pixel_5476/CSA_VREF pixel
Xpixel_5487 pixel_5487/gring pixel_5487/VDD pixel_5487/GND pixel_5487/VREF pixel_5487/ROW_SEL
+ pixel_5487/NB1 pixel_5487/VBIAS pixel_5487/NB2 pixel_5487/AMP_IN pixel_5487/SF_IB
+ pixel_5487/PIX_OUT pixel_5487/CSA_VREF pixel
Xpixel_5498 pixel_5498/gring pixel_5498/VDD pixel_5498/GND pixel_5498/VREF pixel_5498/ROW_SEL
+ pixel_5498/NB1 pixel_5498/VBIAS pixel_5498/NB2 pixel_5498/AMP_IN pixel_5498/SF_IB
+ pixel_5498/PIX_OUT pixel_5498/CSA_VREF pixel
Xpixel_4742 pixel_4742/gring pixel_4742/VDD pixel_4742/GND pixel_4742/VREF pixel_4742/ROW_SEL
+ pixel_4742/NB1 pixel_4742/VBIAS pixel_4742/NB2 pixel_4742/AMP_IN pixel_4742/SF_IB
+ pixel_4742/PIX_OUT pixel_4742/CSA_VREF pixel
Xpixel_4753 pixel_4753/gring pixel_4753/VDD pixel_4753/GND pixel_4753/VREF pixel_4753/ROW_SEL
+ pixel_4753/NB1 pixel_4753/VBIAS pixel_4753/NB2 pixel_4753/AMP_IN pixel_4753/SF_IB
+ pixel_4753/PIX_OUT pixel_4753/CSA_VREF pixel
Xpixel_4764 pixel_4764/gring pixel_4764/VDD pixel_4764/GND pixel_4764/VREF pixel_4764/ROW_SEL
+ pixel_4764/NB1 pixel_4764/VBIAS pixel_4764/NB2 pixel_4764/AMP_IN pixel_4764/SF_IB
+ pixel_4764/PIX_OUT pixel_4764/CSA_VREF pixel
Xpixel_792 pixel_792/gring pixel_792/VDD pixel_792/GND pixel_792/VREF pixel_792/ROW_SEL
+ pixel_792/NB1 pixel_792/VBIAS pixel_792/NB2 pixel_792/AMP_IN pixel_792/SF_IB pixel_792/PIX_OUT
+ pixel_792/CSA_VREF pixel
Xpixel_781 pixel_781/gring pixel_781/VDD pixel_781/GND pixel_781/VREF pixel_781/ROW_SEL
+ pixel_781/NB1 pixel_781/VBIAS pixel_781/NB2 pixel_781/AMP_IN pixel_781/SF_IB pixel_781/PIX_OUT
+ pixel_781/CSA_VREF pixel
Xpixel_770 pixel_770/gring pixel_770/VDD pixel_770/GND pixel_770/VREF pixel_770/ROW_SEL
+ pixel_770/NB1 pixel_770/VBIAS pixel_770/NB2 pixel_770/AMP_IN pixel_770/SF_IB pixel_770/PIX_OUT
+ pixel_770/CSA_VREF pixel
Xpixel_4775 pixel_4775/gring pixel_4775/VDD pixel_4775/GND pixel_4775/VREF pixel_4775/ROW_SEL
+ pixel_4775/NB1 pixel_4775/VBIAS pixel_4775/NB2 pixel_4775/AMP_IN pixel_4775/SF_IB
+ pixel_4775/PIX_OUT pixel_4775/CSA_VREF pixel
Xpixel_4786 pixel_4786/gring pixel_4786/VDD pixel_4786/GND pixel_4786/VREF pixel_4786/ROW_SEL
+ pixel_4786/NB1 pixel_4786/VBIAS pixel_4786/NB2 pixel_4786/AMP_IN pixel_4786/SF_IB
+ pixel_4786/PIX_OUT pixel_4786/CSA_VREF pixel
Xpixel_4797 pixel_4797/gring pixel_4797/VDD pixel_4797/GND pixel_4797/VREF pixel_4797/ROW_SEL
+ pixel_4797/NB1 pixel_4797/VBIAS pixel_4797/NB2 pixel_4797/AMP_IN pixel_4797/SF_IB
+ pixel_4797/PIX_OUT pixel_4797/CSA_VREF pixel
Xpixel_8080 pixel_8080/gring pixel_8080/VDD pixel_8080/GND pixel_8080/VREF pixel_8080/ROW_SEL
+ pixel_8080/NB1 pixel_8080/VBIAS pixel_8080/NB2 pixel_8080/AMP_IN pixel_8080/SF_IB
+ pixel_8080/PIX_OUT pixel_8080/CSA_VREF pixel
Xpixel_8091 pixel_8091/gring pixel_8091/VDD pixel_8091/GND pixel_8091/VREF pixel_8091/ROW_SEL
+ pixel_8091/NB1 pixel_8091/VBIAS pixel_8091/NB2 pixel_8091/AMP_IN pixel_8091/SF_IB
+ pixel_8091/PIX_OUT pixel_8091/CSA_VREF pixel
Xpixel_7390 pixel_7390/gring pixel_7390/VDD pixel_7390/GND pixel_7390/VREF pixel_7390/ROW_SEL
+ pixel_7390/NB1 pixel_7390/VBIAS pixel_7390/NB2 pixel_7390/AMP_IN pixel_7390/SF_IB
+ pixel_7390/PIX_OUT pixel_7390/CSA_VREF pixel
Xpixel_9709 pixel_9709/gring pixel_9709/VDD pixel_9709/GND pixel_9709/VREF pixel_9709/ROW_SEL
+ pixel_9709/NB1 pixel_9709/VBIAS pixel_9709/NB2 pixel_9709/AMP_IN pixel_9709/SF_IB
+ pixel_9709/PIX_OUT pixel_9709/CSA_VREF pixel
Xpixel_4005 pixel_4005/gring pixel_4005/VDD pixel_4005/GND pixel_4005/VREF pixel_4005/ROW_SEL
+ pixel_4005/NB1 pixel_4005/VBIAS pixel_4005/NB2 pixel_4005/AMP_IN pixel_4005/SF_IB
+ pixel_4005/PIX_OUT pixel_4005/CSA_VREF pixel
Xpixel_4016 pixel_4016/gring pixel_4016/VDD pixel_4016/GND pixel_4016/VREF pixel_4016/ROW_SEL
+ pixel_4016/NB1 pixel_4016/VBIAS pixel_4016/NB2 pixel_4016/AMP_IN pixel_4016/SF_IB
+ pixel_4016/PIX_OUT pixel_4016/CSA_VREF pixel
Xpixel_3315 pixel_3315/gring pixel_3315/VDD pixel_3315/GND pixel_3315/VREF pixel_3315/ROW_SEL
+ pixel_3315/NB1 pixel_3315/VBIAS pixel_3315/NB2 pixel_3315/AMP_IN pixel_3315/SF_IB
+ pixel_3315/PIX_OUT pixel_3315/CSA_VREF pixel
Xpixel_3304 pixel_3304/gring pixel_3304/VDD pixel_3304/GND pixel_3304/VREF pixel_3304/ROW_SEL
+ pixel_3304/NB1 pixel_3304/VBIAS pixel_3304/NB2 pixel_3304/AMP_IN pixel_3304/SF_IB
+ pixel_3304/PIX_OUT pixel_3304/CSA_VREF pixel
Xpixel_4027 pixel_4027/gring pixel_4027/VDD pixel_4027/GND pixel_4027/VREF pixel_4027/ROW_SEL
+ pixel_4027/NB1 pixel_4027/VBIAS pixel_4027/NB2 pixel_4027/AMP_IN pixel_4027/SF_IB
+ pixel_4027/PIX_OUT pixel_4027/CSA_VREF pixel
Xpixel_4038 pixel_4038/gring pixel_4038/VDD pixel_4038/GND pixel_4038/VREF pixel_4038/ROW_SEL
+ pixel_4038/NB1 pixel_4038/VBIAS pixel_4038/NB2 pixel_4038/AMP_IN pixel_4038/SF_IB
+ pixel_4038/PIX_OUT pixel_4038/CSA_VREF pixel
Xpixel_4049 pixel_4049/gring pixel_4049/VDD pixel_4049/GND pixel_4049/VREF pixel_4049/ROW_SEL
+ pixel_4049/NB1 pixel_4049/VBIAS pixel_4049/NB2 pixel_4049/AMP_IN pixel_4049/SF_IB
+ pixel_4049/PIX_OUT pixel_4049/CSA_VREF pixel
Xpixel_2603 pixel_2603/gring pixel_2603/VDD pixel_2603/GND pixel_2603/VREF pixel_2603/ROW_SEL
+ pixel_2603/NB1 pixel_2603/VBIAS pixel_2603/NB2 pixel_2603/AMP_IN pixel_2603/SF_IB
+ pixel_2603/PIX_OUT pixel_2603/CSA_VREF pixel
Xpixel_3348 pixel_3348/gring pixel_3348/VDD pixel_3348/GND pixel_3348/VREF pixel_3348/ROW_SEL
+ pixel_3348/NB1 pixel_3348/VBIAS pixel_3348/NB2 pixel_3348/AMP_IN pixel_3348/SF_IB
+ pixel_3348/PIX_OUT pixel_3348/CSA_VREF pixel
Xpixel_3337 pixel_3337/gring pixel_3337/VDD pixel_3337/GND pixel_3337/VREF pixel_3337/ROW_SEL
+ pixel_3337/NB1 pixel_3337/VBIAS pixel_3337/NB2 pixel_3337/AMP_IN pixel_3337/SF_IB
+ pixel_3337/PIX_OUT pixel_3337/CSA_VREF pixel
Xpixel_3326 pixel_3326/gring pixel_3326/VDD pixel_3326/GND pixel_3326/VREF pixel_3326/ROW_SEL
+ pixel_3326/NB1 pixel_3326/VBIAS pixel_3326/NB2 pixel_3326/AMP_IN pixel_3326/SF_IB
+ pixel_3326/PIX_OUT pixel_3326/CSA_VREF pixel
Xpixel_1902 pixel_1902/gring pixel_1902/VDD pixel_1902/GND pixel_1902/VREF pixel_1902/ROW_SEL
+ pixel_1902/NB1 pixel_1902/VBIAS pixel_1902/NB2 pixel_1902/AMP_IN pixel_1902/SF_IB
+ pixel_1902/PIX_OUT pixel_1902/CSA_VREF pixel
Xpixel_2636 pixel_2636/gring pixel_2636/VDD pixel_2636/GND pixel_2636/VREF pixel_2636/ROW_SEL
+ pixel_2636/NB1 pixel_2636/VBIAS pixel_2636/NB2 pixel_2636/AMP_IN pixel_2636/SF_IB
+ pixel_2636/PIX_OUT pixel_2636/CSA_VREF pixel
Xpixel_2625 pixel_2625/gring pixel_2625/VDD pixel_2625/GND pixel_2625/VREF pixel_2625/ROW_SEL
+ pixel_2625/NB1 pixel_2625/VBIAS pixel_2625/NB2 pixel_2625/AMP_IN pixel_2625/SF_IB
+ pixel_2625/PIX_OUT pixel_2625/CSA_VREF pixel
Xpixel_2614 pixel_2614/gring pixel_2614/VDD pixel_2614/GND pixel_2614/VREF pixel_2614/ROW_SEL
+ pixel_2614/NB1 pixel_2614/VBIAS pixel_2614/NB2 pixel_2614/AMP_IN pixel_2614/SF_IB
+ pixel_2614/PIX_OUT pixel_2614/CSA_VREF pixel
Xpixel_3359 pixel_3359/gring pixel_3359/VDD pixel_3359/GND pixel_3359/VREF pixel_3359/ROW_SEL
+ pixel_3359/NB1 pixel_3359/VBIAS pixel_3359/NB2 pixel_3359/AMP_IN pixel_3359/SF_IB
+ pixel_3359/PIX_OUT pixel_3359/CSA_VREF pixel
Xpixel_1935 pixel_1935/gring pixel_1935/VDD pixel_1935/GND pixel_1935/VREF pixel_1935/ROW_SEL
+ pixel_1935/NB1 pixel_1935/VBIAS pixel_1935/NB2 pixel_1935/AMP_IN pixel_1935/SF_IB
+ pixel_1935/PIX_OUT pixel_1935/CSA_VREF pixel
Xpixel_1924 pixel_1924/gring pixel_1924/VDD pixel_1924/GND pixel_1924/VREF pixel_1924/ROW_SEL
+ pixel_1924/NB1 pixel_1924/VBIAS pixel_1924/NB2 pixel_1924/AMP_IN pixel_1924/SF_IB
+ pixel_1924/PIX_OUT pixel_1924/CSA_VREF pixel
Xpixel_1913 pixel_1913/gring pixel_1913/VDD pixel_1913/GND pixel_1913/VREF pixel_1913/ROW_SEL
+ pixel_1913/NB1 pixel_1913/VBIAS pixel_1913/NB2 pixel_1913/AMP_IN pixel_1913/SF_IB
+ pixel_1913/PIX_OUT pixel_1913/CSA_VREF pixel
Xpixel_2669 pixel_2669/gring pixel_2669/VDD pixel_2669/GND pixel_2669/VREF pixel_2669/ROW_SEL
+ pixel_2669/NB1 pixel_2669/VBIAS pixel_2669/NB2 pixel_2669/AMP_IN pixel_2669/SF_IB
+ pixel_2669/PIX_OUT pixel_2669/CSA_VREF pixel
Xpixel_2658 pixel_2658/gring pixel_2658/VDD pixel_2658/GND pixel_2658/VREF pixel_2658/ROW_SEL
+ pixel_2658/NB1 pixel_2658/VBIAS pixel_2658/NB2 pixel_2658/AMP_IN pixel_2658/SF_IB
+ pixel_2658/PIX_OUT pixel_2658/CSA_VREF pixel
Xpixel_2647 pixel_2647/gring pixel_2647/VDD pixel_2647/GND pixel_2647/VREF pixel_2647/ROW_SEL
+ pixel_2647/NB1 pixel_2647/VBIAS pixel_2647/NB2 pixel_2647/AMP_IN pixel_2647/SF_IB
+ pixel_2647/PIX_OUT pixel_2647/CSA_VREF pixel
Xpixel_1968 pixel_1968/gring pixel_1968/VDD pixel_1968/GND pixel_1968/VREF pixel_1968/ROW_SEL
+ pixel_1968/NB1 pixel_1968/VBIAS pixel_1968/NB2 pixel_1968/AMP_IN pixel_1968/SF_IB
+ pixel_1968/PIX_OUT pixel_1968/CSA_VREF pixel
Xpixel_1957 pixel_1957/gring pixel_1957/VDD pixel_1957/GND pixel_1957/VREF pixel_1957/ROW_SEL
+ pixel_1957/NB1 pixel_1957/VBIAS pixel_1957/NB2 pixel_1957/AMP_IN pixel_1957/SF_IB
+ pixel_1957/PIX_OUT pixel_1957/CSA_VREF pixel
Xpixel_1946 pixel_1946/gring pixel_1946/VDD pixel_1946/GND pixel_1946/VREF pixel_1946/ROW_SEL
+ pixel_1946/NB1 pixel_1946/VBIAS pixel_1946/NB2 pixel_1946/AMP_IN pixel_1946/SF_IB
+ pixel_1946/PIX_OUT pixel_1946/CSA_VREF pixel
Xpixel_1979 pixel_1979/gring pixel_1979/VDD pixel_1979/GND pixel_1979/VREF pixel_1979/ROW_SEL
+ pixel_1979/NB1 pixel_1979/VBIAS pixel_1979/NB2 pixel_1979/AMP_IN pixel_1979/SF_IB
+ pixel_1979/PIX_OUT pixel_1979/CSA_VREF pixel
Xpixel_5240 pixel_5240/gring pixel_5240/VDD pixel_5240/GND pixel_5240/VREF pixel_5240/ROW_SEL
+ pixel_5240/NB1 pixel_5240/VBIAS pixel_5240/NB2 pixel_5240/AMP_IN pixel_5240/SF_IB
+ pixel_5240/PIX_OUT pixel_5240/CSA_VREF pixel
Xpixel_5251 pixel_5251/gring pixel_5251/VDD pixel_5251/GND pixel_5251/VREF pixel_5251/ROW_SEL
+ pixel_5251/NB1 pixel_5251/VBIAS pixel_5251/NB2 pixel_5251/AMP_IN pixel_5251/SF_IB
+ pixel_5251/PIX_OUT pixel_5251/CSA_VREF pixel
Xpixel_5262 pixel_5262/gring pixel_5262/VDD pixel_5262/GND pixel_5262/VREF pixel_5262/ROW_SEL
+ pixel_5262/NB1 pixel_5262/VBIAS pixel_5262/NB2 pixel_5262/AMP_IN pixel_5262/SF_IB
+ pixel_5262/PIX_OUT pixel_5262/CSA_VREF pixel
Xpixel_5273 pixel_5273/gring pixel_5273/VDD pixel_5273/GND pixel_5273/VREF pixel_5273/ROW_SEL
+ pixel_5273/NB1 pixel_5273/VBIAS pixel_5273/NB2 pixel_5273/AMP_IN pixel_5273/SF_IB
+ pixel_5273/PIX_OUT pixel_5273/CSA_VREF pixel
Xpixel_5284 pixel_5284/gring pixel_5284/VDD pixel_5284/GND pixel_5284/VREF pixel_5284/ROW_SEL
+ pixel_5284/NB1 pixel_5284/VBIAS pixel_5284/NB2 pixel_5284/AMP_IN pixel_5284/SF_IB
+ pixel_5284/PIX_OUT pixel_5284/CSA_VREF pixel
Xpixel_5295 pixel_5295/gring pixel_5295/VDD pixel_5295/GND pixel_5295/VREF pixel_5295/ROW_SEL
+ pixel_5295/NB1 pixel_5295/VBIAS pixel_5295/NB2 pixel_5295/AMP_IN pixel_5295/SF_IB
+ pixel_5295/PIX_OUT pixel_5295/CSA_VREF pixel
Xpixel_4550 pixel_4550/gring pixel_4550/VDD pixel_4550/GND pixel_4550/VREF pixel_4550/ROW_SEL
+ pixel_4550/NB1 pixel_4550/VBIAS pixel_4550/NB2 pixel_4550/AMP_IN pixel_4550/SF_IB
+ pixel_4550/PIX_OUT pixel_4550/CSA_VREF pixel
Xpixel_4561 pixel_4561/gring pixel_4561/VDD pixel_4561/GND pixel_4561/VREF pixel_4561/ROW_SEL
+ pixel_4561/NB1 pixel_4561/VBIAS pixel_4561/NB2 pixel_4561/AMP_IN pixel_4561/SF_IB
+ pixel_4561/PIX_OUT pixel_4561/CSA_VREF pixel
Xpixel_4572 pixel_4572/gring pixel_4572/VDD pixel_4572/GND pixel_4572/VREF pixel_4572/ROW_SEL
+ pixel_4572/NB1 pixel_4572/VBIAS pixel_4572/NB2 pixel_4572/AMP_IN pixel_4572/SF_IB
+ pixel_4572/PIX_OUT pixel_4572/CSA_VREF pixel
Xpixel_3871 pixel_3871/gring pixel_3871/VDD pixel_3871/GND pixel_3871/VREF pixel_3871/ROW_SEL
+ pixel_3871/NB1 pixel_3871/VBIAS pixel_3871/NB2 pixel_3871/AMP_IN pixel_3871/SF_IB
+ pixel_3871/PIX_OUT pixel_3871/CSA_VREF pixel
Xpixel_3860 pixel_3860/gring pixel_3860/VDD pixel_3860/GND pixel_3860/VREF pixel_3860/ROW_SEL
+ pixel_3860/NB1 pixel_3860/VBIAS pixel_3860/NB2 pixel_3860/AMP_IN pixel_3860/SF_IB
+ pixel_3860/PIX_OUT pixel_3860/CSA_VREF pixel
Xpixel_4583 pixel_4583/gring pixel_4583/VDD pixel_4583/GND pixel_4583/VREF pixel_4583/ROW_SEL
+ pixel_4583/NB1 pixel_4583/VBIAS pixel_4583/NB2 pixel_4583/AMP_IN pixel_4583/SF_IB
+ pixel_4583/PIX_OUT pixel_4583/CSA_VREF pixel
Xpixel_4594 pixel_4594/gring pixel_4594/VDD pixel_4594/GND pixel_4594/VREF pixel_4594/ROW_SEL
+ pixel_4594/NB1 pixel_4594/VBIAS pixel_4594/NB2 pixel_4594/AMP_IN pixel_4594/SF_IB
+ pixel_4594/PIX_OUT pixel_4594/CSA_VREF pixel
Xpixel_3893 pixel_3893/gring pixel_3893/VDD pixel_3893/GND pixel_3893/VREF pixel_3893/ROW_SEL
+ pixel_3893/NB1 pixel_3893/VBIAS pixel_3893/NB2 pixel_3893/AMP_IN pixel_3893/SF_IB
+ pixel_3893/PIX_OUT pixel_3893/CSA_VREF pixel
Xpixel_3882 pixel_3882/gring pixel_3882/VDD pixel_3882/GND pixel_3882/VREF pixel_3882/ROW_SEL
+ pixel_3882/NB1 pixel_3882/VBIAS pixel_3882/NB2 pixel_3882/AMP_IN pixel_3882/SF_IB
+ pixel_3882/PIX_OUT pixel_3882/CSA_VREF pixel
Xpixel_1209 pixel_1209/gring pixel_1209/VDD pixel_1209/GND pixel_1209/VREF pixel_1209/ROW_SEL
+ pixel_1209/NB1 pixel_1209/VBIAS pixel_1209/NB2 pixel_1209/AMP_IN pixel_1209/SF_IB
+ pixel_1209/PIX_OUT pixel_1209/CSA_VREF pixel
Xpixel_9539 pixel_9539/gring pixel_9539/VDD pixel_9539/GND pixel_9539/VREF pixel_9539/ROW_SEL
+ pixel_9539/NB1 pixel_9539/VBIAS pixel_9539/NB2 pixel_9539/AMP_IN pixel_9539/SF_IB
+ pixel_9539/PIX_OUT pixel_9539/CSA_VREF pixel
Xpixel_9528 pixel_9528/gring pixel_9528/VDD pixel_9528/GND pixel_9528/VREF pixel_9528/ROW_SEL
+ pixel_9528/NB1 pixel_9528/VBIAS pixel_9528/NB2 pixel_9528/AMP_IN pixel_9528/SF_IB
+ pixel_9528/PIX_OUT pixel_9528/CSA_VREF pixel
Xpixel_9517 pixel_9517/gring pixel_9517/VDD pixel_9517/GND pixel_9517/VREF pixel_9517/ROW_SEL
+ pixel_9517/NB1 pixel_9517/VBIAS pixel_9517/NB2 pixel_9517/AMP_IN pixel_9517/SF_IB
+ pixel_9517/PIX_OUT pixel_9517/CSA_VREF pixel
Xpixel_9506 pixel_9506/gring pixel_9506/VDD pixel_9506/GND pixel_9506/VREF pixel_9506/ROW_SEL
+ pixel_9506/NB1 pixel_9506/VBIAS pixel_9506/NB2 pixel_9506/AMP_IN pixel_9506/SF_IB
+ pixel_9506/PIX_OUT pixel_9506/CSA_VREF pixel
Xpixel_8827 pixel_8827/gring pixel_8827/VDD pixel_8827/GND pixel_8827/VREF pixel_8827/ROW_SEL
+ pixel_8827/NB1 pixel_8827/VBIAS pixel_8827/NB2 pixel_8827/AMP_IN pixel_8827/SF_IB
+ pixel_8827/PIX_OUT pixel_8827/CSA_VREF pixel
Xpixel_8816 pixel_8816/gring pixel_8816/VDD pixel_8816/GND pixel_8816/VREF pixel_8816/ROW_SEL
+ pixel_8816/NB1 pixel_8816/VBIAS pixel_8816/NB2 pixel_8816/AMP_IN pixel_8816/SF_IB
+ pixel_8816/PIX_OUT pixel_8816/CSA_VREF pixel
Xpixel_8805 pixel_8805/gring pixel_8805/VDD pixel_8805/GND pixel_8805/VREF pixel_8805/ROW_SEL
+ pixel_8805/NB1 pixel_8805/VBIAS pixel_8805/NB2 pixel_8805/AMP_IN pixel_8805/SF_IB
+ pixel_8805/PIX_OUT pixel_8805/CSA_VREF pixel
Xpixel_8849 pixel_8849/gring pixel_8849/VDD pixel_8849/GND pixel_8849/VREF pixel_8849/ROW_SEL
+ pixel_8849/NB1 pixel_8849/VBIAS pixel_8849/NB2 pixel_8849/AMP_IN pixel_8849/SF_IB
+ pixel_8849/PIX_OUT pixel_8849/CSA_VREF pixel
Xpixel_8838 pixel_8838/gring pixel_8838/VDD pixel_8838/GND pixel_8838/VREF pixel_8838/ROW_SEL
+ pixel_8838/NB1 pixel_8838/VBIAS pixel_8838/NB2 pixel_8838/AMP_IN pixel_8838/SF_IB
+ pixel_8838/PIX_OUT pixel_8838/CSA_VREF pixel
Xpixel_3123 pixel_3123/gring pixel_3123/VDD pixel_3123/GND pixel_3123/VREF pixel_3123/ROW_SEL
+ pixel_3123/NB1 pixel_3123/VBIAS pixel_3123/NB2 pixel_3123/AMP_IN pixel_3123/SF_IB
+ pixel_3123/PIX_OUT pixel_3123/CSA_VREF pixel
Xpixel_3112 pixel_3112/gring pixel_3112/VDD pixel_3112/GND pixel_3112/VREF pixel_3112/ROW_SEL
+ pixel_3112/NB1 pixel_3112/VBIAS pixel_3112/NB2 pixel_3112/AMP_IN pixel_3112/SF_IB
+ pixel_3112/PIX_OUT pixel_3112/CSA_VREF pixel
Xpixel_3101 pixel_3101/gring pixel_3101/VDD pixel_3101/GND pixel_3101/VREF pixel_3101/ROW_SEL
+ pixel_3101/NB1 pixel_3101/VBIAS pixel_3101/NB2 pixel_3101/AMP_IN pixel_3101/SF_IB
+ pixel_3101/PIX_OUT pixel_3101/CSA_VREF pixel
Xpixel_2411 pixel_2411/gring pixel_2411/VDD pixel_2411/GND pixel_2411/VREF pixel_2411/ROW_SEL
+ pixel_2411/NB1 pixel_2411/VBIAS pixel_2411/NB2 pixel_2411/AMP_IN pixel_2411/SF_IB
+ pixel_2411/PIX_OUT pixel_2411/CSA_VREF pixel
Xpixel_2400 pixel_2400/gring pixel_2400/VDD pixel_2400/GND pixel_2400/VREF pixel_2400/ROW_SEL
+ pixel_2400/NB1 pixel_2400/VBIAS pixel_2400/NB2 pixel_2400/AMP_IN pixel_2400/SF_IB
+ pixel_2400/PIX_OUT pixel_2400/CSA_VREF pixel
Xpixel_3156 pixel_3156/gring pixel_3156/VDD pixel_3156/GND pixel_3156/VREF pixel_3156/ROW_SEL
+ pixel_3156/NB1 pixel_3156/VBIAS pixel_3156/NB2 pixel_3156/AMP_IN pixel_3156/SF_IB
+ pixel_3156/PIX_OUT pixel_3156/CSA_VREF pixel
Xpixel_3145 pixel_3145/gring pixel_3145/VDD pixel_3145/GND pixel_3145/VREF pixel_3145/ROW_SEL
+ pixel_3145/NB1 pixel_3145/VBIAS pixel_3145/NB2 pixel_3145/AMP_IN pixel_3145/SF_IB
+ pixel_3145/PIX_OUT pixel_3145/CSA_VREF pixel
Xpixel_3134 pixel_3134/gring pixel_3134/VDD pixel_3134/GND pixel_3134/VREF pixel_3134/ROW_SEL
+ pixel_3134/NB1 pixel_3134/VBIAS pixel_3134/NB2 pixel_3134/AMP_IN pixel_3134/SF_IB
+ pixel_3134/PIX_OUT pixel_3134/CSA_VREF pixel
Xpixel_1710 pixel_1710/gring pixel_1710/VDD pixel_1710/GND pixel_1710/VREF pixel_1710/ROW_SEL
+ pixel_1710/NB1 pixel_1710/VBIAS pixel_1710/NB2 pixel_1710/AMP_IN pixel_1710/SF_IB
+ pixel_1710/PIX_OUT pixel_1710/CSA_VREF pixel
Xpixel_2455 pixel_2455/gring pixel_2455/VDD pixel_2455/GND pixel_2455/VREF pixel_2455/ROW_SEL
+ pixel_2455/NB1 pixel_2455/VBIAS pixel_2455/NB2 pixel_2455/AMP_IN pixel_2455/SF_IB
+ pixel_2455/PIX_OUT pixel_2455/CSA_VREF pixel
Xpixel_2444 pixel_2444/gring pixel_2444/VDD pixel_2444/GND pixel_2444/VREF pixel_2444/ROW_SEL
+ pixel_2444/NB1 pixel_2444/VBIAS pixel_2444/NB2 pixel_2444/AMP_IN pixel_2444/SF_IB
+ pixel_2444/PIX_OUT pixel_2444/CSA_VREF pixel
Xpixel_2433 pixel_2433/gring pixel_2433/VDD pixel_2433/GND pixel_2433/VREF pixel_2433/ROW_SEL
+ pixel_2433/NB1 pixel_2433/VBIAS pixel_2433/NB2 pixel_2433/AMP_IN pixel_2433/SF_IB
+ pixel_2433/PIX_OUT pixel_2433/CSA_VREF pixel
Xpixel_2422 pixel_2422/gring pixel_2422/VDD pixel_2422/GND pixel_2422/VREF pixel_2422/ROW_SEL
+ pixel_2422/NB1 pixel_2422/VBIAS pixel_2422/NB2 pixel_2422/AMP_IN pixel_2422/SF_IB
+ pixel_2422/PIX_OUT pixel_2422/CSA_VREF pixel
Xpixel_3189 pixel_3189/gring pixel_3189/VDD pixel_3189/GND pixel_3189/VREF pixel_3189/ROW_SEL
+ pixel_3189/NB1 pixel_3189/VBIAS pixel_3189/NB2 pixel_3189/AMP_IN pixel_3189/SF_IB
+ pixel_3189/PIX_OUT pixel_3189/CSA_VREF pixel
Xpixel_3178 pixel_3178/gring pixel_3178/VDD pixel_3178/GND pixel_3178/VREF pixel_3178/ROW_SEL
+ pixel_3178/NB1 pixel_3178/VBIAS pixel_3178/NB2 pixel_3178/AMP_IN pixel_3178/SF_IB
+ pixel_3178/PIX_OUT pixel_3178/CSA_VREF pixel
Xpixel_3167 pixel_3167/gring pixel_3167/VDD pixel_3167/GND pixel_3167/VREF pixel_3167/ROW_SEL
+ pixel_3167/NB1 pixel_3167/VBIAS pixel_3167/NB2 pixel_3167/AMP_IN pixel_3167/SF_IB
+ pixel_3167/PIX_OUT pixel_3167/CSA_VREF pixel
Xpixel_1743 pixel_1743/gring pixel_1743/VDD pixel_1743/GND pixel_1743/VREF pixel_1743/ROW_SEL
+ pixel_1743/NB1 pixel_1743/VBIAS pixel_1743/NB2 pixel_1743/AMP_IN pixel_1743/SF_IB
+ pixel_1743/PIX_OUT pixel_1743/CSA_VREF pixel
Xpixel_1732 pixel_1732/gring pixel_1732/VDD pixel_1732/GND pixel_1732/VREF pixel_1732/ROW_SEL
+ pixel_1732/NB1 pixel_1732/VBIAS pixel_1732/NB2 pixel_1732/AMP_IN pixel_1732/SF_IB
+ pixel_1732/PIX_OUT pixel_1732/CSA_VREF pixel
Xpixel_1721 pixel_1721/gring pixel_1721/VDD pixel_1721/GND pixel_1721/VREF pixel_1721/ROW_SEL
+ pixel_1721/NB1 pixel_1721/VBIAS pixel_1721/NB2 pixel_1721/AMP_IN pixel_1721/SF_IB
+ pixel_1721/PIX_OUT pixel_1721/CSA_VREF pixel
Xpixel_2488 pixel_2488/gring pixel_2488/VDD pixel_2488/GND pixel_2488/VREF pixel_2488/ROW_SEL
+ pixel_2488/NB1 pixel_2488/VBIAS pixel_2488/NB2 pixel_2488/AMP_IN pixel_2488/SF_IB
+ pixel_2488/PIX_OUT pixel_2488/CSA_VREF pixel
Xpixel_2477 pixel_2477/gring pixel_2477/VDD pixel_2477/GND pixel_2477/VREF pixel_2477/ROW_SEL
+ pixel_2477/NB1 pixel_2477/VBIAS pixel_2477/NB2 pixel_2477/AMP_IN pixel_2477/SF_IB
+ pixel_2477/PIX_OUT pixel_2477/CSA_VREF pixel
Xpixel_2466 pixel_2466/gring pixel_2466/VDD pixel_2466/GND pixel_2466/VREF pixel_2466/ROW_SEL
+ pixel_2466/NB1 pixel_2466/VBIAS pixel_2466/NB2 pixel_2466/AMP_IN pixel_2466/SF_IB
+ pixel_2466/PIX_OUT pixel_2466/CSA_VREF pixel
Xpixel_1776 pixel_1776/gring pixel_1776/VDD pixel_1776/GND pixel_1776/VREF pixel_1776/ROW_SEL
+ pixel_1776/NB1 pixel_1776/VBIAS pixel_1776/NB2 pixel_1776/AMP_IN pixel_1776/SF_IB
+ pixel_1776/PIX_OUT pixel_1776/CSA_VREF pixel
Xpixel_1765 pixel_1765/gring pixel_1765/VDD pixel_1765/GND pixel_1765/VREF pixel_1765/ROW_SEL
+ pixel_1765/NB1 pixel_1765/VBIAS pixel_1765/NB2 pixel_1765/AMP_IN pixel_1765/SF_IB
+ pixel_1765/PIX_OUT pixel_1765/CSA_VREF pixel
Xpixel_1754 pixel_1754/gring pixel_1754/VDD pixel_1754/GND pixel_1754/VREF pixel_1754/ROW_SEL
+ pixel_1754/NB1 pixel_1754/VBIAS pixel_1754/NB2 pixel_1754/AMP_IN pixel_1754/SF_IB
+ pixel_1754/PIX_OUT pixel_1754/CSA_VREF pixel
Xpixel_2499 pixel_2499/gring pixel_2499/VDD pixel_2499/GND pixel_2499/VREF pixel_2499/ROW_SEL
+ pixel_2499/NB1 pixel_2499/VBIAS pixel_2499/NB2 pixel_2499/AMP_IN pixel_2499/SF_IB
+ pixel_2499/PIX_OUT pixel_2499/CSA_VREF pixel
Xpixel_1798 pixel_1798/gring pixel_1798/VDD pixel_1798/GND pixel_1798/VREF pixel_1798/ROW_SEL
+ pixel_1798/NB1 pixel_1798/VBIAS pixel_1798/NB2 pixel_1798/AMP_IN pixel_1798/SF_IB
+ pixel_1798/PIX_OUT pixel_1798/CSA_VREF pixel
Xpixel_1787 pixel_1787/gring pixel_1787/VDD pixel_1787/GND pixel_1787/VREF pixel_1787/ROW_SEL
+ pixel_1787/NB1 pixel_1787/VBIAS pixel_1787/NB2 pixel_1787/AMP_IN pixel_1787/SF_IB
+ pixel_1787/PIX_OUT pixel_1787/CSA_VREF pixel
Xpixel_5070 pixel_5070/gring pixel_5070/VDD pixel_5070/GND pixel_5070/VREF pixel_5070/ROW_SEL
+ pixel_5070/NB1 pixel_5070/VBIAS pixel_5070/NB2 pixel_5070/AMP_IN pixel_5070/SF_IB
+ pixel_5070/PIX_OUT pixel_5070/CSA_VREF pixel
Xpixel_5081 pixel_5081/gring pixel_5081/VDD pixel_5081/GND pixel_5081/VREF pixel_5081/ROW_SEL
+ pixel_5081/NB1 pixel_5081/VBIAS pixel_5081/NB2 pixel_5081/AMP_IN pixel_5081/SF_IB
+ pixel_5081/PIX_OUT pixel_5081/CSA_VREF pixel
Xpixel_5092 pixel_5092/gring pixel_5092/VDD pixel_5092/GND pixel_5092/VREF pixel_5092/ROW_SEL
+ pixel_5092/NB1 pixel_5092/VBIAS pixel_5092/NB2 pixel_5092/AMP_IN pixel_5092/SF_IB
+ pixel_5092/PIX_OUT pixel_5092/CSA_VREF pixel
Xpixel_4380 pixel_4380/gring pixel_4380/VDD pixel_4380/GND pixel_4380/VREF pixel_4380/ROW_SEL
+ pixel_4380/NB1 pixel_4380/VBIAS pixel_4380/NB2 pixel_4380/AMP_IN pixel_4380/SF_IB
+ pixel_4380/PIX_OUT pixel_4380/CSA_VREF pixel
Xpixel_4391 pixel_4391/gring pixel_4391/VDD pixel_4391/GND pixel_4391/VREF pixel_4391/ROW_SEL
+ pixel_4391/NB1 pixel_4391/VBIAS pixel_4391/NB2 pixel_4391/AMP_IN pixel_4391/SF_IB
+ pixel_4391/PIX_OUT pixel_4391/CSA_VREF pixel
Xpixel_3690 pixel_3690/gring pixel_3690/VDD pixel_3690/GND pixel_3690/VREF pixel_3690/ROW_SEL
+ pixel_3690/NB1 pixel_3690/VBIAS pixel_3690/NB2 pixel_3690/AMP_IN pixel_3690/SF_IB
+ pixel_3690/PIX_OUT pixel_3690/CSA_VREF pixel
Xpixel_1039 pixel_1039/gring pixel_1039/VDD pixel_1039/GND pixel_1039/VREF pixel_1039/ROW_SEL
+ pixel_1039/NB1 pixel_1039/VBIAS pixel_1039/NB2 pixel_1039/AMP_IN pixel_1039/SF_IB
+ pixel_1039/PIX_OUT pixel_1039/CSA_VREF pixel
Xpixel_1028 pixel_1028/gring pixel_1028/VDD pixel_1028/GND pixel_1028/VREF pixel_1028/ROW_SEL
+ pixel_1028/NB1 pixel_1028/VBIAS pixel_1028/NB2 pixel_1028/AMP_IN pixel_1028/SF_IB
+ pixel_1028/PIX_OUT pixel_1028/CSA_VREF pixel
Xpixel_1017 pixel_1017/gring pixel_1017/VDD pixel_1017/GND pixel_1017/VREF pixel_1017/ROW_SEL
+ pixel_1017/NB1 pixel_1017/VBIAS pixel_1017/NB2 pixel_1017/AMP_IN pixel_1017/SF_IB
+ pixel_1017/PIX_OUT pixel_1017/CSA_VREF pixel
Xpixel_1006 pixel_1006/gring pixel_1006/VDD pixel_1006/GND pixel_1006/VREF pixel_1006/ROW_SEL
+ pixel_1006/NB1 pixel_1006/VBIAS pixel_1006/NB2 pixel_1006/AMP_IN pixel_1006/SF_IB
+ pixel_1006/PIX_OUT pixel_1006/CSA_VREF pixel
Xpixel_9303 pixel_9303/gring pixel_9303/VDD pixel_9303/GND pixel_9303/VREF pixel_9303/ROW_SEL
+ pixel_9303/NB1 pixel_9303/VBIAS pixel_9303/NB2 pixel_9303/AMP_IN pixel_9303/SF_IB
+ pixel_9303/PIX_OUT pixel_9303/CSA_VREF pixel
Xpixel_8602 pixel_8602/gring pixel_8602/VDD pixel_8602/GND pixel_8602/VREF pixel_8602/ROW_SEL
+ pixel_8602/NB1 pixel_8602/VBIAS pixel_8602/NB2 pixel_8602/AMP_IN pixel_8602/SF_IB
+ pixel_8602/PIX_OUT pixel_8602/CSA_VREF pixel
Xpixel_9347 pixel_9347/gring pixel_9347/VDD pixel_9347/GND pixel_9347/VREF pixel_9347/ROW_SEL
+ pixel_9347/NB1 pixel_9347/VBIAS pixel_9347/NB2 pixel_9347/AMP_IN pixel_9347/SF_IB
+ pixel_9347/PIX_OUT pixel_9347/CSA_VREF pixel
Xpixel_9336 pixel_9336/gring pixel_9336/VDD pixel_9336/GND pixel_9336/VREF pixel_9336/ROW_SEL
+ pixel_9336/NB1 pixel_9336/VBIAS pixel_9336/NB2 pixel_9336/AMP_IN pixel_9336/SF_IB
+ pixel_9336/PIX_OUT pixel_9336/CSA_VREF pixel
Xpixel_9325 pixel_9325/gring pixel_9325/VDD pixel_9325/GND pixel_9325/VREF pixel_9325/ROW_SEL
+ pixel_9325/NB1 pixel_9325/VBIAS pixel_9325/NB2 pixel_9325/AMP_IN pixel_9325/SF_IB
+ pixel_9325/PIX_OUT pixel_9325/CSA_VREF pixel
Xpixel_9314 pixel_9314/gring pixel_9314/VDD pixel_9314/GND pixel_9314/VREF pixel_9314/ROW_SEL
+ pixel_9314/NB1 pixel_9314/VBIAS pixel_9314/NB2 pixel_9314/AMP_IN pixel_9314/SF_IB
+ pixel_9314/PIX_OUT pixel_9314/CSA_VREF pixel
Xpixel_8635 pixel_8635/gring pixel_8635/VDD pixel_8635/GND pixel_8635/VREF pixel_8635/ROW_SEL
+ pixel_8635/NB1 pixel_8635/VBIAS pixel_8635/NB2 pixel_8635/AMP_IN pixel_8635/SF_IB
+ pixel_8635/PIX_OUT pixel_8635/CSA_VREF pixel
Xpixel_8624 pixel_8624/gring pixel_8624/VDD pixel_8624/GND pixel_8624/VREF pixel_8624/ROW_SEL
+ pixel_8624/NB1 pixel_8624/VBIAS pixel_8624/NB2 pixel_8624/AMP_IN pixel_8624/SF_IB
+ pixel_8624/PIX_OUT pixel_8624/CSA_VREF pixel
Xpixel_8613 pixel_8613/gring pixel_8613/VDD pixel_8613/GND pixel_8613/VREF pixel_8613/ROW_SEL
+ pixel_8613/NB1 pixel_8613/VBIAS pixel_8613/NB2 pixel_8613/AMP_IN pixel_8613/SF_IB
+ pixel_8613/PIX_OUT pixel_8613/CSA_VREF pixel
Xpixel_9369 pixel_9369/gring pixel_9369/VDD pixel_9369/GND pixel_9369/VREF pixel_9369/ROW_SEL
+ pixel_9369/NB1 pixel_9369/VBIAS pixel_9369/NB2 pixel_9369/AMP_IN pixel_9369/SF_IB
+ pixel_9369/PIX_OUT pixel_9369/CSA_VREF pixel
Xpixel_9358 pixel_9358/gring pixel_9358/VDD pixel_9358/GND pixel_9358/VREF pixel_9358/ROW_SEL
+ pixel_9358/NB1 pixel_9358/VBIAS pixel_9358/NB2 pixel_9358/AMP_IN pixel_9358/SF_IB
+ pixel_9358/PIX_OUT pixel_9358/CSA_VREF pixel
Xpixel_8679 pixel_8679/gring pixel_8679/VDD pixel_8679/GND pixel_8679/VREF pixel_8679/ROW_SEL
+ pixel_8679/NB1 pixel_8679/VBIAS pixel_8679/NB2 pixel_8679/AMP_IN pixel_8679/SF_IB
+ pixel_8679/PIX_OUT pixel_8679/CSA_VREF pixel
Xpixel_8668 pixel_8668/gring pixel_8668/VDD pixel_8668/GND pixel_8668/VREF pixel_8668/ROW_SEL
+ pixel_8668/NB1 pixel_8668/VBIAS pixel_8668/NB2 pixel_8668/AMP_IN pixel_8668/SF_IB
+ pixel_8668/PIX_OUT pixel_8668/CSA_VREF pixel
Xpixel_8657 pixel_8657/gring pixel_8657/VDD pixel_8657/GND pixel_8657/VREF pixel_8657/ROW_SEL
+ pixel_8657/NB1 pixel_8657/VBIAS pixel_8657/NB2 pixel_8657/AMP_IN pixel_8657/SF_IB
+ pixel_8657/PIX_OUT pixel_8657/CSA_VREF pixel
Xpixel_8646 pixel_8646/gring pixel_8646/VDD pixel_8646/GND pixel_8646/VREF pixel_8646/ROW_SEL
+ pixel_8646/NB1 pixel_8646/VBIAS pixel_8646/NB2 pixel_8646/AMP_IN pixel_8646/SF_IB
+ pixel_8646/PIX_OUT pixel_8646/CSA_VREF pixel
Xpixel_7901 pixel_7901/gring pixel_7901/VDD pixel_7901/GND pixel_7901/VREF pixel_7901/ROW_SEL
+ pixel_7901/NB1 pixel_7901/VBIAS pixel_7901/NB2 pixel_7901/AMP_IN pixel_7901/SF_IB
+ pixel_7901/PIX_OUT pixel_7901/CSA_VREF pixel
Xpixel_7912 pixel_7912/gring pixel_7912/VDD pixel_7912/GND pixel_7912/VREF pixel_7912/ROW_SEL
+ pixel_7912/NB1 pixel_7912/VBIAS pixel_7912/NB2 pixel_7912/AMP_IN pixel_7912/SF_IB
+ pixel_7912/PIX_OUT pixel_7912/CSA_VREF pixel
Xpixel_7923 pixel_7923/gring pixel_7923/VDD pixel_7923/GND pixel_7923/VREF pixel_7923/ROW_SEL
+ pixel_7923/NB1 pixel_7923/VBIAS pixel_7923/NB2 pixel_7923/AMP_IN pixel_7923/SF_IB
+ pixel_7923/PIX_OUT pixel_7923/CSA_VREF pixel
Xpixel_7934 pixel_7934/gring pixel_7934/VDD pixel_7934/GND pixel_7934/VREF pixel_7934/ROW_SEL
+ pixel_7934/NB1 pixel_7934/VBIAS pixel_7934/NB2 pixel_7934/AMP_IN pixel_7934/SF_IB
+ pixel_7934/PIX_OUT pixel_7934/CSA_VREF pixel
Xpixel_7945 pixel_7945/gring pixel_7945/VDD pixel_7945/GND pixel_7945/VREF pixel_7945/ROW_SEL
+ pixel_7945/NB1 pixel_7945/VBIAS pixel_7945/NB2 pixel_7945/AMP_IN pixel_7945/SF_IB
+ pixel_7945/PIX_OUT pixel_7945/CSA_VREF pixel
Xpixel_7956 pixel_7956/gring pixel_7956/VDD pixel_7956/GND pixel_7956/VREF pixel_7956/ROW_SEL
+ pixel_7956/NB1 pixel_7956/VBIAS pixel_7956/NB2 pixel_7956/AMP_IN pixel_7956/SF_IB
+ pixel_7956/PIX_OUT pixel_7956/CSA_VREF pixel
Xpixel_7967 pixel_7967/gring pixel_7967/VDD pixel_7967/GND pixel_7967/VREF pixel_7967/ROW_SEL
+ pixel_7967/NB1 pixel_7967/VBIAS pixel_7967/NB2 pixel_7967/AMP_IN pixel_7967/SF_IB
+ pixel_7967/PIX_OUT pixel_7967/CSA_VREF pixel
Xpixel_7978 pixel_7978/gring pixel_7978/VDD pixel_7978/GND pixel_7978/VREF pixel_7978/ROW_SEL
+ pixel_7978/NB1 pixel_7978/VBIAS pixel_7978/NB2 pixel_7978/AMP_IN pixel_7978/SF_IB
+ pixel_7978/PIX_OUT pixel_7978/CSA_VREF pixel
Xpixel_7989 pixel_7989/gring pixel_7989/VDD pixel_7989/GND pixel_7989/VREF pixel_7989/ROW_SEL
+ pixel_7989/NB1 pixel_7989/VBIAS pixel_7989/NB2 pixel_7989/AMP_IN pixel_7989/SF_IB
+ pixel_7989/PIX_OUT pixel_7989/CSA_VREF pixel
Xpixel_2230 pixel_2230/gring pixel_2230/VDD pixel_2230/GND pixel_2230/VREF pixel_2230/ROW_SEL
+ pixel_2230/NB1 pixel_2230/VBIAS pixel_2230/NB2 pixel_2230/AMP_IN pixel_2230/SF_IB
+ pixel_2230/PIX_OUT pixel_2230/CSA_VREF pixel
Xpixel_2263 pixel_2263/gring pixel_2263/VDD pixel_2263/GND pixel_2263/VREF pixel_2263/ROW_SEL
+ pixel_2263/NB1 pixel_2263/VBIAS pixel_2263/NB2 pixel_2263/AMP_IN pixel_2263/SF_IB
+ pixel_2263/PIX_OUT pixel_2263/CSA_VREF pixel
Xpixel_2252 pixel_2252/gring pixel_2252/VDD pixel_2252/GND pixel_2252/VREF pixel_2252/ROW_SEL
+ pixel_2252/NB1 pixel_2252/VBIAS pixel_2252/NB2 pixel_2252/AMP_IN pixel_2252/SF_IB
+ pixel_2252/PIX_OUT pixel_2252/CSA_VREF pixel
Xpixel_2241 pixel_2241/gring pixel_2241/VDD pixel_2241/GND pixel_2241/VREF pixel_2241/ROW_SEL
+ pixel_2241/NB1 pixel_2241/VBIAS pixel_2241/NB2 pixel_2241/AMP_IN pixel_2241/SF_IB
+ pixel_2241/PIX_OUT pixel_2241/CSA_VREF pixel
Xpixel_1551 pixel_1551/gring pixel_1551/VDD pixel_1551/GND pixel_1551/VREF pixel_1551/ROW_SEL
+ pixel_1551/NB1 pixel_1551/VBIAS pixel_1551/NB2 pixel_1551/AMP_IN pixel_1551/SF_IB
+ pixel_1551/PIX_OUT pixel_1551/CSA_VREF pixel
Xpixel_1540 pixel_1540/gring pixel_1540/VDD pixel_1540/GND pixel_1540/VREF pixel_1540/ROW_SEL
+ pixel_1540/NB1 pixel_1540/VBIAS pixel_1540/NB2 pixel_1540/AMP_IN pixel_1540/SF_IB
+ pixel_1540/PIX_OUT pixel_1540/CSA_VREF pixel
Xpixel_2296 pixel_2296/gring pixel_2296/VDD pixel_2296/GND pixel_2296/VREF pixel_2296/ROW_SEL
+ pixel_2296/NB1 pixel_2296/VBIAS pixel_2296/NB2 pixel_2296/AMP_IN pixel_2296/SF_IB
+ pixel_2296/PIX_OUT pixel_2296/CSA_VREF pixel
Xpixel_2285 pixel_2285/gring pixel_2285/VDD pixel_2285/GND pixel_2285/VREF pixel_2285/ROW_SEL
+ pixel_2285/NB1 pixel_2285/VBIAS pixel_2285/NB2 pixel_2285/AMP_IN pixel_2285/SF_IB
+ pixel_2285/PIX_OUT pixel_2285/CSA_VREF pixel
Xpixel_2274 pixel_2274/gring pixel_2274/VDD pixel_2274/GND pixel_2274/VREF pixel_2274/ROW_SEL
+ pixel_2274/NB1 pixel_2274/VBIAS pixel_2274/NB2 pixel_2274/AMP_IN pixel_2274/SF_IB
+ pixel_2274/PIX_OUT pixel_2274/CSA_VREF pixel
Xpixel_1595 pixel_1595/gring pixel_1595/VDD pixel_1595/GND pixel_1595/VREF pixel_1595/ROW_SEL
+ pixel_1595/NB1 pixel_1595/VBIAS pixel_1595/NB2 pixel_1595/AMP_IN pixel_1595/SF_IB
+ pixel_1595/PIX_OUT pixel_1595/CSA_VREF pixel
Xpixel_1584 pixel_1584/gring pixel_1584/VDD pixel_1584/GND pixel_1584/VREF pixel_1584/ROW_SEL
+ pixel_1584/NB1 pixel_1584/VBIAS pixel_1584/NB2 pixel_1584/AMP_IN pixel_1584/SF_IB
+ pixel_1584/PIX_OUT pixel_1584/CSA_VREF pixel
Xpixel_1573 pixel_1573/gring pixel_1573/VDD pixel_1573/GND pixel_1573/VREF pixel_1573/ROW_SEL
+ pixel_1573/NB1 pixel_1573/VBIAS pixel_1573/NB2 pixel_1573/AMP_IN pixel_1573/SF_IB
+ pixel_1573/PIX_OUT pixel_1573/CSA_VREF pixel
Xpixel_1562 pixel_1562/gring pixel_1562/VDD pixel_1562/GND pixel_1562/VREF pixel_1562/ROW_SEL
+ pixel_1562/NB1 pixel_1562/VBIAS pixel_1562/NB2 pixel_1562/AMP_IN pixel_1562/SF_IB
+ pixel_1562/PIX_OUT pixel_1562/CSA_VREF pixel
Xpixel_9870 pixel_9870/gring pixel_9870/VDD pixel_9870/GND pixel_9870/VREF pixel_9870/ROW_SEL
+ pixel_9870/NB1 pixel_9870/VBIAS pixel_9870/NB2 pixel_9870/AMP_IN pixel_9870/SF_IB
+ pixel_9870/PIX_OUT pixel_9870/CSA_VREF pixel
Xpixel_9881 pixel_9881/gring pixel_9881/VDD pixel_9881/GND pixel_9881/VREF pixel_9881/ROW_SEL
+ pixel_9881/NB1 pixel_9881/VBIAS pixel_9881/NB2 pixel_9881/AMP_IN pixel_9881/SF_IB
+ pixel_9881/PIX_OUT pixel_9881/CSA_VREF pixel
Xpixel_9892 pixel_9892/gring pixel_9892/VDD pixel_9892/GND pixel_9892/VREF pixel_9892/ROW_SEL
+ pixel_9892/NB1 pixel_9892/VBIAS pixel_9892/NB2 pixel_9892/AMP_IN pixel_9892/SF_IB
+ pixel_9892/PIX_OUT pixel_9892/CSA_VREF pixel
Xpixel_7208 pixel_7208/gring pixel_7208/VDD pixel_7208/GND pixel_7208/VREF pixel_7208/ROW_SEL
+ pixel_7208/NB1 pixel_7208/VBIAS pixel_7208/NB2 pixel_7208/AMP_IN pixel_7208/SF_IB
+ pixel_7208/PIX_OUT pixel_7208/CSA_VREF pixel
Xpixel_7219 pixel_7219/gring pixel_7219/VDD pixel_7219/GND pixel_7219/VREF pixel_7219/ROW_SEL
+ pixel_7219/NB1 pixel_7219/VBIAS pixel_7219/NB2 pixel_7219/AMP_IN pixel_7219/SF_IB
+ pixel_7219/PIX_OUT pixel_7219/CSA_VREF pixel
Xpixel_6507 pixel_6507/gring pixel_6507/VDD pixel_6507/GND pixel_6507/VREF pixel_6507/ROW_SEL
+ pixel_6507/NB1 pixel_6507/VBIAS pixel_6507/NB2 pixel_6507/AMP_IN pixel_6507/SF_IB
+ pixel_6507/PIX_OUT pixel_6507/CSA_VREF pixel
Xpixel_6518 pixel_6518/gring pixel_6518/VDD pixel_6518/GND pixel_6518/VREF pixel_6518/ROW_SEL
+ pixel_6518/NB1 pixel_6518/VBIAS pixel_6518/NB2 pixel_6518/AMP_IN pixel_6518/SF_IB
+ pixel_6518/PIX_OUT pixel_6518/CSA_VREF pixel
Xpixel_6529 pixel_6529/gring pixel_6529/VDD pixel_6529/GND pixel_6529/VREF pixel_6529/ROW_SEL
+ pixel_6529/NB1 pixel_6529/VBIAS pixel_6529/NB2 pixel_6529/AMP_IN pixel_6529/SF_IB
+ pixel_6529/PIX_OUT pixel_6529/CSA_VREF pixel
Xpixel_5806 pixel_5806/gring pixel_5806/VDD pixel_5806/GND pixel_5806/VREF pixel_5806/ROW_SEL
+ pixel_5806/NB1 pixel_5806/VBIAS pixel_5806/NB2 pixel_5806/AMP_IN pixel_5806/SF_IB
+ pixel_5806/PIX_OUT pixel_5806/CSA_VREF pixel
Xpixel_5817 pixel_5817/gring pixel_5817/VDD pixel_5817/GND pixel_5817/VREF pixel_5817/ROW_SEL
+ pixel_5817/NB1 pixel_5817/VBIAS pixel_5817/NB2 pixel_5817/AMP_IN pixel_5817/SF_IB
+ pixel_5817/PIX_OUT pixel_5817/CSA_VREF pixel
Xpixel_5828 pixel_5828/gring pixel_5828/VDD pixel_5828/GND pixel_5828/VREF pixel_5828/ROW_SEL
+ pixel_5828/NB1 pixel_5828/VBIAS pixel_5828/NB2 pixel_5828/AMP_IN pixel_5828/SF_IB
+ pixel_5828/PIX_OUT pixel_5828/CSA_VREF pixel
Xpixel_5839 pixel_5839/gring pixel_5839/VDD pixel_5839/GND pixel_5839/VREF pixel_5839/ROW_SEL
+ pixel_5839/NB1 pixel_5839/VBIAS pixel_5839/NB2 pixel_5839/AMP_IN pixel_5839/SF_IB
+ pixel_5839/PIX_OUT pixel_5839/CSA_VREF pixel
Xpixel_9122 pixel_9122/gring pixel_9122/VDD pixel_9122/GND pixel_9122/VREF pixel_9122/ROW_SEL
+ pixel_9122/NB1 pixel_9122/VBIAS pixel_9122/NB2 pixel_9122/AMP_IN pixel_9122/SF_IB
+ pixel_9122/PIX_OUT pixel_9122/CSA_VREF pixel
Xpixel_9111 pixel_9111/gring pixel_9111/VDD pixel_9111/GND pixel_9111/VREF pixel_9111/ROW_SEL
+ pixel_9111/NB1 pixel_9111/VBIAS pixel_9111/NB2 pixel_9111/AMP_IN pixel_9111/SF_IB
+ pixel_9111/PIX_OUT pixel_9111/CSA_VREF pixel
Xpixel_9100 pixel_9100/gring pixel_9100/VDD pixel_9100/GND pixel_9100/VREF pixel_9100/ROW_SEL
+ pixel_9100/NB1 pixel_9100/VBIAS pixel_9100/NB2 pixel_9100/AMP_IN pixel_9100/SF_IB
+ pixel_9100/PIX_OUT pixel_9100/CSA_VREF pixel
Xpixel_8410 pixel_8410/gring pixel_8410/VDD pixel_8410/GND pixel_8410/VREF pixel_8410/ROW_SEL
+ pixel_8410/NB1 pixel_8410/VBIAS pixel_8410/NB2 pixel_8410/AMP_IN pixel_8410/SF_IB
+ pixel_8410/PIX_OUT pixel_8410/CSA_VREF pixel
Xpixel_9155 pixel_9155/gring pixel_9155/VDD pixel_9155/GND pixel_9155/VREF pixel_9155/ROW_SEL
+ pixel_9155/NB1 pixel_9155/VBIAS pixel_9155/NB2 pixel_9155/AMP_IN pixel_9155/SF_IB
+ pixel_9155/PIX_OUT pixel_9155/CSA_VREF pixel
Xpixel_9144 pixel_9144/gring pixel_9144/VDD pixel_9144/GND pixel_9144/VREF pixel_9144/ROW_SEL
+ pixel_9144/NB1 pixel_9144/VBIAS pixel_9144/NB2 pixel_9144/AMP_IN pixel_9144/SF_IB
+ pixel_9144/PIX_OUT pixel_9144/CSA_VREF pixel
Xpixel_9133 pixel_9133/gring pixel_9133/VDD pixel_9133/GND pixel_9133/VREF pixel_9133/ROW_SEL
+ pixel_9133/NB1 pixel_9133/VBIAS pixel_9133/NB2 pixel_9133/AMP_IN pixel_9133/SF_IB
+ pixel_9133/PIX_OUT pixel_9133/CSA_VREF pixel
Xpixel_8432 pixel_8432/gring pixel_8432/VDD pixel_8432/GND pixel_8432/VREF pixel_8432/ROW_SEL
+ pixel_8432/NB1 pixel_8432/VBIAS pixel_8432/NB2 pixel_8432/AMP_IN pixel_8432/SF_IB
+ pixel_8432/PIX_OUT pixel_8432/CSA_VREF pixel
Xpixel_8421 pixel_8421/gring pixel_8421/VDD pixel_8421/GND pixel_8421/VREF pixel_8421/ROW_SEL
+ pixel_8421/NB1 pixel_8421/VBIAS pixel_8421/NB2 pixel_8421/AMP_IN pixel_8421/SF_IB
+ pixel_8421/PIX_OUT pixel_8421/CSA_VREF pixel
Xpixel_9188 pixel_9188/gring pixel_9188/VDD pixel_9188/GND pixel_9188/VREF pixel_9188/ROW_SEL
+ pixel_9188/NB1 pixel_9188/VBIAS pixel_9188/NB2 pixel_9188/AMP_IN pixel_9188/SF_IB
+ pixel_9188/PIX_OUT pixel_9188/CSA_VREF pixel
Xpixel_9177 pixel_9177/gring pixel_9177/VDD pixel_9177/GND pixel_9177/VREF pixel_9177/ROW_SEL
+ pixel_9177/NB1 pixel_9177/VBIAS pixel_9177/NB2 pixel_9177/AMP_IN pixel_9177/SF_IB
+ pixel_9177/PIX_OUT pixel_9177/CSA_VREF pixel
Xpixel_9166 pixel_9166/gring pixel_9166/VDD pixel_9166/GND pixel_9166/VREF pixel_9166/ROW_SEL
+ pixel_9166/NB1 pixel_9166/VBIAS pixel_9166/NB2 pixel_9166/AMP_IN pixel_9166/SF_IB
+ pixel_9166/PIX_OUT pixel_9166/CSA_VREF pixel
Xpixel_8443 pixel_8443/gring pixel_8443/VDD pixel_8443/GND pixel_8443/VREF pixel_8443/ROW_SEL
+ pixel_8443/NB1 pixel_8443/VBIAS pixel_8443/NB2 pixel_8443/AMP_IN pixel_8443/SF_IB
+ pixel_8443/PIX_OUT pixel_8443/CSA_VREF pixel
Xpixel_9199 pixel_9199/gring pixel_9199/VDD pixel_9199/GND pixel_9199/VREF pixel_9199/ROW_SEL
+ pixel_9199/NB1 pixel_9199/VBIAS pixel_9199/NB2 pixel_9199/AMP_IN pixel_9199/SF_IB
+ pixel_9199/PIX_OUT pixel_9199/CSA_VREF pixel
Xpixel_8454 pixel_8454/gring pixel_8454/VDD pixel_8454/GND pixel_8454/VREF pixel_8454/ROW_SEL
+ pixel_8454/NB1 pixel_8454/VBIAS pixel_8454/NB2 pixel_8454/AMP_IN pixel_8454/SF_IB
+ pixel_8454/PIX_OUT pixel_8454/CSA_VREF pixel
Xpixel_8465 pixel_8465/gring pixel_8465/VDD pixel_8465/GND pixel_8465/VREF pixel_8465/ROW_SEL
+ pixel_8465/NB1 pixel_8465/VBIAS pixel_8465/NB2 pixel_8465/AMP_IN pixel_8465/SF_IB
+ pixel_8465/PIX_OUT pixel_8465/CSA_VREF pixel
Xpixel_8476 pixel_8476/gring pixel_8476/VDD pixel_8476/GND pixel_8476/VREF pixel_8476/ROW_SEL
+ pixel_8476/NB1 pixel_8476/VBIAS pixel_8476/NB2 pixel_8476/AMP_IN pixel_8476/SF_IB
+ pixel_8476/PIX_OUT pixel_8476/CSA_VREF pixel
Xpixel_8487 pixel_8487/gring pixel_8487/VDD pixel_8487/GND pixel_8487/VREF pixel_8487/ROW_SEL
+ pixel_8487/NB1 pixel_8487/VBIAS pixel_8487/NB2 pixel_8487/AMP_IN pixel_8487/SF_IB
+ pixel_8487/PIX_OUT pixel_8487/CSA_VREF pixel
Xpixel_7720 pixel_7720/gring pixel_7720/VDD pixel_7720/GND pixel_7720/VREF pixel_7720/ROW_SEL
+ pixel_7720/NB1 pixel_7720/VBIAS pixel_7720/NB2 pixel_7720/AMP_IN pixel_7720/SF_IB
+ pixel_7720/PIX_OUT pixel_7720/CSA_VREF pixel
Xpixel_7731 pixel_7731/gring pixel_7731/VDD pixel_7731/GND pixel_7731/VREF pixel_7731/ROW_SEL
+ pixel_7731/NB1 pixel_7731/VBIAS pixel_7731/NB2 pixel_7731/AMP_IN pixel_7731/SF_IB
+ pixel_7731/PIX_OUT pixel_7731/CSA_VREF pixel
Xpixel_7742 pixel_7742/gring pixel_7742/VDD pixel_7742/GND pixel_7742/VREF pixel_7742/ROW_SEL
+ pixel_7742/NB1 pixel_7742/VBIAS pixel_7742/NB2 pixel_7742/AMP_IN pixel_7742/SF_IB
+ pixel_7742/PIX_OUT pixel_7742/CSA_VREF pixel
Xpixel_8498 pixel_8498/gring pixel_8498/VDD pixel_8498/GND pixel_8498/VREF pixel_8498/ROW_SEL
+ pixel_8498/NB1 pixel_8498/VBIAS pixel_8498/NB2 pixel_8498/AMP_IN pixel_8498/SF_IB
+ pixel_8498/PIX_OUT pixel_8498/CSA_VREF pixel
Xpixel_7753 pixel_7753/gring pixel_7753/VDD pixel_7753/GND pixel_7753/VREF pixel_7753/ROW_SEL
+ pixel_7753/NB1 pixel_7753/VBIAS pixel_7753/NB2 pixel_7753/AMP_IN pixel_7753/SF_IB
+ pixel_7753/PIX_OUT pixel_7753/CSA_VREF pixel
Xpixel_7764 pixel_7764/gring pixel_7764/VDD pixel_7764/GND pixel_7764/VREF pixel_7764/ROW_SEL
+ pixel_7764/NB1 pixel_7764/VBIAS pixel_7764/NB2 pixel_7764/AMP_IN pixel_7764/SF_IB
+ pixel_7764/PIX_OUT pixel_7764/CSA_VREF pixel
Xpixel_7775 pixel_7775/gring pixel_7775/VDD pixel_7775/GND pixel_7775/VREF pixel_7775/ROW_SEL
+ pixel_7775/NB1 pixel_7775/VBIAS pixel_7775/NB2 pixel_7775/AMP_IN pixel_7775/SF_IB
+ pixel_7775/PIX_OUT pixel_7775/CSA_VREF pixel
Xpixel_7786 pixel_7786/gring pixel_7786/VDD pixel_7786/GND pixel_7786/VREF pixel_7786/ROW_SEL
+ pixel_7786/NB1 pixel_7786/VBIAS pixel_7786/NB2 pixel_7786/AMP_IN pixel_7786/SF_IB
+ pixel_7786/PIX_OUT pixel_7786/CSA_VREF pixel
Xpixel_7797 pixel_7797/gring pixel_7797/VDD pixel_7797/GND pixel_7797/VREF pixel_7797/ROW_SEL
+ pixel_7797/NB1 pixel_7797/VBIAS pixel_7797/NB2 pixel_7797/AMP_IN pixel_7797/SF_IB
+ pixel_7797/PIX_OUT pixel_7797/CSA_VREF pixel
Xpixel_2071 pixel_2071/gring pixel_2071/VDD pixel_2071/GND pixel_2071/VREF pixel_2071/ROW_SEL
+ pixel_2071/NB1 pixel_2071/VBIAS pixel_2071/NB2 pixel_2071/AMP_IN pixel_2071/SF_IB
+ pixel_2071/PIX_OUT pixel_2071/CSA_VREF pixel
Xpixel_2060 pixel_2060/gring pixel_2060/VDD pixel_2060/GND pixel_2060/VREF pixel_2060/ROW_SEL
+ pixel_2060/NB1 pixel_2060/VBIAS pixel_2060/NB2 pixel_2060/AMP_IN pixel_2060/SF_IB
+ pixel_2060/PIX_OUT pixel_2060/CSA_VREF pixel
Xpixel_1370 pixel_1370/gring pixel_1370/VDD pixel_1370/GND pixel_1370/VREF pixel_1370/ROW_SEL
+ pixel_1370/NB1 pixel_1370/VBIAS pixel_1370/NB2 pixel_1370/AMP_IN pixel_1370/SF_IB
+ pixel_1370/PIX_OUT pixel_1370/CSA_VREF pixel
Xpixel_2093 pixel_2093/gring pixel_2093/VDD pixel_2093/GND pixel_2093/VREF pixel_2093/ROW_SEL
+ pixel_2093/NB1 pixel_2093/VBIAS pixel_2093/NB2 pixel_2093/AMP_IN pixel_2093/SF_IB
+ pixel_2093/PIX_OUT pixel_2093/CSA_VREF pixel
Xpixel_2082 pixel_2082/gring pixel_2082/VDD pixel_2082/GND pixel_2082/VREF pixel_2082/ROW_SEL
+ pixel_2082/NB1 pixel_2082/VBIAS pixel_2082/NB2 pixel_2082/AMP_IN pixel_2082/SF_IB
+ pixel_2082/PIX_OUT pixel_2082/CSA_VREF pixel
Xpixel_1392 pixel_1392/gring pixel_1392/VDD pixel_1392/GND pixel_1392/VREF pixel_1392/ROW_SEL
+ pixel_1392/NB1 pixel_1392/VBIAS pixel_1392/NB2 pixel_1392/AMP_IN pixel_1392/SF_IB
+ pixel_1392/PIX_OUT pixel_1392/CSA_VREF pixel
Xpixel_1381 pixel_1381/gring pixel_1381/VDD pixel_1381/GND pixel_1381/VREF pixel_1381/ROW_SEL
+ pixel_1381/NB1 pixel_1381/VBIAS pixel_1381/NB2 pixel_1381/AMP_IN pixel_1381/SF_IB
+ pixel_1381/PIX_OUT pixel_1381/CSA_VREF pixel
Xpixel_429 pixel_429/gring pixel_429/VDD pixel_429/GND pixel_429/VREF pixel_429/ROW_SEL
+ pixel_429/NB1 pixel_429/VBIAS pixel_429/NB2 pixel_429/AMP_IN pixel_429/SF_IB pixel_429/PIX_OUT
+ pixel_429/CSA_VREF pixel
Xpixel_418 pixel_418/gring pixel_418/VDD pixel_418/GND pixel_418/VREF pixel_418/ROW_SEL
+ pixel_418/NB1 pixel_418/VBIAS pixel_418/NB2 pixel_418/AMP_IN pixel_418/SF_IB pixel_418/PIX_OUT
+ pixel_418/CSA_VREF pixel
Xpixel_407 pixel_407/gring pixel_407/VDD pixel_407/GND pixel_407/VREF pixel_407/ROW_SEL
+ pixel_407/NB1 pixel_407/VBIAS pixel_407/NB2 pixel_407/AMP_IN pixel_407/SF_IB pixel_407/PIX_OUT
+ pixel_407/CSA_VREF pixel
Xpixel_7005 pixel_7005/gring pixel_7005/VDD pixel_7005/GND pixel_7005/VREF pixel_7005/ROW_SEL
+ pixel_7005/NB1 pixel_7005/VBIAS pixel_7005/NB2 pixel_7005/AMP_IN pixel_7005/SF_IB
+ pixel_7005/PIX_OUT pixel_7005/CSA_VREF pixel
Xpixel_7016 pixel_7016/gring pixel_7016/VDD pixel_7016/GND pixel_7016/VREF pixel_7016/ROW_SEL
+ pixel_7016/NB1 pixel_7016/VBIAS pixel_7016/NB2 pixel_7016/AMP_IN pixel_7016/SF_IB
+ pixel_7016/PIX_OUT pixel_7016/CSA_VREF pixel
Xpixel_7027 pixel_7027/gring pixel_7027/VDD pixel_7027/GND pixel_7027/VREF pixel_7027/ROW_SEL
+ pixel_7027/NB1 pixel_7027/VBIAS pixel_7027/NB2 pixel_7027/AMP_IN pixel_7027/SF_IB
+ pixel_7027/PIX_OUT pixel_7027/CSA_VREF pixel
Xpixel_7038 pixel_7038/gring pixel_7038/VDD pixel_7038/GND pixel_7038/VREF pixel_7038/ROW_SEL
+ pixel_7038/NB1 pixel_7038/VBIAS pixel_7038/NB2 pixel_7038/AMP_IN pixel_7038/SF_IB
+ pixel_7038/PIX_OUT pixel_7038/CSA_VREF pixel
Xpixel_7049 pixel_7049/gring pixel_7049/VDD pixel_7049/GND pixel_7049/VREF pixel_7049/ROW_SEL
+ pixel_7049/NB1 pixel_7049/VBIAS pixel_7049/NB2 pixel_7049/AMP_IN pixel_7049/SF_IB
+ pixel_7049/PIX_OUT pixel_7049/CSA_VREF pixel
Xpixel_6304 pixel_6304/gring pixel_6304/VDD pixel_6304/GND pixel_6304/VREF pixel_6304/ROW_SEL
+ pixel_6304/NB1 pixel_6304/VBIAS pixel_6304/NB2 pixel_6304/AMP_IN pixel_6304/SF_IB
+ pixel_6304/PIX_OUT pixel_6304/CSA_VREF pixel
Xpixel_6315 pixel_6315/gring pixel_6315/VDD pixel_6315/GND pixel_6315/VREF pixel_6315/ROW_SEL
+ pixel_6315/NB1 pixel_6315/VBIAS pixel_6315/NB2 pixel_6315/AMP_IN pixel_6315/SF_IB
+ pixel_6315/PIX_OUT pixel_6315/CSA_VREF pixel
Xpixel_6326 pixel_6326/gring pixel_6326/VDD pixel_6326/GND pixel_6326/VREF pixel_6326/ROW_SEL
+ pixel_6326/NB1 pixel_6326/VBIAS pixel_6326/NB2 pixel_6326/AMP_IN pixel_6326/SF_IB
+ pixel_6326/PIX_OUT pixel_6326/CSA_VREF pixel
Xpixel_6337 pixel_6337/gring pixel_6337/VDD pixel_6337/GND pixel_6337/VREF pixel_6337/ROW_SEL
+ pixel_6337/NB1 pixel_6337/VBIAS pixel_6337/NB2 pixel_6337/AMP_IN pixel_6337/SF_IB
+ pixel_6337/PIX_OUT pixel_6337/CSA_VREF pixel
Xpixel_6348 pixel_6348/gring pixel_6348/VDD pixel_6348/GND pixel_6348/VREF pixel_6348/ROW_SEL
+ pixel_6348/NB1 pixel_6348/VBIAS pixel_6348/NB2 pixel_6348/AMP_IN pixel_6348/SF_IB
+ pixel_6348/PIX_OUT pixel_6348/CSA_VREF pixel
Xpixel_6359 pixel_6359/gring pixel_6359/VDD pixel_6359/GND pixel_6359/VREF pixel_6359/ROW_SEL
+ pixel_6359/NB1 pixel_6359/VBIAS pixel_6359/NB2 pixel_6359/AMP_IN pixel_6359/SF_IB
+ pixel_6359/PIX_OUT pixel_6359/CSA_VREF pixel
Xpixel_5603 pixel_5603/gring pixel_5603/VDD pixel_5603/GND pixel_5603/VREF pixel_5603/ROW_SEL
+ pixel_5603/NB1 pixel_5603/VBIAS pixel_5603/NB2 pixel_5603/AMP_IN pixel_5603/SF_IB
+ pixel_5603/PIX_OUT pixel_5603/CSA_VREF pixel
Xpixel_5614 pixel_5614/gring pixel_5614/VDD pixel_5614/GND pixel_5614/VREF pixel_5614/ROW_SEL
+ pixel_5614/NB1 pixel_5614/VBIAS pixel_5614/NB2 pixel_5614/AMP_IN pixel_5614/SF_IB
+ pixel_5614/PIX_OUT pixel_5614/CSA_VREF pixel
Xpixel_5625 pixel_5625/gring pixel_5625/VDD pixel_5625/GND pixel_5625/VREF pixel_5625/ROW_SEL
+ pixel_5625/NB1 pixel_5625/VBIAS pixel_5625/NB2 pixel_5625/AMP_IN pixel_5625/SF_IB
+ pixel_5625/PIX_OUT pixel_5625/CSA_VREF pixel
Xpixel_5636 pixel_5636/gring pixel_5636/VDD pixel_5636/GND pixel_5636/VREF pixel_5636/ROW_SEL
+ pixel_5636/NB1 pixel_5636/VBIAS pixel_5636/NB2 pixel_5636/AMP_IN pixel_5636/SF_IB
+ pixel_5636/PIX_OUT pixel_5636/CSA_VREF pixel
Xpixel_5647 pixel_5647/gring pixel_5647/VDD pixel_5647/GND pixel_5647/VREF pixel_5647/ROW_SEL
+ pixel_5647/NB1 pixel_5647/VBIAS pixel_5647/NB2 pixel_5647/AMP_IN pixel_5647/SF_IB
+ pixel_5647/PIX_OUT pixel_5647/CSA_VREF pixel
Xpixel_5658 pixel_5658/gring pixel_5658/VDD pixel_5658/GND pixel_5658/VREF pixel_5658/ROW_SEL
+ pixel_5658/NB1 pixel_5658/VBIAS pixel_5658/NB2 pixel_5658/AMP_IN pixel_5658/SF_IB
+ pixel_5658/PIX_OUT pixel_5658/CSA_VREF pixel
Xpixel_4902 pixel_4902/gring pixel_4902/VDD pixel_4902/GND pixel_4902/VREF pixel_4902/ROW_SEL
+ pixel_4902/NB1 pixel_4902/VBIAS pixel_4902/NB2 pixel_4902/AMP_IN pixel_4902/SF_IB
+ pixel_4902/PIX_OUT pixel_4902/CSA_VREF pixel
Xpixel_4913 pixel_4913/gring pixel_4913/VDD pixel_4913/GND pixel_4913/VREF pixel_4913/ROW_SEL
+ pixel_4913/NB1 pixel_4913/VBIAS pixel_4913/NB2 pixel_4913/AMP_IN pixel_4913/SF_IB
+ pixel_4913/PIX_OUT pixel_4913/CSA_VREF pixel
Xpixel_941 pixel_941/gring pixel_941/VDD pixel_941/GND pixel_941/VREF pixel_941/ROW_SEL
+ pixel_941/NB1 pixel_941/VBIAS pixel_941/NB2 pixel_941/AMP_IN pixel_941/SF_IB pixel_941/PIX_OUT
+ pixel_941/CSA_VREF pixel
Xpixel_930 pixel_930/gring pixel_930/VDD pixel_930/GND pixel_930/VREF pixel_930/ROW_SEL
+ pixel_930/NB1 pixel_930/VBIAS pixel_930/NB2 pixel_930/AMP_IN pixel_930/SF_IB pixel_930/PIX_OUT
+ pixel_930/CSA_VREF pixel
Xpixel_5669 pixel_5669/gring pixel_5669/VDD pixel_5669/GND pixel_5669/VREF pixel_5669/ROW_SEL
+ pixel_5669/NB1 pixel_5669/VBIAS pixel_5669/NB2 pixel_5669/AMP_IN pixel_5669/SF_IB
+ pixel_5669/PIX_OUT pixel_5669/CSA_VREF pixel
Xpixel_4924 pixel_4924/gring pixel_4924/VDD pixel_4924/GND pixel_4924/VREF pixel_4924/ROW_SEL
+ pixel_4924/NB1 pixel_4924/VBIAS pixel_4924/NB2 pixel_4924/AMP_IN pixel_4924/SF_IB
+ pixel_4924/PIX_OUT pixel_4924/CSA_VREF pixel
Xpixel_4935 pixel_4935/gring pixel_4935/VDD pixel_4935/GND pixel_4935/VREF pixel_4935/ROW_SEL
+ pixel_4935/NB1 pixel_4935/VBIAS pixel_4935/NB2 pixel_4935/AMP_IN pixel_4935/SF_IB
+ pixel_4935/PIX_OUT pixel_4935/CSA_VREF pixel
Xpixel_4946 pixel_4946/gring pixel_4946/VDD pixel_4946/GND pixel_4946/VREF pixel_4946/ROW_SEL
+ pixel_4946/NB1 pixel_4946/VBIAS pixel_4946/NB2 pixel_4946/AMP_IN pixel_4946/SF_IB
+ pixel_4946/PIX_OUT pixel_4946/CSA_VREF pixel
Xpixel_985 pixel_985/gring pixel_985/VDD pixel_985/GND pixel_985/VREF pixel_985/ROW_SEL
+ pixel_985/NB1 pixel_985/VBIAS pixel_985/NB2 pixel_985/AMP_IN pixel_985/SF_IB pixel_985/PIX_OUT
+ pixel_985/CSA_VREF pixel
Xpixel_974 pixel_974/gring pixel_974/VDD pixel_974/GND pixel_974/VREF pixel_974/ROW_SEL
+ pixel_974/NB1 pixel_974/VBIAS pixel_974/NB2 pixel_974/AMP_IN pixel_974/SF_IB pixel_974/PIX_OUT
+ pixel_974/CSA_VREF pixel
Xpixel_963 pixel_963/gring pixel_963/VDD pixel_963/GND pixel_963/VREF pixel_963/ROW_SEL
+ pixel_963/NB1 pixel_963/VBIAS pixel_963/NB2 pixel_963/AMP_IN pixel_963/SF_IB pixel_963/PIX_OUT
+ pixel_963/CSA_VREF pixel
Xpixel_952 pixel_952/gring pixel_952/VDD pixel_952/GND pixel_952/VREF pixel_952/ROW_SEL
+ pixel_952/NB1 pixel_952/VBIAS pixel_952/NB2 pixel_952/AMP_IN pixel_952/SF_IB pixel_952/PIX_OUT
+ pixel_952/CSA_VREF pixel
Xpixel_4957 pixel_4957/gring pixel_4957/VDD pixel_4957/GND pixel_4957/VREF pixel_4957/ROW_SEL
+ pixel_4957/NB1 pixel_4957/VBIAS pixel_4957/NB2 pixel_4957/AMP_IN pixel_4957/SF_IB
+ pixel_4957/PIX_OUT pixel_4957/CSA_VREF pixel
Xpixel_4968 pixel_4968/gring pixel_4968/VDD pixel_4968/GND pixel_4968/VREF pixel_4968/ROW_SEL
+ pixel_4968/NB1 pixel_4968/VBIAS pixel_4968/NB2 pixel_4968/AMP_IN pixel_4968/SF_IB
+ pixel_4968/PIX_OUT pixel_4968/CSA_VREF pixel
Xpixel_4979 pixel_4979/gring pixel_4979/VDD pixel_4979/GND pixel_4979/VREF pixel_4979/ROW_SEL
+ pixel_4979/NB1 pixel_4979/VBIAS pixel_4979/NB2 pixel_4979/AMP_IN pixel_4979/SF_IB
+ pixel_4979/PIX_OUT pixel_4979/CSA_VREF pixel
Xpixel_996 pixel_996/gring pixel_996/VDD pixel_996/GND pixel_996/VREF pixel_996/ROW_SEL
+ pixel_996/NB1 pixel_996/VBIAS pixel_996/NB2 pixel_996/AMP_IN pixel_996/SF_IB pixel_996/PIX_OUT
+ pixel_996/CSA_VREF pixel
Xpixel_8240 pixel_8240/gring pixel_8240/VDD pixel_8240/GND pixel_8240/VREF pixel_8240/ROW_SEL
+ pixel_8240/NB1 pixel_8240/VBIAS pixel_8240/NB2 pixel_8240/AMP_IN pixel_8240/SF_IB
+ pixel_8240/PIX_OUT pixel_8240/CSA_VREF pixel
Xpixel_8251 pixel_8251/gring pixel_8251/VDD pixel_8251/GND pixel_8251/VREF pixel_8251/ROW_SEL
+ pixel_8251/NB1 pixel_8251/VBIAS pixel_8251/NB2 pixel_8251/AMP_IN pixel_8251/SF_IB
+ pixel_8251/PIX_OUT pixel_8251/CSA_VREF pixel
Xpixel_8262 pixel_8262/gring pixel_8262/VDD pixel_8262/GND pixel_8262/VREF pixel_8262/ROW_SEL
+ pixel_8262/NB1 pixel_8262/VBIAS pixel_8262/NB2 pixel_8262/AMP_IN pixel_8262/SF_IB
+ pixel_8262/PIX_OUT pixel_8262/CSA_VREF pixel
Xpixel_8273 pixel_8273/gring pixel_8273/VDD pixel_8273/GND pixel_8273/VREF pixel_8273/ROW_SEL
+ pixel_8273/NB1 pixel_8273/VBIAS pixel_8273/NB2 pixel_8273/AMP_IN pixel_8273/SF_IB
+ pixel_8273/PIX_OUT pixel_8273/CSA_VREF pixel
Xpixel_8284 pixel_8284/gring pixel_8284/VDD pixel_8284/GND pixel_8284/VREF pixel_8284/ROW_SEL
+ pixel_8284/NB1 pixel_8284/VBIAS pixel_8284/NB2 pixel_8284/AMP_IN pixel_8284/SF_IB
+ pixel_8284/PIX_OUT pixel_8284/CSA_VREF pixel
Xpixel_8295 pixel_8295/gring pixel_8295/VDD pixel_8295/GND pixel_8295/VREF pixel_8295/ROW_SEL
+ pixel_8295/NB1 pixel_8295/VBIAS pixel_8295/NB2 pixel_8295/AMP_IN pixel_8295/SF_IB
+ pixel_8295/PIX_OUT pixel_8295/CSA_VREF pixel
Xpixel_7550 pixel_7550/gring pixel_7550/VDD pixel_7550/GND pixel_7550/VREF pixel_7550/ROW_SEL
+ pixel_7550/NB1 pixel_7550/VBIAS pixel_7550/NB2 pixel_7550/AMP_IN pixel_7550/SF_IB
+ pixel_7550/PIX_OUT pixel_7550/CSA_VREF pixel
Xpixel_7561 pixel_7561/gring pixel_7561/VDD pixel_7561/GND pixel_7561/VREF pixel_7561/ROW_SEL
+ pixel_7561/NB1 pixel_7561/VBIAS pixel_7561/NB2 pixel_7561/AMP_IN pixel_7561/SF_IB
+ pixel_7561/PIX_OUT pixel_7561/CSA_VREF pixel
Xpixel_7572 pixel_7572/gring pixel_7572/VDD pixel_7572/GND pixel_7572/VREF pixel_7572/ROW_SEL
+ pixel_7572/NB1 pixel_7572/VBIAS pixel_7572/NB2 pixel_7572/AMP_IN pixel_7572/SF_IB
+ pixel_7572/PIX_OUT pixel_7572/CSA_VREF pixel
Xpixel_7583 pixel_7583/gring pixel_7583/VDD pixel_7583/GND pixel_7583/VREF pixel_7583/ROW_SEL
+ pixel_7583/NB1 pixel_7583/VBIAS pixel_7583/NB2 pixel_7583/AMP_IN pixel_7583/SF_IB
+ pixel_7583/PIX_OUT pixel_7583/CSA_VREF pixel
Xpixel_7594 pixel_7594/gring pixel_7594/VDD pixel_7594/GND pixel_7594/VREF pixel_7594/ROW_SEL
+ pixel_7594/NB1 pixel_7594/VBIAS pixel_7594/NB2 pixel_7594/AMP_IN pixel_7594/SF_IB
+ pixel_7594/PIX_OUT pixel_7594/CSA_VREF pixel
Xpixel_6860 pixel_6860/gring pixel_6860/VDD pixel_6860/GND pixel_6860/VREF pixel_6860/ROW_SEL
+ pixel_6860/NB1 pixel_6860/VBIAS pixel_6860/NB2 pixel_6860/AMP_IN pixel_6860/SF_IB
+ pixel_6860/PIX_OUT pixel_6860/CSA_VREF pixel
Xpixel_6871 pixel_6871/gring pixel_6871/VDD pixel_6871/GND pixel_6871/VREF pixel_6871/ROW_SEL
+ pixel_6871/NB1 pixel_6871/VBIAS pixel_6871/NB2 pixel_6871/AMP_IN pixel_6871/SF_IB
+ pixel_6871/PIX_OUT pixel_6871/CSA_VREF pixel
Xpixel_6882 pixel_6882/gring pixel_6882/VDD pixel_6882/GND pixel_6882/VREF pixel_6882/ROW_SEL
+ pixel_6882/NB1 pixel_6882/VBIAS pixel_6882/NB2 pixel_6882/AMP_IN pixel_6882/SF_IB
+ pixel_6882/PIX_OUT pixel_6882/CSA_VREF pixel
Xpixel_6893 pixel_6893/gring pixel_6893/VDD pixel_6893/GND pixel_6893/VREF pixel_6893/ROW_SEL
+ pixel_6893/NB1 pixel_6893/VBIAS pixel_6893/NB2 pixel_6893/AMP_IN pixel_6893/SF_IB
+ pixel_6893/PIX_OUT pixel_6893/CSA_VREF pixel
Xpixel_204 pixel_204/gring pixel_204/VDD pixel_204/GND pixel_204/VREF pixel_204/ROW_SEL
+ pixel_204/NB1 pixel_204/VBIAS pixel_204/NB2 pixel_204/AMP_IN pixel_204/SF_IB pixel_204/PIX_OUT
+ pixel_204/CSA_VREF pixel
Xpixel_4209 pixel_4209/gring pixel_4209/VDD pixel_4209/GND pixel_4209/VREF pixel_4209/ROW_SEL
+ pixel_4209/NB1 pixel_4209/VBIAS pixel_4209/NB2 pixel_4209/AMP_IN pixel_4209/SF_IB
+ pixel_4209/PIX_OUT pixel_4209/CSA_VREF pixel
Xpixel_237 pixel_237/gring pixel_237/VDD pixel_237/GND pixel_237/VREF pixel_237/ROW_SEL
+ pixel_237/NB1 pixel_237/VBIAS pixel_237/NB2 pixel_237/AMP_IN pixel_237/SF_IB pixel_237/PIX_OUT
+ pixel_237/CSA_VREF pixel
Xpixel_226 pixel_226/gring pixel_226/VDD pixel_226/GND pixel_226/VREF pixel_226/ROW_SEL
+ pixel_226/NB1 pixel_226/VBIAS pixel_226/NB2 pixel_226/AMP_IN pixel_226/SF_IB pixel_226/PIX_OUT
+ pixel_226/CSA_VREF pixel
Xpixel_215 pixel_215/gring pixel_215/VDD pixel_215/GND pixel_215/VREF pixel_215/ROW_SEL
+ pixel_215/NB1 pixel_215/VBIAS pixel_215/NB2 pixel_215/AMP_IN pixel_215/SF_IB pixel_215/PIX_OUT
+ pixel_215/CSA_VREF pixel
Xpixel_259 pixel_259/gring pixel_259/VDD pixel_259/GND pixel_259/VREF pixel_259/ROW_SEL
+ pixel_259/NB1 pixel_259/VBIAS pixel_259/NB2 pixel_259/AMP_IN pixel_259/SF_IB pixel_259/PIX_OUT
+ pixel_259/CSA_VREF pixel
Xpixel_248 pixel_248/gring pixel_248/VDD pixel_248/GND pixel_248/VREF pixel_248/ROW_SEL
+ pixel_248/NB1 pixel_248/VBIAS pixel_248/NB2 pixel_248/AMP_IN pixel_248/SF_IB pixel_248/PIX_OUT
+ pixel_248/CSA_VREF pixel
Xpixel_3519 pixel_3519/gring pixel_3519/VDD pixel_3519/GND pixel_3519/VREF pixel_3519/ROW_SEL
+ pixel_3519/NB1 pixel_3519/VBIAS pixel_3519/NB2 pixel_3519/AMP_IN pixel_3519/SF_IB
+ pixel_3519/PIX_OUT pixel_3519/CSA_VREF pixel
Xpixel_3508 pixel_3508/gring pixel_3508/VDD pixel_3508/GND pixel_3508/VREF pixel_3508/ROW_SEL
+ pixel_3508/NB1 pixel_3508/VBIAS pixel_3508/NB2 pixel_3508/AMP_IN pixel_3508/SF_IB
+ pixel_3508/PIX_OUT pixel_3508/CSA_VREF pixel
Xpixel_2829 pixel_2829/gring pixel_2829/VDD pixel_2829/GND pixel_2829/VREF pixel_2829/ROW_SEL
+ pixel_2829/NB1 pixel_2829/VBIAS pixel_2829/NB2 pixel_2829/AMP_IN pixel_2829/SF_IB
+ pixel_2829/PIX_OUT pixel_2829/CSA_VREF pixel
Xpixel_2818 pixel_2818/gring pixel_2818/VDD pixel_2818/GND pixel_2818/VREF pixel_2818/ROW_SEL
+ pixel_2818/NB1 pixel_2818/VBIAS pixel_2818/NB2 pixel_2818/AMP_IN pixel_2818/SF_IB
+ pixel_2818/PIX_OUT pixel_2818/CSA_VREF pixel
Xpixel_2807 pixel_2807/gring pixel_2807/VDD pixel_2807/GND pixel_2807/VREF pixel_2807/ROW_SEL
+ pixel_2807/NB1 pixel_2807/VBIAS pixel_2807/NB2 pixel_2807/AMP_IN pixel_2807/SF_IB
+ pixel_2807/PIX_OUT pixel_2807/CSA_VREF pixel
Xpixel_6101 pixel_6101/gring pixel_6101/VDD pixel_6101/GND pixel_6101/VREF pixel_6101/ROW_SEL
+ pixel_6101/NB1 pixel_6101/VBIAS pixel_6101/NB2 pixel_6101/AMP_IN pixel_6101/SF_IB
+ pixel_6101/PIX_OUT pixel_6101/CSA_VREF pixel
Xpixel_6112 pixel_6112/gring pixel_6112/VDD pixel_6112/GND pixel_6112/VREF pixel_6112/ROW_SEL
+ pixel_6112/NB1 pixel_6112/VBIAS pixel_6112/NB2 pixel_6112/AMP_IN pixel_6112/SF_IB
+ pixel_6112/PIX_OUT pixel_6112/CSA_VREF pixel
Xpixel_6123 pixel_6123/gring pixel_6123/VDD pixel_6123/GND pixel_6123/VREF pixel_6123/ROW_SEL
+ pixel_6123/NB1 pixel_6123/VBIAS pixel_6123/NB2 pixel_6123/AMP_IN pixel_6123/SF_IB
+ pixel_6123/PIX_OUT pixel_6123/CSA_VREF pixel
Xpixel_6134 pixel_6134/gring pixel_6134/VDD pixel_6134/GND pixel_6134/VREF pixel_6134/ROW_SEL
+ pixel_6134/NB1 pixel_6134/VBIAS pixel_6134/NB2 pixel_6134/AMP_IN pixel_6134/SF_IB
+ pixel_6134/PIX_OUT pixel_6134/CSA_VREF pixel
Xpixel_6145 pixel_6145/gring pixel_6145/VDD pixel_6145/GND pixel_6145/VREF pixel_6145/ROW_SEL
+ pixel_6145/NB1 pixel_6145/VBIAS pixel_6145/NB2 pixel_6145/AMP_IN pixel_6145/SF_IB
+ pixel_6145/PIX_OUT pixel_6145/CSA_VREF pixel
Xpixel_6156 pixel_6156/gring pixel_6156/VDD pixel_6156/GND pixel_6156/VREF pixel_6156/ROW_SEL
+ pixel_6156/NB1 pixel_6156/VBIAS pixel_6156/NB2 pixel_6156/AMP_IN pixel_6156/SF_IB
+ pixel_6156/PIX_OUT pixel_6156/CSA_VREF pixel
Xpixel_6167 pixel_6167/gring pixel_6167/VDD pixel_6167/GND pixel_6167/VREF pixel_6167/ROW_SEL
+ pixel_6167/NB1 pixel_6167/VBIAS pixel_6167/NB2 pixel_6167/AMP_IN pixel_6167/SF_IB
+ pixel_6167/PIX_OUT pixel_6167/CSA_VREF pixel
Xpixel_5400 pixel_5400/gring pixel_5400/VDD pixel_5400/GND pixel_5400/VREF pixel_5400/ROW_SEL
+ pixel_5400/NB1 pixel_5400/VBIAS pixel_5400/NB2 pixel_5400/AMP_IN pixel_5400/SF_IB
+ pixel_5400/PIX_OUT pixel_5400/CSA_VREF pixel
Xpixel_5411 pixel_5411/gring pixel_5411/VDD pixel_5411/GND pixel_5411/VREF pixel_5411/ROW_SEL
+ pixel_5411/NB1 pixel_5411/VBIAS pixel_5411/NB2 pixel_5411/AMP_IN pixel_5411/SF_IB
+ pixel_5411/PIX_OUT pixel_5411/CSA_VREF pixel
Xpixel_5422 pixel_5422/gring pixel_5422/VDD pixel_5422/GND pixel_5422/VREF pixel_5422/ROW_SEL
+ pixel_5422/NB1 pixel_5422/VBIAS pixel_5422/NB2 pixel_5422/AMP_IN pixel_5422/SF_IB
+ pixel_5422/PIX_OUT pixel_5422/CSA_VREF pixel
Xpixel_5433 pixel_5433/gring pixel_5433/VDD pixel_5433/GND pixel_5433/VREF pixel_5433/ROW_SEL
+ pixel_5433/NB1 pixel_5433/VBIAS pixel_5433/NB2 pixel_5433/AMP_IN pixel_5433/SF_IB
+ pixel_5433/PIX_OUT pixel_5433/CSA_VREF pixel
Xpixel_6178 pixel_6178/gring pixel_6178/VDD pixel_6178/GND pixel_6178/VREF pixel_6178/ROW_SEL
+ pixel_6178/NB1 pixel_6178/VBIAS pixel_6178/NB2 pixel_6178/AMP_IN pixel_6178/SF_IB
+ pixel_6178/PIX_OUT pixel_6178/CSA_VREF pixel
Xpixel_6189 pixel_6189/gring pixel_6189/VDD pixel_6189/GND pixel_6189/VREF pixel_6189/ROW_SEL
+ pixel_6189/NB1 pixel_6189/VBIAS pixel_6189/NB2 pixel_6189/AMP_IN pixel_6189/SF_IB
+ pixel_6189/PIX_OUT pixel_6189/CSA_VREF pixel
Xpixel_5444 pixel_5444/gring pixel_5444/VDD pixel_5444/GND pixel_5444/VREF pixel_5444/ROW_SEL
+ pixel_5444/NB1 pixel_5444/VBIAS pixel_5444/NB2 pixel_5444/AMP_IN pixel_5444/SF_IB
+ pixel_5444/PIX_OUT pixel_5444/CSA_VREF pixel
Xpixel_5455 pixel_5455/gring pixel_5455/VDD pixel_5455/GND pixel_5455/VREF pixel_5455/ROW_SEL
+ pixel_5455/NB1 pixel_5455/VBIAS pixel_5455/NB2 pixel_5455/AMP_IN pixel_5455/SF_IB
+ pixel_5455/PIX_OUT pixel_5455/CSA_VREF pixel
Xpixel_5466 pixel_5466/gring pixel_5466/VDD pixel_5466/GND pixel_5466/VREF pixel_5466/ROW_SEL
+ pixel_5466/NB1 pixel_5466/VBIAS pixel_5466/NB2 pixel_5466/AMP_IN pixel_5466/SF_IB
+ pixel_5466/PIX_OUT pixel_5466/CSA_VREF pixel
Xpixel_4710 pixel_4710/gring pixel_4710/VDD pixel_4710/GND pixel_4710/VREF pixel_4710/ROW_SEL
+ pixel_4710/NB1 pixel_4710/VBIAS pixel_4710/NB2 pixel_4710/AMP_IN pixel_4710/SF_IB
+ pixel_4710/PIX_OUT pixel_4710/CSA_VREF pixel
Xpixel_4721 pixel_4721/gring pixel_4721/VDD pixel_4721/GND pixel_4721/VREF pixel_4721/ROW_SEL
+ pixel_4721/NB1 pixel_4721/VBIAS pixel_4721/NB2 pixel_4721/AMP_IN pixel_4721/SF_IB
+ pixel_4721/PIX_OUT pixel_4721/CSA_VREF pixel
Xpixel_760 pixel_760/gring pixel_760/VDD pixel_760/GND pixel_760/VREF pixel_760/ROW_SEL
+ pixel_760/NB1 pixel_760/VBIAS pixel_760/NB2 pixel_760/AMP_IN pixel_760/SF_IB pixel_760/PIX_OUT
+ pixel_760/CSA_VREF pixel
Xpixel_5477 pixel_5477/gring pixel_5477/VDD pixel_5477/GND pixel_5477/VREF pixel_5477/ROW_SEL
+ pixel_5477/NB1 pixel_5477/VBIAS pixel_5477/NB2 pixel_5477/AMP_IN pixel_5477/SF_IB
+ pixel_5477/PIX_OUT pixel_5477/CSA_VREF pixel
Xpixel_5488 pixel_5488/gring pixel_5488/VDD pixel_5488/GND pixel_5488/VREF pixel_5488/ROW_SEL
+ pixel_5488/NB1 pixel_5488/VBIAS pixel_5488/NB2 pixel_5488/AMP_IN pixel_5488/SF_IB
+ pixel_5488/PIX_OUT pixel_5488/CSA_VREF pixel
Xpixel_5499 pixel_5499/gring pixel_5499/VDD pixel_5499/GND pixel_5499/VREF pixel_5499/ROW_SEL
+ pixel_5499/NB1 pixel_5499/VBIAS pixel_5499/NB2 pixel_5499/AMP_IN pixel_5499/SF_IB
+ pixel_5499/PIX_OUT pixel_5499/CSA_VREF pixel
Xpixel_4732 pixel_4732/gring pixel_4732/VDD pixel_4732/GND pixel_4732/VREF pixel_4732/ROW_SEL
+ pixel_4732/NB1 pixel_4732/VBIAS pixel_4732/NB2 pixel_4732/AMP_IN pixel_4732/SF_IB
+ pixel_4732/PIX_OUT pixel_4732/CSA_VREF pixel
Xpixel_4743 pixel_4743/gring pixel_4743/VDD pixel_4743/GND pixel_4743/VREF pixel_4743/ROW_SEL
+ pixel_4743/NB1 pixel_4743/VBIAS pixel_4743/NB2 pixel_4743/AMP_IN pixel_4743/SF_IB
+ pixel_4743/PIX_OUT pixel_4743/CSA_VREF pixel
Xpixel_4754 pixel_4754/gring pixel_4754/VDD pixel_4754/GND pixel_4754/VREF pixel_4754/ROW_SEL
+ pixel_4754/NB1 pixel_4754/VBIAS pixel_4754/NB2 pixel_4754/AMP_IN pixel_4754/SF_IB
+ pixel_4754/PIX_OUT pixel_4754/CSA_VREF pixel
Xpixel_793 pixel_793/gring pixel_793/VDD pixel_793/GND pixel_793/VREF pixel_793/ROW_SEL
+ pixel_793/NB1 pixel_793/VBIAS pixel_793/NB2 pixel_793/AMP_IN pixel_793/SF_IB pixel_793/PIX_OUT
+ pixel_793/CSA_VREF pixel
Xpixel_782 pixel_782/gring pixel_782/VDD pixel_782/GND pixel_782/VREF pixel_782/ROW_SEL
+ pixel_782/NB1 pixel_782/VBIAS pixel_782/NB2 pixel_782/AMP_IN pixel_782/SF_IB pixel_782/PIX_OUT
+ pixel_782/CSA_VREF pixel
Xpixel_771 pixel_771/gring pixel_771/VDD pixel_771/GND pixel_771/VREF pixel_771/ROW_SEL
+ pixel_771/NB1 pixel_771/VBIAS pixel_771/NB2 pixel_771/AMP_IN pixel_771/SF_IB pixel_771/PIX_OUT
+ pixel_771/CSA_VREF pixel
Xpixel_4765 pixel_4765/gring pixel_4765/VDD pixel_4765/GND pixel_4765/VREF pixel_4765/ROW_SEL
+ pixel_4765/NB1 pixel_4765/VBIAS pixel_4765/NB2 pixel_4765/AMP_IN pixel_4765/SF_IB
+ pixel_4765/PIX_OUT pixel_4765/CSA_VREF pixel
Xpixel_4776 pixel_4776/gring pixel_4776/VDD pixel_4776/GND pixel_4776/VREF pixel_4776/ROW_SEL
+ pixel_4776/NB1 pixel_4776/VBIAS pixel_4776/NB2 pixel_4776/AMP_IN pixel_4776/SF_IB
+ pixel_4776/PIX_OUT pixel_4776/CSA_VREF pixel
Xpixel_4787 pixel_4787/gring pixel_4787/VDD pixel_4787/GND pixel_4787/VREF pixel_4787/ROW_SEL
+ pixel_4787/NB1 pixel_4787/VBIAS pixel_4787/NB2 pixel_4787/AMP_IN pixel_4787/SF_IB
+ pixel_4787/PIX_OUT pixel_4787/CSA_VREF pixel
Xpixel_4798 pixel_4798/gring pixel_4798/VDD pixel_4798/GND pixel_4798/VREF pixel_4798/ROW_SEL
+ pixel_4798/NB1 pixel_4798/VBIAS pixel_4798/NB2 pixel_4798/AMP_IN pixel_4798/SF_IB
+ pixel_4798/PIX_OUT pixel_4798/CSA_VREF pixel
Xpixel_8070 pixel_8070/gring pixel_8070/VDD pixel_8070/GND pixel_8070/VREF pixel_8070/ROW_SEL
+ pixel_8070/NB1 pixel_8070/VBIAS pixel_8070/NB2 pixel_8070/AMP_IN pixel_8070/SF_IB
+ pixel_8070/PIX_OUT pixel_8070/CSA_VREF pixel
Xpixel_8081 pixel_8081/gring pixel_8081/VDD pixel_8081/GND pixel_8081/VREF pixel_8081/ROW_SEL
+ pixel_8081/NB1 pixel_8081/VBIAS pixel_8081/NB2 pixel_8081/AMP_IN pixel_8081/SF_IB
+ pixel_8081/PIX_OUT pixel_8081/CSA_VREF pixel
Xpixel_8092 pixel_8092/gring pixel_8092/VDD pixel_8092/GND pixel_8092/VREF pixel_8092/ROW_SEL
+ pixel_8092/NB1 pixel_8092/VBIAS pixel_8092/NB2 pixel_8092/AMP_IN pixel_8092/SF_IB
+ pixel_8092/PIX_OUT pixel_8092/CSA_VREF pixel
Xpixel_7380 pixel_7380/gring pixel_7380/VDD pixel_7380/GND pixel_7380/VREF pixel_7380/ROW_SEL
+ pixel_7380/NB1 pixel_7380/VBIAS pixel_7380/NB2 pixel_7380/AMP_IN pixel_7380/SF_IB
+ pixel_7380/PIX_OUT pixel_7380/CSA_VREF pixel
Xpixel_7391 pixel_7391/gring pixel_7391/VDD pixel_7391/GND pixel_7391/VREF pixel_7391/ROW_SEL
+ pixel_7391/NB1 pixel_7391/VBIAS pixel_7391/NB2 pixel_7391/AMP_IN pixel_7391/SF_IB
+ pixel_7391/PIX_OUT pixel_7391/CSA_VREF pixel
Xpixel_6690 pixel_6690/gring pixel_6690/VDD pixel_6690/GND pixel_6690/VREF pixel_6690/ROW_SEL
+ pixel_6690/NB1 pixel_6690/VBIAS pixel_6690/NB2 pixel_6690/AMP_IN pixel_6690/SF_IB
+ pixel_6690/PIX_OUT pixel_6690/CSA_VREF pixel
Xpixel_4006 pixel_4006/gring pixel_4006/VDD pixel_4006/GND pixel_4006/VREF pixel_4006/ROW_SEL
+ pixel_4006/NB1 pixel_4006/VBIAS pixel_4006/NB2 pixel_4006/AMP_IN pixel_4006/SF_IB
+ pixel_4006/PIX_OUT pixel_4006/CSA_VREF pixel
Xpixel_4017 pixel_4017/gring pixel_4017/VDD pixel_4017/GND pixel_4017/VREF pixel_4017/ROW_SEL
+ pixel_4017/NB1 pixel_4017/VBIAS pixel_4017/NB2 pixel_4017/AMP_IN pixel_4017/SF_IB
+ pixel_4017/PIX_OUT pixel_4017/CSA_VREF pixel
Xpixel_3305 pixel_3305/gring pixel_3305/VDD pixel_3305/GND pixel_3305/VREF pixel_3305/ROW_SEL
+ pixel_3305/NB1 pixel_3305/VBIAS pixel_3305/NB2 pixel_3305/AMP_IN pixel_3305/SF_IB
+ pixel_3305/PIX_OUT pixel_3305/CSA_VREF pixel
Xpixel_4028 pixel_4028/gring pixel_4028/VDD pixel_4028/GND pixel_4028/VREF pixel_4028/ROW_SEL
+ pixel_4028/NB1 pixel_4028/VBIAS pixel_4028/NB2 pixel_4028/AMP_IN pixel_4028/SF_IB
+ pixel_4028/PIX_OUT pixel_4028/CSA_VREF pixel
Xpixel_4039 pixel_4039/gring pixel_4039/VDD pixel_4039/GND pixel_4039/VREF pixel_4039/ROW_SEL
+ pixel_4039/NB1 pixel_4039/VBIAS pixel_4039/NB2 pixel_4039/AMP_IN pixel_4039/SF_IB
+ pixel_4039/PIX_OUT pixel_4039/CSA_VREF pixel
Xpixel_2604 pixel_2604/gring pixel_2604/VDD pixel_2604/GND pixel_2604/VREF pixel_2604/ROW_SEL
+ pixel_2604/NB1 pixel_2604/VBIAS pixel_2604/NB2 pixel_2604/AMP_IN pixel_2604/SF_IB
+ pixel_2604/PIX_OUT pixel_2604/CSA_VREF pixel
Xpixel_3349 pixel_3349/gring pixel_3349/VDD pixel_3349/GND pixel_3349/VREF pixel_3349/ROW_SEL
+ pixel_3349/NB1 pixel_3349/VBIAS pixel_3349/NB2 pixel_3349/AMP_IN pixel_3349/SF_IB
+ pixel_3349/PIX_OUT pixel_3349/CSA_VREF pixel
Xpixel_3338 pixel_3338/gring pixel_3338/VDD pixel_3338/GND pixel_3338/VREF pixel_3338/ROW_SEL
+ pixel_3338/NB1 pixel_3338/VBIAS pixel_3338/NB2 pixel_3338/AMP_IN pixel_3338/SF_IB
+ pixel_3338/PIX_OUT pixel_3338/CSA_VREF pixel
Xpixel_3327 pixel_3327/gring pixel_3327/VDD pixel_3327/GND pixel_3327/VREF pixel_3327/ROW_SEL
+ pixel_3327/NB1 pixel_3327/VBIAS pixel_3327/NB2 pixel_3327/AMP_IN pixel_3327/SF_IB
+ pixel_3327/PIX_OUT pixel_3327/CSA_VREF pixel
Xpixel_3316 pixel_3316/gring pixel_3316/VDD pixel_3316/GND pixel_3316/VREF pixel_3316/ROW_SEL
+ pixel_3316/NB1 pixel_3316/VBIAS pixel_3316/NB2 pixel_3316/AMP_IN pixel_3316/SF_IB
+ pixel_3316/PIX_OUT pixel_3316/CSA_VREF pixel
Xpixel_2637 pixel_2637/gring pixel_2637/VDD pixel_2637/GND pixel_2637/VREF pixel_2637/ROW_SEL
+ pixel_2637/NB1 pixel_2637/VBIAS pixel_2637/NB2 pixel_2637/AMP_IN pixel_2637/SF_IB
+ pixel_2637/PIX_OUT pixel_2637/CSA_VREF pixel
Xpixel_2626 pixel_2626/gring pixel_2626/VDD pixel_2626/GND pixel_2626/VREF pixel_2626/ROW_SEL
+ pixel_2626/NB1 pixel_2626/VBIAS pixel_2626/NB2 pixel_2626/AMP_IN pixel_2626/SF_IB
+ pixel_2626/PIX_OUT pixel_2626/CSA_VREF pixel
Xpixel_2615 pixel_2615/gring pixel_2615/VDD pixel_2615/GND pixel_2615/VREF pixel_2615/ROW_SEL
+ pixel_2615/NB1 pixel_2615/VBIAS pixel_2615/NB2 pixel_2615/AMP_IN pixel_2615/SF_IB
+ pixel_2615/PIX_OUT pixel_2615/CSA_VREF pixel
Xpixel_1925 pixel_1925/gring pixel_1925/VDD pixel_1925/GND pixel_1925/VREF pixel_1925/ROW_SEL
+ pixel_1925/NB1 pixel_1925/VBIAS pixel_1925/NB2 pixel_1925/AMP_IN pixel_1925/SF_IB
+ pixel_1925/PIX_OUT pixel_1925/CSA_VREF pixel
Xpixel_1914 pixel_1914/gring pixel_1914/VDD pixel_1914/GND pixel_1914/VREF pixel_1914/ROW_SEL
+ pixel_1914/NB1 pixel_1914/VBIAS pixel_1914/NB2 pixel_1914/AMP_IN pixel_1914/SF_IB
+ pixel_1914/PIX_OUT pixel_1914/CSA_VREF pixel
Xpixel_1903 pixel_1903/gring pixel_1903/VDD pixel_1903/GND pixel_1903/VREF pixel_1903/ROW_SEL
+ pixel_1903/NB1 pixel_1903/VBIAS pixel_1903/NB2 pixel_1903/AMP_IN pixel_1903/SF_IB
+ pixel_1903/PIX_OUT pixel_1903/CSA_VREF pixel
Xpixel_2659 pixel_2659/gring pixel_2659/VDD pixel_2659/GND pixel_2659/VREF pixel_2659/ROW_SEL
+ pixel_2659/NB1 pixel_2659/VBIAS pixel_2659/NB2 pixel_2659/AMP_IN pixel_2659/SF_IB
+ pixel_2659/PIX_OUT pixel_2659/CSA_VREF pixel
Xpixel_2648 pixel_2648/gring pixel_2648/VDD pixel_2648/GND pixel_2648/VREF pixel_2648/ROW_SEL
+ pixel_2648/NB1 pixel_2648/VBIAS pixel_2648/NB2 pixel_2648/AMP_IN pixel_2648/SF_IB
+ pixel_2648/PIX_OUT pixel_2648/CSA_VREF pixel
Xpixel_1969 pixel_1969/gring pixel_1969/VDD pixel_1969/GND pixel_1969/VREF pixel_1969/ROW_SEL
+ pixel_1969/NB1 pixel_1969/VBIAS pixel_1969/NB2 pixel_1969/AMP_IN pixel_1969/SF_IB
+ pixel_1969/PIX_OUT pixel_1969/CSA_VREF pixel
Xpixel_1958 pixel_1958/gring pixel_1958/VDD pixel_1958/GND pixel_1958/VREF pixel_1958/ROW_SEL
+ pixel_1958/NB1 pixel_1958/VBIAS pixel_1958/NB2 pixel_1958/AMP_IN pixel_1958/SF_IB
+ pixel_1958/PIX_OUT pixel_1958/CSA_VREF pixel
Xpixel_1947 pixel_1947/gring pixel_1947/VDD pixel_1947/GND pixel_1947/VREF pixel_1947/ROW_SEL
+ pixel_1947/NB1 pixel_1947/VBIAS pixel_1947/NB2 pixel_1947/AMP_IN pixel_1947/SF_IB
+ pixel_1947/PIX_OUT pixel_1947/CSA_VREF pixel
Xpixel_1936 pixel_1936/gring pixel_1936/VDD pixel_1936/GND pixel_1936/VREF pixel_1936/ROW_SEL
+ pixel_1936/NB1 pixel_1936/VBIAS pixel_1936/NB2 pixel_1936/AMP_IN pixel_1936/SF_IB
+ pixel_1936/PIX_OUT pixel_1936/CSA_VREF pixel
Xpixel_5230 pixel_5230/gring pixel_5230/VDD pixel_5230/GND pixel_5230/VREF pixel_5230/ROW_SEL
+ pixel_5230/NB1 pixel_5230/VBIAS pixel_5230/NB2 pixel_5230/AMP_IN pixel_5230/SF_IB
+ pixel_5230/PIX_OUT pixel_5230/CSA_VREF pixel
Xpixel_5241 pixel_5241/gring pixel_5241/VDD pixel_5241/GND pixel_5241/VREF pixel_5241/ROW_SEL
+ pixel_5241/NB1 pixel_5241/VBIAS pixel_5241/NB2 pixel_5241/AMP_IN pixel_5241/SF_IB
+ pixel_5241/PIX_OUT pixel_5241/CSA_VREF pixel
Xpixel_5252 pixel_5252/gring pixel_5252/VDD pixel_5252/GND pixel_5252/VREF pixel_5252/ROW_SEL
+ pixel_5252/NB1 pixel_5252/VBIAS pixel_5252/NB2 pixel_5252/AMP_IN pixel_5252/SF_IB
+ pixel_5252/PIX_OUT pixel_5252/CSA_VREF pixel
Xpixel_5263 pixel_5263/gring pixel_5263/VDD pixel_5263/GND pixel_5263/VREF pixel_5263/ROW_SEL
+ pixel_5263/NB1 pixel_5263/VBIAS pixel_5263/NB2 pixel_5263/AMP_IN pixel_5263/SF_IB
+ pixel_5263/PIX_OUT pixel_5263/CSA_VREF pixel
Xpixel_5274 pixel_5274/gring pixel_5274/VDD pixel_5274/GND pixel_5274/VREF pixel_5274/ROW_SEL
+ pixel_5274/NB1 pixel_5274/VBIAS pixel_5274/NB2 pixel_5274/AMP_IN pixel_5274/SF_IB
+ pixel_5274/PIX_OUT pixel_5274/CSA_VREF pixel
Xpixel_5285 pixel_5285/gring pixel_5285/VDD pixel_5285/GND pixel_5285/VREF pixel_5285/ROW_SEL
+ pixel_5285/NB1 pixel_5285/VBIAS pixel_5285/NB2 pixel_5285/AMP_IN pixel_5285/SF_IB
+ pixel_5285/PIX_OUT pixel_5285/CSA_VREF pixel
Xpixel_5296 pixel_5296/gring pixel_5296/VDD pixel_5296/GND pixel_5296/VREF pixel_5296/ROW_SEL
+ pixel_5296/NB1 pixel_5296/VBIAS pixel_5296/NB2 pixel_5296/AMP_IN pixel_5296/SF_IB
+ pixel_5296/PIX_OUT pixel_5296/CSA_VREF pixel
Xpixel_4540 pixel_4540/gring pixel_4540/VDD pixel_4540/GND pixel_4540/VREF pixel_4540/ROW_SEL
+ pixel_4540/NB1 pixel_4540/VBIAS pixel_4540/NB2 pixel_4540/AMP_IN pixel_4540/SF_IB
+ pixel_4540/PIX_OUT pixel_4540/CSA_VREF pixel
Xpixel_4551 pixel_4551/gring pixel_4551/VDD pixel_4551/GND pixel_4551/VREF pixel_4551/ROW_SEL
+ pixel_4551/NB1 pixel_4551/VBIAS pixel_4551/NB2 pixel_4551/AMP_IN pixel_4551/SF_IB
+ pixel_4551/PIX_OUT pixel_4551/CSA_VREF pixel
Xpixel_4562 pixel_4562/gring pixel_4562/VDD pixel_4562/GND pixel_4562/VREF pixel_4562/ROW_SEL
+ pixel_4562/NB1 pixel_4562/VBIAS pixel_4562/NB2 pixel_4562/AMP_IN pixel_4562/SF_IB
+ pixel_4562/PIX_OUT pixel_4562/CSA_VREF pixel
Xpixel_4573 pixel_4573/gring pixel_4573/VDD pixel_4573/GND pixel_4573/VREF pixel_4573/ROW_SEL
+ pixel_4573/NB1 pixel_4573/VBIAS pixel_4573/NB2 pixel_4573/AMP_IN pixel_4573/SF_IB
+ pixel_4573/PIX_OUT pixel_4573/CSA_VREF pixel
Xpixel_590 pixel_590/gring pixel_590/VDD pixel_590/GND pixel_590/VREF pixel_590/ROW_SEL
+ pixel_590/NB1 pixel_590/VBIAS pixel_590/NB2 pixel_590/AMP_IN pixel_590/SF_IB pixel_590/PIX_OUT
+ pixel_590/CSA_VREF pixel
Xpixel_3861 pixel_3861/gring pixel_3861/VDD pixel_3861/GND pixel_3861/VREF pixel_3861/ROW_SEL
+ pixel_3861/NB1 pixel_3861/VBIAS pixel_3861/NB2 pixel_3861/AMP_IN pixel_3861/SF_IB
+ pixel_3861/PIX_OUT pixel_3861/CSA_VREF pixel
Xpixel_3850 pixel_3850/gring pixel_3850/VDD pixel_3850/GND pixel_3850/VREF pixel_3850/ROW_SEL
+ pixel_3850/NB1 pixel_3850/VBIAS pixel_3850/NB2 pixel_3850/AMP_IN pixel_3850/SF_IB
+ pixel_3850/PIX_OUT pixel_3850/CSA_VREF pixel
Xpixel_4584 pixel_4584/gring pixel_4584/VDD pixel_4584/GND pixel_4584/VREF pixel_4584/ROW_SEL
+ pixel_4584/NB1 pixel_4584/VBIAS pixel_4584/NB2 pixel_4584/AMP_IN pixel_4584/SF_IB
+ pixel_4584/PIX_OUT pixel_4584/CSA_VREF pixel
Xpixel_4595 pixel_4595/gring pixel_4595/VDD pixel_4595/GND pixel_4595/VREF pixel_4595/ROW_SEL
+ pixel_4595/NB1 pixel_4595/VBIAS pixel_4595/NB2 pixel_4595/AMP_IN pixel_4595/SF_IB
+ pixel_4595/PIX_OUT pixel_4595/CSA_VREF pixel
Xpixel_3894 pixel_3894/gring pixel_3894/VDD pixel_3894/GND pixel_3894/VREF pixel_3894/ROW_SEL
+ pixel_3894/NB1 pixel_3894/VBIAS pixel_3894/NB2 pixel_3894/AMP_IN pixel_3894/SF_IB
+ pixel_3894/PIX_OUT pixel_3894/CSA_VREF pixel
Xpixel_3883 pixel_3883/gring pixel_3883/VDD pixel_3883/GND pixel_3883/VREF pixel_3883/ROW_SEL
+ pixel_3883/NB1 pixel_3883/VBIAS pixel_3883/NB2 pixel_3883/AMP_IN pixel_3883/SF_IB
+ pixel_3883/PIX_OUT pixel_3883/CSA_VREF pixel
Xpixel_3872 pixel_3872/gring pixel_3872/VDD pixel_3872/GND pixel_3872/VREF pixel_3872/ROW_SEL
+ pixel_3872/NB1 pixel_3872/VBIAS pixel_3872/NB2 pixel_3872/AMP_IN pixel_3872/SF_IB
+ pixel_3872/PIX_OUT pixel_3872/CSA_VREF pixel
Xpixel_9529 pixel_9529/gring pixel_9529/VDD pixel_9529/GND pixel_9529/VREF pixel_9529/ROW_SEL
+ pixel_9529/NB1 pixel_9529/VBIAS pixel_9529/NB2 pixel_9529/AMP_IN pixel_9529/SF_IB
+ pixel_9529/PIX_OUT pixel_9529/CSA_VREF pixel
Xpixel_9518 pixel_9518/gring pixel_9518/VDD pixel_9518/GND pixel_9518/VREF pixel_9518/ROW_SEL
+ pixel_9518/NB1 pixel_9518/VBIAS pixel_9518/NB2 pixel_9518/AMP_IN pixel_9518/SF_IB
+ pixel_9518/PIX_OUT pixel_9518/CSA_VREF pixel
Xpixel_9507 pixel_9507/gring pixel_9507/VDD pixel_9507/GND pixel_9507/VREF pixel_9507/ROW_SEL
+ pixel_9507/NB1 pixel_9507/VBIAS pixel_9507/NB2 pixel_9507/AMP_IN pixel_9507/SF_IB
+ pixel_9507/PIX_OUT pixel_9507/CSA_VREF pixel
Xpixel_8828 pixel_8828/gring pixel_8828/VDD pixel_8828/GND pixel_8828/VREF pixel_8828/ROW_SEL
+ pixel_8828/NB1 pixel_8828/VBIAS pixel_8828/NB2 pixel_8828/AMP_IN pixel_8828/SF_IB
+ pixel_8828/PIX_OUT pixel_8828/CSA_VREF pixel
Xpixel_8817 pixel_8817/gring pixel_8817/VDD pixel_8817/GND pixel_8817/VREF pixel_8817/ROW_SEL
+ pixel_8817/NB1 pixel_8817/VBIAS pixel_8817/NB2 pixel_8817/AMP_IN pixel_8817/SF_IB
+ pixel_8817/PIX_OUT pixel_8817/CSA_VREF pixel
Xpixel_8806 pixel_8806/gring pixel_8806/VDD pixel_8806/GND pixel_8806/VREF pixel_8806/ROW_SEL
+ pixel_8806/NB1 pixel_8806/VBIAS pixel_8806/NB2 pixel_8806/AMP_IN pixel_8806/SF_IB
+ pixel_8806/PIX_OUT pixel_8806/CSA_VREF pixel
Xpixel_8839 pixel_8839/gring pixel_8839/VDD pixel_8839/GND pixel_8839/VREF pixel_8839/ROW_SEL
+ pixel_8839/NB1 pixel_8839/VBIAS pixel_8839/NB2 pixel_8839/AMP_IN pixel_8839/SF_IB
+ pixel_8839/PIX_OUT pixel_8839/CSA_VREF pixel
Xpixel_3113 pixel_3113/gring pixel_3113/VDD pixel_3113/GND pixel_3113/VREF pixel_3113/ROW_SEL
+ pixel_3113/NB1 pixel_3113/VBIAS pixel_3113/NB2 pixel_3113/AMP_IN pixel_3113/SF_IB
+ pixel_3113/PIX_OUT pixel_3113/CSA_VREF pixel
Xpixel_3102 pixel_3102/gring pixel_3102/VDD pixel_3102/GND pixel_3102/VREF pixel_3102/ROW_SEL
+ pixel_3102/NB1 pixel_3102/VBIAS pixel_3102/NB2 pixel_3102/AMP_IN pixel_3102/SF_IB
+ pixel_3102/PIX_OUT pixel_3102/CSA_VREF pixel
Xpixel_2412 pixel_2412/gring pixel_2412/VDD pixel_2412/GND pixel_2412/VREF pixel_2412/ROW_SEL
+ pixel_2412/NB1 pixel_2412/VBIAS pixel_2412/NB2 pixel_2412/AMP_IN pixel_2412/SF_IB
+ pixel_2412/PIX_OUT pixel_2412/CSA_VREF pixel
Xpixel_2401 pixel_2401/gring pixel_2401/VDD pixel_2401/GND pixel_2401/VREF pixel_2401/ROW_SEL
+ pixel_2401/NB1 pixel_2401/VBIAS pixel_2401/NB2 pixel_2401/AMP_IN pixel_2401/SF_IB
+ pixel_2401/PIX_OUT pixel_2401/CSA_VREF pixel
Xpixel_3157 pixel_3157/gring pixel_3157/VDD pixel_3157/GND pixel_3157/VREF pixel_3157/ROW_SEL
+ pixel_3157/NB1 pixel_3157/VBIAS pixel_3157/NB2 pixel_3157/AMP_IN pixel_3157/SF_IB
+ pixel_3157/PIX_OUT pixel_3157/CSA_VREF pixel
Xpixel_3146 pixel_3146/gring pixel_3146/VDD pixel_3146/GND pixel_3146/VREF pixel_3146/ROW_SEL
+ pixel_3146/NB1 pixel_3146/VBIAS pixel_3146/NB2 pixel_3146/AMP_IN pixel_3146/SF_IB
+ pixel_3146/PIX_OUT pixel_3146/CSA_VREF pixel
Xpixel_3135 pixel_3135/gring pixel_3135/VDD pixel_3135/GND pixel_3135/VREF pixel_3135/ROW_SEL
+ pixel_3135/NB1 pixel_3135/VBIAS pixel_3135/NB2 pixel_3135/AMP_IN pixel_3135/SF_IB
+ pixel_3135/PIX_OUT pixel_3135/CSA_VREF pixel
Xpixel_3124 pixel_3124/gring pixel_3124/VDD pixel_3124/GND pixel_3124/VREF pixel_3124/ROW_SEL
+ pixel_3124/NB1 pixel_3124/VBIAS pixel_3124/NB2 pixel_3124/AMP_IN pixel_3124/SF_IB
+ pixel_3124/PIX_OUT pixel_3124/CSA_VREF pixel
Xpixel_1700 pixel_1700/gring pixel_1700/VDD pixel_1700/GND pixel_1700/VREF pixel_1700/ROW_SEL
+ pixel_1700/NB1 pixel_1700/VBIAS pixel_1700/NB2 pixel_1700/AMP_IN pixel_1700/SF_IB
+ pixel_1700/PIX_OUT pixel_1700/CSA_VREF pixel
Xpixel_2445 pixel_2445/gring pixel_2445/VDD pixel_2445/GND pixel_2445/VREF pixel_2445/ROW_SEL
+ pixel_2445/NB1 pixel_2445/VBIAS pixel_2445/NB2 pixel_2445/AMP_IN pixel_2445/SF_IB
+ pixel_2445/PIX_OUT pixel_2445/CSA_VREF pixel
Xpixel_2434 pixel_2434/gring pixel_2434/VDD pixel_2434/GND pixel_2434/VREF pixel_2434/ROW_SEL
+ pixel_2434/NB1 pixel_2434/VBIAS pixel_2434/NB2 pixel_2434/AMP_IN pixel_2434/SF_IB
+ pixel_2434/PIX_OUT pixel_2434/CSA_VREF pixel
Xpixel_2423 pixel_2423/gring pixel_2423/VDD pixel_2423/GND pixel_2423/VREF pixel_2423/ROW_SEL
+ pixel_2423/NB1 pixel_2423/VBIAS pixel_2423/NB2 pixel_2423/AMP_IN pixel_2423/SF_IB
+ pixel_2423/PIX_OUT pixel_2423/CSA_VREF pixel
Xpixel_3179 pixel_3179/gring pixel_3179/VDD pixel_3179/GND pixel_3179/VREF pixel_3179/ROW_SEL
+ pixel_3179/NB1 pixel_3179/VBIAS pixel_3179/NB2 pixel_3179/AMP_IN pixel_3179/SF_IB
+ pixel_3179/PIX_OUT pixel_3179/CSA_VREF pixel
Xpixel_3168 pixel_3168/gring pixel_3168/VDD pixel_3168/GND pixel_3168/VREF pixel_3168/ROW_SEL
+ pixel_3168/NB1 pixel_3168/VBIAS pixel_3168/NB2 pixel_3168/AMP_IN pixel_3168/SF_IB
+ pixel_3168/PIX_OUT pixel_3168/CSA_VREF pixel
Xpixel_1744 pixel_1744/gring pixel_1744/VDD pixel_1744/GND pixel_1744/VREF pixel_1744/ROW_SEL
+ pixel_1744/NB1 pixel_1744/VBIAS pixel_1744/NB2 pixel_1744/AMP_IN pixel_1744/SF_IB
+ pixel_1744/PIX_OUT pixel_1744/CSA_VREF pixel
Xpixel_1733 pixel_1733/gring pixel_1733/VDD pixel_1733/GND pixel_1733/VREF pixel_1733/ROW_SEL
+ pixel_1733/NB1 pixel_1733/VBIAS pixel_1733/NB2 pixel_1733/AMP_IN pixel_1733/SF_IB
+ pixel_1733/PIX_OUT pixel_1733/CSA_VREF pixel
Xpixel_1722 pixel_1722/gring pixel_1722/VDD pixel_1722/GND pixel_1722/VREF pixel_1722/ROW_SEL
+ pixel_1722/NB1 pixel_1722/VBIAS pixel_1722/NB2 pixel_1722/AMP_IN pixel_1722/SF_IB
+ pixel_1722/PIX_OUT pixel_1722/CSA_VREF pixel
Xpixel_1711 pixel_1711/gring pixel_1711/VDD pixel_1711/GND pixel_1711/VREF pixel_1711/ROW_SEL
+ pixel_1711/NB1 pixel_1711/VBIAS pixel_1711/NB2 pixel_1711/AMP_IN pixel_1711/SF_IB
+ pixel_1711/PIX_OUT pixel_1711/CSA_VREF pixel
Xpixel_2478 pixel_2478/gring pixel_2478/VDD pixel_2478/GND pixel_2478/VREF pixel_2478/ROW_SEL
+ pixel_2478/NB1 pixel_2478/VBIAS pixel_2478/NB2 pixel_2478/AMP_IN pixel_2478/SF_IB
+ pixel_2478/PIX_OUT pixel_2478/CSA_VREF pixel
Xpixel_2467 pixel_2467/gring pixel_2467/VDD pixel_2467/GND pixel_2467/VREF pixel_2467/ROW_SEL
+ pixel_2467/NB1 pixel_2467/VBIAS pixel_2467/NB2 pixel_2467/AMP_IN pixel_2467/SF_IB
+ pixel_2467/PIX_OUT pixel_2467/CSA_VREF pixel
Xpixel_2456 pixel_2456/gring pixel_2456/VDD pixel_2456/GND pixel_2456/VREF pixel_2456/ROW_SEL
+ pixel_2456/NB1 pixel_2456/VBIAS pixel_2456/NB2 pixel_2456/AMP_IN pixel_2456/SF_IB
+ pixel_2456/PIX_OUT pixel_2456/CSA_VREF pixel
Xpixel_1777 pixel_1777/gring pixel_1777/VDD pixel_1777/GND pixel_1777/VREF pixel_1777/ROW_SEL
+ pixel_1777/NB1 pixel_1777/VBIAS pixel_1777/NB2 pixel_1777/AMP_IN pixel_1777/SF_IB
+ pixel_1777/PIX_OUT pixel_1777/CSA_VREF pixel
Xpixel_1766 pixel_1766/gring pixel_1766/VDD pixel_1766/GND pixel_1766/VREF pixel_1766/ROW_SEL
+ pixel_1766/NB1 pixel_1766/VBIAS pixel_1766/NB2 pixel_1766/AMP_IN pixel_1766/SF_IB
+ pixel_1766/PIX_OUT pixel_1766/CSA_VREF pixel
Xpixel_1755 pixel_1755/gring pixel_1755/VDD pixel_1755/GND pixel_1755/VREF pixel_1755/ROW_SEL
+ pixel_1755/NB1 pixel_1755/VBIAS pixel_1755/NB2 pixel_1755/AMP_IN pixel_1755/SF_IB
+ pixel_1755/PIX_OUT pixel_1755/CSA_VREF pixel
Xpixel_2489 pixel_2489/gring pixel_2489/VDD pixel_2489/GND pixel_2489/VREF pixel_2489/ROW_SEL
+ pixel_2489/NB1 pixel_2489/VBIAS pixel_2489/NB2 pixel_2489/AMP_IN pixel_2489/SF_IB
+ pixel_2489/PIX_OUT pixel_2489/CSA_VREF pixel
Xpixel_1799 pixel_1799/gring pixel_1799/VDD pixel_1799/GND pixel_1799/VREF pixel_1799/ROW_SEL
+ pixel_1799/NB1 pixel_1799/VBIAS pixel_1799/NB2 pixel_1799/AMP_IN pixel_1799/SF_IB
+ pixel_1799/PIX_OUT pixel_1799/CSA_VREF pixel
Xpixel_1788 pixel_1788/gring pixel_1788/VDD pixel_1788/GND pixel_1788/VREF pixel_1788/ROW_SEL
+ pixel_1788/NB1 pixel_1788/VBIAS pixel_1788/NB2 pixel_1788/AMP_IN pixel_1788/SF_IB
+ pixel_1788/PIX_OUT pixel_1788/CSA_VREF pixel
Xpixel_5060 pixel_5060/gring pixel_5060/VDD pixel_5060/GND pixel_5060/VREF pixel_5060/ROW_SEL
+ pixel_5060/NB1 pixel_5060/VBIAS pixel_5060/NB2 pixel_5060/AMP_IN pixel_5060/SF_IB
+ pixel_5060/PIX_OUT pixel_5060/CSA_VREF pixel
Xpixel_5071 pixel_5071/gring pixel_5071/VDD pixel_5071/GND pixel_5071/VREF pixel_5071/ROW_SEL
+ pixel_5071/NB1 pixel_5071/VBIAS pixel_5071/NB2 pixel_5071/AMP_IN pixel_5071/SF_IB
+ pixel_5071/PIX_OUT pixel_5071/CSA_VREF pixel
Xpixel_5082 pixel_5082/gring pixel_5082/VDD pixel_5082/GND pixel_5082/VREF pixel_5082/ROW_SEL
+ pixel_5082/NB1 pixel_5082/VBIAS pixel_5082/NB2 pixel_5082/AMP_IN pixel_5082/SF_IB
+ pixel_5082/PIX_OUT pixel_5082/CSA_VREF pixel
Xpixel_5093 pixel_5093/gring pixel_5093/VDD pixel_5093/GND pixel_5093/VREF pixel_5093/ROW_SEL
+ pixel_5093/NB1 pixel_5093/VBIAS pixel_5093/NB2 pixel_5093/AMP_IN pixel_5093/SF_IB
+ pixel_5093/PIX_OUT pixel_5093/CSA_VREF pixel
Xpixel_4370 pixel_4370/gring pixel_4370/VDD pixel_4370/GND pixel_4370/VREF pixel_4370/ROW_SEL
+ pixel_4370/NB1 pixel_4370/VBIAS pixel_4370/NB2 pixel_4370/AMP_IN pixel_4370/SF_IB
+ pixel_4370/PIX_OUT pixel_4370/CSA_VREF pixel
Xpixel_4381 pixel_4381/gring pixel_4381/VDD pixel_4381/GND pixel_4381/VREF pixel_4381/ROW_SEL
+ pixel_4381/NB1 pixel_4381/VBIAS pixel_4381/NB2 pixel_4381/AMP_IN pixel_4381/SF_IB
+ pixel_4381/PIX_OUT pixel_4381/CSA_VREF pixel
Xpixel_4392 pixel_4392/gring pixel_4392/VDD pixel_4392/GND pixel_4392/VREF pixel_4392/ROW_SEL
+ pixel_4392/NB1 pixel_4392/VBIAS pixel_4392/NB2 pixel_4392/AMP_IN pixel_4392/SF_IB
+ pixel_4392/PIX_OUT pixel_4392/CSA_VREF pixel
Xpixel_3691 pixel_3691/gring pixel_3691/VDD pixel_3691/GND pixel_3691/VREF pixel_3691/ROW_SEL
+ pixel_3691/NB1 pixel_3691/VBIAS pixel_3691/NB2 pixel_3691/AMP_IN pixel_3691/SF_IB
+ pixel_3691/PIX_OUT pixel_3691/CSA_VREF pixel
Xpixel_3680 pixel_3680/gring pixel_3680/VDD pixel_3680/GND pixel_3680/VREF pixel_3680/ROW_SEL
+ pixel_3680/NB1 pixel_3680/VBIAS pixel_3680/NB2 pixel_3680/AMP_IN pixel_3680/SF_IB
+ pixel_3680/PIX_OUT pixel_3680/CSA_VREF pixel
Xpixel_2990 pixel_2990/gring pixel_2990/VDD pixel_2990/GND pixel_2990/VREF pixel_2990/ROW_SEL
+ pixel_2990/NB1 pixel_2990/VBIAS pixel_2990/NB2 pixel_2990/AMP_IN pixel_2990/SF_IB
+ pixel_2990/PIX_OUT pixel_2990/CSA_VREF pixel
Xpixel_1029 pixel_1029/gring pixel_1029/VDD pixel_1029/GND pixel_1029/VREF pixel_1029/ROW_SEL
+ pixel_1029/NB1 pixel_1029/VBIAS pixel_1029/NB2 pixel_1029/AMP_IN pixel_1029/SF_IB
+ pixel_1029/PIX_OUT pixel_1029/CSA_VREF pixel
Xpixel_1018 pixel_1018/gring pixel_1018/VDD pixel_1018/GND pixel_1018/VREF pixel_1018/ROW_SEL
+ pixel_1018/NB1 pixel_1018/VBIAS pixel_1018/NB2 pixel_1018/AMP_IN pixel_1018/SF_IB
+ pixel_1018/PIX_OUT pixel_1018/CSA_VREF pixel
Xpixel_1007 pixel_1007/gring pixel_1007/VDD pixel_1007/GND pixel_1007/VREF pixel_1007/ROW_SEL
+ pixel_1007/NB1 pixel_1007/VBIAS pixel_1007/NB2 pixel_1007/AMP_IN pixel_1007/SF_IB
+ pixel_1007/PIX_OUT pixel_1007/CSA_VREF pixel
Xpixel_9304 pixel_9304/gring pixel_9304/VDD pixel_9304/GND pixel_9304/VREF pixel_9304/ROW_SEL
+ pixel_9304/NB1 pixel_9304/VBIAS pixel_9304/NB2 pixel_9304/AMP_IN pixel_9304/SF_IB
+ pixel_9304/PIX_OUT pixel_9304/CSA_VREF pixel
Xpixel_9337 pixel_9337/gring pixel_9337/VDD pixel_9337/GND pixel_9337/VREF pixel_9337/ROW_SEL
+ pixel_9337/NB1 pixel_9337/VBIAS pixel_9337/NB2 pixel_9337/AMP_IN pixel_9337/SF_IB
+ pixel_9337/PIX_OUT pixel_9337/CSA_VREF pixel
Xpixel_9326 pixel_9326/gring pixel_9326/VDD pixel_9326/GND pixel_9326/VREF pixel_9326/ROW_SEL
+ pixel_9326/NB1 pixel_9326/VBIAS pixel_9326/NB2 pixel_9326/AMP_IN pixel_9326/SF_IB
+ pixel_9326/PIX_OUT pixel_9326/CSA_VREF pixel
Xpixel_9315 pixel_9315/gring pixel_9315/VDD pixel_9315/GND pixel_9315/VREF pixel_9315/ROW_SEL
+ pixel_9315/NB1 pixel_9315/VBIAS pixel_9315/NB2 pixel_9315/AMP_IN pixel_9315/SF_IB
+ pixel_9315/PIX_OUT pixel_9315/CSA_VREF pixel
Xpixel_8636 pixel_8636/gring pixel_8636/VDD pixel_8636/GND pixel_8636/VREF pixel_8636/ROW_SEL
+ pixel_8636/NB1 pixel_8636/VBIAS pixel_8636/NB2 pixel_8636/AMP_IN pixel_8636/SF_IB
+ pixel_8636/PIX_OUT pixel_8636/CSA_VREF pixel
Xpixel_8625 pixel_8625/gring pixel_8625/VDD pixel_8625/GND pixel_8625/VREF pixel_8625/ROW_SEL
+ pixel_8625/NB1 pixel_8625/VBIAS pixel_8625/NB2 pixel_8625/AMP_IN pixel_8625/SF_IB
+ pixel_8625/PIX_OUT pixel_8625/CSA_VREF pixel
Xpixel_8614 pixel_8614/gring pixel_8614/VDD pixel_8614/GND pixel_8614/VREF pixel_8614/ROW_SEL
+ pixel_8614/NB1 pixel_8614/VBIAS pixel_8614/NB2 pixel_8614/AMP_IN pixel_8614/SF_IB
+ pixel_8614/PIX_OUT pixel_8614/CSA_VREF pixel
Xpixel_8603 pixel_8603/gring pixel_8603/VDD pixel_8603/GND pixel_8603/VREF pixel_8603/ROW_SEL
+ pixel_8603/NB1 pixel_8603/VBIAS pixel_8603/NB2 pixel_8603/AMP_IN pixel_8603/SF_IB
+ pixel_8603/PIX_OUT pixel_8603/CSA_VREF pixel
Xpixel_9359 pixel_9359/gring pixel_9359/VDD pixel_9359/GND pixel_9359/VREF pixel_9359/ROW_SEL
+ pixel_9359/NB1 pixel_9359/VBIAS pixel_9359/NB2 pixel_9359/AMP_IN pixel_9359/SF_IB
+ pixel_9359/PIX_OUT pixel_9359/CSA_VREF pixel
Xpixel_9348 pixel_9348/gring pixel_9348/VDD pixel_9348/GND pixel_9348/VREF pixel_9348/ROW_SEL
+ pixel_9348/NB1 pixel_9348/VBIAS pixel_9348/NB2 pixel_9348/AMP_IN pixel_9348/SF_IB
+ pixel_9348/PIX_OUT pixel_9348/CSA_VREF pixel
Xpixel_8669 pixel_8669/gring pixel_8669/VDD pixel_8669/GND pixel_8669/VREF pixel_8669/ROW_SEL
+ pixel_8669/NB1 pixel_8669/VBIAS pixel_8669/NB2 pixel_8669/AMP_IN pixel_8669/SF_IB
+ pixel_8669/PIX_OUT pixel_8669/CSA_VREF pixel
Xpixel_8658 pixel_8658/gring pixel_8658/VDD pixel_8658/GND pixel_8658/VREF pixel_8658/ROW_SEL
+ pixel_8658/NB1 pixel_8658/VBIAS pixel_8658/NB2 pixel_8658/AMP_IN pixel_8658/SF_IB
+ pixel_8658/PIX_OUT pixel_8658/CSA_VREF pixel
Xpixel_8647 pixel_8647/gring pixel_8647/VDD pixel_8647/GND pixel_8647/VREF pixel_8647/ROW_SEL
+ pixel_8647/NB1 pixel_8647/VBIAS pixel_8647/NB2 pixel_8647/AMP_IN pixel_8647/SF_IB
+ pixel_8647/PIX_OUT pixel_8647/CSA_VREF pixel
Xpixel_7902 pixel_7902/gring pixel_7902/VDD pixel_7902/GND pixel_7902/VREF pixel_7902/ROW_SEL
+ pixel_7902/NB1 pixel_7902/VBIAS pixel_7902/NB2 pixel_7902/AMP_IN pixel_7902/SF_IB
+ pixel_7902/PIX_OUT pixel_7902/CSA_VREF pixel
Xpixel_7913 pixel_7913/gring pixel_7913/VDD pixel_7913/GND pixel_7913/VREF pixel_7913/ROW_SEL
+ pixel_7913/NB1 pixel_7913/VBIAS pixel_7913/NB2 pixel_7913/AMP_IN pixel_7913/SF_IB
+ pixel_7913/PIX_OUT pixel_7913/CSA_VREF pixel
Xpixel_7924 pixel_7924/gring pixel_7924/VDD pixel_7924/GND pixel_7924/VREF pixel_7924/ROW_SEL
+ pixel_7924/NB1 pixel_7924/VBIAS pixel_7924/NB2 pixel_7924/AMP_IN pixel_7924/SF_IB
+ pixel_7924/PIX_OUT pixel_7924/CSA_VREF pixel
Xpixel_7935 pixel_7935/gring pixel_7935/VDD pixel_7935/GND pixel_7935/VREF pixel_7935/ROW_SEL
+ pixel_7935/NB1 pixel_7935/VBIAS pixel_7935/NB2 pixel_7935/AMP_IN pixel_7935/SF_IB
+ pixel_7935/PIX_OUT pixel_7935/CSA_VREF pixel
Xpixel_7946 pixel_7946/gring pixel_7946/VDD pixel_7946/GND pixel_7946/VREF pixel_7946/ROW_SEL
+ pixel_7946/NB1 pixel_7946/VBIAS pixel_7946/NB2 pixel_7946/AMP_IN pixel_7946/SF_IB
+ pixel_7946/PIX_OUT pixel_7946/CSA_VREF pixel
Xpixel_7957 pixel_7957/gring pixel_7957/VDD pixel_7957/GND pixel_7957/VREF pixel_7957/ROW_SEL
+ pixel_7957/NB1 pixel_7957/VBIAS pixel_7957/NB2 pixel_7957/AMP_IN pixel_7957/SF_IB
+ pixel_7957/PIX_OUT pixel_7957/CSA_VREF pixel
Xpixel_7968 pixel_7968/gring pixel_7968/VDD pixel_7968/GND pixel_7968/VREF pixel_7968/ROW_SEL
+ pixel_7968/NB1 pixel_7968/VBIAS pixel_7968/NB2 pixel_7968/AMP_IN pixel_7968/SF_IB
+ pixel_7968/PIX_OUT pixel_7968/CSA_VREF pixel
Xpixel_7979 pixel_7979/gring pixel_7979/VDD pixel_7979/GND pixel_7979/VREF pixel_7979/ROW_SEL
+ pixel_7979/NB1 pixel_7979/VBIAS pixel_7979/NB2 pixel_7979/AMP_IN pixel_7979/SF_IB
+ pixel_7979/PIX_OUT pixel_7979/CSA_VREF pixel
Xpixel_2220 pixel_2220/gring pixel_2220/VDD pixel_2220/GND pixel_2220/VREF pixel_2220/ROW_SEL
+ pixel_2220/NB1 pixel_2220/VBIAS pixel_2220/NB2 pixel_2220/AMP_IN pixel_2220/SF_IB
+ pixel_2220/PIX_OUT pixel_2220/CSA_VREF pixel
Xpixel_2253 pixel_2253/gring pixel_2253/VDD pixel_2253/GND pixel_2253/VREF pixel_2253/ROW_SEL
+ pixel_2253/NB1 pixel_2253/VBIAS pixel_2253/NB2 pixel_2253/AMP_IN pixel_2253/SF_IB
+ pixel_2253/PIX_OUT pixel_2253/CSA_VREF pixel
Xpixel_2242 pixel_2242/gring pixel_2242/VDD pixel_2242/GND pixel_2242/VREF pixel_2242/ROW_SEL
+ pixel_2242/NB1 pixel_2242/VBIAS pixel_2242/NB2 pixel_2242/AMP_IN pixel_2242/SF_IB
+ pixel_2242/PIX_OUT pixel_2242/CSA_VREF pixel
Xpixel_2231 pixel_2231/gring pixel_2231/VDD pixel_2231/GND pixel_2231/VREF pixel_2231/ROW_SEL
+ pixel_2231/NB1 pixel_2231/VBIAS pixel_2231/NB2 pixel_2231/AMP_IN pixel_2231/SF_IB
+ pixel_2231/PIX_OUT pixel_2231/CSA_VREF pixel
Xpixel_1552 pixel_1552/gring pixel_1552/VDD pixel_1552/GND pixel_1552/VREF pixel_1552/ROW_SEL
+ pixel_1552/NB1 pixel_1552/VBIAS pixel_1552/NB2 pixel_1552/AMP_IN pixel_1552/SF_IB
+ pixel_1552/PIX_OUT pixel_1552/CSA_VREF pixel
Xpixel_1541 pixel_1541/gring pixel_1541/VDD pixel_1541/GND pixel_1541/VREF pixel_1541/ROW_SEL
+ pixel_1541/NB1 pixel_1541/VBIAS pixel_1541/NB2 pixel_1541/AMP_IN pixel_1541/SF_IB
+ pixel_1541/PIX_OUT pixel_1541/CSA_VREF pixel
Xpixel_1530 pixel_1530/gring pixel_1530/VDD pixel_1530/GND pixel_1530/VREF pixel_1530/ROW_SEL
+ pixel_1530/NB1 pixel_1530/VBIAS pixel_1530/NB2 pixel_1530/AMP_IN pixel_1530/SF_IB
+ pixel_1530/PIX_OUT pixel_1530/CSA_VREF pixel
Xpixel_2297 pixel_2297/gring pixel_2297/VDD pixel_2297/GND pixel_2297/VREF pixel_2297/ROW_SEL
+ pixel_2297/NB1 pixel_2297/VBIAS pixel_2297/NB2 pixel_2297/AMP_IN pixel_2297/SF_IB
+ pixel_2297/PIX_OUT pixel_2297/CSA_VREF pixel
Xpixel_2286 pixel_2286/gring pixel_2286/VDD pixel_2286/GND pixel_2286/VREF pixel_2286/ROW_SEL
+ pixel_2286/NB1 pixel_2286/VBIAS pixel_2286/NB2 pixel_2286/AMP_IN pixel_2286/SF_IB
+ pixel_2286/PIX_OUT pixel_2286/CSA_VREF pixel
Xpixel_2275 pixel_2275/gring pixel_2275/VDD pixel_2275/GND pixel_2275/VREF pixel_2275/ROW_SEL
+ pixel_2275/NB1 pixel_2275/VBIAS pixel_2275/NB2 pixel_2275/AMP_IN pixel_2275/SF_IB
+ pixel_2275/PIX_OUT pixel_2275/CSA_VREF pixel
Xpixel_2264 pixel_2264/gring pixel_2264/VDD pixel_2264/GND pixel_2264/VREF pixel_2264/ROW_SEL
+ pixel_2264/NB1 pixel_2264/VBIAS pixel_2264/NB2 pixel_2264/AMP_IN pixel_2264/SF_IB
+ pixel_2264/PIX_OUT pixel_2264/CSA_VREF pixel
Xpixel_1585 pixel_1585/gring pixel_1585/VDD pixel_1585/GND pixel_1585/VREF pixel_1585/ROW_SEL
+ pixel_1585/NB1 pixel_1585/VBIAS pixel_1585/NB2 pixel_1585/AMP_IN pixel_1585/SF_IB
+ pixel_1585/PIX_OUT pixel_1585/CSA_VREF pixel
Xpixel_1574 pixel_1574/gring pixel_1574/VDD pixel_1574/GND pixel_1574/VREF pixel_1574/ROW_SEL
+ pixel_1574/NB1 pixel_1574/VBIAS pixel_1574/NB2 pixel_1574/AMP_IN pixel_1574/SF_IB
+ pixel_1574/PIX_OUT pixel_1574/CSA_VREF pixel
Xpixel_1563 pixel_1563/gring pixel_1563/VDD pixel_1563/GND pixel_1563/VREF pixel_1563/ROW_SEL
+ pixel_1563/NB1 pixel_1563/VBIAS pixel_1563/NB2 pixel_1563/AMP_IN pixel_1563/SF_IB
+ pixel_1563/PIX_OUT pixel_1563/CSA_VREF pixel
Xpixel_1596 pixel_1596/gring pixel_1596/VDD pixel_1596/GND pixel_1596/VREF pixel_1596/ROW_SEL
+ pixel_1596/NB1 pixel_1596/VBIAS pixel_1596/NB2 pixel_1596/AMP_IN pixel_1596/SF_IB
+ pixel_1596/PIX_OUT pixel_1596/CSA_VREF pixel
Xpixel_9860 pixel_9860/gring pixel_9860/VDD pixel_9860/GND pixel_9860/VREF pixel_9860/ROW_SEL
+ pixel_9860/NB1 pixel_9860/VBIAS pixel_9860/NB2 pixel_9860/AMP_IN pixel_9860/SF_IB
+ pixel_9860/PIX_OUT pixel_9860/CSA_VREF pixel
Xpixel_9871 pixel_9871/gring pixel_9871/VDD pixel_9871/GND pixel_9871/VREF pixel_9871/ROW_SEL
+ pixel_9871/NB1 pixel_9871/VBIAS pixel_9871/NB2 pixel_9871/AMP_IN pixel_9871/SF_IB
+ pixel_9871/PIX_OUT pixel_9871/CSA_VREF pixel
Xpixel_9882 pixel_9882/gring pixel_9882/VDD pixel_9882/GND pixel_9882/VREF pixel_9882/ROW_SEL
+ pixel_9882/NB1 pixel_9882/VBIAS pixel_9882/NB2 pixel_9882/AMP_IN pixel_9882/SF_IB
+ pixel_9882/PIX_OUT pixel_9882/CSA_VREF pixel
Xpixel_9893 pixel_9893/gring pixel_9893/VDD pixel_9893/GND pixel_9893/VREF pixel_9893/ROW_SEL
+ pixel_9893/NB1 pixel_9893/VBIAS pixel_9893/NB2 pixel_9893/AMP_IN pixel_9893/SF_IB
+ pixel_9893/PIX_OUT pixel_9893/CSA_VREF pixel
Xpixel_7209 pixel_7209/gring pixel_7209/VDD pixel_7209/GND pixel_7209/VREF pixel_7209/ROW_SEL
+ pixel_7209/NB1 pixel_7209/VBIAS pixel_7209/NB2 pixel_7209/AMP_IN pixel_7209/SF_IB
+ pixel_7209/PIX_OUT pixel_7209/CSA_VREF pixel
Xpixel_6508 pixel_6508/gring pixel_6508/VDD pixel_6508/GND pixel_6508/VREF pixel_6508/ROW_SEL
+ pixel_6508/NB1 pixel_6508/VBIAS pixel_6508/NB2 pixel_6508/AMP_IN pixel_6508/SF_IB
+ pixel_6508/PIX_OUT pixel_6508/CSA_VREF pixel
Xpixel_6519 pixel_6519/gring pixel_6519/VDD pixel_6519/GND pixel_6519/VREF pixel_6519/ROW_SEL
+ pixel_6519/NB1 pixel_6519/VBIAS pixel_6519/NB2 pixel_6519/AMP_IN pixel_6519/SF_IB
+ pixel_6519/PIX_OUT pixel_6519/CSA_VREF pixel
Xpixel_5807 pixel_5807/gring pixel_5807/VDD pixel_5807/GND pixel_5807/VREF pixel_5807/ROW_SEL
+ pixel_5807/NB1 pixel_5807/VBIAS pixel_5807/NB2 pixel_5807/AMP_IN pixel_5807/SF_IB
+ pixel_5807/PIX_OUT pixel_5807/CSA_VREF pixel
Xpixel_5818 pixel_5818/gring pixel_5818/VDD pixel_5818/GND pixel_5818/VREF pixel_5818/ROW_SEL
+ pixel_5818/NB1 pixel_5818/VBIAS pixel_5818/NB2 pixel_5818/AMP_IN pixel_5818/SF_IB
+ pixel_5818/PIX_OUT pixel_5818/CSA_VREF pixel
Xpixel_5829 pixel_5829/gring pixel_5829/VDD pixel_5829/GND pixel_5829/VREF pixel_5829/ROW_SEL
+ pixel_5829/NB1 pixel_5829/VBIAS pixel_5829/NB2 pixel_5829/AMP_IN pixel_5829/SF_IB
+ pixel_5829/PIX_OUT pixel_5829/CSA_VREF pixel
Xpixel_9112 pixel_9112/gring pixel_9112/VDD pixel_9112/GND pixel_9112/VREF pixel_9112/ROW_SEL
+ pixel_9112/NB1 pixel_9112/VBIAS pixel_9112/NB2 pixel_9112/AMP_IN pixel_9112/SF_IB
+ pixel_9112/PIX_OUT pixel_9112/CSA_VREF pixel
Xpixel_9101 pixel_9101/gring pixel_9101/VDD pixel_9101/GND pixel_9101/VREF pixel_9101/ROW_SEL
+ pixel_9101/NB1 pixel_9101/VBIAS pixel_9101/NB2 pixel_9101/AMP_IN pixel_9101/SF_IB
+ pixel_9101/PIX_OUT pixel_9101/CSA_VREF pixel
Xpixel_8411 pixel_8411/gring pixel_8411/VDD pixel_8411/GND pixel_8411/VREF pixel_8411/ROW_SEL
+ pixel_8411/NB1 pixel_8411/VBIAS pixel_8411/NB2 pixel_8411/AMP_IN pixel_8411/SF_IB
+ pixel_8411/PIX_OUT pixel_8411/CSA_VREF pixel
Xpixel_8400 pixel_8400/gring pixel_8400/VDD pixel_8400/GND pixel_8400/VREF pixel_8400/ROW_SEL
+ pixel_8400/NB1 pixel_8400/VBIAS pixel_8400/NB2 pixel_8400/AMP_IN pixel_8400/SF_IB
+ pixel_8400/PIX_OUT pixel_8400/CSA_VREF pixel
Xpixel_9145 pixel_9145/gring pixel_9145/VDD pixel_9145/GND pixel_9145/VREF pixel_9145/ROW_SEL
+ pixel_9145/NB1 pixel_9145/VBIAS pixel_9145/NB2 pixel_9145/AMP_IN pixel_9145/SF_IB
+ pixel_9145/PIX_OUT pixel_9145/CSA_VREF pixel
Xpixel_9134 pixel_9134/gring pixel_9134/VDD pixel_9134/GND pixel_9134/VREF pixel_9134/ROW_SEL
+ pixel_9134/NB1 pixel_9134/VBIAS pixel_9134/NB2 pixel_9134/AMP_IN pixel_9134/SF_IB
+ pixel_9134/PIX_OUT pixel_9134/CSA_VREF pixel
Xpixel_9123 pixel_9123/gring pixel_9123/VDD pixel_9123/GND pixel_9123/VREF pixel_9123/ROW_SEL
+ pixel_9123/NB1 pixel_9123/VBIAS pixel_9123/NB2 pixel_9123/AMP_IN pixel_9123/SF_IB
+ pixel_9123/PIX_OUT pixel_9123/CSA_VREF pixel
Xpixel_8433 pixel_8433/gring pixel_8433/VDD pixel_8433/GND pixel_8433/VREF pixel_8433/ROW_SEL
+ pixel_8433/NB1 pixel_8433/VBIAS pixel_8433/NB2 pixel_8433/AMP_IN pixel_8433/SF_IB
+ pixel_8433/PIX_OUT pixel_8433/CSA_VREF pixel
Xpixel_8422 pixel_8422/gring pixel_8422/VDD pixel_8422/GND pixel_8422/VREF pixel_8422/ROW_SEL
+ pixel_8422/NB1 pixel_8422/VBIAS pixel_8422/NB2 pixel_8422/AMP_IN pixel_8422/SF_IB
+ pixel_8422/PIX_OUT pixel_8422/CSA_VREF pixel
Xpixel_9189 pixel_9189/gring pixel_9189/VDD pixel_9189/GND pixel_9189/VREF pixel_9189/ROW_SEL
+ pixel_9189/NB1 pixel_9189/VBIAS pixel_9189/NB2 pixel_9189/AMP_IN pixel_9189/SF_IB
+ pixel_9189/PIX_OUT pixel_9189/CSA_VREF pixel
Xpixel_9178 pixel_9178/gring pixel_9178/VDD pixel_9178/GND pixel_9178/VREF pixel_9178/ROW_SEL
+ pixel_9178/NB1 pixel_9178/VBIAS pixel_9178/NB2 pixel_9178/AMP_IN pixel_9178/SF_IB
+ pixel_9178/PIX_OUT pixel_9178/CSA_VREF pixel
Xpixel_9167 pixel_9167/gring pixel_9167/VDD pixel_9167/GND pixel_9167/VREF pixel_9167/ROW_SEL
+ pixel_9167/NB1 pixel_9167/VBIAS pixel_9167/NB2 pixel_9167/AMP_IN pixel_9167/SF_IB
+ pixel_9167/PIX_OUT pixel_9167/CSA_VREF pixel
Xpixel_9156 pixel_9156/gring pixel_9156/VDD pixel_9156/GND pixel_9156/VREF pixel_9156/ROW_SEL
+ pixel_9156/NB1 pixel_9156/VBIAS pixel_9156/NB2 pixel_9156/AMP_IN pixel_9156/SF_IB
+ pixel_9156/PIX_OUT pixel_9156/CSA_VREF pixel
Xpixel_8444 pixel_8444/gring pixel_8444/VDD pixel_8444/GND pixel_8444/VREF pixel_8444/ROW_SEL
+ pixel_8444/NB1 pixel_8444/VBIAS pixel_8444/NB2 pixel_8444/AMP_IN pixel_8444/SF_IB
+ pixel_8444/PIX_OUT pixel_8444/CSA_VREF pixel
Xpixel_8455 pixel_8455/gring pixel_8455/VDD pixel_8455/GND pixel_8455/VREF pixel_8455/ROW_SEL
+ pixel_8455/NB1 pixel_8455/VBIAS pixel_8455/NB2 pixel_8455/AMP_IN pixel_8455/SF_IB
+ pixel_8455/PIX_OUT pixel_8455/CSA_VREF pixel
Xpixel_8466 pixel_8466/gring pixel_8466/VDD pixel_8466/GND pixel_8466/VREF pixel_8466/ROW_SEL
+ pixel_8466/NB1 pixel_8466/VBIAS pixel_8466/NB2 pixel_8466/AMP_IN pixel_8466/SF_IB
+ pixel_8466/PIX_OUT pixel_8466/CSA_VREF pixel
Xpixel_8477 pixel_8477/gring pixel_8477/VDD pixel_8477/GND pixel_8477/VREF pixel_8477/ROW_SEL
+ pixel_8477/NB1 pixel_8477/VBIAS pixel_8477/NB2 pixel_8477/AMP_IN pixel_8477/SF_IB
+ pixel_8477/PIX_OUT pixel_8477/CSA_VREF pixel
Xpixel_7710 pixel_7710/gring pixel_7710/VDD pixel_7710/GND pixel_7710/VREF pixel_7710/ROW_SEL
+ pixel_7710/NB1 pixel_7710/VBIAS pixel_7710/NB2 pixel_7710/AMP_IN pixel_7710/SF_IB
+ pixel_7710/PIX_OUT pixel_7710/CSA_VREF pixel
Xpixel_7721 pixel_7721/gring pixel_7721/VDD pixel_7721/GND pixel_7721/VREF pixel_7721/ROW_SEL
+ pixel_7721/NB1 pixel_7721/VBIAS pixel_7721/NB2 pixel_7721/AMP_IN pixel_7721/SF_IB
+ pixel_7721/PIX_OUT pixel_7721/CSA_VREF pixel
Xpixel_7732 pixel_7732/gring pixel_7732/VDD pixel_7732/GND pixel_7732/VREF pixel_7732/ROW_SEL
+ pixel_7732/NB1 pixel_7732/VBIAS pixel_7732/NB2 pixel_7732/AMP_IN pixel_7732/SF_IB
+ pixel_7732/PIX_OUT pixel_7732/CSA_VREF pixel
Xpixel_8488 pixel_8488/gring pixel_8488/VDD pixel_8488/GND pixel_8488/VREF pixel_8488/ROW_SEL
+ pixel_8488/NB1 pixel_8488/VBIAS pixel_8488/NB2 pixel_8488/AMP_IN pixel_8488/SF_IB
+ pixel_8488/PIX_OUT pixel_8488/CSA_VREF pixel
Xpixel_8499 pixel_8499/gring pixel_8499/VDD pixel_8499/GND pixel_8499/VREF pixel_8499/ROW_SEL
+ pixel_8499/NB1 pixel_8499/VBIAS pixel_8499/NB2 pixel_8499/AMP_IN pixel_8499/SF_IB
+ pixel_8499/PIX_OUT pixel_8499/CSA_VREF pixel
Xpixel_7743 pixel_7743/gring pixel_7743/VDD pixel_7743/GND pixel_7743/VREF pixel_7743/ROW_SEL
+ pixel_7743/NB1 pixel_7743/VBIAS pixel_7743/NB2 pixel_7743/AMP_IN pixel_7743/SF_IB
+ pixel_7743/PIX_OUT pixel_7743/CSA_VREF pixel
Xpixel_7754 pixel_7754/gring pixel_7754/VDD pixel_7754/GND pixel_7754/VREF pixel_7754/ROW_SEL
+ pixel_7754/NB1 pixel_7754/VBIAS pixel_7754/NB2 pixel_7754/AMP_IN pixel_7754/SF_IB
+ pixel_7754/PIX_OUT pixel_7754/CSA_VREF pixel
Xpixel_7765 pixel_7765/gring pixel_7765/VDD pixel_7765/GND pixel_7765/VREF pixel_7765/ROW_SEL
+ pixel_7765/NB1 pixel_7765/VBIAS pixel_7765/NB2 pixel_7765/AMP_IN pixel_7765/SF_IB
+ pixel_7765/PIX_OUT pixel_7765/CSA_VREF pixel
Xpixel_7776 pixel_7776/gring pixel_7776/VDD pixel_7776/GND pixel_7776/VREF pixel_7776/ROW_SEL
+ pixel_7776/NB1 pixel_7776/VBIAS pixel_7776/NB2 pixel_7776/AMP_IN pixel_7776/SF_IB
+ pixel_7776/PIX_OUT pixel_7776/CSA_VREF pixel
Xpixel_7787 pixel_7787/gring pixel_7787/VDD pixel_7787/GND pixel_7787/VREF pixel_7787/ROW_SEL
+ pixel_7787/NB1 pixel_7787/VBIAS pixel_7787/NB2 pixel_7787/AMP_IN pixel_7787/SF_IB
+ pixel_7787/PIX_OUT pixel_7787/CSA_VREF pixel
Xpixel_7798 pixel_7798/gring pixel_7798/VDD pixel_7798/GND pixel_7798/VREF pixel_7798/ROW_SEL
+ pixel_7798/NB1 pixel_7798/VBIAS pixel_7798/NB2 pixel_7798/AMP_IN pixel_7798/SF_IB
+ pixel_7798/PIX_OUT pixel_7798/CSA_VREF pixel
Xpixel_2072 pixel_2072/gring pixel_2072/VDD pixel_2072/GND pixel_2072/VREF pixel_2072/ROW_SEL
+ pixel_2072/NB1 pixel_2072/VBIAS pixel_2072/NB2 pixel_2072/AMP_IN pixel_2072/SF_IB
+ pixel_2072/PIX_OUT pixel_2072/CSA_VREF pixel
Xpixel_2061 pixel_2061/gring pixel_2061/VDD pixel_2061/GND pixel_2061/VREF pixel_2061/ROW_SEL
+ pixel_2061/NB1 pixel_2061/VBIAS pixel_2061/NB2 pixel_2061/AMP_IN pixel_2061/SF_IB
+ pixel_2061/PIX_OUT pixel_2061/CSA_VREF pixel
Xpixel_2050 pixel_2050/gring pixel_2050/VDD pixel_2050/GND pixel_2050/VREF pixel_2050/ROW_SEL
+ pixel_2050/NB1 pixel_2050/VBIAS pixel_2050/NB2 pixel_2050/AMP_IN pixel_2050/SF_IB
+ pixel_2050/PIX_OUT pixel_2050/CSA_VREF pixel
Xpixel_1360 pixel_1360/gring pixel_1360/VDD pixel_1360/GND pixel_1360/VREF pixel_1360/ROW_SEL
+ pixel_1360/NB1 pixel_1360/VBIAS pixel_1360/NB2 pixel_1360/AMP_IN pixel_1360/SF_IB
+ pixel_1360/PIX_OUT pixel_1360/CSA_VREF pixel
Xpixel_2094 pixel_2094/gring pixel_2094/VDD pixel_2094/GND pixel_2094/VREF pixel_2094/ROW_SEL
+ pixel_2094/NB1 pixel_2094/VBIAS pixel_2094/NB2 pixel_2094/AMP_IN pixel_2094/SF_IB
+ pixel_2094/PIX_OUT pixel_2094/CSA_VREF pixel
Xpixel_2083 pixel_2083/gring pixel_2083/VDD pixel_2083/GND pixel_2083/VREF pixel_2083/ROW_SEL
+ pixel_2083/NB1 pixel_2083/VBIAS pixel_2083/NB2 pixel_2083/AMP_IN pixel_2083/SF_IB
+ pixel_2083/PIX_OUT pixel_2083/CSA_VREF pixel
Xpixel_1393 pixel_1393/gring pixel_1393/VDD pixel_1393/GND pixel_1393/VREF pixel_1393/ROW_SEL
+ pixel_1393/NB1 pixel_1393/VBIAS pixel_1393/NB2 pixel_1393/AMP_IN pixel_1393/SF_IB
+ pixel_1393/PIX_OUT pixel_1393/CSA_VREF pixel
Xpixel_1382 pixel_1382/gring pixel_1382/VDD pixel_1382/GND pixel_1382/VREF pixel_1382/ROW_SEL
+ pixel_1382/NB1 pixel_1382/VBIAS pixel_1382/NB2 pixel_1382/AMP_IN pixel_1382/SF_IB
+ pixel_1382/PIX_OUT pixel_1382/CSA_VREF pixel
Xpixel_1371 pixel_1371/gring pixel_1371/VDD pixel_1371/GND pixel_1371/VREF pixel_1371/ROW_SEL
+ pixel_1371/NB1 pixel_1371/VBIAS pixel_1371/NB2 pixel_1371/AMP_IN pixel_1371/SF_IB
+ pixel_1371/PIX_OUT pixel_1371/CSA_VREF pixel
Xpixel_9690 pixel_9690/gring pixel_9690/VDD pixel_9690/GND pixel_9690/VREF pixel_9690/ROW_SEL
+ pixel_9690/NB1 pixel_9690/VBIAS pixel_9690/NB2 pixel_9690/AMP_IN pixel_9690/SF_IB
+ pixel_9690/PIX_OUT pixel_9690/CSA_VREF pixel
Xpixel_419 pixel_419/gring pixel_419/VDD pixel_419/GND pixel_419/VREF pixel_419/ROW_SEL
+ pixel_419/NB1 pixel_419/VBIAS pixel_419/NB2 pixel_419/AMP_IN pixel_419/SF_IB pixel_419/PIX_OUT
+ pixel_419/CSA_VREF pixel
Xpixel_408 pixel_408/gring pixel_408/VDD pixel_408/GND pixel_408/VREF pixel_408/ROW_SEL
+ pixel_408/NB1 pixel_408/VBIAS pixel_408/NB2 pixel_408/AMP_IN pixel_408/SF_IB pixel_408/PIX_OUT
+ pixel_408/CSA_VREF pixel
Xpixel_7006 pixel_7006/gring pixel_7006/VDD pixel_7006/GND pixel_7006/VREF pixel_7006/ROW_SEL
+ pixel_7006/NB1 pixel_7006/VBIAS pixel_7006/NB2 pixel_7006/AMP_IN pixel_7006/SF_IB
+ pixel_7006/PIX_OUT pixel_7006/CSA_VREF pixel
Xpixel_7017 pixel_7017/gring pixel_7017/VDD pixel_7017/GND pixel_7017/VREF pixel_7017/ROW_SEL
+ pixel_7017/NB1 pixel_7017/VBIAS pixel_7017/NB2 pixel_7017/AMP_IN pixel_7017/SF_IB
+ pixel_7017/PIX_OUT pixel_7017/CSA_VREF pixel
Xpixel_7028 pixel_7028/gring pixel_7028/VDD pixel_7028/GND pixel_7028/VREF pixel_7028/ROW_SEL
+ pixel_7028/NB1 pixel_7028/VBIAS pixel_7028/NB2 pixel_7028/AMP_IN pixel_7028/SF_IB
+ pixel_7028/PIX_OUT pixel_7028/CSA_VREF pixel
Xpixel_7039 pixel_7039/gring pixel_7039/VDD pixel_7039/GND pixel_7039/VREF pixel_7039/ROW_SEL
+ pixel_7039/NB1 pixel_7039/VBIAS pixel_7039/NB2 pixel_7039/AMP_IN pixel_7039/SF_IB
+ pixel_7039/PIX_OUT pixel_7039/CSA_VREF pixel
Xpixel_6305 pixel_6305/gring pixel_6305/VDD pixel_6305/GND pixel_6305/VREF pixel_6305/ROW_SEL
+ pixel_6305/NB1 pixel_6305/VBIAS pixel_6305/NB2 pixel_6305/AMP_IN pixel_6305/SF_IB
+ pixel_6305/PIX_OUT pixel_6305/CSA_VREF pixel
Xpixel_6316 pixel_6316/gring pixel_6316/VDD pixel_6316/GND pixel_6316/VREF pixel_6316/ROW_SEL
+ pixel_6316/NB1 pixel_6316/VBIAS pixel_6316/NB2 pixel_6316/AMP_IN pixel_6316/SF_IB
+ pixel_6316/PIX_OUT pixel_6316/CSA_VREF pixel
Xpixel_6327 pixel_6327/gring pixel_6327/VDD pixel_6327/GND pixel_6327/VREF pixel_6327/ROW_SEL
+ pixel_6327/NB1 pixel_6327/VBIAS pixel_6327/NB2 pixel_6327/AMP_IN pixel_6327/SF_IB
+ pixel_6327/PIX_OUT pixel_6327/CSA_VREF pixel
Xpixel_6338 pixel_6338/gring pixel_6338/VDD pixel_6338/GND pixel_6338/VREF pixel_6338/ROW_SEL
+ pixel_6338/NB1 pixel_6338/VBIAS pixel_6338/NB2 pixel_6338/AMP_IN pixel_6338/SF_IB
+ pixel_6338/PIX_OUT pixel_6338/CSA_VREF pixel
Xpixel_6349 pixel_6349/gring pixel_6349/VDD pixel_6349/GND pixel_6349/VREF pixel_6349/ROW_SEL
+ pixel_6349/NB1 pixel_6349/VBIAS pixel_6349/NB2 pixel_6349/AMP_IN pixel_6349/SF_IB
+ pixel_6349/PIX_OUT pixel_6349/CSA_VREF pixel
Xpixel_5604 pixel_5604/gring pixel_5604/VDD pixel_5604/GND pixel_5604/VREF pixel_5604/ROW_SEL
+ pixel_5604/NB1 pixel_5604/VBIAS pixel_5604/NB2 pixel_5604/AMP_IN pixel_5604/SF_IB
+ pixel_5604/PIX_OUT pixel_5604/CSA_VREF pixel
Xpixel_5615 pixel_5615/gring pixel_5615/VDD pixel_5615/GND pixel_5615/VREF pixel_5615/ROW_SEL
+ pixel_5615/NB1 pixel_5615/VBIAS pixel_5615/NB2 pixel_5615/AMP_IN pixel_5615/SF_IB
+ pixel_5615/PIX_OUT pixel_5615/CSA_VREF pixel
Xpixel_5626 pixel_5626/gring pixel_5626/VDD pixel_5626/GND pixel_5626/VREF pixel_5626/ROW_SEL
+ pixel_5626/NB1 pixel_5626/VBIAS pixel_5626/NB2 pixel_5626/AMP_IN pixel_5626/SF_IB
+ pixel_5626/PIX_OUT pixel_5626/CSA_VREF pixel
Xpixel_5637 pixel_5637/gring pixel_5637/VDD pixel_5637/GND pixel_5637/VREF pixel_5637/ROW_SEL
+ pixel_5637/NB1 pixel_5637/VBIAS pixel_5637/NB2 pixel_5637/AMP_IN pixel_5637/SF_IB
+ pixel_5637/PIX_OUT pixel_5637/CSA_VREF pixel
Xpixel_5648 pixel_5648/gring pixel_5648/VDD pixel_5648/GND pixel_5648/VREF pixel_5648/ROW_SEL
+ pixel_5648/NB1 pixel_5648/VBIAS pixel_5648/NB2 pixel_5648/AMP_IN pixel_5648/SF_IB
+ pixel_5648/PIX_OUT pixel_5648/CSA_VREF pixel
Xpixel_4903 pixel_4903/gring pixel_4903/VDD pixel_4903/GND pixel_4903/VREF pixel_4903/ROW_SEL
+ pixel_4903/NB1 pixel_4903/VBIAS pixel_4903/NB2 pixel_4903/AMP_IN pixel_4903/SF_IB
+ pixel_4903/PIX_OUT pixel_4903/CSA_VREF pixel
Xpixel_942 pixel_942/gring pixel_942/VDD pixel_942/GND pixel_942/VREF pixel_942/ROW_SEL
+ pixel_942/NB1 pixel_942/VBIAS pixel_942/NB2 pixel_942/AMP_IN pixel_942/SF_IB pixel_942/PIX_OUT
+ pixel_942/CSA_VREF pixel
Xpixel_931 pixel_931/gring pixel_931/VDD pixel_931/GND pixel_931/VREF pixel_931/ROW_SEL
+ pixel_931/NB1 pixel_931/VBIAS pixel_931/NB2 pixel_931/AMP_IN pixel_931/SF_IB pixel_931/PIX_OUT
+ pixel_931/CSA_VREF pixel
Xpixel_920 pixel_920/gring pixel_920/VDD pixel_920/GND pixel_920/VREF pixel_920/ROW_SEL
+ pixel_920/NB1 pixel_920/VBIAS pixel_920/NB2 pixel_920/AMP_IN pixel_920/SF_IB pixel_920/PIX_OUT
+ pixel_920/CSA_VREF pixel
Xpixel_5659 pixel_5659/gring pixel_5659/VDD pixel_5659/GND pixel_5659/VREF pixel_5659/ROW_SEL
+ pixel_5659/NB1 pixel_5659/VBIAS pixel_5659/NB2 pixel_5659/AMP_IN pixel_5659/SF_IB
+ pixel_5659/PIX_OUT pixel_5659/CSA_VREF pixel
Xpixel_4914 pixel_4914/gring pixel_4914/VDD pixel_4914/GND pixel_4914/VREF pixel_4914/ROW_SEL
+ pixel_4914/NB1 pixel_4914/VBIAS pixel_4914/NB2 pixel_4914/AMP_IN pixel_4914/SF_IB
+ pixel_4914/PIX_OUT pixel_4914/CSA_VREF pixel
Xpixel_4925 pixel_4925/gring pixel_4925/VDD pixel_4925/GND pixel_4925/VREF pixel_4925/ROW_SEL
+ pixel_4925/NB1 pixel_4925/VBIAS pixel_4925/NB2 pixel_4925/AMP_IN pixel_4925/SF_IB
+ pixel_4925/PIX_OUT pixel_4925/CSA_VREF pixel
Xpixel_4936 pixel_4936/gring pixel_4936/VDD pixel_4936/GND pixel_4936/VREF pixel_4936/ROW_SEL
+ pixel_4936/NB1 pixel_4936/VBIAS pixel_4936/NB2 pixel_4936/AMP_IN pixel_4936/SF_IB
+ pixel_4936/PIX_OUT pixel_4936/CSA_VREF pixel
Xpixel_4947 pixel_4947/gring pixel_4947/VDD pixel_4947/GND pixel_4947/VREF pixel_4947/ROW_SEL
+ pixel_4947/NB1 pixel_4947/VBIAS pixel_4947/NB2 pixel_4947/AMP_IN pixel_4947/SF_IB
+ pixel_4947/PIX_OUT pixel_4947/CSA_VREF pixel
Xpixel_975 pixel_975/gring pixel_975/VDD pixel_975/GND pixel_975/VREF pixel_975/ROW_SEL
+ pixel_975/NB1 pixel_975/VBIAS pixel_975/NB2 pixel_975/AMP_IN pixel_975/SF_IB pixel_975/PIX_OUT
+ pixel_975/CSA_VREF pixel
Xpixel_964 pixel_964/gring pixel_964/VDD pixel_964/GND pixel_964/VREF pixel_964/ROW_SEL
+ pixel_964/NB1 pixel_964/VBIAS pixel_964/NB2 pixel_964/AMP_IN pixel_964/SF_IB pixel_964/PIX_OUT
+ pixel_964/CSA_VREF pixel
Xpixel_953 pixel_953/gring pixel_953/VDD pixel_953/GND pixel_953/VREF pixel_953/ROW_SEL
+ pixel_953/NB1 pixel_953/VBIAS pixel_953/NB2 pixel_953/AMP_IN pixel_953/SF_IB pixel_953/PIX_OUT
+ pixel_953/CSA_VREF pixel
Xpixel_4958 pixel_4958/gring pixel_4958/VDD pixel_4958/GND pixel_4958/VREF pixel_4958/ROW_SEL
+ pixel_4958/NB1 pixel_4958/VBIAS pixel_4958/NB2 pixel_4958/AMP_IN pixel_4958/SF_IB
+ pixel_4958/PIX_OUT pixel_4958/CSA_VREF pixel
Xpixel_4969 pixel_4969/gring pixel_4969/VDD pixel_4969/GND pixel_4969/VREF pixel_4969/ROW_SEL
+ pixel_4969/NB1 pixel_4969/VBIAS pixel_4969/NB2 pixel_4969/AMP_IN pixel_4969/SF_IB
+ pixel_4969/PIX_OUT pixel_4969/CSA_VREF pixel
Xpixel_997 pixel_997/gring pixel_997/VDD pixel_997/GND pixel_997/VREF pixel_997/ROW_SEL
+ pixel_997/NB1 pixel_997/VBIAS pixel_997/NB2 pixel_997/AMP_IN pixel_997/SF_IB pixel_997/PIX_OUT
+ pixel_997/CSA_VREF pixel
Xpixel_986 pixel_986/gring pixel_986/VDD pixel_986/GND pixel_986/VREF pixel_986/ROW_SEL
+ pixel_986/NB1 pixel_986/VBIAS pixel_986/NB2 pixel_986/AMP_IN pixel_986/SF_IB pixel_986/PIX_OUT
+ pixel_986/CSA_VREF pixel
Xpixel_8230 pixel_8230/gring pixel_8230/VDD pixel_8230/GND pixel_8230/VREF pixel_8230/ROW_SEL
+ pixel_8230/NB1 pixel_8230/VBIAS pixel_8230/NB2 pixel_8230/AMP_IN pixel_8230/SF_IB
+ pixel_8230/PIX_OUT pixel_8230/CSA_VREF pixel
Xpixel_8241 pixel_8241/gring pixel_8241/VDD pixel_8241/GND pixel_8241/VREF pixel_8241/ROW_SEL
+ pixel_8241/NB1 pixel_8241/VBIAS pixel_8241/NB2 pixel_8241/AMP_IN pixel_8241/SF_IB
+ pixel_8241/PIX_OUT pixel_8241/CSA_VREF pixel
Xpixel_8252 pixel_8252/gring pixel_8252/VDD pixel_8252/GND pixel_8252/VREF pixel_8252/ROW_SEL
+ pixel_8252/NB1 pixel_8252/VBIAS pixel_8252/NB2 pixel_8252/AMP_IN pixel_8252/SF_IB
+ pixel_8252/PIX_OUT pixel_8252/CSA_VREF pixel
Xpixel_8263 pixel_8263/gring pixel_8263/VDD pixel_8263/GND pixel_8263/VREF pixel_8263/ROW_SEL
+ pixel_8263/NB1 pixel_8263/VBIAS pixel_8263/NB2 pixel_8263/AMP_IN pixel_8263/SF_IB
+ pixel_8263/PIX_OUT pixel_8263/CSA_VREF pixel
Xpixel_8274 pixel_8274/gring pixel_8274/VDD pixel_8274/GND pixel_8274/VREF pixel_8274/ROW_SEL
+ pixel_8274/NB1 pixel_8274/VBIAS pixel_8274/NB2 pixel_8274/AMP_IN pixel_8274/SF_IB
+ pixel_8274/PIX_OUT pixel_8274/CSA_VREF pixel
Xpixel_8285 pixel_8285/gring pixel_8285/VDD pixel_8285/GND pixel_8285/VREF pixel_8285/ROW_SEL
+ pixel_8285/NB1 pixel_8285/VBIAS pixel_8285/NB2 pixel_8285/AMP_IN pixel_8285/SF_IB
+ pixel_8285/PIX_OUT pixel_8285/CSA_VREF pixel
Xpixel_7540 pixel_7540/gring pixel_7540/VDD pixel_7540/GND pixel_7540/VREF pixel_7540/ROW_SEL
+ pixel_7540/NB1 pixel_7540/VBIAS pixel_7540/NB2 pixel_7540/AMP_IN pixel_7540/SF_IB
+ pixel_7540/PIX_OUT pixel_7540/CSA_VREF pixel
Xpixel_7551 pixel_7551/gring pixel_7551/VDD pixel_7551/GND pixel_7551/VREF pixel_7551/ROW_SEL
+ pixel_7551/NB1 pixel_7551/VBIAS pixel_7551/NB2 pixel_7551/AMP_IN pixel_7551/SF_IB
+ pixel_7551/PIX_OUT pixel_7551/CSA_VREF pixel
Xpixel_8296 pixel_8296/gring pixel_8296/VDD pixel_8296/GND pixel_8296/VREF pixel_8296/ROW_SEL
+ pixel_8296/NB1 pixel_8296/VBIAS pixel_8296/NB2 pixel_8296/AMP_IN pixel_8296/SF_IB
+ pixel_8296/PIX_OUT pixel_8296/CSA_VREF pixel
Xpixel_7562 pixel_7562/gring pixel_7562/VDD pixel_7562/GND pixel_7562/VREF pixel_7562/ROW_SEL
+ pixel_7562/NB1 pixel_7562/VBIAS pixel_7562/NB2 pixel_7562/AMP_IN pixel_7562/SF_IB
+ pixel_7562/PIX_OUT pixel_7562/CSA_VREF pixel
Xpixel_7573 pixel_7573/gring pixel_7573/VDD pixel_7573/GND pixel_7573/VREF pixel_7573/ROW_SEL
+ pixel_7573/NB1 pixel_7573/VBIAS pixel_7573/NB2 pixel_7573/AMP_IN pixel_7573/SF_IB
+ pixel_7573/PIX_OUT pixel_7573/CSA_VREF pixel
Xpixel_7584 pixel_7584/gring pixel_7584/VDD pixel_7584/GND pixel_7584/VREF pixel_7584/ROW_SEL
+ pixel_7584/NB1 pixel_7584/VBIAS pixel_7584/NB2 pixel_7584/AMP_IN pixel_7584/SF_IB
+ pixel_7584/PIX_OUT pixel_7584/CSA_VREF pixel
Xpixel_7595 pixel_7595/gring pixel_7595/VDD pixel_7595/GND pixel_7595/VREF pixel_7595/ROW_SEL
+ pixel_7595/NB1 pixel_7595/VBIAS pixel_7595/NB2 pixel_7595/AMP_IN pixel_7595/SF_IB
+ pixel_7595/PIX_OUT pixel_7595/CSA_VREF pixel
Xpixel_6850 pixel_6850/gring pixel_6850/VDD pixel_6850/GND pixel_6850/VREF pixel_6850/ROW_SEL
+ pixel_6850/NB1 pixel_6850/VBIAS pixel_6850/NB2 pixel_6850/AMP_IN pixel_6850/SF_IB
+ pixel_6850/PIX_OUT pixel_6850/CSA_VREF pixel
Xpixel_6861 pixel_6861/gring pixel_6861/VDD pixel_6861/GND pixel_6861/VREF pixel_6861/ROW_SEL
+ pixel_6861/NB1 pixel_6861/VBIAS pixel_6861/NB2 pixel_6861/AMP_IN pixel_6861/SF_IB
+ pixel_6861/PIX_OUT pixel_6861/CSA_VREF pixel
Xpixel_6872 pixel_6872/gring pixel_6872/VDD pixel_6872/GND pixel_6872/VREF pixel_6872/ROW_SEL
+ pixel_6872/NB1 pixel_6872/VBIAS pixel_6872/NB2 pixel_6872/AMP_IN pixel_6872/SF_IB
+ pixel_6872/PIX_OUT pixel_6872/CSA_VREF pixel
Xpixel_6883 pixel_6883/gring pixel_6883/VDD pixel_6883/GND pixel_6883/VREF pixel_6883/ROW_SEL
+ pixel_6883/NB1 pixel_6883/VBIAS pixel_6883/NB2 pixel_6883/AMP_IN pixel_6883/SF_IB
+ pixel_6883/PIX_OUT pixel_6883/CSA_VREF pixel
Xpixel_6894 pixel_6894/gring pixel_6894/VDD pixel_6894/GND pixel_6894/VREF pixel_6894/ROW_SEL
+ pixel_6894/NB1 pixel_6894/VBIAS pixel_6894/NB2 pixel_6894/AMP_IN pixel_6894/SF_IB
+ pixel_6894/PIX_OUT pixel_6894/CSA_VREF pixel
Xpixel_1190 pixel_1190/gring pixel_1190/VDD pixel_1190/GND pixel_1190/VREF pixel_1190/ROW_SEL
+ pixel_1190/NB1 pixel_1190/VBIAS pixel_1190/NB2 pixel_1190/AMP_IN pixel_1190/SF_IB
+ pixel_1190/PIX_OUT pixel_1190/CSA_VREF pixel
Xpixel_238 pixel_238/gring pixel_238/VDD pixel_238/GND pixel_238/VREF pixel_238/ROW_SEL
+ pixel_238/NB1 pixel_238/VBIAS pixel_238/NB2 pixel_238/AMP_IN pixel_238/SF_IB pixel_238/PIX_OUT
+ pixel_238/CSA_VREF pixel
Xpixel_227 pixel_227/gring pixel_227/VDD pixel_227/GND pixel_227/VREF pixel_227/ROW_SEL
+ pixel_227/NB1 pixel_227/VBIAS pixel_227/NB2 pixel_227/AMP_IN pixel_227/SF_IB pixel_227/PIX_OUT
+ pixel_227/CSA_VREF pixel
Xpixel_216 pixel_216/gring pixel_216/VDD pixel_216/GND pixel_216/VREF pixel_216/ROW_SEL
+ pixel_216/NB1 pixel_216/VBIAS pixel_216/NB2 pixel_216/AMP_IN pixel_216/SF_IB pixel_216/PIX_OUT
+ pixel_216/CSA_VREF pixel
Xpixel_205 pixel_205/gring pixel_205/VDD pixel_205/GND pixel_205/VREF pixel_205/ROW_SEL
+ pixel_205/NB1 pixel_205/VBIAS pixel_205/NB2 pixel_205/AMP_IN pixel_205/SF_IB pixel_205/PIX_OUT
+ pixel_205/CSA_VREF pixel
Xpixel_249 pixel_249/gring pixel_249/VDD pixel_249/GND pixel_249/VREF pixel_249/ROW_SEL
+ pixel_249/NB1 pixel_249/VBIAS pixel_249/NB2 pixel_249/AMP_IN pixel_249/SF_IB pixel_249/PIX_OUT
+ pixel_249/CSA_VREF pixel
Xpixel_3509 pixel_3509/gring pixel_3509/VDD pixel_3509/GND pixel_3509/VREF pixel_3509/ROW_SEL
+ pixel_3509/NB1 pixel_3509/VBIAS pixel_3509/NB2 pixel_3509/AMP_IN pixel_3509/SF_IB
+ pixel_3509/PIX_OUT pixel_3509/CSA_VREF pixel
Xpixel_2819 pixel_2819/gring pixel_2819/VDD pixel_2819/GND pixel_2819/VREF pixel_2819/ROW_SEL
+ pixel_2819/NB1 pixel_2819/VBIAS pixel_2819/NB2 pixel_2819/AMP_IN pixel_2819/SF_IB
+ pixel_2819/PIX_OUT pixel_2819/CSA_VREF pixel
Xpixel_2808 pixel_2808/gring pixel_2808/VDD pixel_2808/GND pixel_2808/VREF pixel_2808/ROW_SEL
+ pixel_2808/NB1 pixel_2808/VBIAS pixel_2808/NB2 pixel_2808/AMP_IN pixel_2808/SF_IB
+ pixel_2808/PIX_OUT pixel_2808/CSA_VREF pixel
Xpixel_6102 pixel_6102/gring pixel_6102/VDD pixel_6102/GND pixel_6102/VREF pixel_6102/ROW_SEL
+ pixel_6102/NB1 pixel_6102/VBIAS pixel_6102/NB2 pixel_6102/AMP_IN pixel_6102/SF_IB
+ pixel_6102/PIX_OUT pixel_6102/CSA_VREF pixel
Xpixel_6113 pixel_6113/gring pixel_6113/VDD pixel_6113/GND pixel_6113/VREF pixel_6113/ROW_SEL
+ pixel_6113/NB1 pixel_6113/VBIAS pixel_6113/NB2 pixel_6113/AMP_IN pixel_6113/SF_IB
+ pixel_6113/PIX_OUT pixel_6113/CSA_VREF pixel
Xpixel_6124 pixel_6124/gring pixel_6124/VDD pixel_6124/GND pixel_6124/VREF pixel_6124/ROW_SEL
+ pixel_6124/NB1 pixel_6124/VBIAS pixel_6124/NB2 pixel_6124/AMP_IN pixel_6124/SF_IB
+ pixel_6124/PIX_OUT pixel_6124/CSA_VREF pixel
Xpixel_6135 pixel_6135/gring pixel_6135/VDD pixel_6135/GND pixel_6135/VREF pixel_6135/ROW_SEL
+ pixel_6135/NB1 pixel_6135/VBIAS pixel_6135/NB2 pixel_6135/AMP_IN pixel_6135/SF_IB
+ pixel_6135/PIX_OUT pixel_6135/CSA_VREF pixel
Xpixel_6146 pixel_6146/gring pixel_6146/VDD pixel_6146/GND pixel_6146/VREF pixel_6146/ROW_SEL
+ pixel_6146/NB1 pixel_6146/VBIAS pixel_6146/NB2 pixel_6146/AMP_IN pixel_6146/SF_IB
+ pixel_6146/PIX_OUT pixel_6146/CSA_VREF pixel
Xpixel_6157 pixel_6157/gring pixel_6157/VDD pixel_6157/GND pixel_6157/VREF pixel_6157/ROW_SEL
+ pixel_6157/NB1 pixel_6157/VBIAS pixel_6157/NB2 pixel_6157/AMP_IN pixel_6157/SF_IB
+ pixel_6157/PIX_OUT pixel_6157/CSA_VREF pixel
Xpixel_6168 pixel_6168/gring pixel_6168/VDD pixel_6168/GND pixel_6168/VREF pixel_6168/ROW_SEL
+ pixel_6168/NB1 pixel_6168/VBIAS pixel_6168/NB2 pixel_6168/AMP_IN pixel_6168/SF_IB
+ pixel_6168/PIX_OUT pixel_6168/CSA_VREF pixel
Xpixel_5401 pixel_5401/gring pixel_5401/VDD pixel_5401/GND pixel_5401/VREF pixel_5401/ROW_SEL
+ pixel_5401/NB1 pixel_5401/VBIAS pixel_5401/NB2 pixel_5401/AMP_IN pixel_5401/SF_IB
+ pixel_5401/PIX_OUT pixel_5401/CSA_VREF pixel
Xpixel_5412 pixel_5412/gring pixel_5412/VDD pixel_5412/GND pixel_5412/VREF pixel_5412/ROW_SEL
+ pixel_5412/NB1 pixel_5412/VBIAS pixel_5412/NB2 pixel_5412/AMP_IN pixel_5412/SF_IB
+ pixel_5412/PIX_OUT pixel_5412/CSA_VREF pixel
Xpixel_5423 pixel_5423/gring pixel_5423/VDD pixel_5423/GND pixel_5423/VREF pixel_5423/ROW_SEL
+ pixel_5423/NB1 pixel_5423/VBIAS pixel_5423/NB2 pixel_5423/AMP_IN pixel_5423/SF_IB
+ pixel_5423/PIX_OUT pixel_5423/CSA_VREF pixel
Xpixel_6179 pixel_6179/gring pixel_6179/VDD pixel_6179/GND pixel_6179/VREF pixel_6179/ROW_SEL
+ pixel_6179/NB1 pixel_6179/VBIAS pixel_6179/NB2 pixel_6179/AMP_IN pixel_6179/SF_IB
+ pixel_6179/PIX_OUT pixel_6179/CSA_VREF pixel
Xpixel_5434 pixel_5434/gring pixel_5434/VDD pixel_5434/GND pixel_5434/VREF pixel_5434/ROW_SEL
+ pixel_5434/NB1 pixel_5434/VBIAS pixel_5434/NB2 pixel_5434/AMP_IN pixel_5434/SF_IB
+ pixel_5434/PIX_OUT pixel_5434/CSA_VREF pixel
Xpixel_5445 pixel_5445/gring pixel_5445/VDD pixel_5445/GND pixel_5445/VREF pixel_5445/ROW_SEL
+ pixel_5445/NB1 pixel_5445/VBIAS pixel_5445/NB2 pixel_5445/AMP_IN pixel_5445/SF_IB
+ pixel_5445/PIX_OUT pixel_5445/CSA_VREF pixel
Xpixel_5456 pixel_5456/gring pixel_5456/VDD pixel_5456/GND pixel_5456/VREF pixel_5456/ROW_SEL
+ pixel_5456/NB1 pixel_5456/VBIAS pixel_5456/NB2 pixel_5456/AMP_IN pixel_5456/SF_IB
+ pixel_5456/PIX_OUT pixel_5456/CSA_VREF pixel
Xpixel_4700 pixel_4700/gring pixel_4700/VDD pixel_4700/GND pixel_4700/VREF pixel_4700/ROW_SEL
+ pixel_4700/NB1 pixel_4700/VBIAS pixel_4700/NB2 pixel_4700/AMP_IN pixel_4700/SF_IB
+ pixel_4700/PIX_OUT pixel_4700/CSA_VREF pixel
Xpixel_4711 pixel_4711/gring pixel_4711/VDD pixel_4711/GND pixel_4711/VREF pixel_4711/ROW_SEL
+ pixel_4711/NB1 pixel_4711/VBIAS pixel_4711/NB2 pixel_4711/AMP_IN pixel_4711/SF_IB
+ pixel_4711/PIX_OUT pixel_4711/CSA_VREF pixel
Xpixel_4722 pixel_4722/gring pixel_4722/VDD pixel_4722/GND pixel_4722/VREF pixel_4722/ROW_SEL
+ pixel_4722/NB1 pixel_4722/VBIAS pixel_4722/NB2 pixel_4722/AMP_IN pixel_4722/SF_IB
+ pixel_4722/PIX_OUT pixel_4722/CSA_VREF pixel
Xpixel_750 pixel_750/gring pixel_750/VDD pixel_750/GND pixel_750/VREF pixel_750/ROW_SEL
+ pixel_750/NB1 pixel_750/VBIAS pixel_750/NB2 pixel_750/AMP_IN pixel_750/SF_IB pixel_750/PIX_OUT
+ pixel_750/CSA_VREF pixel
Xpixel_5467 pixel_5467/gring pixel_5467/VDD pixel_5467/GND pixel_5467/VREF pixel_5467/ROW_SEL
+ pixel_5467/NB1 pixel_5467/VBIAS pixel_5467/NB2 pixel_5467/AMP_IN pixel_5467/SF_IB
+ pixel_5467/PIX_OUT pixel_5467/CSA_VREF pixel
Xpixel_5478 pixel_5478/gring pixel_5478/VDD pixel_5478/GND pixel_5478/VREF pixel_5478/ROW_SEL
+ pixel_5478/NB1 pixel_5478/VBIAS pixel_5478/NB2 pixel_5478/AMP_IN pixel_5478/SF_IB
+ pixel_5478/PIX_OUT pixel_5478/CSA_VREF pixel
Xpixel_5489 pixel_5489/gring pixel_5489/VDD pixel_5489/GND pixel_5489/VREF pixel_5489/ROW_SEL
+ pixel_5489/NB1 pixel_5489/VBIAS pixel_5489/NB2 pixel_5489/AMP_IN pixel_5489/SF_IB
+ pixel_5489/PIX_OUT pixel_5489/CSA_VREF pixel
Xpixel_4733 pixel_4733/gring pixel_4733/VDD pixel_4733/GND pixel_4733/VREF pixel_4733/ROW_SEL
+ pixel_4733/NB1 pixel_4733/VBIAS pixel_4733/NB2 pixel_4733/AMP_IN pixel_4733/SF_IB
+ pixel_4733/PIX_OUT pixel_4733/CSA_VREF pixel
Xpixel_4744 pixel_4744/gring pixel_4744/VDD pixel_4744/GND pixel_4744/VREF pixel_4744/ROW_SEL
+ pixel_4744/NB1 pixel_4744/VBIAS pixel_4744/NB2 pixel_4744/AMP_IN pixel_4744/SF_IB
+ pixel_4744/PIX_OUT pixel_4744/CSA_VREF pixel
Xpixel_4755 pixel_4755/gring pixel_4755/VDD pixel_4755/GND pixel_4755/VREF pixel_4755/ROW_SEL
+ pixel_4755/NB1 pixel_4755/VBIAS pixel_4755/NB2 pixel_4755/AMP_IN pixel_4755/SF_IB
+ pixel_4755/PIX_OUT pixel_4755/CSA_VREF pixel
Xpixel_783 pixel_783/gring pixel_783/VDD pixel_783/GND pixel_783/VREF pixel_783/ROW_SEL
+ pixel_783/NB1 pixel_783/VBIAS pixel_783/NB2 pixel_783/AMP_IN pixel_783/SF_IB pixel_783/PIX_OUT
+ pixel_783/CSA_VREF pixel
Xpixel_772 pixel_772/gring pixel_772/VDD pixel_772/GND pixel_772/VREF pixel_772/ROW_SEL
+ pixel_772/NB1 pixel_772/VBIAS pixel_772/NB2 pixel_772/AMP_IN pixel_772/SF_IB pixel_772/PIX_OUT
+ pixel_772/CSA_VREF pixel
Xpixel_761 pixel_761/gring pixel_761/VDD pixel_761/GND pixel_761/VREF pixel_761/ROW_SEL
+ pixel_761/NB1 pixel_761/VBIAS pixel_761/NB2 pixel_761/AMP_IN pixel_761/SF_IB pixel_761/PIX_OUT
+ pixel_761/CSA_VREF pixel
Xpixel_4766 pixel_4766/gring pixel_4766/VDD pixel_4766/GND pixel_4766/VREF pixel_4766/ROW_SEL
+ pixel_4766/NB1 pixel_4766/VBIAS pixel_4766/NB2 pixel_4766/AMP_IN pixel_4766/SF_IB
+ pixel_4766/PIX_OUT pixel_4766/CSA_VREF pixel
Xpixel_4777 pixel_4777/gring pixel_4777/VDD pixel_4777/GND pixel_4777/VREF pixel_4777/ROW_SEL
+ pixel_4777/NB1 pixel_4777/VBIAS pixel_4777/NB2 pixel_4777/AMP_IN pixel_4777/SF_IB
+ pixel_4777/PIX_OUT pixel_4777/CSA_VREF pixel
Xpixel_4788 pixel_4788/gring pixel_4788/VDD pixel_4788/GND pixel_4788/VREF pixel_4788/ROW_SEL
+ pixel_4788/NB1 pixel_4788/VBIAS pixel_4788/NB2 pixel_4788/AMP_IN pixel_4788/SF_IB
+ pixel_4788/PIX_OUT pixel_4788/CSA_VREF pixel
Xpixel_794 pixel_794/gring pixel_794/VDD pixel_794/GND pixel_794/VREF pixel_794/ROW_SEL
+ pixel_794/NB1 pixel_794/VBIAS pixel_794/NB2 pixel_794/AMP_IN pixel_794/SF_IB pixel_794/PIX_OUT
+ pixel_794/CSA_VREF pixel
Xpixel_4799 pixel_4799/gring pixel_4799/VDD pixel_4799/GND pixel_4799/VREF pixel_4799/ROW_SEL
+ pixel_4799/NB1 pixel_4799/VBIAS pixel_4799/NB2 pixel_4799/AMP_IN pixel_4799/SF_IB
+ pixel_4799/PIX_OUT pixel_4799/CSA_VREF pixel
Xpixel_8060 pixel_8060/gring pixel_8060/VDD pixel_8060/GND pixel_8060/VREF pixel_8060/ROW_SEL
+ pixel_8060/NB1 pixel_8060/VBIAS pixel_8060/NB2 pixel_8060/AMP_IN pixel_8060/SF_IB
+ pixel_8060/PIX_OUT pixel_8060/CSA_VREF pixel
Xpixel_8071 pixel_8071/gring pixel_8071/VDD pixel_8071/GND pixel_8071/VREF pixel_8071/ROW_SEL
+ pixel_8071/NB1 pixel_8071/VBIAS pixel_8071/NB2 pixel_8071/AMP_IN pixel_8071/SF_IB
+ pixel_8071/PIX_OUT pixel_8071/CSA_VREF pixel
Xpixel_8082 pixel_8082/gring pixel_8082/VDD pixel_8082/GND pixel_8082/VREF pixel_8082/ROW_SEL
+ pixel_8082/NB1 pixel_8082/VBIAS pixel_8082/NB2 pixel_8082/AMP_IN pixel_8082/SF_IB
+ pixel_8082/PIX_OUT pixel_8082/CSA_VREF pixel
Xpixel_8093 pixel_8093/gring pixel_8093/VDD pixel_8093/GND pixel_8093/VREF pixel_8093/ROW_SEL
+ pixel_8093/NB1 pixel_8093/VBIAS pixel_8093/NB2 pixel_8093/AMP_IN pixel_8093/SF_IB
+ pixel_8093/PIX_OUT pixel_8093/CSA_VREF pixel
Xpixel_7370 pixel_7370/gring pixel_7370/VDD pixel_7370/GND pixel_7370/VREF pixel_7370/ROW_SEL
+ pixel_7370/NB1 pixel_7370/VBIAS pixel_7370/NB2 pixel_7370/AMP_IN pixel_7370/SF_IB
+ pixel_7370/PIX_OUT pixel_7370/CSA_VREF pixel
Xpixel_7381 pixel_7381/gring pixel_7381/VDD pixel_7381/GND pixel_7381/VREF pixel_7381/ROW_SEL
+ pixel_7381/NB1 pixel_7381/VBIAS pixel_7381/NB2 pixel_7381/AMP_IN pixel_7381/SF_IB
+ pixel_7381/PIX_OUT pixel_7381/CSA_VREF pixel
Xpixel_7392 pixel_7392/gring pixel_7392/VDD pixel_7392/GND pixel_7392/VREF pixel_7392/ROW_SEL
+ pixel_7392/NB1 pixel_7392/VBIAS pixel_7392/NB2 pixel_7392/AMP_IN pixel_7392/SF_IB
+ pixel_7392/PIX_OUT pixel_7392/CSA_VREF pixel
Xpixel_6680 pixel_6680/gring pixel_6680/VDD pixel_6680/GND pixel_6680/VREF pixel_6680/ROW_SEL
+ pixel_6680/NB1 pixel_6680/VBIAS pixel_6680/NB2 pixel_6680/AMP_IN pixel_6680/SF_IB
+ pixel_6680/PIX_OUT pixel_6680/CSA_VREF pixel
Xpixel_6691 pixel_6691/gring pixel_6691/VDD pixel_6691/GND pixel_6691/VREF pixel_6691/ROW_SEL
+ pixel_6691/NB1 pixel_6691/VBIAS pixel_6691/NB2 pixel_6691/AMP_IN pixel_6691/SF_IB
+ pixel_6691/PIX_OUT pixel_6691/CSA_VREF pixel
Xpixel_5990 pixel_5990/gring pixel_5990/VDD pixel_5990/GND pixel_5990/VREF pixel_5990/ROW_SEL
+ pixel_5990/NB1 pixel_5990/VBIAS pixel_5990/NB2 pixel_5990/AMP_IN pixel_5990/SF_IB
+ pixel_5990/PIX_OUT pixel_5990/CSA_VREF pixel
Xpixel_4007 pixel_4007/gring pixel_4007/VDD pixel_4007/GND pixel_4007/VREF pixel_4007/ROW_SEL
+ pixel_4007/NB1 pixel_4007/VBIAS pixel_4007/NB2 pixel_4007/AMP_IN pixel_4007/SF_IB
+ pixel_4007/PIX_OUT pixel_4007/CSA_VREF pixel
Xpixel_3306 pixel_3306/gring pixel_3306/VDD pixel_3306/GND pixel_3306/VREF pixel_3306/ROW_SEL
+ pixel_3306/NB1 pixel_3306/VBIAS pixel_3306/NB2 pixel_3306/AMP_IN pixel_3306/SF_IB
+ pixel_3306/PIX_OUT pixel_3306/CSA_VREF pixel
Xpixel_4018 pixel_4018/gring pixel_4018/VDD pixel_4018/GND pixel_4018/VREF pixel_4018/ROW_SEL
+ pixel_4018/NB1 pixel_4018/VBIAS pixel_4018/NB2 pixel_4018/AMP_IN pixel_4018/SF_IB
+ pixel_4018/PIX_OUT pixel_4018/CSA_VREF pixel
Xpixel_4029 pixel_4029/gring pixel_4029/VDD pixel_4029/GND pixel_4029/VREF pixel_4029/ROW_SEL
+ pixel_4029/NB1 pixel_4029/VBIAS pixel_4029/NB2 pixel_4029/AMP_IN pixel_4029/SF_IB
+ pixel_4029/PIX_OUT pixel_4029/CSA_VREF pixel
Xpixel_3339 pixel_3339/gring pixel_3339/VDD pixel_3339/GND pixel_3339/VREF pixel_3339/ROW_SEL
+ pixel_3339/NB1 pixel_3339/VBIAS pixel_3339/NB2 pixel_3339/AMP_IN pixel_3339/SF_IB
+ pixel_3339/PIX_OUT pixel_3339/CSA_VREF pixel
Xpixel_3328 pixel_3328/gring pixel_3328/VDD pixel_3328/GND pixel_3328/VREF pixel_3328/ROW_SEL
+ pixel_3328/NB1 pixel_3328/VBIAS pixel_3328/NB2 pixel_3328/AMP_IN pixel_3328/SF_IB
+ pixel_3328/PIX_OUT pixel_3328/CSA_VREF pixel
Xpixel_3317 pixel_3317/gring pixel_3317/VDD pixel_3317/GND pixel_3317/VREF pixel_3317/ROW_SEL
+ pixel_3317/NB1 pixel_3317/VBIAS pixel_3317/NB2 pixel_3317/AMP_IN pixel_3317/SF_IB
+ pixel_3317/PIX_OUT pixel_3317/CSA_VREF pixel
Xpixel_2627 pixel_2627/gring pixel_2627/VDD pixel_2627/GND pixel_2627/VREF pixel_2627/ROW_SEL
+ pixel_2627/NB1 pixel_2627/VBIAS pixel_2627/NB2 pixel_2627/AMP_IN pixel_2627/SF_IB
+ pixel_2627/PIX_OUT pixel_2627/CSA_VREF pixel
Xpixel_2616 pixel_2616/gring pixel_2616/VDD pixel_2616/GND pixel_2616/VREF pixel_2616/ROW_SEL
+ pixel_2616/NB1 pixel_2616/VBIAS pixel_2616/NB2 pixel_2616/AMP_IN pixel_2616/SF_IB
+ pixel_2616/PIX_OUT pixel_2616/CSA_VREF pixel
Xpixel_2605 pixel_2605/gring pixel_2605/VDD pixel_2605/GND pixel_2605/VREF pixel_2605/ROW_SEL
+ pixel_2605/NB1 pixel_2605/VBIAS pixel_2605/NB2 pixel_2605/AMP_IN pixel_2605/SF_IB
+ pixel_2605/PIX_OUT pixel_2605/CSA_VREF pixel
Xpixel_1926 pixel_1926/gring pixel_1926/VDD pixel_1926/GND pixel_1926/VREF pixel_1926/ROW_SEL
+ pixel_1926/NB1 pixel_1926/VBIAS pixel_1926/NB2 pixel_1926/AMP_IN pixel_1926/SF_IB
+ pixel_1926/PIX_OUT pixel_1926/CSA_VREF pixel
Xpixel_1915 pixel_1915/gring pixel_1915/VDD pixel_1915/GND pixel_1915/VREF pixel_1915/ROW_SEL
+ pixel_1915/NB1 pixel_1915/VBIAS pixel_1915/NB2 pixel_1915/AMP_IN pixel_1915/SF_IB
+ pixel_1915/PIX_OUT pixel_1915/CSA_VREF pixel
Xpixel_1904 pixel_1904/gring pixel_1904/VDD pixel_1904/GND pixel_1904/VREF pixel_1904/ROW_SEL
+ pixel_1904/NB1 pixel_1904/VBIAS pixel_1904/NB2 pixel_1904/AMP_IN pixel_1904/SF_IB
+ pixel_1904/PIX_OUT pixel_1904/CSA_VREF pixel
Xpixel_2649 pixel_2649/gring pixel_2649/VDD pixel_2649/GND pixel_2649/VREF pixel_2649/ROW_SEL
+ pixel_2649/NB1 pixel_2649/VBIAS pixel_2649/NB2 pixel_2649/AMP_IN pixel_2649/SF_IB
+ pixel_2649/PIX_OUT pixel_2649/CSA_VREF pixel
Xpixel_2638 pixel_2638/gring pixel_2638/VDD pixel_2638/GND pixel_2638/VREF pixel_2638/ROW_SEL
+ pixel_2638/NB1 pixel_2638/VBIAS pixel_2638/NB2 pixel_2638/AMP_IN pixel_2638/SF_IB
+ pixel_2638/PIX_OUT pixel_2638/CSA_VREF pixel
Xpixel_1959 pixel_1959/gring pixel_1959/VDD pixel_1959/GND pixel_1959/VREF pixel_1959/ROW_SEL
+ pixel_1959/NB1 pixel_1959/VBIAS pixel_1959/NB2 pixel_1959/AMP_IN pixel_1959/SF_IB
+ pixel_1959/PIX_OUT pixel_1959/CSA_VREF pixel
Xpixel_1948 pixel_1948/gring pixel_1948/VDD pixel_1948/GND pixel_1948/VREF pixel_1948/ROW_SEL
+ pixel_1948/NB1 pixel_1948/VBIAS pixel_1948/NB2 pixel_1948/AMP_IN pixel_1948/SF_IB
+ pixel_1948/PIX_OUT pixel_1948/CSA_VREF pixel
Xpixel_1937 pixel_1937/gring pixel_1937/VDD pixel_1937/GND pixel_1937/VREF pixel_1937/ROW_SEL
+ pixel_1937/NB1 pixel_1937/VBIAS pixel_1937/NB2 pixel_1937/AMP_IN pixel_1937/SF_IB
+ pixel_1937/PIX_OUT pixel_1937/CSA_VREF pixel
Xpixel_5220 pixel_5220/gring pixel_5220/VDD pixel_5220/GND pixel_5220/VREF pixel_5220/ROW_SEL
+ pixel_5220/NB1 pixel_5220/VBIAS pixel_5220/NB2 pixel_5220/AMP_IN pixel_5220/SF_IB
+ pixel_5220/PIX_OUT pixel_5220/CSA_VREF pixel
Xpixel_5231 pixel_5231/gring pixel_5231/VDD pixel_5231/GND pixel_5231/VREF pixel_5231/ROW_SEL
+ pixel_5231/NB1 pixel_5231/VBIAS pixel_5231/NB2 pixel_5231/AMP_IN pixel_5231/SF_IB
+ pixel_5231/PIX_OUT pixel_5231/CSA_VREF pixel
Xpixel_5242 pixel_5242/gring pixel_5242/VDD pixel_5242/GND pixel_5242/VREF pixel_5242/ROW_SEL
+ pixel_5242/NB1 pixel_5242/VBIAS pixel_5242/NB2 pixel_5242/AMP_IN pixel_5242/SF_IB
+ pixel_5242/PIX_OUT pixel_5242/CSA_VREF pixel
Xpixel_5253 pixel_5253/gring pixel_5253/VDD pixel_5253/GND pixel_5253/VREF pixel_5253/ROW_SEL
+ pixel_5253/NB1 pixel_5253/VBIAS pixel_5253/NB2 pixel_5253/AMP_IN pixel_5253/SF_IB
+ pixel_5253/PIX_OUT pixel_5253/CSA_VREF pixel
Xpixel_5264 pixel_5264/gring pixel_5264/VDD pixel_5264/GND pixel_5264/VREF pixel_5264/ROW_SEL
+ pixel_5264/NB1 pixel_5264/VBIAS pixel_5264/NB2 pixel_5264/AMP_IN pixel_5264/SF_IB
+ pixel_5264/PIX_OUT pixel_5264/CSA_VREF pixel
Xpixel_5275 pixel_5275/gring pixel_5275/VDD pixel_5275/GND pixel_5275/VREF pixel_5275/ROW_SEL
+ pixel_5275/NB1 pixel_5275/VBIAS pixel_5275/NB2 pixel_5275/AMP_IN pixel_5275/SF_IB
+ pixel_5275/PIX_OUT pixel_5275/CSA_VREF pixel
Xpixel_4530 pixel_4530/gring pixel_4530/VDD pixel_4530/GND pixel_4530/VREF pixel_4530/ROW_SEL
+ pixel_4530/NB1 pixel_4530/VBIAS pixel_4530/NB2 pixel_4530/AMP_IN pixel_4530/SF_IB
+ pixel_4530/PIX_OUT pixel_4530/CSA_VREF pixel
Xpixel_5286 pixel_5286/gring pixel_5286/VDD pixel_5286/GND pixel_5286/VREF pixel_5286/ROW_SEL
+ pixel_5286/NB1 pixel_5286/VBIAS pixel_5286/NB2 pixel_5286/AMP_IN pixel_5286/SF_IB
+ pixel_5286/PIX_OUT pixel_5286/CSA_VREF pixel
Xpixel_5297 pixel_5297/gring pixel_5297/VDD pixel_5297/GND pixel_5297/VREF pixel_5297/ROW_SEL
+ pixel_5297/NB1 pixel_5297/VBIAS pixel_5297/NB2 pixel_5297/AMP_IN pixel_5297/SF_IB
+ pixel_5297/PIX_OUT pixel_5297/CSA_VREF pixel
Xpixel_4541 pixel_4541/gring pixel_4541/VDD pixel_4541/GND pixel_4541/VREF pixel_4541/ROW_SEL
+ pixel_4541/NB1 pixel_4541/VBIAS pixel_4541/NB2 pixel_4541/AMP_IN pixel_4541/SF_IB
+ pixel_4541/PIX_OUT pixel_4541/CSA_VREF pixel
Xpixel_4552 pixel_4552/gring pixel_4552/VDD pixel_4552/GND pixel_4552/VREF pixel_4552/ROW_SEL
+ pixel_4552/NB1 pixel_4552/VBIAS pixel_4552/NB2 pixel_4552/AMP_IN pixel_4552/SF_IB
+ pixel_4552/PIX_OUT pixel_4552/CSA_VREF pixel
Xpixel_4563 pixel_4563/gring pixel_4563/VDD pixel_4563/GND pixel_4563/VREF pixel_4563/ROW_SEL
+ pixel_4563/NB1 pixel_4563/VBIAS pixel_4563/NB2 pixel_4563/AMP_IN pixel_4563/SF_IB
+ pixel_4563/PIX_OUT pixel_4563/CSA_VREF pixel
Xpixel_591 pixel_591/gring pixel_591/VDD pixel_591/GND pixel_591/VREF pixel_591/ROW_SEL
+ pixel_591/NB1 pixel_591/VBIAS pixel_591/NB2 pixel_591/AMP_IN pixel_591/SF_IB pixel_591/PIX_OUT
+ pixel_591/CSA_VREF pixel
Xpixel_580 pixel_580/gring pixel_580/VDD pixel_580/GND pixel_580/VREF pixel_580/ROW_SEL
+ pixel_580/NB1 pixel_580/VBIAS pixel_580/NB2 pixel_580/AMP_IN pixel_580/SF_IB pixel_580/PIX_OUT
+ pixel_580/CSA_VREF pixel
Xpixel_3862 pixel_3862/gring pixel_3862/VDD pixel_3862/GND pixel_3862/VREF pixel_3862/ROW_SEL
+ pixel_3862/NB1 pixel_3862/VBIAS pixel_3862/NB2 pixel_3862/AMP_IN pixel_3862/SF_IB
+ pixel_3862/PIX_OUT pixel_3862/CSA_VREF pixel
Xpixel_3851 pixel_3851/gring pixel_3851/VDD pixel_3851/GND pixel_3851/VREF pixel_3851/ROW_SEL
+ pixel_3851/NB1 pixel_3851/VBIAS pixel_3851/NB2 pixel_3851/AMP_IN pixel_3851/SF_IB
+ pixel_3851/PIX_OUT pixel_3851/CSA_VREF pixel
Xpixel_4574 pixel_4574/gring pixel_4574/VDD pixel_4574/GND pixel_4574/VREF pixel_4574/ROW_SEL
+ pixel_4574/NB1 pixel_4574/VBIAS pixel_4574/NB2 pixel_4574/AMP_IN pixel_4574/SF_IB
+ pixel_4574/PIX_OUT pixel_4574/CSA_VREF pixel
Xpixel_4585 pixel_4585/gring pixel_4585/VDD pixel_4585/GND pixel_4585/VREF pixel_4585/ROW_SEL
+ pixel_4585/NB1 pixel_4585/VBIAS pixel_4585/NB2 pixel_4585/AMP_IN pixel_4585/SF_IB
+ pixel_4585/PIX_OUT pixel_4585/CSA_VREF pixel
Xpixel_4596 pixel_4596/gring pixel_4596/VDD pixel_4596/GND pixel_4596/VREF pixel_4596/ROW_SEL
+ pixel_4596/NB1 pixel_4596/VBIAS pixel_4596/NB2 pixel_4596/AMP_IN pixel_4596/SF_IB
+ pixel_4596/PIX_OUT pixel_4596/CSA_VREF pixel
Xpixel_3840 pixel_3840/gring pixel_3840/VDD pixel_3840/GND pixel_3840/VREF pixel_3840/ROW_SEL
+ pixel_3840/NB1 pixel_3840/VBIAS pixel_3840/NB2 pixel_3840/AMP_IN pixel_3840/SF_IB
+ pixel_3840/PIX_OUT pixel_3840/CSA_VREF pixel
Xpixel_3895 pixel_3895/gring pixel_3895/VDD pixel_3895/GND pixel_3895/VREF pixel_3895/ROW_SEL
+ pixel_3895/NB1 pixel_3895/VBIAS pixel_3895/NB2 pixel_3895/AMP_IN pixel_3895/SF_IB
+ pixel_3895/PIX_OUT pixel_3895/CSA_VREF pixel
Xpixel_3884 pixel_3884/gring pixel_3884/VDD pixel_3884/GND pixel_3884/VREF pixel_3884/ROW_SEL
+ pixel_3884/NB1 pixel_3884/VBIAS pixel_3884/NB2 pixel_3884/AMP_IN pixel_3884/SF_IB
+ pixel_3884/PIX_OUT pixel_3884/CSA_VREF pixel
Xpixel_3873 pixel_3873/gring pixel_3873/VDD pixel_3873/GND pixel_3873/VREF pixel_3873/ROW_SEL
+ pixel_3873/NB1 pixel_3873/VBIAS pixel_3873/NB2 pixel_3873/AMP_IN pixel_3873/SF_IB
+ pixel_3873/PIX_OUT pixel_3873/CSA_VREF pixel
Xpixel_9519 pixel_9519/gring pixel_9519/VDD pixel_9519/GND pixel_9519/VREF pixel_9519/ROW_SEL
+ pixel_9519/NB1 pixel_9519/VBIAS pixel_9519/NB2 pixel_9519/AMP_IN pixel_9519/SF_IB
+ pixel_9519/PIX_OUT pixel_9519/CSA_VREF pixel
Xpixel_9508 pixel_9508/gring pixel_9508/VDD pixel_9508/GND pixel_9508/VREF pixel_9508/ROW_SEL
+ pixel_9508/NB1 pixel_9508/VBIAS pixel_9508/NB2 pixel_9508/AMP_IN pixel_9508/SF_IB
+ pixel_9508/PIX_OUT pixel_9508/CSA_VREF pixel
Xpixel_8818 pixel_8818/gring pixel_8818/VDD pixel_8818/GND pixel_8818/VREF pixel_8818/ROW_SEL
+ pixel_8818/NB1 pixel_8818/VBIAS pixel_8818/NB2 pixel_8818/AMP_IN pixel_8818/SF_IB
+ pixel_8818/PIX_OUT pixel_8818/CSA_VREF pixel
Xpixel_8807 pixel_8807/gring pixel_8807/VDD pixel_8807/GND pixel_8807/VREF pixel_8807/ROW_SEL
+ pixel_8807/NB1 pixel_8807/VBIAS pixel_8807/NB2 pixel_8807/AMP_IN pixel_8807/SF_IB
+ pixel_8807/PIX_OUT pixel_8807/CSA_VREF pixel
Xpixel_8829 pixel_8829/gring pixel_8829/VDD pixel_8829/GND pixel_8829/VREF pixel_8829/ROW_SEL
+ pixel_8829/NB1 pixel_8829/VBIAS pixel_8829/NB2 pixel_8829/AMP_IN pixel_8829/SF_IB
+ pixel_8829/PIX_OUT pixel_8829/CSA_VREF pixel
Xpixel_3114 pixel_3114/gring pixel_3114/VDD pixel_3114/GND pixel_3114/VREF pixel_3114/ROW_SEL
+ pixel_3114/NB1 pixel_3114/VBIAS pixel_3114/NB2 pixel_3114/AMP_IN pixel_3114/SF_IB
+ pixel_3114/PIX_OUT pixel_3114/CSA_VREF pixel
Xpixel_3103 pixel_3103/gring pixel_3103/VDD pixel_3103/GND pixel_3103/VREF pixel_3103/ROW_SEL
+ pixel_3103/NB1 pixel_3103/VBIAS pixel_3103/NB2 pixel_3103/AMP_IN pixel_3103/SF_IB
+ pixel_3103/PIX_OUT pixel_3103/CSA_VREF pixel
Xpixel_2402 pixel_2402/gring pixel_2402/VDD pixel_2402/GND pixel_2402/VREF pixel_2402/ROW_SEL
+ pixel_2402/NB1 pixel_2402/VBIAS pixel_2402/NB2 pixel_2402/AMP_IN pixel_2402/SF_IB
+ pixel_2402/PIX_OUT pixel_2402/CSA_VREF pixel
Xpixel_3147 pixel_3147/gring pixel_3147/VDD pixel_3147/GND pixel_3147/VREF pixel_3147/ROW_SEL
+ pixel_3147/NB1 pixel_3147/VBIAS pixel_3147/NB2 pixel_3147/AMP_IN pixel_3147/SF_IB
+ pixel_3147/PIX_OUT pixel_3147/CSA_VREF pixel
Xpixel_3136 pixel_3136/gring pixel_3136/VDD pixel_3136/GND pixel_3136/VREF pixel_3136/ROW_SEL
+ pixel_3136/NB1 pixel_3136/VBIAS pixel_3136/NB2 pixel_3136/AMP_IN pixel_3136/SF_IB
+ pixel_3136/PIX_OUT pixel_3136/CSA_VREF pixel
Xpixel_3125 pixel_3125/gring pixel_3125/VDD pixel_3125/GND pixel_3125/VREF pixel_3125/ROW_SEL
+ pixel_3125/NB1 pixel_3125/VBIAS pixel_3125/NB2 pixel_3125/AMP_IN pixel_3125/SF_IB
+ pixel_3125/PIX_OUT pixel_3125/CSA_VREF pixel
Xpixel_1701 pixel_1701/gring pixel_1701/VDD pixel_1701/GND pixel_1701/VREF pixel_1701/ROW_SEL
+ pixel_1701/NB1 pixel_1701/VBIAS pixel_1701/NB2 pixel_1701/AMP_IN pixel_1701/SF_IB
+ pixel_1701/PIX_OUT pixel_1701/CSA_VREF pixel
Xpixel_2446 pixel_2446/gring pixel_2446/VDD pixel_2446/GND pixel_2446/VREF pixel_2446/ROW_SEL
+ pixel_2446/NB1 pixel_2446/VBIAS pixel_2446/NB2 pixel_2446/AMP_IN pixel_2446/SF_IB
+ pixel_2446/PIX_OUT pixel_2446/CSA_VREF pixel
Xpixel_2435 pixel_2435/gring pixel_2435/VDD pixel_2435/GND pixel_2435/VREF pixel_2435/ROW_SEL
+ pixel_2435/NB1 pixel_2435/VBIAS pixel_2435/NB2 pixel_2435/AMP_IN pixel_2435/SF_IB
+ pixel_2435/PIX_OUT pixel_2435/CSA_VREF pixel
Xpixel_2424 pixel_2424/gring pixel_2424/VDD pixel_2424/GND pixel_2424/VREF pixel_2424/ROW_SEL
+ pixel_2424/NB1 pixel_2424/VBIAS pixel_2424/NB2 pixel_2424/AMP_IN pixel_2424/SF_IB
+ pixel_2424/PIX_OUT pixel_2424/CSA_VREF pixel
Xpixel_2413 pixel_2413/gring pixel_2413/VDD pixel_2413/GND pixel_2413/VREF pixel_2413/ROW_SEL
+ pixel_2413/NB1 pixel_2413/VBIAS pixel_2413/NB2 pixel_2413/AMP_IN pixel_2413/SF_IB
+ pixel_2413/PIX_OUT pixel_2413/CSA_VREF pixel
Xpixel_3169 pixel_3169/gring pixel_3169/VDD pixel_3169/GND pixel_3169/VREF pixel_3169/ROW_SEL
+ pixel_3169/NB1 pixel_3169/VBIAS pixel_3169/NB2 pixel_3169/AMP_IN pixel_3169/SF_IB
+ pixel_3169/PIX_OUT pixel_3169/CSA_VREF pixel
Xpixel_3158 pixel_3158/gring pixel_3158/VDD pixel_3158/GND pixel_3158/VREF pixel_3158/ROW_SEL
+ pixel_3158/NB1 pixel_3158/VBIAS pixel_3158/NB2 pixel_3158/AMP_IN pixel_3158/SF_IB
+ pixel_3158/PIX_OUT pixel_3158/CSA_VREF pixel
Xpixel_1734 pixel_1734/gring pixel_1734/VDD pixel_1734/GND pixel_1734/VREF pixel_1734/ROW_SEL
+ pixel_1734/NB1 pixel_1734/VBIAS pixel_1734/NB2 pixel_1734/AMP_IN pixel_1734/SF_IB
+ pixel_1734/PIX_OUT pixel_1734/CSA_VREF pixel
Xpixel_1723 pixel_1723/gring pixel_1723/VDD pixel_1723/GND pixel_1723/VREF pixel_1723/ROW_SEL
+ pixel_1723/NB1 pixel_1723/VBIAS pixel_1723/NB2 pixel_1723/AMP_IN pixel_1723/SF_IB
+ pixel_1723/PIX_OUT pixel_1723/CSA_VREF pixel
Xpixel_1712 pixel_1712/gring pixel_1712/VDD pixel_1712/GND pixel_1712/VREF pixel_1712/ROW_SEL
+ pixel_1712/NB1 pixel_1712/VBIAS pixel_1712/NB2 pixel_1712/AMP_IN pixel_1712/SF_IB
+ pixel_1712/PIX_OUT pixel_1712/CSA_VREF pixel
Xpixel_2479 pixel_2479/gring pixel_2479/VDD pixel_2479/GND pixel_2479/VREF pixel_2479/ROW_SEL
+ pixel_2479/NB1 pixel_2479/VBIAS pixel_2479/NB2 pixel_2479/AMP_IN pixel_2479/SF_IB
+ pixel_2479/PIX_OUT pixel_2479/CSA_VREF pixel
Xpixel_2468 pixel_2468/gring pixel_2468/VDD pixel_2468/GND pixel_2468/VREF pixel_2468/ROW_SEL
+ pixel_2468/NB1 pixel_2468/VBIAS pixel_2468/NB2 pixel_2468/AMP_IN pixel_2468/SF_IB
+ pixel_2468/PIX_OUT pixel_2468/CSA_VREF pixel
Xpixel_2457 pixel_2457/gring pixel_2457/VDD pixel_2457/GND pixel_2457/VREF pixel_2457/ROW_SEL
+ pixel_2457/NB1 pixel_2457/VBIAS pixel_2457/NB2 pixel_2457/AMP_IN pixel_2457/SF_IB
+ pixel_2457/PIX_OUT pixel_2457/CSA_VREF pixel
Xpixel_1767 pixel_1767/gring pixel_1767/VDD pixel_1767/GND pixel_1767/VREF pixel_1767/ROW_SEL
+ pixel_1767/NB1 pixel_1767/VBIAS pixel_1767/NB2 pixel_1767/AMP_IN pixel_1767/SF_IB
+ pixel_1767/PIX_OUT pixel_1767/CSA_VREF pixel
Xpixel_1756 pixel_1756/gring pixel_1756/VDD pixel_1756/GND pixel_1756/VREF pixel_1756/ROW_SEL
+ pixel_1756/NB1 pixel_1756/VBIAS pixel_1756/NB2 pixel_1756/AMP_IN pixel_1756/SF_IB
+ pixel_1756/PIX_OUT pixel_1756/CSA_VREF pixel
Xpixel_1745 pixel_1745/gring pixel_1745/VDD pixel_1745/GND pixel_1745/VREF pixel_1745/ROW_SEL
+ pixel_1745/NB1 pixel_1745/VBIAS pixel_1745/NB2 pixel_1745/AMP_IN pixel_1745/SF_IB
+ pixel_1745/PIX_OUT pixel_1745/CSA_VREF pixel
Xpixel_1789 pixel_1789/gring pixel_1789/VDD pixel_1789/GND pixel_1789/VREF pixel_1789/ROW_SEL
+ pixel_1789/NB1 pixel_1789/VBIAS pixel_1789/NB2 pixel_1789/AMP_IN pixel_1789/SF_IB
+ pixel_1789/PIX_OUT pixel_1789/CSA_VREF pixel
Xpixel_1778 pixel_1778/gring pixel_1778/VDD pixel_1778/GND pixel_1778/VREF pixel_1778/ROW_SEL
+ pixel_1778/NB1 pixel_1778/VBIAS pixel_1778/NB2 pixel_1778/AMP_IN pixel_1778/SF_IB
+ pixel_1778/PIX_OUT pixel_1778/CSA_VREF pixel
Xpixel_5050 pixel_5050/gring pixel_5050/VDD pixel_5050/GND pixel_5050/VREF pixel_5050/ROW_SEL
+ pixel_5050/NB1 pixel_5050/VBIAS pixel_5050/NB2 pixel_5050/AMP_IN pixel_5050/SF_IB
+ pixel_5050/PIX_OUT pixel_5050/CSA_VREF pixel
Xpixel_5061 pixel_5061/gring pixel_5061/VDD pixel_5061/GND pixel_5061/VREF pixel_5061/ROW_SEL
+ pixel_5061/NB1 pixel_5061/VBIAS pixel_5061/NB2 pixel_5061/AMP_IN pixel_5061/SF_IB
+ pixel_5061/PIX_OUT pixel_5061/CSA_VREF pixel
Xpixel_5072 pixel_5072/gring pixel_5072/VDD pixel_5072/GND pixel_5072/VREF pixel_5072/ROW_SEL
+ pixel_5072/NB1 pixel_5072/VBIAS pixel_5072/NB2 pixel_5072/AMP_IN pixel_5072/SF_IB
+ pixel_5072/PIX_OUT pixel_5072/CSA_VREF pixel
Xpixel_5083 pixel_5083/gring pixel_5083/VDD pixel_5083/GND pixel_5083/VREF pixel_5083/ROW_SEL
+ pixel_5083/NB1 pixel_5083/VBIAS pixel_5083/NB2 pixel_5083/AMP_IN pixel_5083/SF_IB
+ pixel_5083/PIX_OUT pixel_5083/CSA_VREF pixel
Xpixel_5094 pixel_5094/gring pixel_5094/VDD pixel_5094/GND pixel_5094/VREF pixel_5094/ROW_SEL
+ pixel_5094/NB1 pixel_5094/VBIAS pixel_5094/NB2 pixel_5094/AMP_IN pixel_5094/SF_IB
+ pixel_5094/PIX_OUT pixel_5094/CSA_VREF pixel
Xpixel_4360 pixel_4360/gring pixel_4360/VDD pixel_4360/GND pixel_4360/VREF pixel_4360/ROW_SEL
+ pixel_4360/NB1 pixel_4360/VBIAS pixel_4360/NB2 pixel_4360/AMP_IN pixel_4360/SF_IB
+ pixel_4360/PIX_OUT pixel_4360/CSA_VREF pixel
Xpixel_4371 pixel_4371/gring pixel_4371/VDD pixel_4371/GND pixel_4371/VREF pixel_4371/ROW_SEL
+ pixel_4371/NB1 pixel_4371/VBIAS pixel_4371/NB2 pixel_4371/AMP_IN pixel_4371/SF_IB
+ pixel_4371/PIX_OUT pixel_4371/CSA_VREF pixel
Xpixel_3670 pixel_3670/gring pixel_3670/VDD pixel_3670/GND pixel_3670/VREF pixel_3670/ROW_SEL
+ pixel_3670/NB1 pixel_3670/VBIAS pixel_3670/NB2 pixel_3670/AMP_IN pixel_3670/SF_IB
+ pixel_3670/PIX_OUT pixel_3670/CSA_VREF pixel
Xpixel_4382 pixel_4382/gring pixel_4382/VDD pixel_4382/GND pixel_4382/VREF pixel_4382/ROW_SEL
+ pixel_4382/NB1 pixel_4382/VBIAS pixel_4382/NB2 pixel_4382/AMP_IN pixel_4382/SF_IB
+ pixel_4382/PIX_OUT pixel_4382/CSA_VREF pixel
Xpixel_4393 pixel_4393/gring pixel_4393/VDD pixel_4393/GND pixel_4393/VREF pixel_4393/ROW_SEL
+ pixel_4393/NB1 pixel_4393/VBIAS pixel_4393/NB2 pixel_4393/AMP_IN pixel_4393/SF_IB
+ pixel_4393/PIX_OUT pixel_4393/CSA_VREF pixel
Xpixel_3692 pixel_3692/gring pixel_3692/VDD pixel_3692/GND pixel_3692/VREF pixel_3692/ROW_SEL
+ pixel_3692/NB1 pixel_3692/VBIAS pixel_3692/NB2 pixel_3692/AMP_IN pixel_3692/SF_IB
+ pixel_3692/PIX_OUT pixel_3692/CSA_VREF pixel
Xpixel_3681 pixel_3681/gring pixel_3681/VDD pixel_3681/GND pixel_3681/VREF pixel_3681/ROW_SEL
+ pixel_3681/NB1 pixel_3681/VBIAS pixel_3681/NB2 pixel_3681/AMP_IN pixel_3681/SF_IB
+ pixel_3681/PIX_OUT pixel_3681/CSA_VREF pixel
Xpixel_2991 pixel_2991/gring pixel_2991/VDD pixel_2991/GND pixel_2991/VREF pixel_2991/ROW_SEL
+ pixel_2991/NB1 pixel_2991/VBIAS pixel_2991/NB2 pixel_2991/AMP_IN pixel_2991/SF_IB
+ pixel_2991/PIX_OUT pixel_2991/CSA_VREF pixel
Xpixel_2980 pixel_2980/gring pixel_2980/VDD pixel_2980/GND pixel_2980/VREF pixel_2980/ROW_SEL
+ pixel_2980/NB1 pixel_2980/VBIAS pixel_2980/NB2 pixel_2980/AMP_IN pixel_2980/SF_IB
+ pixel_2980/PIX_OUT pixel_2980/CSA_VREF pixel
Xpixel_1019 pixel_1019/gring pixel_1019/VDD pixel_1019/GND pixel_1019/VREF pixel_1019/ROW_SEL
+ pixel_1019/NB1 pixel_1019/VBIAS pixel_1019/NB2 pixel_1019/AMP_IN pixel_1019/SF_IB
+ pixel_1019/PIX_OUT pixel_1019/CSA_VREF pixel
Xpixel_1008 pixel_1008/gring pixel_1008/VDD pixel_1008/GND pixel_1008/VREF pixel_1008/ROW_SEL
+ pixel_1008/NB1 pixel_1008/VBIAS pixel_1008/NB2 pixel_1008/AMP_IN pixel_1008/SF_IB
+ pixel_1008/PIX_OUT pixel_1008/CSA_VREF pixel
Xpixel_9338 pixel_9338/gring pixel_9338/VDD pixel_9338/GND pixel_9338/VREF pixel_9338/ROW_SEL
+ pixel_9338/NB1 pixel_9338/VBIAS pixel_9338/NB2 pixel_9338/AMP_IN pixel_9338/SF_IB
+ pixel_9338/PIX_OUT pixel_9338/CSA_VREF pixel
Xpixel_9327 pixel_9327/gring pixel_9327/VDD pixel_9327/GND pixel_9327/VREF pixel_9327/ROW_SEL
+ pixel_9327/NB1 pixel_9327/VBIAS pixel_9327/NB2 pixel_9327/AMP_IN pixel_9327/SF_IB
+ pixel_9327/PIX_OUT pixel_9327/CSA_VREF pixel
Xpixel_9316 pixel_9316/gring pixel_9316/VDD pixel_9316/GND pixel_9316/VREF pixel_9316/ROW_SEL
+ pixel_9316/NB1 pixel_9316/VBIAS pixel_9316/NB2 pixel_9316/AMP_IN pixel_9316/SF_IB
+ pixel_9316/PIX_OUT pixel_9316/CSA_VREF pixel
Xpixel_9305 pixel_9305/gring pixel_9305/VDD pixel_9305/GND pixel_9305/VREF pixel_9305/ROW_SEL
+ pixel_9305/NB1 pixel_9305/VBIAS pixel_9305/NB2 pixel_9305/AMP_IN pixel_9305/SF_IB
+ pixel_9305/PIX_OUT pixel_9305/CSA_VREF pixel
Xpixel_8626 pixel_8626/gring pixel_8626/VDD pixel_8626/GND pixel_8626/VREF pixel_8626/ROW_SEL
+ pixel_8626/NB1 pixel_8626/VBIAS pixel_8626/NB2 pixel_8626/AMP_IN pixel_8626/SF_IB
+ pixel_8626/PIX_OUT pixel_8626/CSA_VREF pixel
Xpixel_8615 pixel_8615/gring pixel_8615/VDD pixel_8615/GND pixel_8615/VREF pixel_8615/ROW_SEL
+ pixel_8615/NB1 pixel_8615/VBIAS pixel_8615/NB2 pixel_8615/AMP_IN pixel_8615/SF_IB
+ pixel_8615/PIX_OUT pixel_8615/CSA_VREF pixel
Xpixel_8604 pixel_8604/gring pixel_8604/VDD pixel_8604/GND pixel_8604/VREF pixel_8604/ROW_SEL
+ pixel_8604/NB1 pixel_8604/VBIAS pixel_8604/NB2 pixel_8604/AMP_IN pixel_8604/SF_IB
+ pixel_8604/PIX_OUT pixel_8604/CSA_VREF pixel
Xpixel_9349 pixel_9349/gring pixel_9349/VDD pixel_9349/GND pixel_9349/VREF pixel_9349/ROW_SEL
+ pixel_9349/NB1 pixel_9349/VBIAS pixel_9349/NB2 pixel_9349/AMP_IN pixel_9349/SF_IB
+ pixel_9349/PIX_OUT pixel_9349/CSA_VREF pixel
Xpixel_8659 pixel_8659/gring pixel_8659/VDD pixel_8659/GND pixel_8659/VREF pixel_8659/ROW_SEL
+ pixel_8659/NB1 pixel_8659/VBIAS pixel_8659/NB2 pixel_8659/AMP_IN pixel_8659/SF_IB
+ pixel_8659/PIX_OUT pixel_8659/CSA_VREF pixel
Xpixel_8648 pixel_8648/gring pixel_8648/VDD pixel_8648/GND pixel_8648/VREF pixel_8648/ROW_SEL
+ pixel_8648/NB1 pixel_8648/VBIAS pixel_8648/NB2 pixel_8648/AMP_IN pixel_8648/SF_IB
+ pixel_8648/PIX_OUT pixel_8648/CSA_VREF pixel
Xpixel_8637 pixel_8637/gring pixel_8637/VDD pixel_8637/GND pixel_8637/VREF pixel_8637/ROW_SEL
+ pixel_8637/NB1 pixel_8637/VBIAS pixel_8637/NB2 pixel_8637/AMP_IN pixel_8637/SF_IB
+ pixel_8637/PIX_OUT pixel_8637/CSA_VREF pixel
Xpixel_7903 pixel_7903/gring pixel_7903/VDD pixel_7903/GND pixel_7903/VREF pixel_7903/ROW_SEL
+ pixel_7903/NB1 pixel_7903/VBIAS pixel_7903/NB2 pixel_7903/AMP_IN pixel_7903/SF_IB
+ pixel_7903/PIX_OUT pixel_7903/CSA_VREF pixel
Xpixel_7914 pixel_7914/gring pixel_7914/VDD pixel_7914/GND pixel_7914/VREF pixel_7914/ROW_SEL
+ pixel_7914/NB1 pixel_7914/VBIAS pixel_7914/NB2 pixel_7914/AMP_IN pixel_7914/SF_IB
+ pixel_7914/PIX_OUT pixel_7914/CSA_VREF pixel
Xpixel_7925 pixel_7925/gring pixel_7925/VDD pixel_7925/GND pixel_7925/VREF pixel_7925/ROW_SEL
+ pixel_7925/NB1 pixel_7925/VBIAS pixel_7925/NB2 pixel_7925/AMP_IN pixel_7925/SF_IB
+ pixel_7925/PIX_OUT pixel_7925/CSA_VREF pixel
Xpixel_7936 pixel_7936/gring pixel_7936/VDD pixel_7936/GND pixel_7936/VREF pixel_7936/ROW_SEL
+ pixel_7936/NB1 pixel_7936/VBIAS pixel_7936/NB2 pixel_7936/AMP_IN pixel_7936/SF_IB
+ pixel_7936/PIX_OUT pixel_7936/CSA_VREF pixel
Xpixel_7947 pixel_7947/gring pixel_7947/VDD pixel_7947/GND pixel_7947/VREF pixel_7947/ROW_SEL
+ pixel_7947/NB1 pixel_7947/VBIAS pixel_7947/NB2 pixel_7947/AMP_IN pixel_7947/SF_IB
+ pixel_7947/PIX_OUT pixel_7947/CSA_VREF pixel
Xpixel_7958 pixel_7958/gring pixel_7958/VDD pixel_7958/GND pixel_7958/VREF pixel_7958/ROW_SEL
+ pixel_7958/NB1 pixel_7958/VBIAS pixel_7958/NB2 pixel_7958/AMP_IN pixel_7958/SF_IB
+ pixel_7958/PIX_OUT pixel_7958/CSA_VREF pixel
Xpixel_7969 pixel_7969/gring pixel_7969/VDD pixel_7969/GND pixel_7969/VREF pixel_7969/ROW_SEL
+ pixel_7969/NB1 pixel_7969/VBIAS pixel_7969/NB2 pixel_7969/AMP_IN pixel_7969/SF_IB
+ pixel_7969/PIX_OUT pixel_7969/CSA_VREF pixel
Xpixel_2221 pixel_2221/gring pixel_2221/VDD pixel_2221/GND pixel_2221/VREF pixel_2221/ROW_SEL
+ pixel_2221/NB1 pixel_2221/VBIAS pixel_2221/NB2 pixel_2221/AMP_IN pixel_2221/SF_IB
+ pixel_2221/PIX_OUT pixel_2221/CSA_VREF pixel
Xpixel_2210 pixel_2210/gring pixel_2210/VDD pixel_2210/GND pixel_2210/VREF pixel_2210/ROW_SEL
+ pixel_2210/NB1 pixel_2210/VBIAS pixel_2210/NB2 pixel_2210/AMP_IN pixel_2210/SF_IB
+ pixel_2210/PIX_OUT pixel_2210/CSA_VREF pixel
Xpixel_2254 pixel_2254/gring pixel_2254/VDD pixel_2254/GND pixel_2254/VREF pixel_2254/ROW_SEL
+ pixel_2254/NB1 pixel_2254/VBIAS pixel_2254/NB2 pixel_2254/AMP_IN pixel_2254/SF_IB
+ pixel_2254/PIX_OUT pixel_2254/CSA_VREF pixel
Xpixel_2243 pixel_2243/gring pixel_2243/VDD pixel_2243/GND pixel_2243/VREF pixel_2243/ROW_SEL
+ pixel_2243/NB1 pixel_2243/VBIAS pixel_2243/NB2 pixel_2243/AMP_IN pixel_2243/SF_IB
+ pixel_2243/PIX_OUT pixel_2243/CSA_VREF pixel
Xpixel_2232 pixel_2232/gring pixel_2232/VDD pixel_2232/GND pixel_2232/VREF pixel_2232/ROW_SEL
+ pixel_2232/NB1 pixel_2232/VBIAS pixel_2232/NB2 pixel_2232/AMP_IN pixel_2232/SF_IB
+ pixel_2232/PIX_OUT pixel_2232/CSA_VREF pixel
Xpixel_1542 pixel_1542/gring pixel_1542/VDD pixel_1542/GND pixel_1542/VREF pixel_1542/ROW_SEL
+ pixel_1542/NB1 pixel_1542/VBIAS pixel_1542/NB2 pixel_1542/AMP_IN pixel_1542/SF_IB
+ pixel_1542/PIX_OUT pixel_1542/CSA_VREF pixel
Xpixel_1531 pixel_1531/gring pixel_1531/VDD pixel_1531/GND pixel_1531/VREF pixel_1531/ROW_SEL
+ pixel_1531/NB1 pixel_1531/VBIAS pixel_1531/NB2 pixel_1531/AMP_IN pixel_1531/SF_IB
+ pixel_1531/PIX_OUT pixel_1531/CSA_VREF pixel
Xpixel_1520 pixel_1520/gring pixel_1520/VDD pixel_1520/GND pixel_1520/VREF pixel_1520/ROW_SEL
+ pixel_1520/NB1 pixel_1520/VBIAS pixel_1520/NB2 pixel_1520/AMP_IN pixel_1520/SF_IB
+ pixel_1520/PIX_OUT pixel_1520/CSA_VREF pixel
Xpixel_2287 pixel_2287/gring pixel_2287/VDD pixel_2287/GND pixel_2287/VREF pixel_2287/ROW_SEL
+ pixel_2287/NB1 pixel_2287/VBIAS pixel_2287/NB2 pixel_2287/AMP_IN pixel_2287/SF_IB
+ pixel_2287/PIX_OUT pixel_2287/CSA_VREF pixel
Xpixel_2276 pixel_2276/gring pixel_2276/VDD pixel_2276/GND pixel_2276/VREF pixel_2276/ROW_SEL
+ pixel_2276/NB1 pixel_2276/VBIAS pixel_2276/NB2 pixel_2276/AMP_IN pixel_2276/SF_IB
+ pixel_2276/PIX_OUT pixel_2276/CSA_VREF pixel
Xpixel_2265 pixel_2265/gring pixel_2265/VDD pixel_2265/GND pixel_2265/VREF pixel_2265/ROW_SEL
+ pixel_2265/NB1 pixel_2265/VBIAS pixel_2265/NB2 pixel_2265/AMP_IN pixel_2265/SF_IB
+ pixel_2265/PIX_OUT pixel_2265/CSA_VREF pixel
Xpixel_1586 pixel_1586/gring pixel_1586/VDD pixel_1586/GND pixel_1586/VREF pixel_1586/ROW_SEL
+ pixel_1586/NB1 pixel_1586/VBIAS pixel_1586/NB2 pixel_1586/AMP_IN pixel_1586/SF_IB
+ pixel_1586/PIX_OUT pixel_1586/CSA_VREF pixel
Xpixel_1575 pixel_1575/gring pixel_1575/VDD pixel_1575/GND pixel_1575/VREF pixel_1575/ROW_SEL
+ pixel_1575/NB1 pixel_1575/VBIAS pixel_1575/NB2 pixel_1575/AMP_IN pixel_1575/SF_IB
+ pixel_1575/PIX_OUT pixel_1575/CSA_VREF pixel
Xpixel_1564 pixel_1564/gring pixel_1564/VDD pixel_1564/GND pixel_1564/VREF pixel_1564/ROW_SEL
+ pixel_1564/NB1 pixel_1564/VBIAS pixel_1564/NB2 pixel_1564/AMP_IN pixel_1564/SF_IB
+ pixel_1564/PIX_OUT pixel_1564/CSA_VREF pixel
Xpixel_1553 pixel_1553/gring pixel_1553/VDD pixel_1553/GND pixel_1553/VREF pixel_1553/ROW_SEL
+ pixel_1553/NB1 pixel_1553/VBIAS pixel_1553/NB2 pixel_1553/AMP_IN pixel_1553/SF_IB
+ pixel_1553/PIX_OUT pixel_1553/CSA_VREF pixel
Xpixel_2298 pixel_2298/gring pixel_2298/VDD pixel_2298/GND pixel_2298/VREF pixel_2298/ROW_SEL
+ pixel_2298/NB1 pixel_2298/VBIAS pixel_2298/NB2 pixel_2298/AMP_IN pixel_2298/SF_IB
+ pixel_2298/PIX_OUT pixel_2298/CSA_VREF pixel
Xpixel_1597 pixel_1597/gring pixel_1597/VDD pixel_1597/GND pixel_1597/VREF pixel_1597/ROW_SEL
+ pixel_1597/NB1 pixel_1597/VBIAS pixel_1597/NB2 pixel_1597/AMP_IN pixel_1597/SF_IB
+ pixel_1597/PIX_OUT pixel_1597/CSA_VREF pixel
Xpixel_9850 pixel_9850/gring pixel_9850/VDD pixel_9850/GND pixel_9850/VREF pixel_9850/ROW_SEL
+ pixel_9850/NB1 pixel_9850/VBIAS pixel_9850/NB2 pixel_9850/AMP_IN pixel_9850/SF_IB
+ pixel_9850/PIX_OUT pixel_9850/CSA_VREF pixel
Xpixel_9861 pixel_9861/gring pixel_9861/VDD pixel_9861/GND pixel_9861/VREF pixel_9861/ROW_SEL
+ pixel_9861/NB1 pixel_9861/VBIAS pixel_9861/NB2 pixel_9861/AMP_IN pixel_9861/SF_IB
+ pixel_9861/PIX_OUT pixel_9861/CSA_VREF pixel
Xpixel_9872 pixel_9872/gring pixel_9872/VDD pixel_9872/GND pixel_9872/VREF pixel_9872/ROW_SEL
+ pixel_9872/NB1 pixel_9872/VBIAS pixel_9872/NB2 pixel_9872/AMP_IN pixel_9872/SF_IB
+ pixel_9872/PIX_OUT pixel_9872/CSA_VREF pixel
Xpixel_9883 pixel_9883/gring pixel_9883/VDD pixel_9883/GND pixel_9883/VREF pixel_9883/ROW_SEL
+ pixel_9883/NB1 pixel_9883/VBIAS pixel_9883/NB2 pixel_9883/AMP_IN pixel_9883/SF_IB
+ pixel_9883/PIX_OUT pixel_9883/CSA_VREF pixel
Xpixel_9894 pixel_9894/gring pixel_9894/VDD pixel_9894/GND pixel_9894/VREF pixel_9894/ROW_SEL
+ pixel_9894/NB1 pixel_9894/VBIAS pixel_9894/NB2 pixel_9894/AMP_IN pixel_9894/SF_IB
+ pixel_9894/PIX_OUT pixel_9894/CSA_VREF pixel
Xpixel_4190 pixel_4190/gring pixel_4190/VDD pixel_4190/GND pixel_4190/VREF pixel_4190/ROW_SEL
+ pixel_4190/NB1 pixel_4190/VBIAS pixel_4190/NB2 pixel_4190/AMP_IN pixel_4190/SF_IB
+ pixel_4190/PIX_OUT pixel_4190/CSA_VREF pixel
Xpixel_6509 pixel_6509/gring pixel_6509/VDD pixel_6509/GND pixel_6509/VREF pixel_6509/ROW_SEL
+ pixel_6509/NB1 pixel_6509/VBIAS pixel_6509/NB2 pixel_6509/AMP_IN pixel_6509/SF_IB
+ pixel_6509/PIX_OUT pixel_6509/CSA_VREF pixel
Xpixel_5808 pixel_5808/gring pixel_5808/VDD pixel_5808/GND pixel_5808/VREF pixel_5808/ROW_SEL
+ pixel_5808/NB1 pixel_5808/VBIAS pixel_5808/NB2 pixel_5808/AMP_IN pixel_5808/SF_IB
+ pixel_5808/PIX_OUT pixel_5808/CSA_VREF pixel
Xpixel_5819 pixel_5819/gring pixel_5819/VDD pixel_5819/GND pixel_5819/VREF pixel_5819/ROW_SEL
+ pixel_5819/NB1 pixel_5819/VBIAS pixel_5819/NB2 pixel_5819/AMP_IN pixel_5819/SF_IB
+ pixel_5819/PIX_OUT pixel_5819/CSA_VREF pixel
Xpixel_9113 pixel_9113/gring pixel_9113/VDD pixel_9113/GND pixel_9113/VREF pixel_9113/ROW_SEL
+ pixel_9113/NB1 pixel_9113/VBIAS pixel_9113/NB2 pixel_9113/AMP_IN pixel_9113/SF_IB
+ pixel_9113/PIX_OUT pixel_9113/CSA_VREF pixel
Xpixel_9102 pixel_9102/gring pixel_9102/VDD pixel_9102/GND pixel_9102/VREF pixel_9102/ROW_SEL
+ pixel_9102/NB1 pixel_9102/VBIAS pixel_9102/NB2 pixel_9102/AMP_IN pixel_9102/SF_IB
+ pixel_9102/PIX_OUT pixel_9102/CSA_VREF pixel
Xpixel_8401 pixel_8401/gring pixel_8401/VDD pixel_8401/GND pixel_8401/VREF pixel_8401/ROW_SEL
+ pixel_8401/NB1 pixel_8401/VBIAS pixel_8401/NB2 pixel_8401/AMP_IN pixel_8401/SF_IB
+ pixel_8401/PIX_OUT pixel_8401/CSA_VREF pixel
Xpixel_9146 pixel_9146/gring pixel_9146/VDD pixel_9146/GND pixel_9146/VREF pixel_9146/ROW_SEL
+ pixel_9146/NB1 pixel_9146/VBIAS pixel_9146/NB2 pixel_9146/AMP_IN pixel_9146/SF_IB
+ pixel_9146/PIX_OUT pixel_9146/CSA_VREF pixel
Xpixel_9135 pixel_9135/gring pixel_9135/VDD pixel_9135/GND pixel_9135/VREF pixel_9135/ROW_SEL
+ pixel_9135/NB1 pixel_9135/VBIAS pixel_9135/NB2 pixel_9135/AMP_IN pixel_9135/SF_IB
+ pixel_9135/PIX_OUT pixel_9135/CSA_VREF pixel
Xpixel_9124 pixel_9124/gring pixel_9124/VDD pixel_9124/GND pixel_9124/VREF pixel_9124/ROW_SEL
+ pixel_9124/NB1 pixel_9124/VBIAS pixel_9124/NB2 pixel_9124/AMP_IN pixel_9124/SF_IB
+ pixel_9124/PIX_OUT pixel_9124/CSA_VREF pixel
Xpixel_8434 pixel_8434/gring pixel_8434/VDD pixel_8434/GND pixel_8434/VREF pixel_8434/ROW_SEL
+ pixel_8434/NB1 pixel_8434/VBIAS pixel_8434/NB2 pixel_8434/AMP_IN pixel_8434/SF_IB
+ pixel_8434/PIX_OUT pixel_8434/CSA_VREF pixel
Xpixel_8423 pixel_8423/gring pixel_8423/VDD pixel_8423/GND pixel_8423/VREF pixel_8423/ROW_SEL
+ pixel_8423/NB1 pixel_8423/VBIAS pixel_8423/NB2 pixel_8423/AMP_IN pixel_8423/SF_IB
+ pixel_8423/PIX_OUT pixel_8423/CSA_VREF pixel
Xpixel_8412 pixel_8412/gring pixel_8412/VDD pixel_8412/GND pixel_8412/VREF pixel_8412/ROW_SEL
+ pixel_8412/NB1 pixel_8412/VBIAS pixel_8412/NB2 pixel_8412/AMP_IN pixel_8412/SF_IB
+ pixel_8412/PIX_OUT pixel_8412/CSA_VREF pixel
Xpixel_9179 pixel_9179/gring pixel_9179/VDD pixel_9179/GND pixel_9179/VREF pixel_9179/ROW_SEL
+ pixel_9179/NB1 pixel_9179/VBIAS pixel_9179/NB2 pixel_9179/AMP_IN pixel_9179/SF_IB
+ pixel_9179/PIX_OUT pixel_9179/CSA_VREF pixel
Xpixel_9168 pixel_9168/gring pixel_9168/VDD pixel_9168/GND pixel_9168/VREF pixel_9168/ROW_SEL
+ pixel_9168/NB1 pixel_9168/VBIAS pixel_9168/NB2 pixel_9168/AMP_IN pixel_9168/SF_IB
+ pixel_9168/PIX_OUT pixel_9168/CSA_VREF pixel
Xpixel_9157 pixel_9157/gring pixel_9157/VDD pixel_9157/GND pixel_9157/VREF pixel_9157/ROW_SEL
+ pixel_9157/NB1 pixel_9157/VBIAS pixel_9157/NB2 pixel_9157/AMP_IN pixel_9157/SF_IB
+ pixel_9157/PIX_OUT pixel_9157/CSA_VREF pixel
Xpixel_7700 pixel_7700/gring pixel_7700/VDD pixel_7700/GND pixel_7700/VREF pixel_7700/ROW_SEL
+ pixel_7700/NB1 pixel_7700/VBIAS pixel_7700/NB2 pixel_7700/AMP_IN pixel_7700/SF_IB
+ pixel_7700/PIX_OUT pixel_7700/CSA_VREF pixel
Xpixel_8445 pixel_8445/gring pixel_8445/VDD pixel_8445/GND pixel_8445/VREF pixel_8445/ROW_SEL
+ pixel_8445/NB1 pixel_8445/VBIAS pixel_8445/NB2 pixel_8445/AMP_IN pixel_8445/SF_IB
+ pixel_8445/PIX_OUT pixel_8445/CSA_VREF pixel
Xpixel_8456 pixel_8456/gring pixel_8456/VDD pixel_8456/GND pixel_8456/VREF pixel_8456/ROW_SEL
+ pixel_8456/NB1 pixel_8456/VBIAS pixel_8456/NB2 pixel_8456/AMP_IN pixel_8456/SF_IB
+ pixel_8456/PIX_OUT pixel_8456/CSA_VREF pixel
Xpixel_8467 pixel_8467/gring pixel_8467/VDD pixel_8467/GND pixel_8467/VREF pixel_8467/ROW_SEL
+ pixel_8467/NB1 pixel_8467/VBIAS pixel_8467/NB2 pixel_8467/AMP_IN pixel_8467/SF_IB
+ pixel_8467/PIX_OUT pixel_8467/CSA_VREF pixel
Xpixel_8478 pixel_8478/gring pixel_8478/VDD pixel_8478/GND pixel_8478/VREF pixel_8478/ROW_SEL
+ pixel_8478/NB1 pixel_8478/VBIAS pixel_8478/NB2 pixel_8478/AMP_IN pixel_8478/SF_IB
+ pixel_8478/PIX_OUT pixel_8478/CSA_VREF pixel
Xpixel_7711 pixel_7711/gring pixel_7711/VDD pixel_7711/GND pixel_7711/VREF pixel_7711/ROW_SEL
+ pixel_7711/NB1 pixel_7711/VBIAS pixel_7711/NB2 pixel_7711/AMP_IN pixel_7711/SF_IB
+ pixel_7711/PIX_OUT pixel_7711/CSA_VREF pixel
Xpixel_7722 pixel_7722/gring pixel_7722/VDD pixel_7722/GND pixel_7722/VREF pixel_7722/ROW_SEL
+ pixel_7722/NB1 pixel_7722/VBIAS pixel_7722/NB2 pixel_7722/AMP_IN pixel_7722/SF_IB
+ pixel_7722/PIX_OUT pixel_7722/CSA_VREF pixel
Xpixel_7733 pixel_7733/gring pixel_7733/VDD pixel_7733/GND pixel_7733/VREF pixel_7733/ROW_SEL
+ pixel_7733/NB1 pixel_7733/VBIAS pixel_7733/NB2 pixel_7733/AMP_IN pixel_7733/SF_IB
+ pixel_7733/PIX_OUT pixel_7733/CSA_VREF pixel
Xpixel_8489 pixel_8489/gring pixel_8489/VDD pixel_8489/GND pixel_8489/VREF pixel_8489/ROW_SEL
+ pixel_8489/NB1 pixel_8489/VBIAS pixel_8489/NB2 pixel_8489/AMP_IN pixel_8489/SF_IB
+ pixel_8489/PIX_OUT pixel_8489/CSA_VREF pixel
Xpixel_7744 pixel_7744/gring pixel_7744/VDD pixel_7744/GND pixel_7744/VREF pixel_7744/ROW_SEL
+ pixel_7744/NB1 pixel_7744/VBIAS pixel_7744/NB2 pixel_7744/AMP_IN pixel_7744/SF_IB
+ pixel_7744/PIX_OUT pixel_7744/CSA_VREF pixel
Xpixel_7755 pixel_7755/gring pixel_7755/VDD pixel_7755/GND pixel_7755/VREF pixel_7755/ROW_SEL
+ pixel_7755/NB1 pixel_7755/VBIAS pixel_7755/NB2 pixel_7755/AMP_IN pixel_7755/SF_IB
+ pixel_7755/PIX_OUT pixel_7755/CSA_VREF pixel
Xpixel_7766 pixel_7766/gring pixel_7766/VDD pixel_7766/GND pixel_7766/VREF pixel_7766/ROW_SEL
+ pixel_7766/NB1 pixel_7766/VBIAS pixel_7766/NB2 pixel_7766/AMP_IN pixel_7766/SF_IB
+ pixel_7766/PIX_OUT pixel_7766/CSA_VREF pixel
Xpixel_7777 pixel_7777/gring pixel_7777/VDD pixel_7777/GND pixel_7777/VREF pixel_7777/ROW_SEL
+ pixel_7777/NB1 pixel_7777/VBIAS pixel_7777/NB2 pixel_7777/AMP_IN pixel_7777/SF_IB
+ pixel_7777/PIX_OUT pixel_7777/CSA_VREF pixel
Xpixel_7788 pixel_7788/gring pixel_7788/VDD pixel_7788/GND pixel_7788/VREF pixel_7788/ROW_SEL
+ pixel_7788/NB1 pixel_7788/VBIAS pixel_7788/NB2 pixel_7788/AMP_IN pixel_7788/SF_IB
+ pixel_7788/PIX_OUT pixel_7788/CSA_VREF pixel
Xpixel_7799 pixel_7799/gring pixel_7799/VDD pixel_7799/GND pixel_7799/VREF pixel_7799/ROW_SEL
+ pixel_7799/NB1 pixel_7799/VBIAS pixel_7799/NB2 pixel_7799/AMP_IN pixel_7799/SF_IB
+ pixel_7799/PIX_OUT pixel_7799/CSA_VREF pixel
Xpixel_2062 pixel_2062/gring pixel_2062/VDD pixel_2062/GND pixel_2062/VREF pixel_2062/ROW_SEL
+ pixel_2062/NB1 pixel_2062/VBIAS pixel_2062/NB2 pixel_2062/AMP_IN pixel_2062/SF_IB
+ pixel_2062/PIX_OUT pixel_2062/CSA_VREF pixel
Xpixel_2051 pixel_2051/gring pixel_2051/VDD pixel_2051/GND pixel_2051/VREF pixel_2051/ROW_SEL
+ pixel_2051/NB1 pixel_2051/VBIAS pixel_2051/NB2 pixel_2051/AMP_IN pixel_2051/SF_IB
+ pixel_2051/PIX_OUT pixel_2051/CSA_VREF pixel
Xpixel_2040 pixel_2040/gring pixel_2040/VDD pixel_2040/GND pixel_2040/VREF pixel_2040/ROW_SEL
+ pixel_2040/NB1 pixel_2040/VBIAS pixel_2040/NB2 pixel_2040/AMP_IN pixel_2040/SF_IB
+ pixel_2040/PIX_OUT pixel_2040/CSA_VREF pixel
Xpixel_1361 pixel_1361/gring pixel_1361/VDD pixel_1361/GND pixel_1361/VREF pixel_1361/ROW_SEL
+ pixel_1361/NB1 pixel_1361/VBIAS pixel_1361/NB2 pixel_1361/AMP_IN pixel_1361/SF_IB
+ pixel_1361/PIX_OUT pixel_1361/CSA_VREF pixel
Xpixel_1350 pixel_1350/gring pixel_1350/VDD pixel_1350/GND pixel_1350/VREF pixel_1350/ROW_SEL
+ pixel_1350/NB1 pixel_1350/VBIAS pixel_1350/NB2 pixel_1350/AMP_IN pixel_1350/SF_IB
+ pixel_1350/PIX_OUT pixel_1350/CSA_VREF pixel
Xpixel_2095 pixel_2095/gring pixel_2095/VDD pixel_2095/GND pixel_2095/VREF pixel_2095/ROW_SEL
+ pixel_2095/NB1 pixel_2095/VBIAS pixel_2095/NB2 pixel_2095/AMP_IN pixel_2095/SF_IB
+ pixel_2095/PIX_OUT pixel_2095/CSA_VREF pixel
Xpixel_2084 pixel_2084/gring pixel_2084/VDD pixel_2084/GND pixel_2084/VREF pixel_2084/ROW_SEL
+ pixel_2084/NB1 pixel_2084/VBIAS pixel_2084/NB2 pixel_2084/AMP_IN pixel_2084/SF_IB
+ pixel_2084/PIX_OUT pixel_2084/CSA_VREF pixel
Xpixel_2073 pixel_2073/gring pixel_2073/VDD pixel_2073/GND pixel_2073/VREF pixel_2073/ROW_SEL
+ pixel_2073/NB1 pixel_2073/VBIAS pixel_2073/NB2 pixel_2073/AMP_IN pixel_2073/SF_IB
+ pixel_2073/PIX_OUT pixel_2073/CSA_VREF pixel
Xpixel_1394 pixel_1394/gring pixel_1394/VDD pixel_1394/GND pixel_1394/VREF pixel_1394/ROW_SEL
+ pixel_1394/NB1 pixel_1394/VBIAS pixel_1394/NB2 pixel_1394/AMP_IN pixel_1394/SF_IB
+ pixel_1394/PIX_OUT pixel_1394/CSA_VREF pixel
Xpixel_1383 pixel_1383/gring pixel_1383/VDD pixel_1383/GND pixel_1383/VREF pixel_1383/ROW_SEL
+ pixel_1383/NB1 pixel_1383/VBIAS pixel_1383/NB2 pixel_1383/AMP_IN pixel_1383/SF_IB
+ pixel_1383/PIX_OUT pixel_1383/CSA_VREF pixel
Xpixel_1372 pixel_1372/gring pixel_1372/VDD pixel_1372/GND pixel_1372/VREF pixel_1372/ROW_SEL
+ pixel_1372/NB1 pixel_1372/VBIAS pixel_1372/NB2 pixel_1372/AMP_IN pixel_1372/SF_IB
+ pixel_1372/PIX_OUT pixel_1372/CSA_VREF pixel
Xpixel_9691 pixel_9691/gring pixel_9691/VDD pixel_9691/GND pixel_9691/VREF pixel_9691/ROW_SEL
+ pixel_9691/NB1 pixel_9691/VBIAS pixel_9691/NB2 pixel_9691/AMP_IN pixel_9691/SF_IB
+ pixel_9691/PIX_OUT pixel_9691/CSA_VREF pixel
Xpixel_9680 pixel_9680/gring pixel_9680/VDD pixel_9680/GND pixel_9680/VREF pixel_9680/ROW_SEL
+ pixel_9680/NB1 pixel_9680/VBIAS pixel_9680/NB2 pixel_9680/AMP_IN pixel_9680/SF_IB
+ pixel_9680/PIX_OUT pixel_9680/CSA_VREF pixel
Xpixel_8990 pixel_8990/gring pixel_8990/VDD pixel_8990/GND pixel_8990/VREF pixel_8990/ROW_SEL
+ pixel_8990/NB1 pixel_8990/VBIAS pixel_8990/NB2 pixel_8990/AMP_IN pixel_8990/SF_IB
+ pixel_8990/PIX_OUT pixel_8990/CSA_VREF pixel
Xpixel_409 pixel_409/gring pixel_409/VDD pixel_409/GND pixel_409/VREF pixel_409/ROW_SEL
+ pixel_409/NB1 pixel_409/VBIAS pixel_409/NB2 pixel_409/AMP_IN pixel_409/SF_IB pixel_409/PIX_OUT
+ pixel_409/CSA_VREF pixel
Xpixel_7007 pixel_7007/gring pixel_7007/VDD pixel_7007/GND pixel_7007/VREF pixel_7007/ROW_SEL
+ pixel_7007/NB1 pixel_7007/VBIAS pixel_7007/NB2 pixel_7007/AMP_IN pixel_7007/SF_IB
+ pixel_7007/PIX_OUT pixel_7007/CSA_VREF pixel
Xpixel_7018 pixel_7018/gring pixel_7018/VDD pixel_7018/GND pixel_7018/VREF pixel_7018/ROW_SEL
+ pixel_7018/NB1 pixel_7018/VBIAS pixel_7018/NB2 pixel_7018/AMP_IN pixel_7018/SF_IB
+ pixel_7018/PIX_OUT pixel_7018/CSA_VREF pixel
Xpixel_7029 pixel_7029/gring pixel_7029/VDD pixel_7029/GND pixel_7029/VREF pixel_7029/ROW_SEL
+ pixel_7029/NB1 pixel_7029/VBIAS pixel_7029/NB2 pixel_7029/AMP_IN pixel_7029/SF_IB
+ pixel_7029/PIX_OUT pixel_7029/CSA_VREF pixel
Xpixel_6306 pixel_6306/gring pixel_6306/VDD pixel_6306/GND pixel_6306/VREF pixel_6306/ROW_SEL
+ pixel_6306/NB1 pixel_6306/VBIAS pixel_6306/NB2 pixel_6306/AMP_IN pixel_6306/SF_IB
+ pixel_6306/PIX_OUT pixel_6306/CSA_VREF pixel
Xpixel_6317 pixel_6317/gring pixel_6317/VDD pixel_6317/GND pixel_6317/VREF pixel_6317/ROW_SEL
+ pixel_6317/NB1 pixel_6317/VBIAS pixel_6317/NB2 pixel_6317/AMP_IN pixel_6317/SF_IB
+ pixel_6317/PIX_OUT pixel_6317/CSA_VREF pixel
Xpixel_6328 pixel_6328/gring pixel_6328/VDD pixel_6328/GND pixel_6328/VREF pixel_6328/ROW_SEL
+ pixel_6328/NB1 pixel_6328/VBIAS pixel_6328/NB2 pixel_6328/AMP_IN pixel_6328/SF_IB
+ pixel_6328/PIX_OUT pixel_6328/CSA_VREF pixel
Xpixel_6339 pixel_6339/gring pixel_6339/VDD pixel_6339/GND pixel_6339/VREF pixel_6339/ROW_SEL
+ pixel_6339/NB1 pixel_6339/VBIAS pixel_6339/NB2 pixel_6339/AMP_IN pixel_6339/SF_IB
+ pixel_6339/PIX_OUT pixel_6339/CSA_VREF pixel
Xpixel_5605 pixel_5605/gring pixel_5605/VDD pixel_5605/GND pixel_5605/VREF pixel_5605/ROW_SEL
+ pixel_5605/NB1 pixel_5605/VBIAS pixel_5605/NB2 pixel_5605/AMP_IN pixel_5605/SF_IB
+ pixel_5605/PIX_OUT pixel_5605/CSA_VREF pixel
Xpixel_5616 pixel_5616/gring pixel_5616/VDD pixel_5616/GND pixel_5616/VREF pixel_5616/ROW_SEL
+ pixel_5616/NB1 pixel_5616/VBIAS pixel_5616/NB2 pixel_5616/AMP_IN pixel_5616/SF_IB
+ pixel_5616/PIX_OUT pixel_5616/CSA_VREF pixel
Xpixel_5627 pixel_5627/gring pixel_5627/VDD pixel_5627/GND pixel_5627/VREF pixel_5627/ROW_SEL
+ pixel_5627/NB1 pixel_5627/VBIAS pixel_5627/NB2 pixel_5627/AMP_IN pixel_5627/SF_IB
+ pixel_5627/PIX_OUT pixel_5627/CSA_VREF pixel
Xpixel_5638 pixel_5638/gring pixel_5638/VDD pixel_5638/GND pixel_5638/VREF pixel_5638/ROW_SEL
+ pixel_5638/NB1 pixel_5638/VBIAS pixel_5638/NB2 pixel_5638/AMP_IN pixel_5638/SF_IB
+ pixel_5638/PIX_OUT pixel_5638/CSA_VREF pixel
Xpixel_5649 pixel_5649/gring pixel_5649/VDD pixel_5649/GND pixel_5649/VREF pixel_5649/ROW_SEL
+ pixel_5649/NB1 pixel_5649/VBIAS pixel_5649/NB2 pixel_5649/AMP_IN pixel_5649/SF_IB
+ pixel_5649/PIX_OUT pixel_5649/CSA_VREF pixel
Xpixel_4904 pixel_4904/gring pixel_4904/VDD pixel_4904/GND pixel_4904/VREF pixel_4904/ROW_SEL
+ pixel_4904/NB1 pixel_4904/VBIAS pixel_4904/NB2 pixel_4904/AMP_IN pixel_4904/SF_IB
+ pixel_4904/PIX_OUT pixel_4904/CSA_VREF pixel
Xpixel_932 pixel_932/gring pixel_932/VDD pixel_932/GND pixel_932/VREF pixel_932/ROW_SEL
+ pixel_932/NB1 pixel_932/VBIAS pixel_932/NB2 pixel_932/AMP_IN pixel_932/SF_IB pixel_932/PIX_OUT
+ pixel_932/CSA_VREF pixel
Xpixel_921 pixel_921/gring pixel_921/VDD pixel_921/GND pixel_921/VREF pixel_921/ROW_SEL
+ pixel_921/NB1 pixel_921/VBIAS pixel_921/NB2 pixel_921/AMP_IN pixel_921/SF_IB pixel_921/PIX_OUT
+ pixel_921/CSA_VREF pixel
Xpixel_910 pixel_910/gring pixel_910/VDD pixel_910/GND pixel_910/VREF pixel_910/ROW_SEL
+ pixel_910/NB1 pixel_910/VBIAS pixel_910/NB2 pixel_910/AMP_IN pixel_910/SF_IB pixel_910/PIX_OUT
+ pixel_910/CSA_VREF pixel
Xpixel_4915 pixel_4915/gring pixel_4915/VDD pixel_4915/GND pixel_4915/VREF pixel_4915/ROW_SEL
+ pixel_4915/NB1 pixel_4915/VBIAS pixel_4915/NB2 pixel_4915/AMP_IN pixel_4915/SF_IB
+ pixel_4915/PIX_OUT pixel_4915/CSA_VREF pixel
Xpixel_4926 pixel_4926/gring pixel_4926/VDD pixel_4926/GND pixel_4926/VREF pixel_4926/ROW_SEL
+ pixel_4926/NB1 pixel_4926/VBIAS pixel_4926/NB2 pixel_4926/AMP_IN pixel_4926/SF_IB
+ pixel_4926/PIX_OUT pixel_4926/CSA_VREF pixel
Xpixel_4937 pixel_4937/gring pixel_4937/VDD pixel_4937/GND pixel_4937/VREF pixel_4937/ROW_SEL
+ pixel_4937/NB1 pixel_4937/VBIAS pixel_4937/NB2 pixel_4937/AMP_IN pixel_4937/SF_IB
+ pixel_4937/PIX_OUT pixel_4937/CSA_VREF pixel
Xpixel_976 pixel_976/gring pixel_976/VDD pixel_976/GND pixel_976/VREF pixel_976/ROW_SEL
+ pixel_976/NB1 pixel_976/VBIAS pixel_976/NB2 pixel_976/AMP_IN pixel_976/SF_IB pixel_976/PIX_OUT
+ pixel_976/CSA_VREF pixel
Xpixel_965 pixel_965/gring pixel_965/VDD pixel_965/GND pixel_965/VREF pixel_965/ROW_SEL
+ pixel_965/NB1 pixel_965/VBIAS pixel_965/NB2 pixel_965/AMP_IN pixel_965/SF_IB pixel_965/PIX_OUT
+ pixel_965/CSA_VREF pixel
Xpixel_954 pixel_954/gring pixel_954/VDD pixel_954/GND pixel_954/VREF pixel_954/ROW_SEL
+ pixel_954/NB1 pixel_954/VBIAS pixel_954/NB2 pixel_954/AMP_IN pixel_954/SF_IB pixel_954/PIX_OUT
+ pixel_954/CSA_VREF pixel
Xpixel_943 pixel_943/gring pixel_943/VDD pixel_943/GND pixel_943/VREF pixel_943/ROW_SEL
+ pixel_943/NB1 pixel_943/VBIAS pixel_943/NB2 pixel_943/AMP_IN pixel_943/SF_IB pixel_943/PIX_OUT
+ pixel_943/CSA_VREF pixel
Xpixel_4948 pixel_4948/gring pixel_4948/VDD pixel_4948/GND pixel_4948/VREF pixel_4948/ROW_SEL
+ pixel_4948/NB1 pixel_4948/VBIAS pixel_4948/NB2 pixel_4948/AMP_IN pixel_4948/SF_IB
+ pixel_4948/PIX_OUT pixel_4948/CSA_VREF pixel
Xpixel_4959 pixel_4959/gring pixel_4959/VDD pixel_4959/GND pixel_4959/VREF pixel_4959/ROW_SEL
+ pixel_4959/NB1 pixel_4959/VBIAS pixel_4959/NB2 pixel_4959/AMP_IN pixel_4959/SF_IB
+ pixel_4959/PIX_OUT pixel_4959/CSA_VREF pixel
Xpixel_998 pixel_998/gring pixel_998/VDD pixel_998/GND pixel_998/VREF pixel_998/ROW_SEL
+ pixel_998/NB1 pixel_998/VBIAS pixel_998/NB2 pixel_998/AMP_IN pixel_998/SF_IB pixel_998/PIX_OUT
+ pixel_998/CSA_VREF pixel
Xpixel_987 pixel_987/gring pixel_987/VDD pixel_987/GND pixel_987/VREF pixel_987/ROW_SEL
+ pixel_987/NB1 pixel_987/VBIAS pixel_987/NB2 pixel_987/AMP_IN pixel_987/SF_IB pixel_987/PIX_OUT
+ pixel_987/CSA_VREF pixel
Xpixel_8220 pixel_8220/gring pixel_8220/VDD pixel_8220/GND pixel_8220/VREF pixel_8220/ROW_SEL
+ pixel_8220/NB1 pixel_8220/VBIAS pixel_8220/NB2 pixel_8220/AMP_IN pixel_8220/SF_IB
+ pixel_8220/PIX_OUT pixel_8220/CSA_VREF pixel
Xpixel_8231 pixel_8231/gring pixel_8231/VDD pixel_8231/GND pixel_8231/VREF pixel_8231/ROW_SEL
+ pixel_8231/NB1 pixel_8231/VBIAS pixel_8231/NB2 pixel_8231/AMP_IN pixel_8231/SF_IB
+ pixel_8231/PIX_OUT pixel_8231/CSA_VREF pixel
Xpixel_8242 pixel_8242/gring pixel_8242/VDD pixel_8242/GND pixel_8242/VREF pixel_8242/ROW_SEL
+ pixel_8242/NB1 pixel_8242/VBIAS pixel_8242/NB2 pixel_8242/AMP_IN pixel_8242/SF_IB
+ pixel_8242/PIX_OUT pixel_8242/CSA_VREF pixel
Xpixel_8253 pixel_8253/gring pixel_8253/VDD pixel_8253/GND pixel_8253/VREF pixel_8253/ROW_SEL
+ pixel_8253/NB1 pixel_8253/VBIAS pixel_8253/NB2 pixel_8253/AMP_IN pixel_8253/SF_IB
+ pixel_8253/PIX_OUT pixel_8253/CSA_VREF pixel
Xpixel_8264 pixel_8264/gring pixel_8264/VDD pixel_8264/GND pixel_8264/VREF pixel_8264/ROW_SEL
+ pixel_8264/NB1 pixel_8264/VBIAS pixel_8264/NB2 pixel_8264/AMP_IN pixel_8264/SF_IB
+ pixel_8264/PIX_OUT pixel_8264/CSA_VREF pixel
Xpixel_8275 pixel_8275/gring pixel_8275/VDD pixel_8275/GND pixel_8275/VREF pixel_8275/ROW_SEL
+ pixel_8275/NB1 pixel_8275/VBIAS pixel_8275/NB2 pixel_8275/AMP_IN pixel_8275/SF_IB
+ pixel_8275/PIX_OUT pixel_8275/CSA_VREF pixel
Xpixel_8286 pixel_8286/gring pixel_8286/VDD pixel_8286/GND pixel_8286/VREF pixel_8286/ROW_SEL
+ pixel_8286/NB1 pixel_8286/VBIAS pixel_8286/NB2 pixel_8286/AMP_IN pixel_8286/SF_IB
+ pixel_8286/PIX_OUT pixel_8286/CSA_VREF pixel
Xpixel_7530 pixel_7530/gring pixel_7530/VDD pixel_7530/GND pixel_7530/VREF pixel_7530/ROW_SEL
+ pixel_7530/NB1 pixel_7530/VBIAS pixel_7530/NB2 pixel_7530/AMP_IN pixel_7530/SF_IB
+ pixel_7530/PIX_OUT pixel_7530/CSA_VREF pixel
Xpixel_7541 pixel_7541/gring pixel_7541/VDD pixel_7541/GND pixel_7541/VREF pixel_7541/ROW_SEL
+ pixel_7541/NB1 pixel_7541/VBIAS pixel_7541/NB2 pixel_7541/AMP_IN pixel_7541/SF_IB
+ pixel_7541/PIX_OUT pixel_7541/CSA_VREF pixel
Xpixel_8297 pixel_8297/gring pixel_8297/VDD pixel_8297/GND pixel_8297/VREF pixel_8297/ROW_SEL
+ pixel_8297/NB1 pixel_8297/VBIAS pixel_8297/NB2 pixel_8297/AMP_IN pixel_8297/SF_IB
+ pixel_8297/PIX_OUT pixel_8297/CSA_VREF pixel
Xpixel_7552 pixel_7552/gring pixel_7552/VDD pixel_7552/GND pixel_7552/VREF pixel_7552/ROW_SEL
+ pixel_7552/NB1 pixel_7552/VBIAS pixel_7552/NB2 pixel_7552/AMP_IN pixel_7552/SF_IB
+ pixel_7552/PIX_OUT pixel_7552/CSA_VREF pixel
Xpixel_7563 pixel_7563/gring pixel_7563/VDD pixel_7563/GND pixel_7563/VREF pixel_7563/ROW_SEL
+ pixel_7563/NB1 pixel_7563/VBIAS pixel_7563/NB2 pixel_7563/AMP_IN pixel_7563/SF_IB
+ pixel_7563/PIX_OUT pixel_7563/CSA_VREF pixel
Xpixel_7574 pixel_7574/gring pixel_7574/VDD pixel_7574/GND pixel_7574/VREF pixel_7574/ROW_SEL
+ pixel_7574/NB1 pixel_7574/VBIAS pixel_7574/NB2 pixel_7574/AMP_IN pixel_7574/SF_IB
+ pixel_7574/PIX_OUT pixel_7574/CSA_VREF pixel
Xpixel_6840 pixel_6840/gring pixel_6840/VDD pixel_6840/GND pixel_6840/VREF pixel_6840/ROW_SEL
+ pixel_6840/NB1 pixel_6840/VBIAS pixel_6840/NB2 pixel_6840/AMP_IN pixel_6840/SF_IB
+ pixel_6840/PIX_OUT pixel_6840/CSA_VREF pixel
Xpixel_7585 pixel_7585/gring pixel_7585/VDD pixel_7585/GND pixel_7585/VREF pixel_7585/ROW_SEL
+ pixel_7585/NB1 pixel_7585/VBIAS pixel_7585/NB2 pixel_7585/AMP_IN pixel_7585/SF_IB
+ pixel_7585/PIX_OUT pixel_7585/CSA_VREF pixel
Xpixel_7596 pixel_7596/gring pixel_7596/VDD pixel_7596/GND pixel_7596/VREF pixel_7596/ROW_SEL
+ pixel_7596/NB1 pixel_7596/VBIAS pixel_7596/NB2 pixel_7596/AMP_IN pixel_7596/SF_IB
+ pixel_7596/PIX_OUT pixel_7596/CSA_VREF pixel
Xpixel_6851 pixel_6851/gring pixel_6851/VDD pixel_6851/GND pixel_6851/VREF pixel_6851/ROW_SEL
+ pixel_6851/NB1 pixel_6851/VBIAS pixel_6851/NB2 pixel_6851/AMP_IN pixel_6851/SF_IB
+ pixel_6851/PIX_OUT pixel_6851/CSA_VREF pixel
Xpixel_6862 pixel_6862/gring pixel_6862/VDD pixel_6862/GND pixel_6862/VREF pixel_6862/ROW_SEL
+ pixel_6862/NB1 pixel_6862/VBIAS pixel_6862/NB2 pixel_6862/AMP_IN pixel_6862/SF_IB
+ pixel_6862/PIX_OUT pixel_6862/CSA_VREF pixel
Xpixel_6873 pixel_6873/gring pixel_6873/VDD pixel_6873/GND pixel_6873/VREF pixel_6873/ROW_SEL
+ pixel_6873/NB1 pixel_6873/VBIAS pixel_6873/NB2 pixel_6873/AMP_IN pixel_6873/SF_IB
+ pixel_6873/PIX_OUT pixel_6873/CSA_VREF pixel
Xpixel_6884 pixel_6884/gring pixel_6884/VDD pixel_6884/GND pixel_6884/VREF pixel_6884/ROW_SEL
+ pixel_6884/NB1 pixel_6884/VBIAS pixel_6884/NB2 pixel_6884/AMP_IN pixel_6884/SF_IB
+ pixel_6884/PIX_OUT pixel_6884/CSA_VREF pixel
Xpixel_6895 pixel_6895/gring pixel_6895/VDD pixel_6895/GND pixel_6895/VREF pixel_6895/ROW_SEL
+ pixel_6895/NB1 pixel_6895/VBIAS pixel_6895/NB2 pixel_6895/AMP_IN pixel_6895/SF_IB
+ pixel_6895/PIX_OUT pixel_6895/CSA_VREF pixel
Xpixel_1191 pixel_1191/gring pixel_1191/VDD pixel_1191/GND pixel_1191/VREF pixel_1191/ROW_SEL
+ pixel_1191/NB1 pixel_1191/VBIAS pixel_1191/NB2 pixel_1191/AMP_IN pixel_1191/SF_IB
+ pixel_1191/PIX_OUT pixel_1191/CSA_VREF pixel
Xpixel_1180 pixel_1180/gring pixel_1180/VDD pixel_1180/GND pixel_1180/VREF pixel_1180/ROW_SEL
+ pixel_1180/NB1 pixel_1180/VBIAS pixel_1180/NB2 pixel_1180/AMP_IN pixel_1180/SF_IB
+ pixel_1180/PIX_OUT pixel_1180/CSA_VREF pixel
Xpixel_228 pixel_228/gring pixel_228/VDD pixel_228/GND pixel_228/VREF pixel_228/ROW_SEL
+ pixel_228/NB1 pixel_228/VBIAS pixel_228/NB2 pixel_228/AMP_IN pixel_228/SF_IB pixel_228/PIX_OUT
+ pixel_228/CSA_VREF pixel
Xpixel_217 pixel_217/gring pixel_217/VDD pixel_217/GND pixel_217/VREF pixel_217/ROW_SEL
+ pixel_217/NB1 pixel_217/VBIAS pixel_217/NB2 pixel_217/AMP_IN pixel_217/SF_IB pixel_217/PIX_OUT
+ pixel_217/CSA_VREF pixel
Xpixel_206 pixel_206/gring pixel_206/VDD pixel_206/GND pixel_206/VREF pixel_206/ROW_SEL
+ pixel_206/NB1 pixel_206/VBIAS pixel_206/NB2 pixel_206/AMP_IN pixel_206/SF_IB pixel_206/PIX_OUT
+ pixel_206/CSA_VREF pixel
Xpixel_239 pixel_239/gring pixel_239/VDD pixel_239/GND pixel_239/VREF pixel_239/ROW_SEL
+ pixel_239/NB1 pixel_239/VBIAS pixel_239/NB2 pixel_239/AMP_IN pixel_239/SF_IB pixel_239/PIX_OUT
+ pixel_239/CSA_VREF pixel
Xpixel_2809 pixel_2809/gring pixel_2809/VDD pixel_2809/GND pixel_2809/VREF pixel_2809/ROW_SEL
+ pixel_2809/NB1 pixel_2809/VBIAS pixel_2809/NB2 pixel_2809/AMP_IN pixel_2809/SF_IB
+ pixel_2809/PIX_OUT pixel_2809/CSA_VREF pixel
Xpixel_6103 pixel_6103/gring pixel_6103/VDD pixel_6103/GND pixel_6103/VREF pixel_6103/ROW_SEL
+ pixel_6103/NB1 pixel_6103/VBIAS pixel_6103/NB2 pixel_6103/AMP_IN pixel_6103/SF_IB
+ pixel_6103/PIX_OUT pixel_6103/CSA_VREF pixel
Xpixel_6114 pixel_6114/gring pixel_6114/VDD pixel_6114/GND pixel_6114/VREF pixel_6114/ROW_SEL
+ pixel_6114/NB1 pixel_6114/VBIAS pixel_6114/NB2 pixel_6114/AMP_IN pixel_6114/SF_IB
+ pixel_6114/PIX_OUT pixel_6114/CSA_VREF pixel
Xpixel_6125 pixel_6125/gring pixel_6125/VDD pixel_6125/GND pixel_6125/VREF pixel_6125/ROW_SEL
+ pixel_6125/NB1 pixel_6125/VBIAS pixel_6125/NB2 pixel_6125/AMP_IN pixel_6125/SF_IB
+ pixel_6125/PIX_OUT pixel_6125/CSA_VREF pixel
Xpixel_6136 pixel_6136/gring pixel_6136/VDD pixel_6136/GND pixel_6136/VREF pixel_6136/ROW_SEL
+ pixel_6136/NB1 pixel_6136/VBIAS pixel_6136/NB2 pixel_6136/AMP_IN pixel_6136/SF_IB
+ pixel_6136/PIX_OUT pixel_6136/CSA_VREF pixel
Xpixel_6147 pixel_6147/gring pixel_6147/VDD pixel_6147/GND pixel_6147/VREF pixel_6147/ROW_SEL
+ pixel_6147/NB1 pixel_6147/VBIAS pixel_6147/NB2 pixel_6147/AMP_IN pixel_6147/SF_IB
+ pixel_6147/PIX_OUT pixel_6147/CSA_VREF pixel
Xpixel_6158 pixel_6158/gring pixel_6158/VDD pixel_6158/GND pixel_6158/VREF pixel_6158/ROW_SEL
+ pixel_6158/NB1 pixel_6158/VBIAS pixel_6158/NB2 pixel_6158/AMP_IN pixel_6158/SF_IB
+ pixel_6158/PIX_OUT pixel_6158/CSA_VREF pixel
Xpixel_5402 pixel_5402/gring pixel_5402/VDD pixel_5402/GND pixel_5402/VREF pixel_5402/ROW_SEL
+ pixel_5402/NB1 pixel_5402/VBIAS pixel_5402/NB2 pixel_5402/AMP_IN pixel_5402/SF_IB
+ pixel_5402/PIX_OUT pixel_5402/CSA_VREF pixel
Xpixel_5413 pixel_5413/gring pixel_5413/VDD pixel_5413/GND pixel_5413/VREF pixel_5413/ROW_SEL
+ pixel_5413/NB1 pixel_5413/VBIAS pixel_5413/NB2 pixel_5413/AMP_IN pixel_5413/SF_IB
+ pixel_5413/PIX_OUT pixel_5413/CSA_VREF pixel
Xpixel_5424 pixel_5424/gring pixel_5424/VDD pixel_5424/GND pixel_5424/VREF pixel_5424/ROW_SEL
+ pixel_5424/NB1 pixel_5424/VBIAS pixel_5424/NB2 pixel_5424/AMP_IN pixel_5424/SF_IB
+ pixel_5424/PIX_OUT pixel_5424/CSA_VREF pixel
Xpixel_6169 pixel_6169/gring pixel_6169/VDD pixel_6169/GND pixel_6169/VREF pixel_6169/ROW_SEL
+ pixel_6169/NB1 pixel_6169/VBIAS pixel_6169/NB2 pixel_6169/AMP_IN pixel_6169/SF_IB
+ pixel_6169/PIX_OUT pixel_6169/CSA_VREF pixel
Xpixel_5435 pixel_5435/gring pixel_5435/VDD pixel_5435/GND pixel_5435/VREF pixel_5435/ROW_SEL
+ pixel_5435/NB1 pixel_5435/VBIAS pixel_5435/NB2 pixel_5435/AMP_IN pixel_5435/SF_IB
+ pixel_5435/PIX_OUT pixel_5435/CSA_VREF pixel
Xpixel_5446 pixel_5446/gring pixel_5446/VDD pixel_5446/GND pixel_5446/VREF pixel_5446/ROW_SEL
+ pixel_5446/NB1 pixel_5446/VBIAS pixel_5446/NB2 pixel_5446/AMP_IN pixel_5446/SF_IB
+ pixel_5446/PIX_OUT pixel_5446/CSA_VREF pixel
Xpixel_5457 pixel_5457/gring pixel_5457/VDD pixel_5457/GND pixel_5457/VREF pixel_5457/ROW_SEL
+ pixel_5457/NB1 pixel_5457/VBIAS pixel_5457/NB2 pixel_5457/AMP_IN pixel_5457/SF_IB
+ pixel_5457/PIX_OUT pixel_5457/CSA_VREF pixel
Xpixel_4701 pixel_4701/gring pixel_4701/VDD pixel_4701/GND pixel_4701/VREF pixel_4701/ROW_SEL
+ pixel_4701/NB1 pixel_4701/VBIAS pixel_4701/NB2 pixel_4701/AMP_IN pixel_4701/SF_IB
+ pixel_4701/PIX_OUT pixel_4701/CSA_VREF pixel
Xpixel_4712 pixel_4712/gring pixel_4712/VDD pixel_4712/GND pixel_4712/VREF pixel_4712/ROW_SEL
+ pixel_4712/NB1 pixel_4712/VBIAS pixel_4712/NB2 pixel_4712/AMP_IN pixel_4712/SF_IB
+ pixel_4712/PIX_OUT pixel_4712/CSA_VREF pixel
Xpixel_751 pixel_751/gring pixel_751/VDD pixel_751/GND pixel_751/VREF pixel_751/ROW_SEL
+ pixel_751/NB1 pixel_751/VBIAS pixel_751/NB2 pixel_751/AMP_IN pixel_751/SF_IB pixel_751/PIX_OUT
+ pixel_751/CSA_VREF pixel
Xpixel_740 pixel_740/gring pixel_740/VDD pixel_740/GND pixel_740/VREF pixel_740/ROW_SEL
+ pixel_740/NB1 pixel_740/VBIAS pixel_740/NB2 pixel_740/AMP_IN pixel_740/SF_IB pixel_740/PIX_OUT
+ pixel_740/CSA_VREF pixel
Xpixel_5468 pixel_5468/gring pixel_5468/VDD pixel_5468/GND pixel_5468/VREF pixel_5468/ROW_SEL
+ pixel_5468/NB1 pixel_5468/VBIAS pixel_5468/NB2 pixel_5468/AMP_IN pixel_5468/SF_IB
+ pixel_5468/PIX_OUT pixel_5468/CSA_VREF pixel
Xpixel_5479 pixel_5479/gring pixel_5479/VDD pixel_5479/GND pixel_5479/VREF pixel_5479/ROW_SEL
+ pixel_5479/NB1 pixel_5479/VBIAS pixel_5479/NB2 pixel_5479/AMP_IN pixel_5479/SF_IB
+ pixel_5479/PIX_OUT pixel_5479/CSA_VREF pixel
Xpixel_4723 pixel_4723/gring pixel_4723/VDD pixel_4723/GND pixel_4723/VREF pixel_4723/ROW_SEL
+ pixel_4723/NB1 pixel_4723/VBIAS pixel_4723/NB2 pixel_4723/AMP_IN pixel_4723/SF_IB
+ pixel_4723/PIX_OUT pixel_4723/CSA_VREF pixel
Xpixel_4734 pixel_4734/gring pixel_4734/VDD pixel_4734/GND pixel_4734/VREF pixel_4734/ROW_SEL
+ pixel_4734/NB1 pixel_4734/VBIAS pixel_4734/NB2 pixel_4734/AMP_IN pixel_4734/SF_IB
+ pixel_4734/PIX_OUT pixel_4734/CSA_VREF pixel
Xpixel_4745 pixel_4745/gring pixel_4745/VDD pixel_4745/GND pixel_4745/VREF pixel_4745/ROW_SEL
+ pixel_4745/NB1 pixel_4745/VBIAS pixel_4745/NB2 pixel_4745/AMP_IN pixel_4745/SF_IB
+ pixel_4745/PIX_OUT pixel_4745/CSA_VREF pixel
Xpixel_784 pixel_784/gring pixel_784/VDD pixel_784/GND pixel_784/VREF pixel_784/ROW_SEL
+ pixel_784/NB1 pixel_784/VBIAS pixel_784/NB2 pixel_784/AMP_IN pixel_784/SF_IB pixel_784/PIX_OUT
+ pixel_784/CSA_VREF pixel
Xpixel_773 pixel_773/gring pixel_773/VDD pixel_773/GND pixel_773/VREF pixel_773/ROW_SEL
+ pixel_773/NB1 pixel_773/VBIAS pixel_773/NB2 pixel_773/AMP_IN pixel_773/SF_IB pixel_773/PIX_OUT
+ pixel_773/CSA_VREF pixel
Xpixel_762 pixel_762/gring pixel_762/VDD pixel_762/GND pixel_762/VREF pixel_762/ROW_SEL
+ pixel_762/NB1 pixel_762/VBIAS pixel_762/NB2 pixel_762/AMP_IN pixel_762/SF_IB pixel_762/PIX_OUT
+ pixel_762/CSA_VREF pixel
Xpixel_4756 pixel_4756/gring pixel_4756/VDD pixel_4756/GND pixel_4756/VREF pixel_4756/ROW_SEL
+ pixel_4756/NB1 pixel_4756/VBIAS pixel_4756/NB2 pixel_4756/AMP_IN pixel_4756/SF_IB
+ pixel_4756/PIX_OUT pixel_4756/CSA_VREF pixel
Xpixel_4767 pixel_4767/gring pixel_4767/VDD pixel_4767/GND pixel_4767/VREF pixel_4767/ROW_SEL
+ pixel_4767/NB1 pixel_4767/VBIAS pixel_4767/NB2 pixel_4767/AMP_IN pixel_4767/SF_IB
+ pixel_4767/PIX_OUT pixel_4767/CSA_VREF pixel
Xpixel_4778 pixel_4778/gring pixel_4778/VDD pixel_4778/GND pixel_4778/VREF pixel_4778/ROW_SEL
+ pixel_4778/NB1 pixel_4778/VBIAS pixel_4778/NB2 pixel_4778/AMP_IN pixel_4778/SF_IB
+ pixel_4778/PIX_OUT pixel_4778/CSA_VREF pixel
Xpixel_4789 pixel_4789/gring pixel_4789/VDD pixel_4789/GND pixel_4789/VREF pixel_4789/ROW_SEL
+ pixel_4789/NB1 pixel_4789/VBIAS pixel_4789/NB2 pixel_4789/AMP_IN pixel_4789/SF_IB
+ pixel_4789/PIX_OUT pixel_4789/CSA_VREF pixel
Xpixel_795 pixel_795/gring pixel_795/VDD pixel_795/GND pixel_795/VREF pixel_795/ROW_SEL
+ pixel_795/NB1 pixel_795/VBIAS pixel_795/NB2 pixel_795/AMP_IN pixel_795/SF_IB pixel_795/PIX_OUT
+ pixel_795/CSA_VREF pixel
Xpixel_8050 pixel_8050/gring pixel_8050/VDD pixel_8050/GND pixel_8050/VREF pixel_8050/ROW_SEL
+ pixel_8050/NB1 pixel_8050/VBIAS pixel_8050/NB2 pixel_8050/AMP_IN pixel_8050/SF_IB
+ pixel_8050/PIX_OUT pixel_8050/CSA_VREF pixel
Xpixel_8061 pixel_8061/gring pixel_8061/VDD pixel_8061/GND pixel_8061/VREF pixel_8061/ROW_SEL
+ pixel_8061/NB1 pixel_8061/VBIAS pixel_8061/NB2 pixel_8061/AMP_IN pixel_8061/SF_IB
+ pixel_8061/PIX_OUT pixel_8061/CSA_VREF pixel
Xpixel_8072 pixel_8072/gring pixel_8072/VDD pixel_8072/GND pixel_8072/VREF pixel_8072/ROW_SEL
+ pixel_8072/NB1 pixel_8072/VBIAS pixel_8072/NB2 pixel_8072/AMP_IN pixel_8072/SF_IB
+ pixel_8072/PIX_OUT pixel_8072/CSA_VREF pixel
Xpixel_8083 pixel_8083/gring pixel_8083/VDD pixel_8083/GND pixel_8083/VREF pixel_8083/ROW_SEL
+ pixel_8083/NB1 pixel_8083/VBIAS pixel_8083/NB2 pixel_8083/AMP_IN pixel_8083/SF_IB
+ pixel_8083/PIX_OUT pixel_8083/CSA_VREF pixel
Xpixel_8094 pixel_8094/gring pixel_8094/VDD pixel_8094/GND pixel_8094/VREF pixel_8094/ROW_SEL
+ pixel_8094/NB1 pixel_8094/VBIAS pixel_8094/NB2 pixel_8094/AMP_IN pixel_8094/SF_IB
+ pixel_8094/PIX_OUT pixel_8094/CSA_VREF pixel
Xpixel_7360 pixel_7360/gring pixel_7360/VDD pixel_7360/GND pixel_7360/VREF pixel_7360/ROW_SEL
+ pixel_7360/NB1 pixel_7360/VBIAS pixel_7360/NB2 pixel_7360/AMP_IN pixel_7360/SF_IB
+ pixel_7360/PIX_OUT pixel_7360/CSA_VREF pixel
Xpixel_7371 pixel_7371/gring pixel_7371/VDD pixel_7371/GND pixel_7371/VREF pixel_7371/ROW_SEL
+ pixel_7371/NB1 pixel_7371/VBIAS pixel_7371/NB2 pixel_7371/AMP_IN pixel_7371/SF_IB
+ pixel_7371/PIX_OUT pixel_7371/CSA_VREF pixel
Xpixel_7382 pixel_7382/gring pixel_7382/VDD pixel_7382/GND pixel_7382/VREF pixel_7382/ROW_SEL
+ pixel_7382/NB1 pixel_7382/VBIAS pixel_7382/NB2 pixel_7382/AMP_IN pixel_7382/SF_IB
+ pixel_7382/PIX_OUT pixel_7382/CSA_VREF pixel
Xpixel_7393 pixel_7393/gring pixel_7393/VDD pixel_7393/GND pixel_7393/VREF pixel_7393/ROW_SEL
+ pixel_7393/NB1 pixel_7393/VBIAS pixel_7393/NB2 pixel_7393/AMP_IN pixel_7393/SF_IB
+ pixel_7393/PIX_OUT pixel_7393/CSA_VREF pixel
Xpixel_6670 pixel_6670/gring pixel_6670/VDD pixel_6670/GND pixel_6670/VREF pixel_6670/ROW_SEL
+ pixel_6670/NB1 pixel_6670/VBIAS pixel_6670/NB2 pixel_6670/AMP_IN pixel_6670/SF_IB
+ pixel_6670/PIX_OUT pixel_6670/CSA_VREF pixel
Xpixel_6681 pixel_6681/gring pixel_6681/VDD pixel_6681/GND pixel_6681/VREF pixel_6681/ROW_SEL
+ pixel_6681/NB1 pixel_6681/VBIAS pixel_6681/NB2 pixel_6681/AMP_IN pixel_6681/SF_IB
+ pixel_6681/PIX_OUT pixel_6681/CSA_VREF pixel
Xpixel_6692 pixel_6692/gring pixel_6692/VDD pixel_6692/GND pixel_6692/VREF pixel_6692/ROW_SEL
+ pixel_6692/NB1 pixel_6692/VBIAS pixel_6692/NB2 pixel_6692/AMP_IN pixel_6692/SF_IB
+ pixel_6692/PIX_OUT pixel_6692/CSA_VREF pixel
Xpixel_5980 pixel_5980/gring pixel_5980/VDD pixel_5980/GND pixel_5980/VREF pixel_5980/ROW_SEL
+ pixel_5980/NB1 pixel_5980/VBIAS pixel_5980/NB2 pixel_5980/AMP_IN pixel_5980/SF_IB
+ pixel_5980/PIX_OUT pixel_5980/CSA_VREF pixel
Xpixel_5991 pixel_5991/gring pixel_5991/VDD pixel_5991/GND pixel_5991/VREF pixel_5991/ROW_SEL
+ pixel_5991/NB1 pixel_5991/VBIAS pixel_5991/NB2 pixel_5991/AMP_IN pixel_5991/SF_IB
+ pixel_5991/PIX_OUT pixel_5991/CSA_VREF pixel
Xpixel_4008 pixel_4008/gring pixel_4008/VDD pixel_4008/GND pixel_4008/VREF pixel_4008/ROW_SEL
+ pixel_4008/NB1 pixel_4008/VBIAS pixel_4008/NB2 pixel_4008/AMP_IN pixel_4008/SF_IB
+ pixel_4008/PIX_OUT pixel_4008/CSA_VREF pixel
Xpixel_4019 pixel_4019/gring pixel_4019/VDD pixel_4019/GND pixel_4019/VREF pixel_4019/ROW_SEL
+ pixel_4019/NB1 pixel_4019/VBIAS pixel_4019/NB2 pixel_4019/AMP_IN pixel_4019/SF_IB
+ pixel_4019/PIX_OUT pixel_4019/CSA_VREF pixel
Xpixel_3329 pixel_3329/gring pixel_3329/VDD pixel_3329/GND pixel_3329/VREF pixel_3329/ROW_SEL
+ pixel_3329/NB1 pixel_3329/VBIAS pixel_3329/NB2 pixel_3329/AMP_IN pixel_3329/SF_IB
+ pixel_3329/PIX_OUT pixel_3329/CSA_VREF pixel
Xpixel_3318 pixel_3318/gring pixel_3318/VDD pixel_3318/GND pixel_3318/VREF pixel_3318/ROW_SEL
+ pixel_3318/NB1 pixel_3318/VBIAS pixel_3318/NB2 pixel_3318/AMP_IN pixel_3318/SF_IB
+ pixel_3318/PIX_OUT pixel_3318/CSA_VREF pixel
Xpixel_3307 pixel_3307/gring pixel_3307/VDD pixel_3307/GND pixel_3307/VREF pixel_3307/ROW_SEL
+ pixel_3307/NB1 pixel_3307/VBIAS pixel_3307/NB2 pixel_3307/AMP_IN pixel_3307/SF_IB
+ pixel_3307/PIX_OUT pixel_3307/CSA_VREF pixel
Xpixel_2628 pixel_2628/gring pixel_2628/VDD pixel_2628/GND pixel_2628/VREF pixel_2628/ROW_SEL
+ pixel_2628/NB1 pixel_2628/VBIAS pixel_2628/NB2 pixel_2628/AMP_IN pixel_2628/SF_IB
+ pixel_2628/PIX_OUT pixel_2628/CSA_VREF pixel
Xpixel_2617 pixel_2617/gring pixel_2617/VDD pixel_2617/GND pixel_2617/VREF pixel_2617/ROW_SEL
+ pixel_2617/NB1 pixel_2617/VBIAS pixel_2617/NB2 pixel_2617/AMP_IN pixel_2617/SF_IB
+ pixel_2617/PIX_OUT pixel_2617/CSA_VREF pixel
Xpixel_2606 pixel_2606/gring pixel_2606/VDD pixel_2606/GND pixel_2606/VREF pixel_2606/ROW_SEL
+ pixel_2606/NB1 pixel_2606/VBIAS pixel_2606/NB2 pixel_2606/AMP_IN pixel_2606/SF_IB
+ pixel_2606/PIX_OUT pixel_2606/CSA_VREF pixel
Xpixel_1916 pixel_1916/gring pixel_1916/VDD pixel_1916/GND pixel_1916/VREF pixel_1916/ROW_SEL
+ pixel_1916/NB1 pixel_1916/VBIAS pixel_1916/NB2 pixel_1916/AMP_IN pixel_1916/SF_IB
+ pixel_1916/PIX_OUT pixel_1916/CSA_VREF pixel
Xpixel_1905 pixel_1905/gring pixel_1905/VDD pixel_1905/GND pixel_1905/VREF pixel_1905/ROW_SEL
+ pixel_1905/NB1 pixel_1905/VBIAS pixel_1905/NB2 pixel_1905/AMP_IN pixel_1905/SF_IB
+ pixel_1905/PIX_OUT pixel_1905/CSA_VREF pixel
Xpixel_2639 pixel_2639/gring pixel_2639/VDD pixel_2639/GND pixel_2639/VREF pixel_2639/ROW_SEL
+ pixel_2639/NB1 pixel_2639/VBIAS pixel_2639/NB2 pixel_2639/AMP_IN pixel_2639/SF_IB
+ pixel_2639/PIX_OUT pixel_2639/CSA_VREF pixel
Xpixel_1949 pixel_1949/gring pixel_1949/VDD pixel_1949/GND pixel_1949/VREF pixel_1949/ROW_SEL
+ pixel_1949/NB1 pixel_1949/VBIAS pixel_1949/NB2 pixel_1949/AMP_IN pixel_1949/SF_IB
+ pixel_1949/PIX_OUT pixel_1949/CSA_VREF pixel
Xpixel_1938 pixel_1938/gring pixel_1938/VDD pixel_1938/GND pixel_1938/VREF pixel_1938/ROW_SEL
+ pixel_1938/NB1 pixel_1938/VBIAS pixel_1938/NB2 pixel_1938/AMP_IN pixel_1938/SF_IB
+ pixel_1938/PIX_OUT pixel_1938/CSA_VREF pixel
Xpixel_1927 pixel_1927/gring pixel_1927/VDD pixel_1927/GND pixel_1927/VREF pixel_1927/ROW_SEL
+ pixel_1927/NB1 pixel_1927/VBIAS pixel_1927/NB2 pixel_1927/AMP_IN pixel_1927/SF_IB
+ pixel_1927/PIX_OUT pixel_1927/CSA_VREF pixel
Xpixel_5210 pixel_5210/gring pixel_5210/VDD pixel_5210/GND pixel_5210/VREF pixel_5210/ROW_SEL
+ pixel_5210/NB1 pixel_5210/VBIAS pixel_5210/NB2 pixel_5210/AMP_IN pixel_5210/SF_IB
+ pixel_5210/PIX_OUT pixel_5210/CSA_VREF pixel
Xpixel_5221 pixel_5221/gring pixel_5221/VDD pixel_5221/GND pixel_5221/VREF pixel_5221/ROW_SEL
+ pixel_5221/NB1 pixel_5221/VBIAS pixel_5221/NB2 pixel_5221/AMP_IN pixel_5221/SF_IB
+ pixel_5221/PIX_OUT pixel_5221/CSA_VREF pixel
Xpixel_5232 pixel_5232/gring pixel_5232/VDD pixel_5232/GND pixel_5232/VREF pixel_5232/ROW_SEL
+ pixel_5232/NB1 pixel_5232/VBIAS pixel_5232/NB2 pixel_5232/AMP_IN pixel_5232/SF_IB
+ pixel_5232/PIX_OUT pixel_5232/CSA_VREF pixel
Xpixel_5243 pixel_5243/gring pixel_5243/VDD pixel_5243/GND pixel_5243/VREF pixel_5243/ROW_SEL
+ pixel_5243/NB1 pixel_5243/VBIAS pixel_5243/NB2 pixel_5243/AMP_IN pixel_5243/SF_IB
+ pixel_5243/PIX_OUT pixel_5243/CSA_VREF pixel
Xpixel_5254 pixel_5254/gring pixel_5254/VDD pixel_5254/GND pixel_5254/VREF pixel_5254/ROW_SEL
+ pixel_5254/NB1 pixel_5254/VBIAS pixel_5254/NB2 pixel_5254/AMP_IN pixel_5254/SF_IB
+ pixel_5254/PIX_OUT pixel_5254/CSA_VREF pixel
Xpixel_5265 pixel_5265/gring pixel_5265/VDD pixel_5265/GND pixel_5265/VREF pixel_5265/ROW_SEL
+ pixel_5265/NB1 pixel_5265/VBIAS pixel_5265/NB2 pixel_5265/AMP_IN pixel_5265/SF_IB
+ pixel_5265/PIX_OUT pixel_5265/CSA_VREF pixel
Xpixel_4520 pixel_4520/gring pixel_4520/VDD pixel_4520/GND pixel_4520/VREF pixel_4520/ROW_SEL
+ pixel_4520/NB1 pixel_4520/VBIAS pixel_4520/NB2 pixel_4520/AMP_IN pixel_4520/SF_IB
+ pixel_4520/PIX_OUT pixel_4520/CSA_VREF pixel
Xpixel_5276 pixel_5276/gring pixel_5276/VDD pixel_5276/GND pixel_5276/VREF pixel_5276/ROW_SEL
+ pixel_5276/NB1 pixel_5276/VBIAS pixel_5276/NB2 pixel_5276/AMP_IN pixel_5276/SF_IB
+ pixel_5276/PIX_OUT pixel_5276/CSA_VREF pixel
Xpixel_5287 pixel_5287/gring pixel_5287/VDD pixel_5287/GND pixel_5287/VREF pixel_5287/ROW_SEL
+ pixel_5287/NB1 pixel_5287/VBIAS pixel_5287/NB2 pixel_5287/AMP_IN pixel_5287/SF_IB
+ pixel_5287/PIX_OUT pixel_5287/CSA_VREF pixel
Xpixel_5298 pixel_5298/gring pixel_5298/VDD pixel_5298/GND pixel_5298/VREF pixel_5298/ROW_SEL
+ pixel_5298/NB1 pixel_5298/VBIAS pixel_5298/NB2 pixel_5298/AMP_IN pixel_5298/SF_IB
+ pixel_5298/PIX_OUT pixel_5298/CSA_VREF pixel
Xpixel_4531 pixel_4531/gring pixel_4531/VDD pixel_4531/GND pixel_4531/VREF pixel_4531/ROW_SEL
+ pixel_4531/NB1 pixel_4531/VBIAS pixel_4531/NB2 pixel_4531/AMP_IN pixel_4531/SF_IB
+ pixel_4531/PIX_OUT pixel_4531/CSA_VREF pixel
Xpixel_4542 pixel_4542/gring pixel_4542/VDD pixel_4542/GND pixel_4542/VREF pixel_4542/ROW_SEL
+ pixel_4542/NB1 pixel_4542/VBIAS pixel_4542/NB2 pixel_4542/AMP_IN pixel_4542/SF_IB
+ pixel_4542/PIX_OUT pixel_4542/CSA_VREF pixel
Xpixel_4553 pixel_4553/gring pixel_4553/VDD pixel_4553/GND pixel_4553/VREF pixel_4553/ROW_SEL
+ pixel_4553/NB1 pixel_4553/VBIAS pixel_4553/NB2 pixel_4553/AMP_IN pixel_4553/SF_IB
+ pixel_4553/PIX_OUT pixel_4553/CSA_VREF pixel
Xpixel_4564 pixel_4564/gring pixel_4564/VDD pixel_4564/GND pixel_4564/VREF pixel_4564/ROW_SEL
+ pixel_4564/NB1 pixel_4564/VBIAS pixel_4564/NB2 pixel_4564/AMP_IN pixel_4564/SF_IB
+ pixel_4564/PIX_OUT pixel_4564/CSA_VREF pixel
Xpixel_592 pixel_592/gring pixel_592/VDD pixel_592/GND pixel_592/VREF pixel_592/ROW_SEL
+ pixel_592/NB1 pixel_592/VBIAS pixel_592/NB2 pixel_592/AMP_IN pixel_592/SF_IB pixel_592/PIX_OUT
+ pixel_592/CSA_VREF pixel
Xpixel_581 pixel_581/gring pixel_581/VDD pixel_581/GND pixel_581/VREF pixel_581/ROW_SEL
+ pixel_581/NB1 pixel_581/VBIAS pixel_581/NB2 pixel_581/AMP_IN pixel_581/SF_IB pixel_581/PIX_OUT
+ pixel_581/CSA_VREF pixel
Xpixel_570 pixel_570/gring pixel_570/VDD pixel_570/GND pixel_570/VREF pixel_570/ROW_SEL
+ pixel_570/NB1 pixel_570/VBIAS pixel_570/NB2 pixel_570/AMP_IN pixel_570/SF_IB pixel_570/PIX_OUT
+ pixel_570/CSA_VREF pixel
Xpixel_3852 pixel_3852/gring pixel_3852/VDD pixel_3852/GND pixel_3852/VREF pixel_3852/ROW_SEL
+ pixel_3852/NB1 pixel_3852/VBIAS pixel_3852/NB2 pixel_3852/AMP_IN pixel_3852/SF_IB
+ pixel_3852/PIX_OUT pixel_3852/CSA_VREF pixel
Xpixel_4575 pixel_4575/gring pixel_4575/VDD pixel_4575/GND pixel_4575/VREF pixel_4575/ROW_SEL
+ pixel_4575/NB1 pixel_4575/VBIAS pixel_4575/NB2 pixel_4575/AMP_IN pixel_4575/SF_IB
+ pixel_4575/PIX_OUT pixel_4575/CSA_VREF pixel
Xpixel_4586 pixel_4586/gring pixel_4586/VDD pixel_4586/GND pixel_4586/VREF pixel_4586/ROW_SEL
+ pixel_4586/NB1 pixel_4586/VBIAS pixel_4586/NB2 pixel_4586/AMP_IN pixel_4586/SF_IB
+ pixel_4586/PIX_OUT pixel_4586/CSA_VREF pixel
Xpixel_4597 pixel_4597/gring pixel_4597/VDD pixel_4597/GND pixel_4597/VREF pixel_4597/ROW_SEL
+ pixel_4597/NB1 pixel_4597/VBIAS pixel_4597/NB2 pixel_4597/AMP_IN pixel_4597/SF_IB
+ pixel_4597/PIX_OUT pixel_4597/CSA_VREF pixel
Xpixel_3830 pixel_3830/gring pixel_3830/VDD pixel_3830/GND pixel_3830/VREF pixel_3830/ROW_SEL
+ pixel_3830/NB1 pixel_3830/VBIAS pixel_3830/NB2 pixel_3830/AMP_IN pixel_3830/SF_IB
+ pixel_3830/PIX_OUT pixel_3830/CSA_VREF pixel
Xpixel_3841 pixel_3841/gring pixel_3841/VDD pixel_3841/GND pixel_3841/VREF pixel_3841/ROW_SEL
+ pixel_3841/NB1 pixel_3841/VBIAS pixel_3841/NB2 pixel_3841/AMP_IN pixel_3841/SF_IB
+ pixel_3841/PIX_OUT pixel_3841/CSA_VREF pixel
Xpixel_3885 pixel_3885/gring pixel_3885/VDD pixel_3885/GND pixel_3885/VREF pixel_3885/ROW_SEL
+ pixel_3885/NB1 pixel_3885/VBIAS pixel_3885/NB2 pixel_3885/AMP_IN pixel_3885/SF_IB
+ pixel_3885/PIX_OUT pixel_3885/CSA_VREF pixel
Xpixel_3874 pixel_3874/gring pixel_3874/VDD pixel_3874/GND pixel_3874/VREF pixel_3874/ROW_SEL
+ pixel_3874/NB1 pixel_3874/VBIAS pixel_3874/NB2 pixel_3874/AMP_IN pixel_3874/SF_IB
+ pixel_3874/PIX_OUT pixel_3874/CSA_VREF pixel
Xpixel_3863 pixel_3863/gring pixel_3863/VDD pixel_3863/GND pixel_3863/VREF pixel_3863/ROW_SEL
+ pixel_3863/NB1 pixel_3863/VBIAS pixel_3863/NB2 pixel_3863/AMP_IN pixel_3863/SF_IB
+ pixel_3863/PIX_OUT pixel_3863/CSA_VREF pixel
Xpixel_3896 pixel_3896/gring pixel_3896/VDD pixel_3896/GND pixel_3896/VREF pixel_3896/ROW_SEL
+ pixel_3896/NB1 pixel_3896/VBIAS pixel_3896/NB2 pixel_3896/AMP_IN pixel_3896/SF_IB
+ pixel_3896/PIX_OUT pixel_3896/CSA_VREF pixel
Xpixel_7190 pixel_7190/gring pixel_7190/VDD pixel_7190/GND pixel_7190/VREF pixel_7190/ROW_SEL
+ pixel_7190/NB1 pixel_7190/VBIAS pixel_7190/NB2 pixel_7190/AMP_IN pixel_7190/SF_IB
+ pixel_7190/PIX_OUT pixel_7190/CSA_VREF pixel
Xpixel_9509 pixel_9509/gring pixel_9509/VDD pixel_9509/GND pixel_9509/VREF pixel_9509/ROW_SEL
+ pixel_9509/NB1 pixel_9509/VBIAS pixel_9509/NB2 pixel_9509/AMP_IN pixel_9509/SF_IB
+ pixel_9509/PIX_OUT pixel_9509/CSA_VREF pixel
Xpixel_8808 pixel_8808/gring pixel_8808/VDD pixel_8808/GND pixel_8808/VREF pixel_8808/ROW_SEL
+ pixel_8808/NB1 pixel_8808/VBIAS pixel_8808/NB2 pixel_8808/AMP_IN pixel_8808/SF_IB
+ pixel_8808/PIX_OUT pixel_8808/CSA_VREF pixel
Xpixel_8819 pixel_8819/gring pixel_8819/VDD pixel_8819/GND pixel_8819/VREF pixel_8819/ROW_SEL
+ pixel_8819/NB1 pixel_8819/VBIAS pixel_8819/NB2 pixel_8819/AMP_IN pixel_8819/SF_IB
+ pixel_8819/PIX_OUT pixel_8819/CSA_VREF pixel
Xpixel_3104 pixel_3104/gring pixel_3104/VDD pixel_3104/GND pixel_3104/VREF pixel_3104/ROW_SEL
+ pixel_3104/NB1 pixel_3104/VBIAS pixel_3104/NB2 pixel_3104/AMP_IN pixel_3104/SF_IB
+ pixel_3104/PIX_OUT pixel_3104/CSA_VREF pixel
Xpixel_2403 pixel_2403/gring pixel_2403/VDD pixel_2403/GND pixel_2403/VREF pixel_2403/ROW_SEL
+ pixel_2403/NB1 pixel_2403/VBIAS pixel_2403/NB2 pixel_2403/AMP_IN pixel_2403/SF_IB
+ pixel_2403/PIX_OUT pixel_2403/CSA_VREF pixel
Xpixel_3148 pixel_3148/gring pixel_3148/VDD pixel_3148/GND pixel_3148/VREF pixel_3148/ROW_SEL
+ pixel_3148/NB1 pixel_3148/VBIAS pixel_3148/NB2 pixel_3148/AMP_IN pixel_3148/SF_IB
+ pixel_3148/PIX_OUT pixel_3148/CSA_VREF pixel
Xpixel_3137 pixel_3137/gring pixel_3137/VDD pixel_3137/GND pixel_3137/VREF pixel_3137/ROW_SEL
+ pixel_3137/NB1 pixel_3137/VBIAS pixel_3137/NB2 pixel_3137/AMP_IN pixel_3137/SF_IB
+ pixel_3137/PIX_OUT pixel_3137/CSA_VREF pixel
Xpixel_3126 pixel_3126/gring pixel_3126/VDD pixel_3126/GND pixel_3126/VREF pixel_3126/ROW_SEL
+ pixel_3126/NB1 pixel_3126/VBIAS pixel_3126/NB2 pixel_3126/AMP_IN pixel_3126/SF_IB
+ pixel_3126/PIX_OUT pixel_3126/CSA_VREF pixel
Xpixel_3115 pixel_3115/gring pixel_3115/VDD pixel_3115/GND pixel_3115/VREF pixel_3115/ROW_SEL
+ pixel_3115/NB1 pixel_3115/VBIAS pixel_3115/NB2 pixel_3115/AMP_IN pixel_3115/SF_IB
+ pixel_3115/PIX_OUT pixel_3115/CSA_VREF pixel
Xpixel_2436 pixel_2436/gring pixel_2436/VDD pixel_2436/GND pixel_2436/VREF pixel_2436/ROW_SEL
+ pixel_2436/NB1 pixel_2436/VBIAS pixel_2436/NB2 pixel_2436/AMP_IN pixel_2436/SF_IB
+ pixel_2436/PIX_OUT pixel_2436/CSA_VREF pixel
Xpixel_2425 pixel_2425/gring pixel_2425/VDD pixel_2425/GND pixel_2425/VREF pixel_2425/ROW_SEL
+ pixel_2425/NB1 pixel_2425/VBIAS pixel_2425/NB2 pixel_2425/AMP_IN pixel_2425/SF_IB
+ pixel_2425/PIX_OUT pixel_2425/CSA_VREF pixel
Xpixel_2414 pixel_2414/gring pixel_2414/VDD pixel_2414/GND pixel_2414/VREF pixel_2414/ROW_SEL
+ pixel_2414/NB1 pixel_2414/VBIAS pixel_2414/NB2 pixel_2414/AMP_IN pixel_2414/SF_IB
+ pixel_2414/PIX_OUT pixel_2414/CSA_VREF pixel
Xpixel_3159 pixel_3159/gring pixel_3159/VDD pixel_3159/GND pixel_3159/VREF pixel_3159/ROW_SEL
+ pixel_3159/NB1 pixel_3159/VBIAS pixel_3159/NB2 pixel_3159/AMP_IN pixel_3159/SF_IB
+ pixel_3159/PIX_OUT pixel_3159/CSA_VREF pixel
Xpixel_1735 pixel_1735/gring pixel_1735/VDD pixel_1735/GND pixel_1735/VREF pixel_1735/ROW_SEL
+ pixel_1735/NB1 pixel_1735/VBIAS pixel_1735/NB2 pixel_1735/AMP_IN pixel_1735/SF_IB
+ pixel_1735/PIX_OUT pixel_1735/CSA_VREF pixel
Xpixel_1724 pixel_1724/gring pixel_1724/VDD pixel_1724/GND pixel_1724/VREF pixel_1724/ROW_SEL
+ pixel_1724/NB1 pixel_1724/VBIAS pixel_1724/NB2 pixel_1724/AMP_IN pixel_1724/SF_IB
+ pixel_1724/PIX_OUT pixel_1724/CSA_VREF pixel
Xpixel_1713 pixel_1713/gring pixel_1713/VDD pixel_1713/GND pixel_1713/VREF pixel_1713/ROW_SEL
+ pixel_1713/NB1 pixel_1713/VBIAS pixel_1713/NB2 pixel_1713/AMP_IN pixel_1713/SF_IB
+ pixel_1713/PIX_OUT pixel_1713/CSA_VREF pixel
Xpixel_1702 pixel_1702/gring pixel_1702/VDD pixel_1702/GND pixel_1702/VREF pixel_1702/ROW_SEL
+ pixel_1702/NB1 pixel_1702/VBIAS pixel_1702/NB2 pixel_1702/AMP_IN pixel_1702/SF_IB
+ pixel_1702/PIX_OUT pixel_1702/CSA_VREF pixel
Xpixel_2469 pixel_2469/gring pixel_2469/VDD pixel_2469/GND pixel_2469/VREF pixel_2469/ROW_SEL
+ pixel_2469/NB1 pixel_2469/VBIAS pixel_2469/NB2 pixel_2469/AMP_IN pixel_2469/SF_IB
+ pixel_2469/PIX_OUT pixel_2469/CSA_VREF pixel
Xpixel_2458 pixel_2458/gring pixel_2458/VDD pixel_2458/GND pixel_2458/VREF pixel_2458/ROW_SEL
+ pixel_2458/NB1 pixel_2458/VBIAS pixel_2458/NB2 pixel_2458/AMP_IN pixel_2458/SF_IB
+ pixel_2458/PIX_OUT pixel_2458/CSA_VREF pixel
Xpixel_2447 pixel_2447/gring pixel_2447/VDD pixel_2447/GND pixel_2447/VREF pixel_2447/ROW_SEL
+ pixel_2447/NB1 pixel_2447/VBIAS pixel_2447/NB2 pixel_2447/AMP_IN pixel_2447/SF_IB
+ pixel_2447/PIX_OUT pixel_2447/CSA_VREF pixel
Xpixel_1768 pixel_1768/gring pixel_1768/VDD pixel_1768/GND pixel_1768/VREF pixel_1768/ROW_SEL
+ pixel_1768/NB1 pixel_1768/VBIAS pixel_1768/NB2 pixel_1768/AMP_IN pixel_1768/SF_IB
+ pixel_1768/PIX_OUT pixel_1768/CSA_VREF pixel
Xpixel_1757 pixel_1757/gring pixel_1757/VDD pixel_1757/GND pixel_1757/VREF pixel_1757/ROW_SEL
+ pixel_1757/NB1 pixel_1757/VBIAS pixel_1757/NB2 pixel_1757/AMP_IN pixel_1757/SF_IB
+ pixel_1757/PIX_OUT pixel_1757/CSA_VREF pixel
Xpixel_1746 pixel_1746/gring pixel_1746/VDD pixel_1746/GND pixel_1746/VREF pixel_1746/ROW_SEL
+ pixel_1746/NB1 pixel_1746/VBIAS pixel_1746/NB2 pixel_1746/AMP_IN pixel_1746/SF_IB
+ pixel_1746/PIX_OUT pixel_1746/CSA_VREF pixel
Xpixel_1779 pixel_1779/gring pixel_1779/VDD pixel_1779/GND pixel_1779/VREF pixel_1779/ROW_SEL
+ pixel_1779/NB1 pixel_1779/VBIAS pixel_1779/NB2 pixel_1779/AMP_IN pixel_1779/SF_IB
+ pixel_1779/PIX_OUT pixel_1779/CSA_VREF pixel
Xpixel_5040 pixel_5040/gring pixel_5040/VDD pixel_5040/GND pixel_5040/VREF pixel_5040/ROW_SEL
+ pixel_5040/NB1 pixel_5040/VBIAS pixel_5040/NB2 pixel_5040/AMP_IN pixel_5040/SF_IB
+ pixel_5040/PIX_OUT pixel_5040/CSA_VREF pixel
Xpixel_5051 pixel_5051/gring pixel_5051/VDD pixel_5051/GND pixel_5051/VREF pixel_5051/ROW_SEL
+ pixel_5051/NB1 pixel_5051/VBIAS pixel_5051/NB2 pixel_5051/AMP_IN pixel_5051/SF_IB
+ pixel_5051/PIX_OUT pixel_5051/CSA_VREF pixel
Xpixel_5062 pixel_5062/gring pixel_5062/VDD pixel_5062/GND pixel_5062/VREF pixel_5062/ROW_SEL
+ pixel_5062/NB1 pixel_5062/VBIAS pixel_5062/NB2 pixel_5062/AMP_IN pixel_5062/SF_IB
+ pixel_5062/PIX_OUT pixel_5062/CSA_VREF pixel
Xpixel_5073 pixel_5073/gring pixel_5073/VDD pixel_5073/GND pixel_5073/VREF pixel_5073/ROW_SEL
+ pixel_5073/NB1 pixel_5073/VBIAS pixel_5073/NB2 pixel_5073/AMP_IN pixel_5073/SF_IB
+ pixel_5073/PIX_OUT pixel_5073/CSA_VREF pixel
Xpixel_5084 pixel_5084/gring pixel_5084/VDD pixel_5084/GND pixel_5084/VREF pixel_5084/ROW_SEL
+ pixel_5084/NB1 pixel_5084/VBIAS pixel_5084/NB2 pixel_5084/AMP_IN pixel_5084/SF_IB
+ pixel_5084/PIX_OUT pixel_5084/CSA_VREF pixel
Xpixel_5095 pixel_5095/gring pixel_5095/VDD pixel_5095/GND pixel_5095/VREF pixel_5095/ROW_SEL
+ pixel_5095/NB1 pixel_5095/VBIAS pixel_5095/NB2 pixel_5095/AMP_IN pixel_5095/SF_IB
+ pixel_5095/PIX_OUT pixel_5095/CSA_VREF pixel
Xpixel_4350 pixel_4350/gring pixel_4350/VDD pixel_4350/GND pixel_4350/VREF pixel_4350/ROW_SEL
+ pixel_4350/NB1 pixel_4350/VBIAS pixel_4350/NB2 pixel_4350/AMP_IN pixel_4350/SF_IB
+ pixel_4350/PIX_OUT pixel_4350/CSA_VREF pixel
Xpixel_4361 pixel_4361/gring pixel_4361/VDD pixel_4361/GND pixel_4361/VREF pixel_4361/ROW_SEL
+ pixel_4361/NB1 pixel_4361/VBIAS pixel_4361/NB2 pixel_4361/AMP_IN pixel_4361/SF_IB
+ pixel_4361/PIX_OUT pixel_4361/CSA_VREF pixel
Xpixel_4372 pixel_4372/gring pixel_4372/VDD pixel_4372/GND pixel_4372/VREF pixel_4372/ROW_SEL
+ pixel_4372/NB1 pixel_4372/VBIAS pixel_4372/NB2 pixel_4372/AMP_IN pixel_4372/SF_IB
+ pixel_4372/PIX_OUT pixel_4372/CSA_VREF pixel
Xpixel_3660 pixel_3660/gring pixel_3660/VDD pixel_3660/GND pixel_3660/VREF pixel_3660/ROW_SEL
+ pixel_3660/NB1 pixel_3660/VBIAS pixel_3660/NB2 pixel_3660/AMP_IN pixel_3660/SF_IB
+ pixel_3660/PIX_OUT pixel_3660/CSA_VREF pixel
Xpixel_4383 pixel_4383/gring pixel_4383/VDD pixel_4383/GND pixel_4383/VREF pixel_4383/ROW_SEL
+ pixel_4383/NB1 pixel_4383/VBIAS pixel_4383/NB2 pixel_4383/AMP_IN pixel_4383/SF_IB
+ pixel_4383/PIX_OUT pixel_4383/CSA_VREF pixel
Xpixel_4394 pixel_4394/gring pixel_4394/VDD pixel_4394/GND pixel_4394/VREF pixel_4394/ROW_SEL
+ pixel_4394/NB1 pixel_4394/VBIAS pixel_4394/NB2 pixel_4394/AMP_IN pixel_4394/SF_IB
+ pixel_4394/PIX_OUT pixel_4394/CSA_VREF pixel
Xpixel_3693 pixel_3693/gring pixel_3693/VDD pixel_3693/GND pixel_3693/VREF pixel_3693/ROW_SEL
+ pixel_3693/NB1 pixel_3693/VBIAS pixel_3693/NB2 pixel_3693/AMP_IN pixel_3693/SF_IB
+ pixel_3693/PIX_OUT pixel_3693/CSA_VREF pixel
Xpixel_3682 pixel_3682/gring pixel_3682/VDD pixel_3682/GND pixel_3682/VREF pixel_3682/ROW_SEL
+ pixel_3682/NB1 pixel_3682/VBIAS pixel_3682/NB2 pixel_3682/AMP_IN pixel_3682/SF_IB
+ pixel_3682/PIX_OUT pixel_3682/CSA_VREF pixel
Xpixel_3671 pixel_3671/gring pixel_3671/VDD pixel_3671/GND pixel_3671/VREF pixel_3671/ROW_SEL
+ pixel_3671/NB1 pixel_3671/VBIAS pixel_3671/NB2 pixel_3671/AMP_IN pixel_3671/SF_IB
+ pixel_3671/PIX_OUT pixel_3671/CSA_VREF pixel
Xpixel_2992 pixel_2992/gring pixel_2992/VDD pixel_2992/GND pixel_2992/VREF pixel_2992/ROW_SEL
+ pixel_2992/NB1 pixel_2992/VBIAS pixel_2992/NB2 pixel_2992/AMP_IN pixel_2992/SF_IB
+ pixel_2992/PIX_OUT pixel_2992/CSA_VREF pixel
Xpixel_2981 pixel_2981/gring pixel_2981/VDD pixel_2981/GND pixel_2981/VREF pixel_2981/ROW_SEL
+ pixel_2981/NB1 pixel_2981/VBIAS pixel_2981/NB2 pixel_2981/AMP_IN pixel_2981/SF_IB
+ pixel_2981/PIX_OUT pixel_2981/CSA_VREF pixel
Xpixel_2970 pixel_2970/gring pixel_2970/VDD pixel_2970/GND pixel_2970/VREF pixel_2970/ROW_SEL
+ pixel_2970/NB1 pixel_2970/VBIAS pixel_2970/NB2 pixel_2970/AMP_IN pixel_2970/SF_IB
+ pixel_2970/PIX_OUT pixel_2970/CSA_VREF pixel
Xpixel_1009 pixel_1009/gring pixel_1009/VDD pixel_1009/GND pixel_1009/VREF pixel_1009/ROW_SEL
+ pixel_1009/NB1 pixel_1009/VBIAS pixel_1009/NB2 pixel_1009/AMP_IN pixel_1009/SF_IB
+ pixel_1009/PIX_OUT pixel_1009/CSA_VREF pixel
Xpixel_9328 pixel_9328/gring pixel_9328/VDD pixel_9328/GND pixel_9328/VREF pixel_9328/ROW_SEL
+ pixel_9328/NB1 pixel_9328/VBIAS pixel_9328/NB2 pixel_9328/AMP_IN pixel_9328/SF_IB
+ pixel_9328/PIX_OUT pixel_9328/CSA_VREF pixel
Xpixel_9317 pixel_9317/gring pixel_9317/VDD pixel_9317/GND pixel_9317/VREF pixel_9317/ROW_SEL
+ pixel_9317/NB1 pixel_9317/VBIAS pixel_9317/NB2 pixel_9317/AMP_IN pixel_9317/SF_IB
+ pixel_9317/PIX_OUT pixel_9317/CSA_VREF pixel
Xpixel_9306 pixel_9306/gring pixel_9306/VDD pixel_9306/GND pixel_9306/VREF pixel_9306/ROW_SEL
+ pixel_9306/NB1 pixel_9306/VBIAS pixel_9306/NB2 pixel_9306/AMP_IN pixel_9306/SF_IB
+ pixel_9306/PIX_OUT pixel_9306/CSA_VREF pixel
Xpixel_8627 pixel_8627/gring pixel_8627/VDD pixel_8627/GND pixel_8627/VREF pixel_8627/ROW_SEL
+ pixel_8627/NB1 pixel_8627/VBIAS pixel_8627/NB2 pixel_8627/AMP_IN pixel_8627/SF_IB
+ pixel_8627/PIX_OUT pixel_8627/CSA_VREF pixel
Xpixel_8616 pixel_8616/gring pixel_8616/VDD pixel_8616/GND pixel_8616/VREF pixel_8616/ROW_SEL
+ pixel_8616/NB1 pixel_8616/VBIAS pixel_8616/NB2 pixel_8616/AMP_IN pixel_8616/SF_IB
+ pixel_8616/PIX_OUT pixel_8616/CSA_VREF pixel
Xpixel_8605 pixel_8605/gring pixel_8605/VDD pixel_8605/GND pixel_8605/VREF pixel_8605/ROW_SEL
+ pixel_8605/NB1 pixel_8605/VBIAS pixel_8605/NB2 pixel_8605/AMP_IN pixel_8605/SF_IB
+ pixel_8605/PIX_OUT pixel_8605/CSA_VREF pixel
Xpixel_9339 pixel_9339/gring pixel_9339/VDD pixel_9339/GND pixel_9339/VREF pixel_9339/ROW_SEL
+ pixel_9339/NB1 pixel_9339/VBIAS pixel_9339/NB2 pixel_9339/AMP_IN pixel_9339/SF_IB
+ pixel_9339/PIX_OUT pixel_9339/CSA_VREF pixel
Xpixel_8649 pixel_8649/gring pixel_8649/VDD pixel_8649/GND pixel_8649/VREF pixel_8649/ROW_SEL
+ pixel_8649/NB1 pixel_8649/VBIAS pixel_8649/NB2 pixel_8649/AMP_IN pixel_8649/SF_IB
+ pixel_8649/PIX_OUT pixel_8649/CSA_VREF pixel
Xpixel_8638 pixel_8638/gring pixel_8638/VDD pixel_8638/GND pixel_8638/VREF pixel_8638/ROW_SEL
+ pixel_8638/NB1 pixel_8638/VBIAS pixel_8638/NB2 pixel_8638/AMP_IN pixel_8638/SF_IB
+ pixel_8638/PIX_OUT pixel_8638/CSA_VREF pixel
Xpixel_7904 pixel_7904/gring pixel_7904/VDD pixel_7904/GND pixel_7904/VREF pixel_7904/ROW_SEL
+ pixel_7904/NB1 pixel_7904/VBIAS pixel_7904/NB2 pixel_7904/AMP_IN pixel_7904/SF_IB
+ pixel_7904/PIX_OUT pixel_7904/CSA_VREF pixel
Xpixel_7915 pixel_7915/gring pixel_7915/VDD pixel_7915/GND pixel_7915/VREF pixel_7915/ROW_SEL
+ pixel_7915/NB1 pixel_7915/VBIAS pixel_7915/NB2 pixel_7915/AMP_IN pixel_7915/SF_IB
+ pixel_7915/PIX_OUT pixel_7915/CSA_VREF pixel
Xpixel_7926 pixel_7926/gring pixel_7926/VDD pixel_7926/GND pixel_7926/VREF pixel_7926/ROW_SEL
+ pixel_7926/NB1 pixel_7926/VBIAS pixel_7926/NB2 pixel_7926/AMP_IN pixel_7926/SF_IB
+ pixel_7926/PIX_OUT pixel_7926/CSA_VREF pixel
Xpixel_7937 pixel_7937/gring pixel_7937/VDD pixel_7937/GND pixel_7937/VREF pixel_7937/ROW_SEL
+ pixel_7937/NB1 pixel_7937/VBIAS pixel_7937/NB2 pixel_7937/AMP_IN pixel_7937/SF_IB
+ pixel_7937/PIX_OUT pixel_7937/CSA_VREF pixel
Xpixel_7948 pixel_7948/gring pixel_7948/VDD pixel_7948/GND pixel_7948/VREF pixel_7948/ROW_SEL
+ pixel_7948/NB1 pixel_7948/VBIAS pixel_7948/NB2 pixel_7948/AMP_IN pixel_7948/SF_IB
+ pixel_7948/PIX_OUT pixel_7948/CSA_VREF pixel
Xpixel_7959 pixel_7959/gring pixel_7959/VDD pixel_7959/GND pixel_7959/VREF pixel_7959/ROW_SEL
+ pixel_7959/NB1 pixel_7959/VBIAS pixel_7959/NB2 pixel_7959/AMP_IN pixel_7959/SF_IB
+ pixel_7959/PIX_OUT pixel_7959/CSA_VREF pixel
Xpixel_2211 pixel_2211/gring pixel_2211/VDD pixel_2211/GND pixel_2211/VREF pixel_2211/ROW_SEL
+ pixel_2211/NB1 pixel_2211/VBIAS pixel_2211/NB2 pixel_2211/AMP_IN pixel_2211/SF_IB
+ pixel_2211/PIX_OUT pixel_2211/CSA_VREF pixel
Xpixel_2200 pixel_2200/gring pixel_2200/VDD pixel_2200/GND pixel_2200/VREF pixel_2200/ROW_SEL
+ pixel_2200/NB1 pixel_2200/VBIAS pixel_2200/NB2 pixel_2200/AMP_IN pixel_2200/SF_IB
+ pixel_2200/PIX_OUT pixel_2200/CSA_VREF pixel
Xpixel_1510 pixel_1510/gring pixel_1510/VDD pixel_1510/GND pixel_1510/VREF pixel_1510/ROW_SEL
+ pixel_1510/NB1 pixel_1510/VBIAS pixel_1510/NB2 pixel_1510/AMP_IN pixel_1510/SF_IB
+ pixel_1510/PIX_OUT pixel_1510/CSA_VREF pixel
Xpixel_2244 pixel_2244/gring pixel_2244/VDD pixel_2244/GND pixel_2244/VREF pixel_2244/ROW_SEL
+ pixel_2244/NB1 pixel_2244/VBIAS pixel_2244/NB2 pixel_2244/AMP_IN pixel_2244/SF_IB
+ pixel_2244/PIX_OUT pixel_2244/CSA_VREF pixel
Xpixel_2233 pixel_2233/gring pixel_2233/VDD pixel_2233/GND pixel_2233/VREF pixel_2233/ROW_SEL
+ pixel_2233/NB1 pixel_2233/VBIAS pixel_2233/NB2 pixel_2233/AMP_IN pixel_2233/SF_IB
+ pixel_2233/PIX_OUT pixel_2233/CSA_VREF pixel
Xpixel_2222 pixel_2222/gring pixel_2222/VDD pixel_2222/GND pixel_2222/VREF pixel_2222/ROW_SEL
+ pixel_2222/NB1 pixel_2222/VBIAS pixel_2222/NB2 pixel_2222/AMP_IN pixel_2222/SF_IB
+ pixel_2222/PIX_OUT pixel_2222/CSA_VREF pixel
Xpixel_1543 pixel_1543/gring pixel_1543/VDD pixel_1543/GND pixel_1543/VREF pixel_1543/ROW_SEL
+ pixel_1543/NB1 pixel_1543/VBIAS pixel_1543/NB2 pixel_1543/AMP_IN pixel_1543/SF_IB
+ pixel_1543/PIX_OUT pixel_1543/CSA_VREF pixel
Xpixel_1532 pixel_1532/gring pixel_1532/VDD pixel_1532/GND pixel_1532/VREF pixel_1532/ROW_SEL
+ pixel_1532/NB1 pixel_1532/VBIAS pixel_1532/NB2 pixel_1532/AMP_IN pixel_1532/SF_IB
+ pixel_1532/PIX_OUT pixel_1532/CSA_VREF pixel
Xpixel_1521 pixel_1521/gring pixel_1521/VDD pixel_1521/GND pixel_1521/VREF pixel_1521/ROW_SEL
+ pixel_1521/NB1 pixel_1521/VBIAS pixel_1521/NB2 pixel_1521/AMP_IN pixel_1521/SF_IB
+ pixel_1521/PIX_OUT pixel_1521/CSA_VREF pixel
Xpixel_2288 pixel_2288/gring pixel_2288/VDD pixel_2288/GND pixel_2288/VREF pixel_2288/ROW_SEL
+ pixel_2288/NB1 pixel_2288/VBIAS pixel_2288/NB2 pixel_2288/AMP_IN pixel_2288/SF_IB
+ pixel_2288/PIX_OUT pixel_2288/CSA_VREF pixel
Xpixel_2277 pixel_2277/gring pixel_2277/VDD pixel_2277/GND pixel_2277/VREF pixel_2277/ROW_SEL
+ pixel_2277/NB1 pixel_2277/VBIAS pixel_2277/NB2 pixel_2277/AMP_IN pixel_2277/SF_IB
+ pixel_2277/PIX_OUT pixel_2277/CSA_VREF pixel
Xpixel_2266 pixel_2266/gring pixel_2266/VDD pixel_2266/GND pixel_2266/VREF pixel_2266/ROW_SEL
+ pixel_2266/NB1 pixel_2266/VBIAS pixel_2266/NB2 pixel_2266/AMP_IN pixel_2266/SF_IB
+ pixel_2266/PIX_OUT pixel_2266/CSA_VREF pixel
Xpixel_2255 pixel_2255/gring pixel_2255/VDD pixel_2255/GND pixel_2255/VREF pixel_2255/ROW_SEL
+ pixel_2255/NB1 pixel_2255/VBIAS pixel_2255/NB2 pixel_2255/AMP_IN pixel_2255/SF_IB
+ pixel_2255/PIX_OUT pixel_2255/CSA_VREF pixel
Xpixel_1576 pixel_1576/gring pixel_1576/VDD pixel_1576/GND pixel_1576/VREF pixel_1576/ROW_SEL
+ pixel_1576/NB1 pixel_1576/VBIAS pixel_1576/NB2 pixel_1576/AMP_IN pixel_1576/SF_IB
+ pixel_1576/PIX_OUT pixel_1576/CSA_VREF pixel
Xpixel_1565 pixel_1565/gring pixel_1565/VDD pixel_1565/GND pixel_1565/VREF pixel_1565/ROW_SEL
+ pixel_1565/NB1 pixel_1565/VBIAS pixel_1565/NB2 pixel_1565/AMP_IN pixel_1565/SF_IB
+ pixel_1565/PIX_OUT pixel_1565/CSA_VREF pixel
Xpixel_1554 pixel_1554/gring pixel_1554/VDD pixel_1554/GND pixel_1554/VREF pixel_1554/ROW_SEL
+ pixel_1554/NB1 pixel_1554/VBIAS pixel_1554/NB2 pixel_1554/AMP_IN pixel_1554/SF_IB
+ pixel_1554/PIX_OUT pixel_1554/CSA_VREF pixel
Xpixel_2299 pixel_2299/gring pixel_2299/VDD pixel_2299/GND pixel_2299/VREF pixel_2299/ROW_SEL
+ pixel_2299/NB1 pixel_2299/VBIAS pixel_2299/NB2 pixel_2299/AMP_IN pixel_2299/SF_IB
+ pixel_2299/PIX_OUT pixel_2299/CSA_VREF pixel
Xpixel_1598 pixel_1598/gring pixel_1598/VDD pixel_1598/GND pixel_1598/VREF pixel_1598/ROW_SEL
+ pixel_1598/NB1 pixel_1598/VBIAS pixel_1598/NB2 pixel_1598/AMP_IN pixel_1598/SF_IB
+ pixel_1598/PIX_OUT pixel_1598/CSA_VREF pixel
Xpixel_1587 pixel_1587/gring pixel_1587/VDD pixel_1587/GND pixel_1587/VREF pixel_1587/ROW_SEL
+ pixel_1587/NB1 pixel_1587/VBIAS pixel_1587/NB2 pixel_1587/AMP_IN pixel_1587/SF_IB
+ pixel_1587/PIX_OUT pixel_1587/CSA_VREF pixel
Xpixel_9840 pixel_9840/gring pixel_9840/VDD pixel_9840/GND pixel_9840/VREF pixel_9840/ROW_SEL
+ pixel_9840/NB1 pixel_9840/VBIAS pixel_9840/NB2 pixel_9840/AMP_IN pixel_9840/SF_IB
+ pixel_9840/PIX_OUT pixel_9840/CSA_VREF pixel
Xpixel_9851 pixel_9851/gring pixel_9851/VDD pixel_9851/GND pixel_9851/VREF pixel_9851/ROW_SEL
+ pixel_9851/NB1 pixel_9851/VBIAS pixel_9851/NB2 pixel_9851/AMP_IN pixel_9851/SF_IB
+ pixel_9851/PIX_OUT pixel_9851/CSA_VREF pixel
Xpixel_9862 pixel_9862/gring pixel_9862/VDD pixel_9862/GND pixel_9862/VREF pixel_9862/ROW_SEL
+ pixel_9862/NB1 pixel_9862/VBIAS pixel_9862/NB2 pixel_9862/AMP_IN pixel_9862/SF_IB
+ pixel_9862/PIX_OUT pixel_9862/CSA_VREF pixel
Xpixel_9873 pixel_9873/gring pixel_9873/VDD pixel_9873/GND pixel_9873/VREF pixel_9873/ROW_SEL
+ pixel_9873/NB1 pixel_9873/VBIAS pixel_9873/NB2 pixel_9873/AMP_IN pixel_9873/SF_IB
+ pixel_9873/PIX_OUT pixel_9873/CSA_VREF pixel
Xpixel_9884 pixel_9884/gring pixel_9884/VDD pixel_9884/GND pixel_9884/VREF pixel_9884/ROW_SEL
+ pixel_9884/NB1 pixel_9884/VBIAS pixel_9884/NB2 pixel_9884/AMP_IN pixel_9884/SF_IB
+ pixel_9884/PIX_OUT pixel_9884/CSA_VREF pixel
Xpixel_9895 pixel_9895/gring pixel_9895/VDD pixel_9895/GND pixel_9895/VREF pixel_9895/ROW_SEL
+ pixel_9895/NB1 pixel_9895/VBIAS pixel_9895/NB2 pixel_9895/AMP_IN pixel_9895/SF_IB
+ pixel_9895/PIX_OUT pixel_9895/CSA_VREF pixel
Xpixel_4180 pixel_4180/gring pixel_4180/VDD pixel_4180/GND pixel_4180/VREF pixel_4180/ROW_SEL
+ pixel_4180/NB1 pixel_4180/VBIAS pixel_4180/NB2 pixel_4180/AMP_IN pixel_4180/SF_IB
+ pixel_4180/PIX_OUT pixel_4180/CSA_VREF pixel
Xpixel_4191 pixel_4191/gring pixel_4191/VDD pixel_4191/GND pixel_4191/VREF pixel_4191/ROW_SEL
+ pixel_4191/NB1 pixel_4191/VBIAS pixel_4191/NB2 pixel_4191/AMP_IN pixel_4191/SF_IB
+ pixel_4191/PIX_OUT pixel_4191/CSA_VREF pixel
Xpixel_3490 pixel_3490/gring pixel_3490/VDD pixel_3490/GND pixel_3490/VREF pixel_3490/ROW_SEL
+ pixel_3490/NB1 pixel_3490/VBIAS pixel_3490/NB2 pixel_3490/AMP_IN pixel_3490/SF_IB
+ pixel_3490/PIX_OUT pixel_3490/CSA_VREF pixel
Xpixel_5809 pixel_5809/gring pixel_5809/VDD pixel_5809/GND pixel_5809/VREF pixel_5809/ROW_SEL
+ pixel_5809/NB1 pixel_5809/VBIAS pixel_5809/NB2 pixel_5809/AMP_IN pixel_5809/SF_IB
+ pixel_5809/PIX_OUT pixel_5809/CSA_VREF pixel
Xpixel_9103 pixel_9103/gring pixel_9103/VDD pixel_9103/GND pixel_9103/VREF pixel_9103/ROW_SEL
+ pixel_9103/NB1 pixel_9103/VBIAS pixel_9103/NB2 pixel_9103/AMP_IN pixel_9103/SF_IB
+ pixel_9103/PIX_OUT pixel_9103/CSA_VREF pixel
Xpixel_8402 pixel_8402/gring pixel_8402/VDD pixel_8402/GND pixel_8402/VREF pixel_8402/ROW_SEL
+ pixel_8402/NB1 pixel_8402/VBIAS pixel_8402/NB2 pixel_8402/AMP_IN pixel_8402/SF_IB
+ pixel_8402/PIX_OUT pixel_8402/CSA_VREF pixel
Xpixel_9136 pixel_9136/gring pixel_9136/VDD pixel_9136/GND pixel_9136/VREF pixel_9136/ROW_SEL
+ pixel_9136/NB1 pixel_9136/VBIAS pixel_9136/NB2 pixel_9136/AMP_IN pixel_9136/SF_IB
+ pixel_9136/PIX_OUT pixel_9136/CSA_VREF pixel
Xpixel_9125 pixel_9125/gring pixel_9125/VDD pixel_9125/GND pixel_9125/VREF pixel_9125/ROW_SEL
+ pixel_9125/NB1 pixel_9125/VBIAS pixel_9125/NB2 pixel_9125/AMP_IN pixel_9125/SF_IB
+ pixel_9125/PIX_OUT pixel_9125/CSA_VREF pixel
Xpixel_9114 pixel_9114/gring pixel_9114/VDD pixel_9114/GND pixel_9114/VREF pixel_9114/ROW_SEL
+ pixel_9114/NB1 pixel_9114/VBIAS pixel_9114/NB2 pixel_9114/AMP_IN pixel_9114/SF_IB
+ pixel_9114/PIX_OUT pixel_9114/CSA_VREF pixel
Xpixel_8435 pixel_8435/gring pixel_8435/VDD pixel_8435/GND pixel_8435/VREF pixel_8435/ROW_SEL
+ pixel_8435/NB1 pixel_8435/VBIAS pixel_8435/NB2 pixel_8435/AMP_IN pixel_8435/SF_IB
+ pixel_8435/PIX_OUT pixel_8435/CSA_VREF pixel
Xpixel_8424 pixel_8424/gring pixel_8424/VDD pixel_8424/GND pixel_8424/VREF pixel_8424/ROW_SEL
+ pixel_8424/NB1 pixel_8424/VBIAS pixel_8424/NB2 pixel_8424/AMP_IN pixel_8424/SF_IB
+ pixel_8424/PIX_OUT pixel_8424/CSA_VREF pixel
Xpixel_8413 pixel_8413/gring pixel_8413/VDD pixel_8413/GND pixel_8413/VREF pixel_8413/ROW_SEL
+ pixel_8413/NB1 pixel_8413/VBIAS pixel_8413/NB2 pixel_8413/AMP_IN pixel_8413/SF_IB
+ pixel_8413/PIX_OUT pixel_8413/CSA_VREF pixel
Xpixel_9169 pixel_9169/gring pixel_9169/VDD pixel_9169/GND pixel_9169/VREF pixel_9169/ROW_SEL
+ pixel_9169/NB1 pixel_9169/VBIAS pixel_9169/NB2 pixel_9169/AMP_IN pixel_9169/SF_IB
+ pixel_9169/PIX_OUT pixel_9169/CSA_VREF pixel
Xpixel_9158 pixel_9158/gring pixel_9158/VDD pixel_9158/GND pixel_9158/VREF pixel_9158/ROW_SEL
+ pixel_9158/NB1 pixel_9158/VBIAS pixel_9158/NB2 pixel_9158/AMP_IN pixel_9158/SF_IB
+ pixel_9158/PIX_OUT pixel_9158/CSA_VREF pixel
Xpixel_9147 pixel_9147/gring pixel_9147/VDD pixel_9147/GND pixel_9147/VREF pixel_9147/ROW_SEL
+ pixel_9147/NB1 pixel_9147/VBIAS pixel_9147/NB2 pixel_9147/AMP_IN pixel_9147/SF_IB
+ pixel_9147/PIX_OUT pixel_9147/CSA_VREF pixel
Xpixel_8446 pixel_8446/gring pixel_8446/VDD pixel_8446/GND pixel_8446/VREF pixel_8446/ROW_SEL
+ pixel_8446/NB1 pixel_8446/VBIAS pixel_8446/NB2 pixel_8446/AMP_IN pixel_8446/SF_IB
+ pixel_8446/PIX_OUT pixel_8446/CSA_VREF pixel
Xpixel_8457 pixel_8457/gring pixel_8457/VDD pixel_8457/GND pixel_8457/VREF pixel_8457/ROW_SEL
+ pixel_8457/NB1 pixel_8457/VBIAS pixel_8457/NB2 pixel_8457/AMP_IN pixel_8457/SF_IB
+ pixel_8457/PIX_OUT pixel_8457/CSA_VREF pixel
Xpixel_8468 pixel_8468/gring pixel_8468/VDD pixel_8468/GND pixel_8468/VREF pixel_8468/ROW_SEL
+ pixel_8468/NB1 pixel_8468/VBIAS pixel_8468/NB2 pixel_8468/AMP_IN pixel_8468/SF_IB
+ pixel_8468/PIX_OUT pixel_8468/CSA_VREF pixel
Xpixel_7701 pixel_7701/gring pixel_7701/VDD pixel_7701/GND pixel_7701/VREF pixel_7701/ROW_SEL
+ pixel_7701/NB1 pixel_7701/VBIAS pixel_7701/NB2 pixel_7701/AMP_IN pixel_7701/SF_IB
+ pixel_7701/PIX_OUT pixel_7701/CSA_VREF pixel
Xpixel_7712 pixel_7712/gring pixel_7712/VDD pixel_7712/GND pixel_7712/VREF pixel_7712/ROW_SEL
+ pixel_7712/NB1 pixel_7712/VBIAS pixel_7712/NB2 pixel_7712/AMP_IN pixel_7712/SF_IB
+ pixel_7712/PIX_OUT pixel_7712/CSA_VREF pixel
Xpixel_7723 pixel_7723/gring pixel_7723/VDD pixel_7723/GND pixel_7723/VREF pixel_7723/ROW_SEL
+ pixel_7723/NB1 pixel_7723/VBIAS pixel_7723/NB2 pixel_7723/AMP_IN pixel_7723/SF_IB
+ pixel_7723/PIX_OUT pixel_7723/CSA_VREF pixel
Xpixel_8479 pixel_8479/gring pixel_8479/VDD pixel_8479/GND pixel_8479/VREF pixel_8479/ROW_SEL
+ pixel_8479/NB1 pixel_8479/VBIAS pixel_8479/NB2 pixel_8479/AMP_IN pixel_8479/SF_IB
+ pixel_8479/PIX_OUT pixel_8479/CSA_VREF pixel
Xpixel_7734 pixel_7734/gring pixel_7734/VDD pixel_7734/GND pixel_7734/VREF pixel_7734/ROW_SEL
+ pixel_7734/NB1 pixel_7734/VBIAS pixel_7734/NB2 pixel_7734/AMP_IN pixel_7734/SF_IB
+ pixel_7734/PIX_OUT pixel_7734/CSA_VREF pixel
Xpixel_7745 pixel_7745/gring pixel_7745/VDD pixel_7745/GND pixel_7745/VREF pixel_7745/ROW_SEL
+ pixel_7745/NB1 pixel_7745/VBIAS pixel_7745/NB2 pixel_7745/AMP_IN pixel_7745/SF_IB
+ pixel_7745/PIX_OUT pixel_7745/CSA_VREF pixel
Xpixel_7756 pixel_7756/gring pixel_7756/VDD pixel_7756/GND pixel_7756/VREF pixel_7756/ROW_SEL
+ pixel_7756/NB1 pixel_7756/VBIAS pixel_7756/NB2 pixel_7756/AMP_IN pixel_7756/SF_IB
+ pixel_7756/PIX_OUT pixel_7756/CSA_VREF pixel
Xpixel_7767 pixel_7767/gring pixel_7767/VDD pixel_7767/GND pixel_7767/VREF pixel_7767/ROW_SEL
+ pixel_7767/NB1 pixel_7767/VBIAS pixel_7767/NB2 pixel_7767/AMP_IN pixel_7767/SF_IB
+ pixel_7767/PIX_OUT pixel_7767/CSA_VREF pixel
Xpixel_7778 pixel_7778/gring pixel_7778/VDD pixel_7778/GND pixel_7778/VREF pixel_7778/ROW_SEL
+ pixel_7778/NB1 pixel_7778/VBIAS pixel_7778/NB2 pixel_7778/AMP_IN pixel_7778/SF_IB
+ pixel_7778/PIX_OUT pixel_7778/CSA_VREF pixel
Xpixel_7789 pixel_7789/gring pixel_7789/VDD pixel_7789/GND pixel_7789/VREF pixel_7789/ROW_SEL
+ pixel_7789/NB1 pixel_7789/VBIAS pixel_7789/NB2 pixel_7789/AMP_IN pixel_7789/SF_IB
+ pixel_7789/PIX_OUT pixel_7789/CSA_VREF pixel
Xpixel_2063 pixel_2063/gring pixel_2063/VDD pixel_2063/GND pixel_2063/VREF pixel_2063/ROW_SEL
+ pixel_2063/NB1 pixel_2063/VBIAS pixel_2063/NB2 pixel_2063/AMP_IN pixel_2063/SF_IB
+ pixel_2063/PIX_OUT pixel_2063/CSA_VREF pixel
Xpixel_2052 pixel_2052/gring pixel_2052/VDD pixel_2052/GND pixel_2052/VREF pixel_2052/ROW_SEL
+ pixel_2052/NB1 pixel_2052/VBIAS pixel_2052/NB2 pixel_2052/AMP_IN pixel_2052/SF_IB
+ pixel_2052/PIX_OUT pixel_2052/CSA_VREF pixel
Xpixel_2041 pixel_2041/gring pixel_2041/VDD pixel_2041/GND pixel_2041/VREF pixel_2041/ROW_SEL
+ pixel_2041/NB1 pixel_2041/VBIAS pixel_2041/NB2 pixel_2041/AMP_IN pixel_2041/SF_IB
+ pixel_2041/PIX_OUT pixel_2041/CSA_VREF pixel
Xpixel_2030 pixel_2030/gring pixel_2030/VDD pixel_2030/GND pixel_2030/VREF pixel_2030/ROW_SEL
+ pixel_2030/NB1 pixel_2030/VBIAS pixel_2030/NB2 pixel_2030/AMP_IN pixel_2030/SF_IB
+ pixel_2030/PIX_OUT pixel_2030/CSA_VREF pixel
Xpixel_1351 pixel_1351/gring pixel_1351/VDD pixel_1351/GND pixel_1351/VREF pixel_1351/ROW_SEL
+ pixel_1351/NB1 pixel_1351/VBIAS pixel_1351/NB2 pixel_1351/AMP_IN pixel_1351/SF_IB
+ pixel_1351/PIX_OUT pixel_1351/CSA_VREF pixel
Xpixel_1340 pixel_1340/gring pixel_1340/VDD pixel_1340/GND pixel_1340/VREF pixel_1340/ROW_SEL
+ pixel_1340/NB1 pixel_1340/VBIAS pixel_1340/NB2 pixel_1340/AMP_IN pixel_1340/SF_IB
+ pixel_1340/PIX_OUT pixel_1340/CSA_VREF pixel
Xpixel_2096 pixel_2096/gring pixel_2096/VDD pixel_2096/GND pixel_2096/VREF pixel_2096/ROW_SEL
+ pixel_2096/NB1 pixel_2096/VBIAS pixel_2096/NB2 pixel_2096/AMP_IN pixel_2096/SF_IB
+ pixel_2096/PIX_OUT pixel_2096/CSA_VREF pixel
Xpixel_2085 pixel_2085/gring pixel_2085/VDD pixel_2085/GND pixel_2085/VREF pixel_2085/ROW_SEL
+ pixel_2085/NB1 pixel_2085/VBIAS pixel_2085/NB2 pixel_2085/AMP_IN pixel_2085/SF_IB
+ pixel_2085/PIX_OUT pixel_2085/CSA_VREF pixel
Xpixel_2074 pixel_2074/gring pixel_2074/VDD pixel_2074/GND pixel_2074/VREF pixel_2074/ROW_SEL
+ pixel_2074/NB1 pixel_2074/VBIAS pixel_2074/NB2 pixel_2074/AMP_IN pixel_2074/SF_IB
+ pixel_2074/PIX_OUT pixel_2074/CSA_VREF pixel
Xpixel_1384 pixel_1384/gring pixel_1384/VDD pixel_1384/GND pixel_1384/VREF pixel_1384/ROW_SEL
+ pixel_1384/NB1 pixel_1384/VBIAS pixel_1384/NB2 pixel_1384/AMP_IN pixel_1384/SF_IB
+ pixel_1384/PIX_OUT pixel_1384/CSA_VREF pixel
Xpixel_1373 pixel_1373/gring pixel_1373/VDD pixel_1373/GND pixel_1373/VREF pixel_1373/ROW_SEL
+ pixel_1373/NB1 pixel_1373/VBIAS pixel_1373/NB2 pixel_1373/AMP_IN pixel_1373/SF_IB
+ pixel_1373/PIX_OUT pixel_1373/CSA_VREF pixel
Xpixel_1362 pixel_1362/gring pixel_1362/VDD pixel_1362/GND pixel_1362/VREF pixel_1362/ROW_SEL
+ pixel_1362/NB1 pixel_1362/VBIAS pixel_1362/NB2 pixel_1362/AMP_IN pixel_1362/SF_IB
+ pixel_1362/PIX_OUT pixel_1362/CSA_VREF pixel
Xpixel_1395 pixel_1395/gring pixel_1395/VDD pixel_1395/GND pixel_1395/VREF pixel_1395/ROW_SEL
+ pixel_1395/NB1 pixel_1395/VBIAS pixel_1395/NB2 pixel_1395/AMP_IN pixel_1395/SF_IB
+ pixel_1395/PIX_OUT pixel_1395/CSA_VREF pixel
Xpixel_9692 pixel_9692/gring pixel_9692/VDD pixel_9692/GND pixel_9692/VREF pixel_9692/ROW_SEL
+ pixel_9692/NB1 pixel_9692/VBIAS pixel_9692/NB2 pixel_9692/AMP_IN pixel_9692/SF_IB
+ pixel_9692/PIX_OUT pixel_9692/CSA_VREF pixel
Xpixel_9670 pixel_9670/gring pixel_9670/VDD pixel_9670/GND pixel_9670/VREF pixel_9670/ROW_SEL
+ pixel_9670/NB1 pixel_9670/VBIAS pixel_9670/NB2 pixel_9670/AMP_IN pixel_9670/SF_IB
+ pixel_9670/PIX_OUT pixel_9670/CSA_VREF pixel
Xpixel_9681 pixel_9681/gring pixel_9681/VDD pixel_9681/GND pixel_9681/VREF pixel_9681/ROW_SEL
+ pixel_9681/NB1 pixel_9681/VBIAS pixel_9681/NB2 pixel_9681/AMP_IN pixel_9681/SF_IB
+ pixel_9681/PIX_OUT pixel_9681/CSA_VREF pixel
Xpixel_8991 pixel_8991/gring pixel_8991/VDD pixel_8991/GND pixel_8991/VREF pixel_8991/ROW_SEL
+ pixel_8991/NB1 pixel_8991/VBIAS pixel_8991/NB2 pixel_8991/AMP_IN pixel_8991/SF_IB
+ pixel_8991/PIX_OUT pixel_8991/CSA_VREF pixel
Xpixel_8980 pixel_8980/gring pixel_8980/VDD pixel_8980/GND pixel_8980/VREF pixel_8980/ROW_SEL
+ pixel_8980/NB1 pixel_8980/VBIAS pixel_8980/NB2 pixel_8980/AMP_IN pixel_8980/SF_IB
+ pixel_8980/PIX_OUT pixel_8980/CSA_VREF pixel
Xpixel_7008 pixel_7008/gring pixel_7008/VDD pixel_7008/GND pixel_7008/VREF pixel_7008/ROW_SEL
+ pixel_7008/NB1 pixel_7008/VBIAS pixel_7008/NB2 pixel_7008/AMP_IN pixel_7008/SF_IB
+ pixel_7008/PIX_OUT pixel_7008/CSA_VREF pixel
Xpixel_7019 pixel_7019/gring pixel_7019/VDD pixel_7019/GND pixel_7019/VREF pixel_7019/ROW_SEL
+ pixel_7019/NB1 pixel_7019/VBIAS pixel_7019/NB2 pixel_7019/AMP_IN pixel_7019/SF_IB
+ pixel_7019/PIX_OUT pixel_7019/CSA_VREF pixel
Xpixel_6307 pixel_6307/gring pixel_6307/VDD pixel_6307/GND pixel_6307/VREF pixel_6307/ROW_SEL
+ pixel_6307/NB1 pixel_6307/VBIAS pixel_6307/NB2 pixel_6307/AMP_IN pixel_6307/SF_IB
+ pixel_6307/PIX_OUT pixel_6307/CSA_VREF pixel
Xpixel_6318 pixel_6318/gring pixel_6318/VDD pixel_6318/GND pixel_6318/VREF pixel_6318/ROW_SEL
+ pixel_6318/NB1 pixel_6318/VBIAS pixel_6318/NB2 pixel_6318/AMP_IN pixel_6318/SF_IB
+ pixel_6318/PIX_OUT pixel_6318/CSA_VREF pixel
Xpixel_6329 pixel_6329/gring pixel_6329/VDD pixel_6329/GND pixel_6329/VREF pixel_6329/ROW_SEL
+ pixel_6329/NB1 pixel_6329/VBIAS pixel_6329/NB2 pixel_6329/AMP_IN pixel_6329/SF_IB
+ pixel_6329/PIX_OUT pixel_6329/CSA_VREF pixel
Xpixel_5606 pixel_5606/gring pixel_5606/VDD pixel_5606/GND pixel_5606/VREF pixel_5606/ROW_SEL
+ pixel_5606/NB1 pixel_5606/VBIAS pixel_5606/NB2 pixel_5606/AMP_IN pixel_5606/SF_IB
+ pixel_5606/PIX_OUT pixel_5606/CSA_VREF pixel
Xpixel_900 pixel_900/gring pixel_900/VDD pixel_900/GND pixel_900/VREF pixel_900/ROW_SEL
+ pixel_900/NB1 pixel_900/VBIAS pixel_900/NB2 pixel_900/AMP_IN pixel_900/SF_IB pixel_900/PIX_OUT
+ pixel_900/CSA_VREF pixel
Xpixel_5617 pixel_5617/gring pixel_5617/VDD pixel_5617/GND pixel_5617/VREF pixel_5617/ROW_SEL
+ pixel_5617/NB1 pixel_5617/VBIAS pixel_5617/NB2 pixel_5617/AMP_IN pixel_5617/SF_IB
+ pixel_5617/PIX_OUT pixel_5617/CSA_VREF pixel
Xpixel_5628 pixel_5628/gring pixel_5628/VDD pixel_5628/GND pixel_5628/VREF pixel_5628/ROW_SEL
+ pixel_5628/NB1 pixel_5628/VBIAS pixel_5628/NB2 pixel_5628/AMP_IN pixel_5628/SF_IB
+ pixel_5628/PIX_OUT pixel_5628/CSA_VREF pixel
Xpixel_5639 pixel_5639/gring pixel_5639/VDD pixel_5639/GND pixel_5639/VREF pixel_5639/ROW_SEL
+ pixel_5639/NB1 pixel_5639/VBIAS pixel_5639/NB2 pixel_5639/AMP_IN pixel_5639/SF_IB
+ pixel_5639/PIX_OUT pixel_5639/CSA_VREF pixel
Xpixel_933 pixel_933/gring pixel_933/VDD pixel_933/GND pixel_933/VREF pixel_933/ROW_SEL
+ pixel_933/NB1 pixel_933/VBIAS pixel_933/NB2 pixel_933/AMP_IN pixel_933/SF_IB pixel_933/PIX_OUT
+ pixel_933/CSA_VREF pixel
Xpixel_922 pixel_922/gring pixel_922/VDD pixel_922/GND pixel_922/VREF pixel_922/ROW_SEL
+ pixel_922/NB1 pixel_922/VBIAS pixel_922/NB2 pixel_922/AMP_IN pixel_922/SF_IB pixel_922/PIX_OUT
+ pixel_922/CSA_VREF pixel
Xpixel_911 pixel_911/gring pixel_911/VDD pixel_911/GND pixel_911/VREF pixel_911/ROW_SEL
+ pixel_911/NB1 pixel_911/VBIAS pixel_911/NB2 pixel_911/AMP_IN pixel_911/SF_IB pixel_911/PIX_OUT
+ pixel_911/CSA_VREF pixel
Xpixel_4905 pixel_4905/gring pixel_4905/VDD pixel_4905/GND pixel_4905/VREF pixel_4905/ROW_SEL
+ pixel_4905/NB1 pixel_4905/VBIAS pixel_4905/NB2 pixel_4905/AMP_IN pixel_4905/SF_IB
+ pixel_4905/PIX_OUT pixel_4905/CSA_VREF pixel
Xpixel_4916 pixel_4916/gring pixel_4916/VDD pixel_4916/GND pixel_4916/VREF pixel_4916/ROW_SEL
+ pixel_4916/NB1 pixel_4916/VBIAS pixel_4916/NB2 pixel_4916/AMP_IN pixel_4916/SF_IB
+ pixel_4916/PIX_OUT pixel_4916/CSA_VREF pixel
Xpixel_4927 pixel_4927/gring pixel_4927/VDD pixel_4927/GND pixel_4927/VREF pixel_4927/ROW_SEL
+ pixel_4927/NB1 pixel_4927/VBIAS pixel_4927/NB2 pixel_4927/AMP_IN pixel_4927/SF_IB
+ pixel_4927/PIX_OUT pixel_4927/CSA_VREF pixel
Xpixel_4938 pixel_4938/gring pixel_4938/VDD pixel_4938/GND pixel_4938/VREF pixel_4938/ROW_SEL
+ pixel_4938/NB1 pixel_4938/VBIAS pixel_4938/NB2 pixel_4938/AMP_IN pixel_4938/SF_IB
+ pixel_4938/PIX_OUT pixel_4938/CSA_VREF pixel
Xpixel_966 pixel_966/gring pixel_966/VDD pixel_966/GND pixel_966/VREF pixel_966/ROW_SEL
+ pixel_966/NB1 pixel_966/VBIAS pixel_966/NB2 pixel_966/AMP_IN pixel_966/SF_IB pixel_966/PIX_OUT
+ pixel_966/CSA_VREF pixel
Xpixel_955 pixel_955/gring pixel_955/VDD pixel_955/GND pixel_955/VREF pixel_955/ROW_SEL
+ pixel_955/NB1 pixel_955/VBIAS pixel_955/NB2 pixel_955/AMP_IN pixel_955/SF_IB pixel_955/PIX_OUT
+ pixel_955/CSA_VREF pixel
Xpixel_944 pixel_944/gring pixel_944/VDD pixel_944/GND pixel_944/VREF pixel_944/ROW_SEL
+ pixel_944/NB1 pixel_944/VBIAS pixel_944/NB2 pixel_944/AMP_IN pixel_944/SF_IB pixel_944/PIX_OUT
+ pixel_944/CSA_VREF pixel
Xpixel_4949 pixel_4949/gring pixel_4949/VDD pixel_4949/GND pixel_4949/VREF pixel_4949/ROW_SEL
+ pixel_4949/NB1 pixel_4949/VBIAS pixel_4949/NB2 pixel_4949/AMP_IN pixel_4949/SF_IB
+ pixel_4949/PIX_OUT pixel_4949/CSA_VREF pixel
Xpixel_999 pixel_999/gring pixel_999/VDD pixel_999/GND pixel_999/VREF pixel_999/ROW_SEL
+ pixel_999/NB1 pixel_999/VBIAS pixel_999/NB2 pixel_999/AMP_IN pixel_999/SF_IB pixel_999/PIX_OUT
+ pixel_999/CSA_VREF pixel
Xpixel_988 pixel_988/gring pixel_988/VDD pixel_988/GND pixel_988/VREF pixel_988/ROW_SEL
+ pixel_988/NB1 pixel_988/VBIAS pixel_988/NB2 pixel_988/AMP_IN pixel_988/SF_IB pixel_988/PIX_OUT
+ pixel_988/CSA_VREF pixel
Xpixel_977 pixel_977/gring pixel_977/VDD pixel_977/GND pixel_977/VREF pixel_977/ROW_SEL
+ pixel_977/NB1 pixel_977/VBIAS pixel_977/NB2 pixel_977/AMP_IN pixel_977/SF_IB pixel_977/PIX_OUT
+ pixel_977/CSA_VREF pixel
Xpixel_8210 pixel_8210/gring pixel_8210/VDD pixel_8210/GND pixel_8210/VREF pixel_8210/ROW_SEL
+ pixel_8210/NB1 pixel_8210/VBIAS pixel_8210/NB2 pixel_8210/AMP_IN pixel_8210/SF_IB
+ pixel_8210/PIX_OUT pixel_8210/CSA_VREF pixel
Xpixel_8221 pixel_8221/gring pixel_8221/VDD pixel_8221/GND pixel_8221/VREF pixel_8221/ROW_SEL
+ pixel_8221/NB1 pixel_8221/VBIAS pixel_8221/NB2 pixel_8221/AMP_IN pixel_8221/SF_IB
+ pixel_8221/PIX_OUT pixel_8221/CSA_VREF pixel
Xpixel_8232 pixel_8232/gring pixel_8232/VDD pixel_8232/GND pixel_8232/VREF pixel_8232/ROW_SEL
+ pixel_8232/NB1 pixel_8232/VBIAS pixel_8232/NB2 pixel_8232/AMP_IN pixel_8232/SF_IB
+ pixel_8232/PIX_OUT pixel_8232/CSA_VREF pixel
Xpixel_8243 pixel_8243/gring pixel_8243/VDD pixel_8243/GND pixel_8243/VREF pixel_8243/ROW_SEL
+ pixel_8243/NB1 pixel_8243/VBIAS pixel_8243/NB2 pixel_8243/AMP_IN pixel_8243/SF_IB
+ pixel_8243/PIX_OUT pixel_8243/CSA_VREF pixel
Xpixel_8254 pixel_8254/gring pixel_8254/VDD pixel_8254/GND pixel_8254/VREF pixel_8254/ROW_SEL
+ pixel_8254/NB1 pixel_8254/VBIAS pixel_8254/NB2 pixel_8254/AMP_IN pixel_8254/SF_IB
+ pixel_8254/PIX_OUT pixel_8254/CSA_VREF pixel
Xpixel_8265 pixel_8265/gring pixel_8265/VDD pixel_8265/GND pixel_8265/VREF pixel_8265/ROW_SEL
+ pixel_8265/NB1 pixel_8265/VBIAS pixel_8265/NB2 pixel_8265/AMP_IN pixel_8265/SF_IB
+ pixel_8265/PIX_OUT pixel_8265/CSA_VREF pixel
Xpixel_8276 pixel_8276/gring pixel_8276/VDD pixel_8276/GND pixel_8276/VREF pixel_8276/ROW_SEL
+ pixel_8276/NB1 pixel_8276/VBIAS pixel_8276/NB2 pixel_8276/AMP_IN pixel_8276/SF_IB
+ pixel_8276/PIX_OUT pixel_8276/CSA_VREF pixel
Xpixel_7520 pixel_7520/gring pixel_7520/VDD pixel_7520/GND pixel_7520/VREF pixel_7520/ROW_SEL
+ pixel_7520/NB1 pixel_7520/VBIAS pixel_7520/NB2 pixel_7520/AMP_IN pixel_7520/SF_IB
+ pixel_7520/PIX_OUT pixel_7520/CSA_VREF pixel
Xpixel_7531 pixel_7531/gring pixel_7531/VDD pixel_7531/GND pixel_7531/VREF pixel_7531/ROW_SEL
+ pixel_7531/NB1 pixel_7531/VBIAS pixel_7531/NB2 pixel_7531/AMP_IN pixel_7531/SF_IB
+ pixel_7531/PIX_OUT pixel_7531/CSA_VREF pixel
Xpixel_7542 pixel_7542/gring pixel_7542/VDD pixel_7542/GND pixel_7542/VREF pixel_7542/ROW_SEL
+ pixel_7542/NB1 pixel_7542/VBIAS pixel_7542/NB2 pixel_7542/AMP_IN pixel_7542/SF_IB
+ pixel_7542/PIX_OUT pixel_7542/CSA_VREF pixel
Xpixel_8287 pixel_8287/gring pixel_8287/VDD pixel_8287/GND pixel_8287/VREF pixel_8287/ROW_SEL
+ pixel_8287/NB1 pixel_8287/VBIAS pixel_8287/NB2 pixel_8287/AMP_IN pixel_8287/SF_IB
+ pixel_8287/PIX_OUT pixel_8287/CSA_VREF pixel
Xpixel_8298 pixel_8298/gring pixel_8298/VDD pixel_8298/GND pixel_8298/VREF pixel_8298/ROW_SEL
+ pixel_8298/NB1 pixel_8298/VBIAS pixel_8298/NB2 pixel_8298/AMP_IN pixel_8298/SF_IB
+ pixel_8298/PIX_OUT pixel_8298/CSA_VREF pixel
Xpixel_7553 pixel_7553/gring pixel_7553/VDD pixel_7553/GND pixel_7553/VREF pixel_7553/ROW_SEL
+ pixel_7553/NB1 pixel_7553/VBIAS pixel_7553/NB2 pixel_7553/AMP_IN pixel_7553/SF_IB
+ pixel_7553/PIX_OUT pixel_7553/CSA_VREF pixel
Xpixel_7564 pixel_7564/gring pixel_7564/VDD pixel_7564/GND pixel_7564/VREF pixel_7564/ROW_SEL
+ pixel_7564/NB1 pixel_7564/VBIAS pixel_7564/NB2 pixel_7564/AMP_IN pixel_7564/SF_IB
+ pixel_7564/PIX_OUT pixel_7564/CSA_VREF pixel
Xpixel_7575 pixel_7575/gring pixel_7575/VDD pixel_7575/GND pixel_7575/VREF pixel_7575/ROW_SEL
+ pixel_7575/NB1 pixel_7575/VBIAS pixel_7575/NB2 pixel_7575/AMP_IN pixel_7575/SF_IB
+ pixel_7575/PIX_OUT pixel_7575/CSA_VREF pixel
Xpixel_6830 pixel_6830/gring pixel_6830/VDD pixel_6830/GND pixel_6830/VREF pixel_6830/ROW_SEL
+ pixel_6830/NB1 pixel_6830/VBIAS pixel_6830/NB2 pixel_6830/AMP_IN pixel_6830/SF_IB
+ pixel_6830/PIX_OUT pixel_6830/CSA_VREF pixel
Xpixel_7586 pixel_7586/gring pixel_7586/VDD pixel_7586/GND pixel_7586/VREF pixel_7586/ROW_SEL
+ pixel_7586/NB1 pixel_7586/VBIAS pixel_7586/NB2 pixel_7586/AMP_IN pixel_7586/SF_IB
+ pixel_7586/PIX_OUT pixel_7586/CSA_VREF pixel
Xpixel_7597 pixel_7597/gring pixel_7597/VDD pixel_7597/GND pixel_7597/VREF pixel_7597/ROW_SEL
+ pixel_7597/NB1 pixel_7597/VBIAS pixel_7597/NB2 pixel_7597/AMP_IN pixel_7597/SF_IB
+ pixel_7597/PIX_OUT pixel_7597/CSA_VREF pixel
Xpixel_6841 pixel_6841/gring pixel_6841/VDD pixel_6841/GND pixel_6841/VREF pixel_6841/ROW_SEL
+ pixel_6841/NB1 pixel_6841/VBIAS pixel_6841/NB2 pixel_6841/AMP_IN pixel_6841/SF_IB
+ pixel_6841/PIX_OUT pixel_6841/CSA_VREF pixel
Xpixel_6852 pixel_6852/gring pixel_6852/VDD pixel_6852/GND pixel_6852/VREF pixel_6852/ROW_SEL
+ pixel_6852/NB1 pixel_6852/VBIAS pixel_6852/NB2 pixel_6852/AMP_IN pixel_6852/SF_IB
+ pixel_6852/PIX_OUT pixel_6852/CSA_VREF pixel
Xpixel_6863 pixel_6863/gring pixel_6863/VDD pixel_6863/GND pixel_6863/VREF pixel_6863/ROW_SEL
+ pixel_6863/NB1 pixel_6863/VBIAS pixel_6863/NB2 pixel_6863/AMP_IN pixel_6863/SF_IB
+ pixel_6863/PIX_OUT pixel_6863/CSA_VREF pixel
Xpixel_6874 pixel_6874/gring pixel_6874/VDD pixel_6874/GND pixel_6874/VREF pixel_6874/ROW_SEL
+ pixel_6874/NB1 pixel_6874/VBIAS pixel_6874/NB2 pixel_6874/AMP_IN pixel_6874/SF_IB
+ pixel_6874/PIX_OUT pixel_6874/CSA_VREF pixel
Xpixel_6885 pixel_6885/gring pixel_6885/VDD pixel_6885/GND pixel_6885/VREF pixel_6885/ROW_SEL
+ pixel_6885/NB1 pixel_6885/VBIAS pixel_6885/NB2 pixel_6885/AMP_IN pixel_6885/SF_IB
+ pixel_6885/PIX_OUT pixel_6885/CSA_VREF pixel
Xpixel_6896 pixel_6896/gring pixel_6896/VDD pixel_6896/GND pixel_6896/VREF pixel_6896/ROW_SEL
+ pixel_6896/NB1 pixel_6896/VBIAS pixel_6896/NB2 pixel_6896/AMP_IN pixel_6896/SF_IB
+ pixel_6896/PIX_OUT pixel_6896/CSA_VREF pixel
Xpixel_1192 pixel_1192/gring pixel_1192/VDD pixel_1192/GND pixel_1192/VREF pixel_1192/ROW_SEL
+ pixel_1192/NB1 pixel_1192/VBIAS pixel_1192/NB2 pixel_1192/AMP_IN pixel_1192/SF_IB
+ pixel_1192/PIX_OUT pixel_1192/CSA_VREF pixel
Xpixel_1181 pixel_1181/gring pixel_1181/VDD pixel_1181/GND pixel_1181/VREF pixel_1181/ROW_SEL
+ pixel_1181/NB1 pixel_1181/VBIAS pixel_1181/NB2 pixel_1181/AMP_IN pixel_1181/SF_IB
+ pixel_1181/PIX_OUT pixel_1181/CSA_VREF pixel
Xpixel_1170 pixel_1170/gring pixel_1170/VDD pixel_1170/GND pixel_1170/VREF pixel_1170/ROW_SEL
+ pixel_1170/NB1 pixel_1170/VBIAS pixel_1170/NB2 pixel_1170/AMP_IN pixel_1170/SF_IB
+ pixel_1170/PIX_OUT pixel_1170/CSA_VREF pixel
Xpixel_229 pixel_229/gring pixel_229/VDD pixel_229/GND pixel_229/VREF pixel_229/ROW_SEL
+ pixel_229/NB1 pixel_229/VBIAS pixel_229/NB2 pixel_229/AMP_IN pixel_229/SF_IB pixel_229/PIX_OUT
+ pixel_229/CSA_VREF pixel
Xpixel_218 pixel_218/gring pixel_218/VDD pixel_218/GND pixel_218/VREF pixel_218/ROW_SEL
+ pixel_218/NB1 pixel_218/VBIAS pixel_218/NB2 pixel_218/AMP_IN pixel_218/SF_IB pixel_218/PIX_OUT
+ pixel_218/CSA_VREF pixel
Xpixel_207 pixel_207/gring pixel_207/VDD pixel_207/GND pixel_207/VREF pixel_207/ROW_SEL
+ pixel_207/NB1 pixel_207/VBIAS pixel_207/NB2 pixel_207/AMP_IN pixel_207/SF_IB pixel_207/PIX_OUT
+ pixel_207/CSA_VREF pixel
Xpixel_6104 pixel_6104/gring pixel_6104/VDD pixel_6104/GND pixel_6104/VREF pixel_6104/ROW_SEL
+ pixel_6104/NB1 pixel_6104/VBIAS pixel_6104/NB2 pixel_6104/AMP_IN pixel_6104/SF_IB
+ pixel_6104/PIX_OUT pixel_6104/CSA_VREF pixel
Xpixel_6115 pixel_6115/gring pixel_6115/VDD pixel_6115/GND pixel_6115/VREF pixel_6115/ROW_SEL
+ pixel_6115/NB1 pixel_6115/VBIAS pixel_6115/NB2 pixel_6115/AMP_IN pixel_6115/SF_IB
+ pixel_6115/PIX_OUT pixel_6115/CSA_VREF pixel
Xpixel_6126 pixel_6126/gring pixel_6126/VDD pixel_6126/GND pixel_6126/VREF pixel_6126/ROW_SEL
+ pixel_6126/NB1 pixel_6126/VBIAS pixel_6126/NB2 pixel_6126/AMP_IN pixel_6126/SF_IB
+ pixel_6126/PIX_OUT pixel_6126/CSA_VREF pixel
Xpixel_6137 pixel_6137/gring pixel_6137/VDD pixel_6137/GND pixel_6137/VREF pixel_6137/ROW_SEL
+ pixel_6137/NB1 pixel_6137/VBIAS pixel_6137/NB2 pixel_6137/AMP_IN pixel_6137/SF_IB
+ pixel_6137/PIX_OUT pixel_6137/CSA_VREF pixel
Xpixel_6148 pixel_6148/gring pixel_6148/VDD pixel_6148/GND pixel_6148/VREF pixel_6148/ROW_SEL
+ pixel_6148/NB1 pixel_6148/VBIAS pixel_6148/NB2 pixel_6148/AMP_IN pixel_6148/SF_IB
+ pixel_6148/PIX_OUT pixel_6148/CSA_VREF pixel
Xpixel_6159 pixel_6159/gring pixel_6159/VDD pixel_6159/GND pixel_6159/VREF pixel_6159/ROW_SEL
+ pixel_6159/NB1 pixel_6159/VBIAS pixel_6159/NB2 pixel_6159/AMP_IN pixel_6159/SF_IB
+ pixel_6159/PIX_OUT pixel_6159/CSA_VREF pixel
Xpixel_5403 pixel_5403/gring pixel_5403/VDD pixel_5403/GND pixel_5403/VREF pixel_5403/ROW_SEL
+ pixel_5403/NB1 pixel_5403/VBIAS pixel_5403/NB2 pixel_5403/AMP_IN pixel_5403/SF_IB
+ pixel_5403/PIX_OUT pixel_5403/CSA_VREF pixel
Xpixel_5414 pixel_5414/gring pixel_5414/VDD pixel_5414/GND pixel_5414/VREF pixel_5414/ROW_SEL
+ pixel_5414/NB1 pixel_5414/VBIAS pixel_5414/NB2 pixel_5414/AMP_IN pixel_5414/SF_IB
+ pixel_5414/PIX_OUT pixel_5414/CSA_VREF pixel
Xpixel_5425 pixel_5425/gring pixel_5425/VDD pixel_5425/GND pixel_5425/VREF pixel_5425/ROW_SEL
+ pixel_5425/NB1 pixel_5425/VBIAS pixel_5425/NB2 pixel_5425/AMP_IN pixel_5425/SF_IB
+ pixel_5425/PIX_OUT pixel_5425/CSA_VREF pixel
Xpixel_5436 pixel_5436/gring pixel_5436/VDD pixel_5436/GND pixel_5436/VREF pixel_5436/ROW_SEL
+ pixel_5436/NB1 pixel_5436/VBIAS pixel_5436/NB2 pixel_5436/AMP_IN pixel_5436/SF_IB
+ pixel_5436/PIX_OUT pixel_5436/CSA_VREF pixel
Xpixel_5447 pixel_5447/gring pixel_5447/VDD pixel_5447/GND pixel_5447/VREF pixel_5447/ROW_SEL
+ pixel_5447/NB1 pixel_5447/VBIAS pixel_5447/NB2 pixel_5447/AMP_IN pixel_5447/SF_IB
+ pixel_5447/PIX_OUT pixel_5447/CSA_VREF pixel
Xpixel_4702 pixel_4702/gring pixel_4702/VDD pixel_4702/GND pixel_4702/VREF pixel_4702/ROW_SEL
+ pixel_4702/NB1 pixel_4702/VBIAS pixel_4702/NB2 pixel_4702/AMP_IN pixel_4702/SF_IB
+ pixel_4702/PIX_OUT pixel_4702/CSA_VREF pixel
Xpixel_4713 pixel_4713/gring pixel_4713/VDD pixel_4713/GND pixel_4713/VREF pixel_4713/ROW_SEL
+ pixel_4713/NB1 pixel_4713/VBIAS pixel_4713/NB2 pixel_4713/AMP_IN pixel_4713/SF_IB
+ pixel_4713/PIX_OUT pixel_4713/CSA_VREF pixel
Xpixel_741 pixel_741/gring pixel_741/VDD pixel_741/GND pixel_741/VREF pixel_741/ROW_SEL
+ pixel_741/NB1 pixel_741/VBIAS pixel_741/NB2 pixel_741/AMP_IN pixel_741/SF_IB pixel_741/PIX_OUT
+ pixel_741/CSA_VREF pixel
Xpixel_730 pixel_730/gring pixel_730/VDD pixel_730/GND pixel_730/VREF pixel_730/ROW_SEL
+ pixel_730/NB1 pixel_730/VBIAS pixel_730/NB2 pixel_730/AMP_IN pixel_730/SF_IB pixel_730/PIX_OUT
+ pixel_730/CSA_VREF pixel
Xpixel_5458 pixel_5458/gring pixel_5458/VDD pixel_5458/GND pixel_5458/VREF pixel_5458/ROW_SEL
+ pixel_5458/NB1 pixel_5458/VBIAS pixel_5458/NB2 pixel_5458/AMP_IN pixel_5458/SF_IB
+ pixel_5458/PIX_OUT pixel_5458/CSA_VREF pixel
Xpixel_5469 pixel_5469/gring pixel_5469/VDD pixel_5469/GND pixel_5469/VREF pixel_5469/ROW_SEL
+ pixel_5469/NB1 pixel_5469/VBIAS pixel_5469/NB2 pixel_5469/AMP_IN pixel_5469/SF_IB
+ pixel_5469/PIX_OUT pixel_5469/CSA_VREF pixel
Xpixel_4724 pixel_4724/gring pixel_4724/VDD pixel_4724/GND pixel_4724/VREF pixel_4724/ROW_SEL
+ pixel_4724/NB1 pixel_4724/VBIAS pixel_4724/NB2 pixel_4724/AMP_IN pixel_4724/SF_IB
+ pixel_4724/PIX_OUT pixel_4724/CSA_VREF pixel
Xpixel_4735 pixel_4735/gring pixel_4735/VDD pixel_4735/GND pixel_4735/VREF pixel_4735/ROW_SEL
+ pixel_4735/NB1 pixel_4735/VBIAS pixel_4735/NB2 pixel_4735/AMP_IN pixel_4735/SF_IB
+ pixel_4735/PIX_OUT pixel_4735/CSA_VREF pixel
Xpixel_4746 pixel_4746/gring pixel_4746/VDD pixel_4746/GND pixel_4746/VREF pixel_4746/ROW_SEL
+ pixel_4746/NB1 pixel_4746/VBIAS pixel_4746/NB2 pixel_4746/AMP_IN pixel_4746/SF_IB
+ pixel_4746/PIX_OUT pixel_4746/CSA_VREF pixel
Xpixel_774 pixel_774/gring pixel_774/VDD pixel_774/GND pixel_774/VREF pixel_774/ROW_SEL
+ pixel_774/NB1 pixel_774/VBIAS pixel_774/NB2 pixel_774/AMP_IN pixel_774/SF_IB pixel_774/PIX_OUT
+ pixel_774/CSA_VREF pixel
Xpixel_763 pixel_763/gring pixel_763/VDD pixel_763/GND pixel_763/VREF pixel_763/ROW_SEL
+ pixel_763/NB1 pixel_763/VBIAS pixel_763/NB2 pixel_763/AMP_IN pixel_763/SF_IB pixel_763/PIX_OUT
+ pixel_763/CSA_VREF pixel
Xpixel_752 pixel_752/gring pixel_752/VDD pixel_752/GND pixel_752/VREF pixel_752/ROW_SEL
+ pixel_752/NB1 pixel_752/VBIAS pixel_752/NB2 pixel_752/AMP_IN pixel_752/SF_IB pixel_752/PIX_OUT
+ pixel_752/CSA_VREF pixel
Xpixel_4757 pixel_4757/gring pixel_4757/VDD pixel_4757/GND pixel_4757/VREF pixel_4757/ROW_SEL
+ pixel_4757/NB1 pixel_4757/VBIAS pixel_4757/NB2 pixel_4757/AMP_IN pixel_4757/SF_IB
+ pixel_4757/PIX_OUT pixel_4757/CSA_VREF pixel
Xpixel_4768 pixel_4768/gring pixel_4768/VDD pixel_4768/GND pixel_4768/VREF pixel_4768/ROW_SEL
+ pixel_4768/NB1 pixel_4768/VBIAS pixel_4768/NB2 pixel_4768/AMP_IN pixel_4768/SF_IB
+ pixel_4768/PIX_OUT pixel_4768/CSA_VREF pixel
Xpixel_4779 pixel_4779/gring pixel_4779/VDD pixel_4779/GND pixel_4779/VREF pixel_4779/ROW_SEL
+ pixel_4779/NB1 pixel_4779/VBIAS pixel_4779/NB2 pixel_4779/AMP_IN pixel_4779/SF_IB
+ pixel_4779/PIX_OUT pixel_4779/CSA_VREF pixel
Xpixel_796 pixel_796/gring pixel_796/VDD pixel_796/GND pixel_796/VREF pixel_796/ROW_SEL
+ pixel_796/NB1 pixel_796/VBIAS pixel_796/NB2 pixel_796/AMP_IN pixel_796/SF_IB pixel_796/PIX_OUT
+ pixel_796/CSA_VREF pixel
Xpixel_785 pixel_785/gring pixel_785/VDD pixel_785/GND pixel_785/VREF pixel_785/ROW_SEL
+ pixel_785/NB1 pixel_785/VBIAS pixel_785/NB2 pixel_785/AMP_IN pixel_785/SF_IB pixel_785/PIX_OUT
+ pixel_785/CSA_VREF pixel
Xpixel_8040 pixel_8040/gring pixel_8040/VDD pixel_8040/GND pixel_8040/VREF pixel_8040/ROW_SEL
+ pixel_8040/NB1 pixel_8040/VBIAS pixel_8040/NB2 pixel_8040/AMP_IN pixel_8040/SF_IB
+ pixel_8040/PIX_OUT pixel_8040/CSA_VREF pixel
Xpixel_8051 pixel_8051/gring pixel_8051/VDD pixel_8051/GND pixel_8051/VREF pixel_8051/ROW_SEL
+ pixel_8051/NB1 pixel_8051/VBIAS pixel_8051/NB2 pixel_8051/AMP_IN pixel_8051/SF_IB
+ pixel_8051/PIX_OUT pixel_8051/CSA_VREF pixel
Xpixel_8062 pixel_8062/gring pixel_8062/VDD pixel_8062/GND pixel_8062/VREF pixel_8062/ROW_SEL
+ pixel_8062/NB1 pixel_8062/VBIAS pixel_8062/NB2 pixel_8062/AMP_IN pixel_8062/SF_IB
+ pixel_8062/PIX_OUT pixel_8062/CSA_VREF pixel
Xpixel_8073 pixel_8073/gring pixel_8073/VDD pixel_8073/GND pixel_8073/VREF pixel_8073/ROW_SEL
+ pixel_8073/NB1 pixel_8073/VBIAS pixel_8073/NB2 pixel_8073/AMP_IN pixel_8073/SF_IB
+ pixel_8073/PIX_OUT pixel_8073/CSA_VREF pixel
Xpixel_8084 pixel_8084/gring pixel_8084/VDD pixel_8084/GND pixel_8084/VREF pixel_8084/ROW_SEL
+ pixel_8084/NB1 pixel_8084/VBIAS pixel_8084/NB2 pixel_8084/AMP_IN pixel_8084/SF_IB
+ pixel_8084/PIX_OUT pixel_8084/CSA_VREF pixel
Xpixel_8095 pixel_8095/gring pixel_8095/VDD pixel_8095/GND pixel_8095/VREF pixel_8095/ROW_SEL
+ pixel_8095/NB1 pixel_8095/VBIAS pixel_8095/NB2 pixel_8095/AMP_IN pixel_8095/SF_IB
+ pixel_8095/PIX_OUT pixel_8095/CSA_VREF pixel
Xpixel_7350 pixel_7350/gring pixel_7350/VDD pixel_7350/GND pixel_7350/VREF pixel_7350/ROW_SEL
+ pixel_7350/NB1 pixel_7350/VBIAS pixel_7350/NB2 pixel_7350/AMP_IN pixel_7350/SF_IB
+ pixel_7350/PIX_OUT pixel_7350/CSA_VREF pixel
Xpixel_7361 pixel_7361/gring pixel_7361/VDD pixel_7361/GND pixel_7361/VREF pixel_7361/ROW_SEL
+ pixel_7361/NB1 pixel_7361/VBIAS pixel_7361/NB2 pixel_7361/AMP_IN pixel_7361/SF_IB
+ pixel_7361/PIX_OUT pixel_7361/CSA_VREF pixel
Xpixel_7372 pixel_7372/gring pixel_7372/VDD pixel_7372/GND pixel_7372/VREF pixel_7372/ROW_SEL
+ pixel_7372/NB1 pixel_7372/VBIAS pixel_7372/NB2 pixel_7372/AMP_IN pixel_7372/SF_IB
+ pixel_7372/PIX_OUT pixel_7372/CSA_VREF pixel
Xpixel_7383 pixel_7383/gring pixel_7383/VDD pixel_7383/GND pixel_7383/VREF pixel_7383/ROW_SEL
+ pixel_7383/NB1 pixel_7383/VBIAS pixel_7383/NB2 pixel_7383/AMP_IN pixel_7383/SF_IB
+ pixel_7383/PIX_OUT pixel_7383/CSA_VREF pixel
Xpixel_7394 pixel_7394/gring pixel_7394/VDD pixel_7394/GND pixel_7394/VREF pixel_7394/ROW_SEL
+ pixel_7394/NB1 pixel_7394/VBIAS pixel_7394/NB2 pixel_7394/AMP_IN pixel_7394/SF_IB
+ pixel_7394/PIX_OUT pixel_7394/CSA_VREF pixel
Xpixel_6660 pixel_6660/gring pixel_6660/VDD pixel_6660/GND pixel_6660/VREF pixel_6660/ROW_SEL
+ pixel_6660/NB1 pixel_6660/VBIAS pixel_6660/NB2 pixel_6660/AMP_IN pixel_6660/SF_IB
+ pixel_6660/PIX_OUT pixel_6660/CSA_VREF pixel
Xpixel_6671 pixel_6671/gring pixel_6671/VDD pixel_6671/GND pixel_6671/VREF pixel_6671/ROW_SEL
+ pixel_6671/NB1 pixel_6671/VBIAS pixel_6671/NB2 pixel_6671/AMP_IN pixel_6671/SF_IB
+ pixel_6671/PIX_OUT pixel_6671/CSA_VREF pixel
Xpixel_6682 pixel_6682/gring pixel_6682/VDD pixel_6682/GND pixel_6682/VREF pixel_6682/ROW_SEL
+ pixel_6682/NB1 pixel_6682/VBIAS pixel_6682/NB2 pixel_6682/AMP_IN pixel_6682/SF_IB
+ pixel_6682/PIX_OUT pixel_6682/CSA_VREF pixel
Xpixel_6693 pixel_6693/gring pixel_6693/VDD pixel_6693/GND pixel_6693/VREF pixel_6693/ROW_SEL
+ pixel_6693/NB1 pixel_6693/VBIAS pixel_6693/NB2 pixel_6693/AMP_IN pixel_6693/SF_IB
+ pixel_6693/PIX_OUT pixel_6693/CSA_VREF pixel
Xpixel_5970 pixel_5970/gring pixel_5970/VDD pixel_5970/GND pixel_5970/VREF pixel_5970/ROW_SEL
+ pixel_5970/NB1 pixel_5970/VBIAS pixel_5970/NB2 pixel_5970/AMP_IN pixel_5970/SF_IB
+ pixel_5970/PIX_OUT pixel_5970/CSA_VREF pixel
Xpixel_5981 pixel_5981/gring pixel_5981/VDD pixel_5981/GND pixel_5981/VREF pixel_5981/ROW_SEL
+ pixel_5981/NB1 pixel_5981/VBIAS pixel_5981/NB2 pixel_5981/AMP_IN pixel_5981/SF_IB
+ pixel_5981/PIX_OUT pixel_5981/CSA_VREF pixel
Xpixel_5992 pixel_5992/gring pixel_5992/VDD pixel_5992/GND pixel_5992/VREF pixel_5992/ROW_SEL
+ pixel_5992/NB1 pixel_5992/VBIAS pixel_5992/NB2 pixel_5992/AMP_IN pixel_5992/SF_IB
+ pixel_5992/PIX_OUT pixel_5992/CSA_VREF pixel
Xpixel_4009 pixel_4009/gring pixel_4009/VDD pixel_4009/GND pixel_4009/VREF pixel_4009/ROW_SEL
+ pixel_4009/NB1 pixel_4009/VBIAS pixel_4009/NB2 pixel_4009/AMP_IN pixel_4009/SF_IB
+ pixel_4009/PIX_OUT pixel_4009/CSA_VREF pixel
Xpixel_3319 pixel_3319/gring pixel_3319/VDD pixel_3319/GND pixel_3319/VREF pixel_3319/ROW_SEL
+ pixel_3319/NB1 pixel_3319/VBIAS pixel_3319/NB2 pixel_3319/AMP_IN pixel_3319/SF_IB
+ pixel_3319/PIX_OUT pixel_3319/CSA_VREF pixel
Xpixel_3308 pixel_3308/gring pixel_3308/VDD pixel_3308/GND pixel_3308/VREF pixel_3308/ROW_SEL
+ pixel_3308/NB1 pixel_3308/VBIAS pixel_3308/NB2 pixel_3308/AMP_IN pixel_3308/SF_IB
+ pixel_3308/PIX_OUT pixel_3308/CSA_VREF pixel
Xpixel_2618 pixel_2618/gring pixel_2618/VDD pixel_2618/GND pixel_2618/VREF pixel_2618/ROW_SEL
+ pixel_2618/NB1 pixel_2618/VBIAS pixel_2618/NB2 pixel_2618/AMP_IN pixel_2618/SF_IB
+ pixel_2618/PIX_OUT pixel_2618/CSA_VREF pixel
Xpixel_2607 pixel_2607/gring pixel_2607/VDD pixel_2607/GND pixel_2607/VREF pixel_2607/ROW_SEL
+ pixel_2607/NB1 pixel_2607/VBIAS pixel_2607/NB2 pixel_2607/AMP_IN pixel_2607/SF_IB
+ pixel_2607/PIX_OUT pixel_2607/CSA_VREF pixel
Xpixel_1917 pixel_1917/gring pixel_1917/VDD pixel_1917/GND pixel_1917/VREF pixel_1917/ROW_SEL
+ pixel_1917/NB1 pixel_1917/VBIAS pixel_1917/NB2 pixel_1917/AMP_IN pixel_1917/SF_IB
+ pixel_1917/PIX_OUT pixel_1917/CSA_VREF pixel
Xpixel_1906 pixel_1906/gring pixel_1906/VDD pixel_1906/GND pixel_1906/VREF pixel_1906/ROW_SEL
+ pixel_1906/NB1 pixel_1906/VBIAS pixel_1906/NB2 pixel_1906/AMP_IN pixel_1906/SF_IB
+ pixel_1906/PIX_OUT pixel_1906/CSA_VREF pixel
Xpixel_2629 pixel_2629/gring pixel_2629/VDD pixel_2629/GND pixel_2629/VREF pixel_2629/ROW_SEL
+ pixel_2629/NB1 pixel_2629/VBIAS pixel_2629/NB2 pixel_2629/AMP_IN pixel_2629/SF_IB
+ pixel_2629/PIX_OUT pixel_2629/CSA_VREF pixel
Xpixel_1939 pixel_1939/gring pixel_1939/VDD pixel_1939/GND pixel_1939/VREF pixel_1939/ROW_SEL
+ pixel_1939/NB1 pixel_1939/VBIAS pixel_1939/NB2 pixel_1939/AMP_IN pixel_1939/SF_IB
+ pixel_1939/PIX_OUT pixel_1939/CSA_VREF pixel
Xpixel_1928 pixel_1928/gring pixel_1928/VDD pixel_1928/GND pixel_1928/VREF pixel_1928/ROW_SEL
+ pixel_1928/NB1 pixel_1928/VBIAS pixel_1928/NB2 pixel_1928/AMP_IN pixel_1928/SF_IB
+ pixel_1928/PIX_OUT pixel_1928/CSA_VREF pixel
Xpixel_5200 pixel_5200/gring pixel_5200/VDD pixel_5200/GND pixel_5200/VREF pixel_5200/ROW_SEL
+ pixel_5200/NB1 pixel_5200/VBIAS pixel_5200/NB2 pixel_5200/AMP_IN pixel_5200/SF_IB
+ pixel_5200/PIX_OUT pixel_5200/CSA_VREF pixel
Xpixel_5211 pixel_5211/gring pixel_5211/VDD pixel_5211/GND pixel_5211/VREF pixel_5211/ROW_SEL
+ pixel_5211/NB1 pixel_5211/VBIAS pixel_5211/NB2 pixel_5211/AMP_IN pixel_5211/SF_IB
+ pixel_5211/PIX_OUT pixel_5211/CSA_VREF pixel
Xpixel_5222 pixel_5222/gring pixel_5222/VDD pixel_5222/GND pixel_5222/VREF pixel_5222/ROW_SEL
+ pixel_5222/NB1 pixel_5222/VBIAS pixel_5222/NB2 pixel_5222/AMP_IN pixel_5222/SF_IB
+ pixel_5222/PIX_OUT pixel_5222/CSA_VREF pixel
Xpixel_5233 pixel_5233/gring pixel_5233/VDD pixel_5233/GND pixel_5233/VREF pixel_5233/ROW_SEL
+ pixel_5233/NB1 pixel_5233/VBIAS pixel_5233/NB2 pixel_5233/AMP_IN pixel_5233/SF_IB
+ pixel_5233/PIX_OUT pixel_5233/CSA_VREF pixel
Xpixel_5244 pixel_5244/gring pixel_5244/VDD pixel_5244/GND pixel_5244/VREF pixel_5244/ROW_SEL
+ pixel_5244/NB1 pixel_5244/VBIAS pixel_5244/NB2 pixel_5244/AMP_IN pixel_5244/SF_IB
+ pixel_5244/PIX_OUT pixel_5244/CSA_VREF pixel
Xpixel_5255 pixel_5255/gring pixel_5255/VDD pixel_5255/GND pixel_5255/VREF pixel_5255/ROW_SEL
+ pixel_5255/NB1 pixel_5255/VBIAS pixel_5255/NB2 pixel_5255/AMP_IN pixel_5255/SF_IB
+ pixel_5255/PIX_OUT pixel_5255/CSA_VREF pixel
Xpixel_5266 pixel_5266/gring pixel_5266/VDD pixel_5266/GND pixel_5266/VREF pixel_5266/ROW_SEL
+ pixel_5266/NB1 pixel_5266/VBIAS pixel_5266/NB2 pixel_5266/AMP_IN pixel_5266/SF_IB
+ pixel_5266/PIX_OUT pixel_5266/CSA_VREF pixel
Xpixel_4510 pixel_4510/gring pixel_4510/VDD pixel_4510/GND pixel_4510/VREF pixel_4510/ROW_SEL
+ pixel_4510/NB1 pixel_4510/VBIAS pixel_4510/NB2 pixel_4510/AMP_IN pixel_4510/SF_IB
+ pixel_4510/PIX_OUT pixel_4510/CSA_VREF pixel
Xpixel_4521 pixel_4521/gring pixel_4521/VDD pixel_4521/GND pixel_4521/VREF pixel_4521/ROW_SEL
+ pixel_4521/NB1 pixel_4521/VBIAS pixel_4521/NB2 pixel_4521/AMP_IN pixel_4521/SF_IB
+ pixel_4521/PIX_OUT pixel_4521/CSA_VREF pixel
Xpixel_5277 pixel_5277/gring pixel_5277/VDD pixel_5277/GND pixel_5277/VREF pixel_5277/ROW_SEL
+ pixel_5277/NB1 pixel_5277/VBIAS pixel_5277/NB2 pixel_5277/AMP_IN pixel_5277/SF_IB
+ pixel_5277/PIX_OUT pixel_5277/CSA_VREF pixel
Xpixel_5288 pixel_5288/gring pixel_5288/VDD pixel_5288/GND pixel_5288/VREF pixel_5288/ROW_SEL
+ pixel_5288/NB1 pixel_5288/VBIAS pixel_5288/NB2 pixel_5288/AMP_IN pixel_5288/SF_IB
+ pixel_5288/PIX_OUT pixel_5288/CSA_VREF pixel
Xpixel_5299 pixel_5299/gring pixel_5299/VDD pixel_5299/GND pixel_5299/VREF pixel_5299/ROW_SEL
+ pixel_5299/NB1 pixel_5299/VBIAS pixel_5299/NB2 pixel_5299/AMP_IN pixel_5299/SF_IB
+ pixel_5299/PIX_OUT pixel_5299/CSA_VREF pixel
Xpixel_4532 pixel_4532/gring pixel_4532/VDD pixel_4532/GND pixel_4532/VREF pixel_4532/ROW_SEL
+ pixel_4532/NB1 pixel_4532/VBIAS pixel_4532/NB2 pixel_4532/AMP_IN pixel_4532/SF_IB
+ pixel_4532/PIX_OUT pixel_4532/CSA_VREF pixel
Xpixel_4543 pixel_4543/gring pixel_4543/VDD pixel_4543/GND pixel_4543/VREF pixel_4543/ROW_SEL
+ pixel_4543/NB1 pixel_4543/VBIAS pixel_4543/NB2 pixel_4543/AMP_IN pixel_4543/SF_IB
+ pixel_4543/PIX_OUT pixel_4543/CSA_VREF pixel
Xpixel_4554 pixel_4554/gring pixel_4554/VDD pixel_4554/GND pixel_4554/VREF pixel_4554/ROW_SEL
+ pixel_4554/NB1 pixel_4554/VBIAS pixel_4554/NB2 pixel_4554/AMP_IN pixel_4554/SF_IB
+ pixel_4554/PIX_OUT pixel_4554/CSA_VREF pixel
Xpixel_593 pixel_593/gring pixel_593/VDD pixel_593/GND pixel_593/VREF pixel_593/ROW_SEL
+ pixel_593/NB1 pixel_593/VBIAS pixel_593/NB2 pixel_593/AMP_IN pixel_593/SF_IB pixel_593/PIX_OUT
+ pixel_593/CSA_VREF pixel
Xpixel_582 pixel_582/gring pixel_582/VDD pixel_582/GND pixel_582/VREF pixel_582/ROW_SEL
+ pixel_582/NB1 pixel_582/VBIAS pixel_582/NB2 pixel_582/AMP_IN pixel_582/SF_IB pixel_582/PIX_OUT
+ pixel_582/CSA_VREF pixel
Xpixel_571 pixel_571/gring pixel_571/VDD pixel_571/GND pixel_571/VREF pixel_571/ROW_SEL
+ pixel_571/NB1 pixel_571/VBIAS pixel_571/NB2 pixel_571/AMP_IN pixel_571/SF_IB pixel_571/PIX_OUT
+ pixel_571/CSA_VREF pixel
Xpixel_560 pixel_560/gring pixel_560/VDD pixel_560/GND pixel_560/VREF pixel_560/ROW_SEL
+ pixel_560/NB1 pixel_560/VBIAS pixel_560/NB2 pixel_560/AMP_IN pixel_560/SF_IB pixel_560/PIX_OUT
+ pixel_560/CSA_VREF pixel
Xpixel_3853 pixel_3853/gring pixel_3853/VDD pixel_3853/GND pixel_3853/VREF pixel_3853/ROW_SEL
+ pixel_3853/NB1 pixel_3853/VBIAS pixel_3853/NB2 pixel_3853/AMP_IN pixel_3853/SF_IB
+ pixel_3853/PIX_OUT pixel_3853/CSA_VREF pixel
Xpixel_4565 pixel_4565/gring pixel_4565/VDD pixel_4565/GND pixel_4565/VREF pixel_4565/ROW_SEL
+ pixel_4565/NB1 pixel_4565/VBIAS pixel_4565/NB2 pixel_4565/AMP_IN pixel_4565/SF_IB
+ pixel_4565/PIX_OUT pixel_4565/CSA_VREF pixel
Xpixel_4576 pixel_4576/gring pixel_4576/VDD pixel_4576/GND pixel_4576/VREF pixel_4576/ROW_SEL
+ pixel_4576/NB1 pixel_4576/VBIAS pixel_4576/NB2 pixel_4576/AMP_IN pixel_4576/SF_IB
+ pixel_4576/PIX_OUT pixel_4576/CSA_VREF pixel
Xpixel_4587 pixel_4587/gring pixel_4587/VDD pixel_4587/GND pixel_4587/VREF pixel_4587/ROW_SEL
+ pixel_4587/NB1 pixel_4587/VBIAS pixel_4587/NB2 pixel_4587/AMP_IN pixel_4587/SF_IB
+ pixel_4587/PIX_OUT pixel_4587/CSA_VREF pixel
Xpixel_3820 pixel_3820/gring pixel_3820/VDD pixel_3820/GND pixel_3820/VREF pixel_3820/ROW_SEL
+ pixel_3820/NB1 pixel_3820/VBIAS pixel_3820/NB2 pixel_3820/AMP_IN pixel_3820/SF_IB
+ pixel_3820/PIX_OUT pixel_3820/CSA_VREF pixel
Xpixel_3831 pixel_3831/gring pixel_3831/VDD pixel_3831/GND pixel_3831/VREF pixel_3831/ROW_SEL
+ pixel_3831/NB1 pixel_3831/VBIAS pixel_3831/NB2 pixel_3831/AMP_IN pixel_3831/SF_IB
+ pixel_3831/PIX_OUT pixel_3831/CSA_VREF pixel
Xpixel_3842 pixel_3842/gring pixel_3842/VDD pixel_3842/GND pixel_3842/VREF pixel_3842/ROW_SEL
+ pixel_3842/NB1 pixel_3842/VBIAS pixel_3842/NB2 pixel_3842/AMP_IN pixel_3842/SF_IB
+ pixel_3842/PIX_OUT pixel_3842/CSA_VREF pixel
Xpixel_3886 pixel_3886/gring pixel_3886/VDD pixel_3886/GND pixel_3886/VREF pixel_3886/ROW_SEL
+ pixel_3886/NB1 pixel_3886/VBIAS pixel_3886/NB2 pixel_3886/AMP_IN pixel_3886/SF_IB
+ pixel_3886/PIX_OUT pixel_3886/CSA_VREF pixel
Xpixel_3875 pixel_3875/gring pixel_3875/VDD pixel_3875/GND pixel_3875/VREF pixel_3875/ROW_SEL
+ pixel_3875/NB1 pixel_3875/VBIAS pixel_3875/NB2 pixel_3875/AMP_IN pixel_3875/SF_IB
+ pixel_3875/PIX_OUT pixel_3875/CSA_VREF pixel
Xpixel_3864 pixel_3864/gring pixel_3864/VDD pixel_3864/GND pixel_3864/VREF pixel_3864/ROW_SEL
+ pixel_3864/NB1 pixel_3864/VBIAS pixel_3864/NB2 pixel_3864/AMP_IN pixel_3864/SF_IB
+ pixel_3864/PIX_OUT pixel_3864/CSA_VREF pixel
Xpixel_4598 pixel_4598/gring pixel_4598/VDD pixel_4598/GND pixel_4598/VREF pixel_4598/ROW_SEL
+ pixel_4598/NB1 pixel_4598/VBIAS pixel_4598/NB2 pixel_4598/AMP_IN pixel_4598/SF_IB
+ pixel_4598/PIX_OUT pixel_4598/CSA_VREF pixel
Xpixel_3897 pixel_3897/gring pixel_3897/VDD pixel_3897/GND pixel_3897/VREF pixel_3897/ROW_SEL
+ pixel_3897/NB1 pixel_3897/VBIAS pixel_3897/NB2 pixel_3897/AMP_IN pixel_3897/SF_IB
+ pixel_3897/PIX_OUT pixel_3897/CSA_VREF pixel
Xpixel_7180 pixel_7180/gring pixel_7180/VDD pixel_7180/GND pixel_7180/VREF pixel_7180/ROW_SEL
+ pixel_7180/NB1 pixel_7180/VBIAS pixel_7180/NB2 pixel_7180/AMP_IN pixel_7180/SF_IB
+ pixel_7180/PIX_OUT pixel_7180/CSA_VREF pixel
Xpixel_7191 pixel_7191/gring pixel_7191/VDD pixel_7191/GND pixel_7191/VREF pixel_7191/ROW_SEL
+ pixel_7191/NB1 pixel_7191/VBIAS pixel_7191/NB2 pixel_7191/AMP_IN pixel_7191/SF_IB
+ pixel_7191/PIX_OUT pixel_7191/CSA_VREF pixel
Xpixel_6490 pixel_6490/gring pixel_6490/VDD pixel_6490/GND pixel_6490/VREF pixel_6490/ROW_SEL
+ pixel_6490/NB1 pixel_6490/VBIAS pixel_6490/NB2 pixel_6490/AMP_IN pixel_6490/SF_IB
+ pixel_6490/PIX_OUT pixel_6490/CSA_VREF pixel
Xpixel_8809 pixel_8809/gring pixel_8809/VDD pixel_8809/GND pixel_8809/VREF pixel_8809/ROW_SEL
+ pixel_8809/NB1 pixel_8809/VBIAS pixel_8809/NB2 pixel_8809/AMP_IN pixel_8809/SF_IB
+ pixel_8809/PIX_OUT pixel_8809/CSA_VREF pixel
Xpixel_3105 pixel_3105/gring pixel_3105/VDD pixel_3105/GND pixel_3105/VREF pixel_3105/ROW_SEL
+ pixel_3105/NB1 pixel_3105/VBIAS pixel_3105/NB2 pixel_3105/AMP_IN pixel_3105/SF_IB
+ pixel_3105/PIX_OUT pixel_3105/CSA_VREF pixel
Xpixel_3138 pixel_3138/gring pixel_3138/VDD pixel_3138/GND pixel_3138/VREF pixel_3138/ROW_SEL
+ pixel_3138/NB1 pixel_3138/VBIAS pixel_3138/NB2 pixel_3138/AMP_IN pixel_3138/SF_IB
+ pixel_3138/PIX_OUT pixel_3138/CSA_VREF pixel
Xpixel_3127 pixel_3127/gring pixel_3127/VDD pixel_3127/GND pixel_3127/VREF pixel_3127/ROW_SEL
+ pixel_3127/NB1 pixel_3127/VBIAS pixel_3127/NB2 pixel_3127/AMP_IN pixel_3127/SF_IB
+ pixel_3127/PIX_OUT pixel_3127/CSA_VREF pixel
Xpixel_3116 pixel_3116/gring pixel_3116/VDD pixel_3116/GND pixel_3116/VREF pixel_3116/ROW_SEL
+ pixel_3116/NB1 pixel_3116/VBIAS pixel_3116/NB2 pixel_3116/AMP_IN pixel_3116/SF_IB
+ pixel_3116/PIX_OUT pixel_3116/CSA_VREF pixel
Xpixel_2437 pixel_2437/gring pixel_2437/VDD pixel_2437/GND pixel_2437/VREF pixel_2437/ROW_SEL
+ pixel_2437/NB1 pixel_2437/VBIAS pixel_2437/NB2 pixel_2437/AMP_IN pixel_2437/SF_IB
+ pixel_2437/PIX_OUT pixel_2437/CSA_VREF pixel
Xpixel_2426 pixel_2426/gring pixel_2426/VDD pixel_2426/GND pixel_2426/VREF pixel_2426/ROW_SEL
+ pixel_2426/NB1 pixel_2426/VBIAS pixel_2426/NB2 pixel_2426/AMP_IN pixel_2426/SF_IB
+ pixel_2426/PIX_OUT pixel_2426/CSA_VREF pixel
Xpixel_2415 pixel_2415/gring pixel_2415/VDD pixel_2415/GND pixel_2415/VREF pixel_2415/ROW_SEL
+ pixel_2415/NB1 pixel_2415/VBIAS pixel_2415/NB2 pixel_2415/AMP_IN pixel_2415/SF_IB
+ pixel_2415/PIX_OUT pixel_2415/CSA_VREF pixel
Xpixel_2404 pixel_2404/gring pixel_2404/VDD pixel_2404/GND pixel_2404/VREF pixel_2404/ROW_SEL
+ pixel_2404/NB1 pixel_2404/VBIAS pixel_2404/NB2 pixel_2404/AMP_IN pixel_2404/SF_IB
+ pixel_2404/PIX_OUT pixel_2404/CSA_VREF pixel
Xpixel_3149 pixel_3149/gring pixel_3149/VDD pixel_3149/GND pixel_3149/VREF pixel_3149/ROW_SEL
+ pixel_3149/NB1 pixel_3149/VBIAS pixel_3149/NB2 pixel_3149/AMP_IN pixel_3149/SF_IB
+ pixel_3149/PIX_OUT pixel_3149/CSA_VREF pixel
Xpixel_1725 pixel_1725/gring pixel_1725/VDD pixel_1725/GND pixel_1725/VREF pixel_1725/ROW_SEL
+ pixel_1725/NB1 pixel_1725/VBIAS pixel_1725/NB2 pixel_1725/AMP_IN pixel_1725/SF_IB
+ pixel_1725/PIX_OUT pixel_1725/CSA_VREF pixel
Xpixel_1714 pixel_1714/gring pixel_1714/VDD pixel_1714/GND pixel_1714/VREF pixel_1714/ROW_SEL
+ pixel_1714/NB1 pixel_1714/VBIAS pixel_1714/NB2 pixel_1714/AMP_IN pixel_1714/SF_IB
+ pixel_1714/PIX_OUT pixel_1714/CSA_VREF pixel
Xpixel_1703 pixel_1703/gring pixel_1703/VDD pixel_1703/GND pixel_1703/VREF pixel_1703/ROW_SEL
+ pixel_1703/NB1 pixel_1703/VBIAS pixel_1703/NB2 pixel_1703/AMP_IN pixel_1703/SF_IB
+ pixel_1703/PIX_OUT pixel_1703/CSA_VREF pixel
Xpixel_2459 pixel_2459/gring pixel_2459/VDD pixel_2459/GND pixel_2459/VREF pixel_2459/ROW_SEL
+ pixel_2459/NB1 pixel_2459/VBIAS pixel_2459/NB2 pixel_2459/AMP_IN pixel_2459/SF_IB
+ pixel_2459/PIX_OUT pixel_2459/CSA_VREF pixel
Xpixel_2448 pixel_2448/gring pixel_2448/VDD pixel_2448/GND pixel_2448/VREF pixel_2448/ROW_SEL
+ pixel_2448/NB1 pixel_2448/VBIAS pixel_2448/NB2 pixel_2448/AMP_IN pixel_2448/SF_IB
+ pixel_2448/PIX_OUT pixel_2448/CSA_VREF pixel
Xpixel_1758 pixel_1758/gring pixel_1758/VDD pixel_1758/GND pixel_1758/VREF pixel_1758/ROW_SEL
+ pixel_1758/NB1 pixel_1758/VBIAS pixel_1758/NB2 pixel_1758/AMP_IN pixel_1758/SF_IB
+ pixel_1758/PIX_OUT pixel_1758/CSA_VREF pixel
Xpixel_1747 pixel_1747/gring pixel_1747/VDD pixel_1747/GND pixel_1747/VREF pixel_1747/ROW_SEL
+ pixel_1747/NB1 pixel_1747/VBIAS pixel_1747/NB2 pixel_1747/AMP_IN pixel_1747/SF_IB
+ pixel_1747/PIX_OUT pixel_1747/CSA_VREF pixel
Xpixel_1736 pixel_1736/gring pixel_1736/VDD pixel_1736/GND pixel_1736/VREF pixel_1736/ROW_SEL
+ pixel_1736/NB1 pixel_1736/VBIAS pixel_1736/NB2 pixel_1736/AMP_IN pixel_1736/SF_IB
+ pixel_1736/PIX_OUT pixel_1736/CSA_VREF pixel
Xpixel_1769 pixel_1769/gring pixel_1769/VDD pixel_1769/GND pixel_1769/VREF pixel_1769/ROW_SEL
+ pixel_1769/NB1 pixel_1769/VBIAS pixel_1769/NB2 pixel_1769/AMP_IN pixel_1769/SF_IB
+ pixel_1769/PIX_OUT pixel_1769/CSA_VREF pixel
Xpixel_5030 pixel_5030/gring pixel_5030/VDD pixel_5030/GND pixel_5030/VREF pixel_5030/ROW_SEL
+ pixel_5030/NB1 pixel_5030/VBIAS pixel_5030/NB2 pixel_5030/AMP_IN pixel_5030/SF_IB
+ pixel_5030/PIX_OUT pixel_5030/CSA_VREF pixel
Xpixel_5041 pixel_5041/gring pixel_5041/VDD pixel_5041/GND pixel_5041/VREF pixel_5041/ROW_SEL
+ pixel_5041/NB1 pixel_5041/VBIAS pixel_5041/NB2 pixel_5041/AMP_IN pixel_5041/SF_IB
+ pixel_5041/PIX_OUT pixel_5041/CSA_VREF pixel
Xpixel_5052 pixel_5052/gring pixel_5052/VDD pixel_5052/GND pixel_5052/VREF pixel_5052/ROW_SEL
+ pixel_5052/NB1 pixel_5052/VBIAS pixel_5052/NB2 pixel_5052/AMP_IN pixel_5052/SF_IB
+ pixel_5052/PIX_OUT pixel_5052/CSA_VREF pixel
Xpixel_5063 pixel_5063/gring pixel_5063/VDD pixel_5063/GND pixel_5063/VREF pixel_5063/ROW_SEL
+ pixel_5063/NB1 pixel_5063/VBIAS pixel_5063/NB2 pixel_5063/AMP_IN pixel_5063/SF_IB
+ pixel_5063/PIX_OUT pixel_5063/CSA_VREF pixel
Xpixel_5074 pixel_5074/gring pixel_5074/VDD pixel_5074/GND pixel_5074/VREF pixel_5074/ROW_SEL
+ pixel_5074/NB1 pixel_5074/VBIAS pixel_5074/NB2 pixel_5074/AMP_IN pixel_5074/SF_IB
+ pixel_5074/PIX_OUT pixel_5074/CSA_VREF pixel
Xpixel_5085 pixel_5085/gring pixel_5085/VDD pixel_5085/GND pixel_5085/VREF pixel_5085/ROW_SEL
+ pixel_5085/NB1 pixel_5085/VBIAS pixel_5085/NB2 pixel_5085/AMP_IN pixel_5085/SF_IB
+ pixel_5085/PIX_OUT pixel_5085/CSA_VREF pixel
Xpixel_5096 pixel_5096/gring pixel_5096/VDD pixel_5096/GND pixel_5096/VREF pixel_5096/ROW_SEL
+ pixel_5096/NB1 pixel_5096/VBIAS pixel_5096/NB2 pixel_5096/AMP_IN pixel_5096/SF_IB
+ pixel_5096/PIX_OUT pixel_5096/CSA_VREF pixel
Xpixel_4340 pixel_4340/gring pixel_4340/VDD pixel_4340/GND pixel_4340/VREF pixel_4340/ROW_SEL
+ pixel_4340/NB1 pixel_4340/VBIAS pixel_4340/NB2 pixel_4340/AMP_IN pixel_4340/SF_IB
+ pixel_4340/PIX_OUT pixel_4340/CSA_VREF pixel
Xpixel_4351 pixel_4351/gring pixel_4351/VDD pixel_4351/GND pixel_4351/VREF pixel_4351/ROW_SEL
+ pixel_4351/NB1 pixel_4351/VBIAS pixel_4351/NB2 pixel_4351/AMP_IN pixel_4351/SF_IB
+ pixel_4351/PIX_OUT pixel_4351/CSA_VREF pixel
Xpixel_4362 pixel_4362/gring pixel_4362/VDD pixel_4362/GND pixel_4362/VREF pixel_4362/ROW_SEL
+ pixel_4362/NB1 pixel_4362/VBIAS pixel_4362/NB2 pixel_4362/AMP_IN pixel_4362/SF_IB
+ pixel_4362/PIX_OUT pixel_4362/CSA_VREF pixel
Xpixel_390 pixel_390/gring pixel_390/VDD pixel_390/GND pixel_390/VREF pixel_390/ROW_SEL
+ pixel_390/NB1 pixel_390/VBIAS pixel_390/NB2 pixel_390/AMP_IN pixel_390/SF_IB pixel_390/PIX_OUT
+ pixel_390/CSA_VREF pixel
Xpixel_3661 pixel_3661/gring pixel_3661/VDD pixel_3661/GND pixel_3661/VREF pixel_3661/ROW_SEL
+ pixel_3661/NB1 pixel_3661/VBIAS pixel_3661/NB2 pixel_3661/AMP_IN pixel_3661/SF_IB
+ pixel_3661/PIX_OUT pixel_3661/CSA_VREF pixel
Xpixel_3650 pixel_3650/gring pixel_3650/VDD pixel_3650/GND pixel_3650/VREF pixel_3650/ROW_SEL
+ pixel_3650/NB1 pixel_3650/VBIAS pixel_3650/NB2 pixel_3650/AMP_IN pixel_3650/SF_IB
+ pixel_3650/PIX_OUT pixel_3650/CSA_VREF pixel
Xpixel_4373 pixel_4373/gring pixel_4373/VDD pixel_4373/GND pixel_4373/VREF pixel_4373/ROW_SEL
+ pixel_4373/NB1 pixel_4373/VBIAS pixel_4373/NB2 pixel_4373/AMP_IN pixel_4373/SF_IB
+ pixel_4373/PIX_OUT pixel_4373/CSA_VREF pixel
Xpixel_4384 pixel_4384/gring pixel_4384/VDD pixel_4384/GND pixel_4384/VREF pixel_4384/ROW_SEL
+ pixel_4384/NB1 pixel_4384/VBIAS pixel_4384/NB2 pixel_4384/AMP_IN pixel_4384/SF_IB
+ pixel_4384/PIX_OUT pixel_4384/CSA_VREF pixel
Xpixel_4395 pixel_4395/gring pixel_4395/VDD pixel_4395/GND pixel_4395/VREF pixel_4395/ROW_SEL
+ pixel_4395/NB1 pixel_4395/VBIAS pixel_4395/NB2 pixel_4395/AMP_IN pixel_4395/SF_IB
+ pixel_4395/PIX_OUT pixel_4395/CSA_VREF pixel
Xpixel_3694 pixel_3694/gring pixel_3694/VDD pixel_3694/GND pixel_3694/VREF pixel_3694/ROW_SEL
+ pixel_3694/NB1 pixel_3694/VBIAS pixel_3694/NB2 pixel_3694/AMP_IN pixel_3694/SF_IB
+ pixel_3694/PIX_OUT pixel_3694/CSA_VREF pixel
Xpixel_3683 pixel_3683/gring pixel_3683/VDD pixel_3683/GND pixel_3683/VREF pixel_3683/ROW_SEL
+ pixel_3683/NB1 pixel_3683/VBIAS pixel_3683/NB2 pixel_3683/AMP_IN pixel_3683/SF_IB
+ pixel_3683/PIX_OUT pixel_3683/CSA_VREF pixel
Xpixel_3672 pixel_3672/gring pixel_3672/VDD pixel_3672/GND pixel_3672/VREF pixel_3672/ROW_SEL
+ pixel_3672/NB1 pixel_3672/VBIAS pixel_3672/NB2 pixel_3672/AMP_IN pixel_3672/SF_IB
+ pixel_3672/PIX_OUT pixel_3672/CSA_VREF pixel
Xpixel_2982 pixel_2982/gring pixel_2982/VDD pixel_2982/GND pixel_2982/VREF pixel_2982/ROW_SEL
+ pixel_2982/NB1 pixel_2982/VBIAS pixel_2982/NB2 pixel_2982/AMP_IN pixel_2982/SF_IB
+ pixel_2982/PIX_OUT pixel_2982/CSA_VREF pixel
Xpixel_2971 pixel_2971/gring pixel_2971/VDD pixel_2971/GND pixel_2971/VREF pixel_2971/ROW_SEL
+ pixel_2971/NB1 pixel_2971/VBIAS pixel_2971/NB2 pixel_2971/AMP_IN pixel_2971/SF_IB
+ pixel_2971/PIX_OUT pixel_2971/CSA_VREF pixel
Xpixel_2960 pixel_2960/gring pixel_2960/VDD pixel_2960/GND pixel_2960/VREF pixel_2960/ROW_SEL
+ pixel_2960/NB1 pixel_2960/VBIAS pixel_2960/NB2 pixel_2960/AMP_IN pixel_2960/SF_IB
+ pixel_2960/PIX_OUT pixel_2960/CSA_VREF pixel
Xpixel_2993 pixel_2993/gring pixel_2993/VDD pixel_2993/GND pixel_2993/VREF pixel_2993/ROW_SEL
+ pixel_2993/NB1 pixel_2993/VBIAS pixel_2993/NB2 pixel_2993/AMP_IN pixel_2993/SF_IB
+ pixel_2993/PIX_OUT pixel_2993/CSA_VREF pixel
Xpixel_9329 pixel_9329/gring pixel_9329/VDD pixel_9329/GND pixel_9329/VREF pixel_9329/ROW_SEL
+ pixel_9329/NB1 pixel_9329/VBIAS pixel_9329/NB2 pixel_9329/AMP_IN pixel_9329/SF_IB
+ pixel_9329/PIX_OUT pixel_9329/CSA_VREF pixel
Xpixel_9318 pixel_9318/gring pixel_9318/VDD pixel_9318/GND pixel_9318/VREF pixel_9318/ROW_SEL
+ pixel_9318/NB1 pixel_9318/VBIAS pixel_9318/NB2 pixel_9318/AMP_IN pixel_9318/SF_IB
+ pixel_9318/PIX_OUT pixel_9318/CSA_VREF pixel
Xpixel_9307 pixel_9307/gring pixel_9307/VDD pixel_9307/GND pixel_9307/VREF pixel_9307/ROW_SEL
+ pixel_9307/NB1 pixel_9307/VBIAS pixel_9307/NB2 pixel_9307/AMP_IN pixel_9307/SF_IB
+ pixel_9307/PIX_OUT pixel_9307/CSA_VREF pixel
Xpixel_8617 pixel_8617/gring pixel_8617/VDD pixel_8617/GND pixel_8617/VREF pixel_8617/ROW_SEL
+ pixel_8617/NB1 pixel_8617/VBIAS pixel_8617/NB2 pixel_8617/AMP_IN pixel_8617/SF_IB
+ pixel_8617/PIX_OUT pixel_8617/CSA_VREF pixel
Xpixel_8606 pixel_8606/gring pixel_8606/VDD pixel_8606/GND pixel_8606/VREF pixel_8606/ROW_SEL
+ pixel_8606/NB1 pixel_8606/VBIAS pixel_8606/NB2 pixel_8606/AMP_IN pixel_8606/SF_IB
+ pixel_8606/PIX_OUT pixel_8606/CSA_VREF pixel
Xpixel_8639 pixel_8639/gring pixel_8639/VDD pixel_8639/GND pixel_8639/VREF pixel_8639/ROW_SEL
+ pixel_8639/NB1 pixel_8639/VBIAS pixel_8639/NB2 pixel_8639/AMP_IN pixel_8639/SF_IB
+ pixel_8639/PIX_OUT pixel_8639/CSA_VREF pixel
Xpixel_8628 pixel_8628/gring pixel_8628/VDD pixel_8628/GND pixel_8628/VREF pixel_8628/ROW_SEL
+ pixel_8628/NB1 pixel_8628/VBIAS pixel_8628/NB2 pixel_8628/AMP_IN pixel_8628/SF_IB
+ pixel_8628/PIX_OUT pixel_8628/CSA_VREF pixel
Xpixel_7905 pixel_7905/gring pixel_7905/VDD pixel_7905/GND pixel_7905/VREF pixel_7905/ROW_SEL
+ pixel_7905/NB1 pixel_7905/VBIAS pixel_7905/NB2 pixel_7905/AMP_IN pixel_7905/SF_IB
+ pixel_7905/PIX_OUT pixel_7905/CSA_VREF pixel
Xpixel_7916 pixel_7916/gring pixel_7916/VDD pixel_7916/GND pixel_7916/VREF pixel_7916/ROW_SEL
+ pixel_7916/NB1 pixel_7916/VBIAS pixel_7916/NB2 pixel_7916/AMP_IN pixel_7916/SF_IB
+ pixel_7916/PIX_OUT pixel_7916/CSA_VREF pixel
Xpixel_7927 pixel_7927/gring pixel_7927/VDD pixel_7927/GND pixel_7927/VREF pixel_7927/ROW_SEL
+ pixel_7927/NB1 pixel_7927/VBIAS pixel_7927/NB2 pixel_7927/AMP_IN pixel_7927/SF_IB
+ pixel_7927/PIX_OUT pixel_7927/CSA_VREF pixel
Xpixel_7938 pixel_7938/gring pixel_7938/VDD pixel_7938/GND pixel_7938/VREF pixel_7938/ROW_SEL
+ pixel_7938/NB1 pixel_7938/VBIAS pixel_7938/NB2 pixel_7938/AMP_IN pixel_7938/SF_IB
+ pixel_7938/PIX_OUT pixel_7938/CSA_VREF pixel
Xpixel_7949 pixel_7949/gring pixel_7949/VDD pixel_7949/GND pixel_7949/VREF pixel_7949/ROW_SEL
+ pixel_7949/NB1 pixel_7949/VBIAS pixel_7949/NB2 pixel_7949/AMP_IN pixel_7949/SF_IB
+ pixel_7949/PIX_OUT pixel_7949/CSA_VREF pixel
Xpixel_2212 pixel_2212/gring pixel_2212/VDD pixel_2212/GND pixel_2212/VREF pixel_2212/ROW_SEL
+ pixel_2212/NB1 pixel_2212/VBIAS pixel_2212/NB2 pixel_2212/AMP_IN pixel_2212/SF_IB
+ pixel_2212/PIX_OUT pixel_2212/CSA_VREF pixel
Xpixel_2201 pixel_2201/gring pixel_2201/VDD pixel_2201/GND pixel_2201/VREF pixel_2201/ROW_SEL
+ pixel_2201/NB1 pixel_2201/VBIAS pixel_2201/NB2 pixel_2201/AMP_IN pixel_2201/SF_IB
+ pixel_2201/PIX_OUT pixel_2201/CSA_VREF pixel
Xpixel_1500 pixel_1500/gring pixel_1500/VDD pixel_1500/GND pixel_1500/VREF pixel_1500/ROW_SEL
+ pixel_1500/NB1 pixel_1500/VBIAS pixel_1500/NB2 pixel_1500/AMP_IN pixel_1500/SF_IB
+ pixel_1500/PIX_OUT pixel_1500/CSA_VREF pixel
Xpixel_2245 pixel_2245/gring pixel_2245/VDD pixel_2245/GND pixel_2245/VREF pixel_2245/ROW_SEL
+ pixel_2245/NB1 pixel_2245/VBIAS pixel_2245/NB2 pixel_2245/AMP_IN pixel_2245/SF_IB
+ pixel_2245/PIX_OUT pixel_2245/CSA_VREF pixel
Xpixel_2234 pixel_2234/gring pixel_2234/VDD pixel_2234/GND pixel_2234/VREF pixel_2234/ROW_SEL
+ pixel_2234/NB1 pixel_2234/VBIAS pixel_2234/NB2 pixel_2234/AMP_IN pixel_2234/SF_IB
+ pixel_2234/PIX_OUT pixel_2234/CSA_VREF pixel
Xpixel_2223 pixel_2223/gring pixel_2223/VDD pixel_2223/GND pixel_2223/VREF pixel_2223/ROW_SEL
+ pixel_2223/NB1 pixel_2223/VBIAS pixel_2223/NB2 pixel_2223/AMP_IN pixel_2223/SF_IB
+ pixel_2223/PIX_OUT pixel_2223/CSA_VREF pixel
Xpixel_1533 pixel_1533/gring pixel_1533/VDD pixel_1533/GND pixel_1533/VREF pixel_1533/ROW_SEL
+ pixel_1533/NB1 pixel_1533/VBIAS pixel_1533/NB2 pixel_1533/AMP_IN pixel_1533/SF_IB
+ pixel_1533/PIX_OUT pixel_1533/CSA_VREF pixel
Xpixel_1522 pixel_1522/gring pixel_1522/VDD pixel_1522/GND pixel_1522/VREF pixel_1522/ROW_SEL
+ pixel_1522/NB1 pixel_1522/VBIAS pixel_1522/NB2 pixel_1522/AMP_IN pixel_1522/SF_IB
+ pixel_1522/PIX_OUT pixel_1522/CSA_VREF pixel
Xpixel_1511 pixel_1511/gring pixel_1511/VDD pixel_1511/GND pixel_1511/VREF pixel_1511/ROW_SEL
+ pixel_1511/NB1 pixel_1511/VBIAS pixel_1511/NB2 pixel_1511/AMP_IN pixel_1511/SF_IB
+ pixel_1511/PIX_OUT pixel_1511/CSA_VREF pixel
Xpixel_2278 pixel_2278/gring pixel_2278/VDD pixel_2278/GND pixel_2278/VREF pixel_2278/ROW_SEL
+ pixel_2278/NB1 pixel_2278/VBIAS pixel_2278/NB2 pixel_2278/AMP_IN pixel_2278/SF_IB
+ pixel_2278/PIX_OUT pixel_2278/CSA_VREF pixel
Xpixel_2267 pixel_2267/gring pixel_2267/VDD pixel_2267/GND pixel_2267/VREF pixel_2267/ROW_SEL
+ pixel_2267/NB1 pixel_2267/VBIAS pixel_2267/NB2 pixel_2267/AMP_IN pixel_2267/SF_IB
+ pixel_2267/PIX_OUT pixel_2267/CSA_VREF pixel
Xpixel_2256 pixel_2256/gring pixel_2256/VDD pixel_2256/GND pixel_2256/VREF pixel_2256/ROW_SEL
+ pixel_2256/NB1 pixel_2256/VBIAS pixel_2256/NB2 pixel_2256/AMP_IN pixel_2256/SF_IB
+ pixel_2256/PIX_OUT pixel_2256/CSA_VREF pixel
Xpixel_1577 pixel_1577/gring pixel_1577/VDD pixel_1577/GND pixel_1577/VREF pixel_1577/ROW_SEL
+ pixel_1577/NB1 pixel_1577/VBIAS pixel_1577/NB2 pixel_1577/AMP_IN pixel_1577/SF_IB
+ pixel_1577/PIX_OUT pixel_1577/CSA_VREF pixel
Xpixel_1566 pixel_1566/gring pixel_1566/VDD pixel_1566/GND pixel_1566/VREF pixel_1566/ROW_SEL
+ pixel_1566/NB1 pixel_1566/VBIAS pixel_1566/NB2 pixel_1566/AMP_IN pixel_1566/SF_IB
+ pixel_1566/PIX_OUT pixel_1566/CSA_VREF pixel
Xpixel_1555 pixel_1555/gring pixel_1555/VDD pixel_1555/GND pixel_1555/VREF pixel_1555/ROW_SEL
+ pixel_1555/NB1 pixel_1555/VBIAS pixel_1555/NB2 pixel_1555/AMP_IN pixel_1555/SF_IB
+ pixel_1555/PIX_OUT pixel_1555/CSA_VREF pixel
Xpixel_1544 pixel_1544/gring pixel_1544/VDD pixel_1544/GND pixel_1544/VREF pixel_1544/ROW_SEL
+ pixel_1544/NB1 pixel_1544/VBIAS pixel_1544/NB2 pixel_1544/AMP_IN pixel_1544/SF_IB
+ pixel_1544/PIX_OUT pixel_1544/CSA_VREF pixel
Xpixel_2289 pixel_2289/gring pixel_2289/VDD pixel_2289/GND pixel_2289/VREF pixel_2289/ROW_SEL
+ pixel_2289/NB1 pixel_2289/VBIAS pixel_2289/NB2 pixel_2289/AMP_IN pixel_2289/SF_IB
+ pixel_2289/PIX_OUT pixel_2289/CSA_VREF pixel
Xpixel_1599 pixel_1599/gring pixel_1599/VDD pixel_1599/GND pixel_1599/VREF pixel_1599/ROW_SEL
+ pixel_1599/NB1 pixel_1599/VBIAS pixel_1599/NB2 pixel_1599/AMP_IN pixel_1599/SF_IB
+ pixel_1599/PIX_OUT pixel_1599/CSA_VREF pixel
Xpixel_1588 pixel_1588/gring pixel_1588/VDD pixel_1588/GND pixel_1588/VREF pixel_1588/ROW_SEL
+ pixel_1588/NB1 pixel_1588/VBIAS pixel_1588/NB2 pixel_1588/AMP_IN pixel_1588/SF_IB
+ pixel_1588/PIX_OUT pixel_1588/CSA_VREF pixel
Xpixel_9841 pixel_9841/gring pixel_9841/VDD pixel_9841/GND pixel_9841/VREF pixel_9841/ROW_SEL
+ pixel_9841/NB1 pixel_9841/VBIAS pixel_9841/NB2 pixel_9841/AMP_IN pixel_9841/SF_IB
+ pixel_9841/PIX_OUT pixel_9841/CSA_VREF pixel
Xpixel_9830 pixel_9830/gring pixel_9830/VDD pixel_9830/GND pixel_9830/VREF pixel_9830/ROW_SEL
+ pixel_9830/NB1 pixel_9830/VBIAS pixel_9830/NB2 pixel_9830/AMP_IN pixel_9830/SF_IB
+ pixel_9830/PIX_OUT pixel_9830/CSA_VREF pixel
Xpixel_9852 pixel_9852/gring pixel_9852/VDD pixel_9852/GND pixel_9852/VREF pixel_9852/ROW_SEL
+ pixel_9852/NB1 pixel_9852/VBIAS pixel_9852/NB2 pixel_9852/AMP_IN pixel_9852/SF_IB
+ pixel_9852/PIX_OUT pixel_9852/CSA_VREF pixel
Xpixel_9863 pixel_9863/gring pixel_9863/VDD pixel_9863/GND pixel_9863/VREF pixel_9863/ROW_SEL
+ pixel_9863/NB1 pixel_9863/VBIAS pixel_9863/NB2 pixel_9863/AMP_IN pixel_9863/SF_IB
+ pixel_9863/PIX_OUT pixel_9863/CSA_VREF pixel
Xpixel_9874 pixel_9874/gring pixel_9874/VDD pixel_9874/GND pixel_9874/VREF pixel_9874/ROW_SEL
+ pixel_9874/NB1 pixel_9874/VBIAS pixel_9874/NB2 pixel_9874/AMP_IN pixel_9874/SF_IB
+ pixel_9874/PIX_OUT pixel_9874/CSA_VREF pixel
Xpixel_9885 pixel_9885/gring pixel_9885/VDD pixel_9885/GND pixel_9885/VREF pixel_9885/ROW_SEL
+ pixel_9885/NB1 pixel_9885/VBIAS pixel_9885/NB2 pixel_9885/AMP_IN pixel_9885/SF_IB
+ pixel_9885/PIX_OUT pixel_9885/CSA_VREF pixel
Xpixel_9896 pixel_9896/gring pixel_9896/VDD pixel_9896/GND pixel_9896/VREF pixel_9896/ROW_SEL
+ pixel_9896/NB1 pixel_9896/VBIAS pixel_9896/NB2 pixel_9896/AMP_IN pixel_9896/SF_IB
+ pixel_9896/PIX_OUT pixel_9896/CSA_VREF pixel
Xpixel_4170 pixel_4170/gring pixel_4170/VDD pixel_4170/GND pixel_4170/VREF pixel_4170/ROW_SEL
+ pixel_4170/NB1 pixel_4170/VBIAS pixel_4170/NB2 pixel_4170/AMP_IN pixel_4170/SF_IB
+ pixel_4170/PIX_OUT pixel_4170/CSA_VREF pixel
Xpixel_4181 pixel_4181/gring pixel_4181/VDD pixel_4181/GND pixel_4181/VREF pixel_4181/ROW_SEL
+ pixel_4181/NB1 pixel_4181/VBIAS pixel_4181/NB2 pixel_4181/AMP_IN pixel_4181/SF_IB
+ pixel_4181/PIX_OUT pixel_4181/CSA_VREF pixel
Xpixel_4192 pixel_4192/gring pixel_4192/VDD pixel_4192/GND pixel_4192/VREF pixel_4192/ROW_SEL
+ pixel_4192/NB1 pixel_4192/VBIAS pixel_4192/NB2 pixel_4192/AMP_IN pixel_4192/SF_IB
+ pixel_4192/PIX_OUT pixel_4192/CSA_VREF pixel
Xpixel_3491 pixel_3491/gring pixel_3491/VDD pixel_3491/GND pixel_3491/VREF pixel_3491/ROW_SEL
+ pixel_3491/NB1 pixel_3491/VBIAS pixel_3491/NB2 pixel_3491/AMP_IN pixel_3491/SF_IB
+ pixel_3491/PIX_OUT pixel_3491/CSA_VREF pixel
Xpixel_3480 pixel_3480/gring pixel_3480/VDD pixel_3480/GND pixel_3480/VREF pixel_3480/ROW_SEL
+ pixel_3480/NB1 pixel_3480/VBIAS pixel_3480/NB2 pixel_3480/AMP_IN pixel_3480/SF_IB
+ pixel_3480/PIX_OUT pixel_3480/CSA_VREF pixel
Xpixel_2790 pixel_2790/gring pixel_2790/VDD pixel_2790/GND pixel_2790/VREF pixel_2790/ROW_SEL
+ pixel_2790/NB1 pixel_2790/VBIAS pixel_2790/NB2 pixel_2790/AMP_IN pixel_2790/SF_IB
+ pixel_2790/PIX_OUT pixel_2790/CSA_VREF pixel
Xpixel_9104 pixel_9104/gring pixel_9104/VDD pixel_9104/GND pixel_9104/VREF pixel_9104/ROW_SEL
+ pixel_9104/NB1 pixel_9104/VBIAS pixel_9104/NB2 pixel_9104/AMP_IN pixel_9104/SF_IB
+ pixel_9104/PIX_OUT pixel_9104/CSA_VREF pixel
Xpixel_9137 pixel_9137/gring pixel_9137/VDD pixel_9137/GND pixel_9137/VREF pixel_9137/ROW_SEL
+ pixel_9137/NB1 pixel_9137/VBIAS pixel_9137/NB2 pixel_9137/AMP_IN pixel_9137/SF_IB
+ pixel_9137/PIX_OUT pixel_9137/CSA_VREF pixel
Xpixel_9126 pixel_9126/gring pixel_9126/VDD pixel_9126/GND pixel_9126/VREF pixel_9126/ROW_SEL
+ pixel_9126/NB1 pixel_9126/VBIAS pixel_9126/NB2 pixel_9126/AMP_IN pixel_9126/SF_IB
+ pixel_9126/PIX_OUT pixel_9126/CSA_VREF pixel
Xpixel_9115 pixel_9115/gring pixel_9115/VDD pixel_9115/GND pixel_9115/VREF pixel_9115/ROW_SEL
+ pixel_9115/NB1 pixel_9115/VBIAS pixel_9115/NB2 pixel_9115/AMP_IN pixel_9115/SF_IB
+ pixel_9115/PIX_OUT pixel_9115/CSA_VREF pixel
Xpixel_8425 pixel_8425/gring pixel_8425/VDD pixel_8425/GND pixel_8425/VREF pixel_8425/ROW_SEL
+ pixel_8425/NB1 pixel_8425/VBIAS pixel_8425/NB2 pixel_8425/AMP_IN pixel_8425/SF_IB
+ pixel_8425/PIX_OUT pixel_8425/CSA_VREF pixel
Xpixel_8414 pixel_8414/gring pixel_8414/VDD pixel_8414/GND pixel_8414/VREF pixel_8414/ROW_SEL
+ pixel_8414/NB1 pixel_8414/VBIAS pixel_8414/NB2 pixel_8414/AMP_IN pixel_8414/SF_IB
+ pixel_8414/PIX_OUT pixel_8414/CSA_VREF pixel
Xpixel_8403 pixel_8403/gring pixel_8403/VDD pixel_8403/GND pixel_8403/VREF pixel_8403/ROW_SEL
+ pixel_8403/NB1 pixel_8403/VBIAS pixel_8403/NB2 pixel_8403/AMP_IN pixel_8403/SF_IB
+ pixel_8403/PIX_OUT pixel_8403/CSA_VREF pixel
Xpixel_9159 pixel_9159/gring pixel_9159/VDD pixel_9159/GND pixel_9159/VREF pixel_9159/ROW_SEL
+ pixel_9159/NB1 pixel_9159/VBIAS pixel_9159/NB2 pixel_9159/AMP_IN pixel_9159/SF_IB
+ pixel_9159/PIX_OUT pixel_9159/CSA_VREF pixel
Xpixel_9148 pixel_9148/gring pixel_9148/VDD pixel_9148/GND pixel_9148/VREF pixel_9148/ROW_SEL
+ pixel_9148/NB1 pixel_9148/VBIAS pixel_9148/NB2 pixel_9148/AMP_IN pixel_9148/SF_IB
+ pixel_9148/PIX_OUT pixel_9148/CSA_VREF pixel
Xpixel_8436 pixel_8436/gring pixel_8436/VDD pixel_8436/GND pixel_8436/VREF pixel_8436/ROW_SEL
+ pixel_8436/NB1 pixel_8436/VBIAS pixel_8436/NB2 pixel_8436/AMP_IN pixel_8436/SF_IB
+ pixel_8436/PIX_OUT pixel_8436/CSA_VREF pixel
Xpixel_8447 pixel_8447/gring pixel_8447/VDD pixel_8447/GND pixel_8447/VREF pixel_8447/ROW_SEL
+ pixel_8447/NB1 pixel_8447/VBIAS pixel_8447/NB2 pixel_8447/AMP_IN pixel_8447/SF_IB
+ pixel_8447/PIX_OUT pixel_8447/CSA_VREF pixel
Xpixel_8458 pixel_8458/gring pixel_8458/VDD pixel_8458/GND pixel_8458/VREF pixel_8458/ROW_SEL
+ pixel_8458/NB1 pixel_8458/VBIAS pixel_8458/NB2 pixel_8458/AMP_IN pixel_8458/SF_IB
+ pixel_8458/PIX_OUT pixel_8458/CSA_VREF pixel
Xpixel_8469 pixel_8469/gring pixel_8469/VDD pixel_8469/GND pixel_8469/VREF pixel_8469/ROW_SEL
+ pixel_8469/NB1 pixel_8469/VBIAS pixel_8469/NB2 pixel_8469/AMP_IN pixel_8469/SF_IB
+ pixel_8469/PIX_OUT pixel_8469/CSA_VREF pixel
Xpixel_7702 pixel_7702/gring pixel_7702/VDD pixel_7702/GND pixel_7702/VREF pixel_7702/ROW_SEL
+ pixel_7702/NB1 pixel_7702/VBIAS pixel_7702/NB2 pixel_7702/AMP_IN pixel_7702/SF_IB
+ pixel_7702/PIX_OUT pixel_7702/CSA_VREF pixel
Xpixel_7713 pixel_7713/gring pixel_7713/VDD pixel_7713/GND pixel_7713/VREF pixel_7713/ROW_SEL
+ pixel_7713/NB1 pixel_7713/VBIAS pixel_7713/NB2 pixel_7713/AMP_IN pixel_7713/SF_IB
+ pixel_7713/PIX_OUT pixel_7713/CSA_VREF pixel
Xpixel_7724 pixel_7724/gring pixel_7724/VDD pixel_7724/GND pixel_7724/VREF pixel_7724/ROW_SEL
+ pixel_7724/NB1 pixel_7724/VBIAS pixel_7724/NB2 pixel_7724/AMP_IN pixel_7724/SF_IB
+ pixel_7724/PIX_OUT pixel_7724/CSA_VREF pixel
Xpixel_7735 pixel_7735/gring pixel_7735/VDD pixel_7735/GND pixel_7735/VREF pixel_7735/ROW_SEL
+ pixel_7735/NB1 pixel_7735/VBIAS pixel_7735/NB2 pixel_7735/AMP_IN pixel_7735/SF_IB
+ pixel_7735/PIX_OUT pixel_7735/CSA_VREF pixel
Xpixel_7746 pixel_7746/gring pixel_7746/VDD pixel_7746/GND pixel_7746/VREF pixel_7746/ROW_SEL
+ pixel_7746/NB1 pixel_7746/VBIAS pixel_7746/NB2 pixel_7746/AMP_IN pixel_7746/SF_IB
+ pixel_7746/PIX_OUT pixel_7746/CSA_VREF pixel
Xpixel_7757 pixel_7757/gring pixel_7757/VDD pixel_7757/GND pixel_7757/VREF pixel_7757/ROW_SEL
+ pixel_7757/NB1 pixel_7757/VBIAS pixel_7757/NB2 pixel_7757/AMP_IN pixel_7757/SF_IB
+ pixel_7757/PIX_OUT pixel_7757/CSA_VREF pixel
Xpixel_7768 pixel_7768/gring pixel_7768/VDD pixel_7768/GND pixel_7768/VREF pixel_7768/ROW_SEL
+ pixel_7768/NB1 pixel_7768/VBIAS pixel_7768/NB2 pixel_7768/AMP_IN pixel_7768/SF_IB
+ pixel_7768/PIX_OUT pixel_7768/CSA_VREF pixel
Xpixel_7779 pixel_7779/gring pixel_7779/VDD pixel_7779/GND pixel_7779/VREF pixel_7779/ROW_SEL
+ pixel_7779/NB1 pixel_7779/VBIAS pixel_7779/NB2 pixel_7779/AMP_IN pixel_7779/SF_IB
+ pixel_7779/PIX_OUT pixel_7779/CSA_VREF pixel
Xpixel_2020 pixel_2020/gring pixel_2020/VDD pixel_2020/GND pixel_2020/VREF pixel_2020/ROW_SEL
+ pixel_2020/NB1 pixel_2020/VBIAS pixel_2020/NB2 pixel_2020/AMP_IN pixel_2020/SF_IB
+ pixel_2020/PIX_OUT pixel_2020/CSA_VREF pixel
Xpixel_2053 pixel_2053/gring pixel_2053/VDD pixel_2053/GND pixel_2053/VREF pixel_2053/ROW_SEL
+ pixel_2053/NB1 pixel_2053/VBIAS pixel_2053/NB2 pixel_2053/AMP_IN pixel_2053/SF_IB
+ pixel_2053/PIX_OUT pixel_2053/CSA_VREF pixel
Xpixel_2042 pixel_2042/gring pixel_2042/VDD pixel_2042/GND pixel_2042/VREF pixel_2042/ROW_SEL
+ pixel_2042/NB1 pixel_2042/VBIAS pixel_2042/NB2 pixel_2042/AMP_IN pixel_2042/SF_IB
+ pixel_2042/PIX_OUT pixel_2042/CSA_VREF pixel
Xpixel_2031 pixel_2031/gring pixel_2031/VDD pixel_2031/GND pixel_2031/VREF pixel_2031/ROW_SEL
+ pixel_2031/NB1 pixel_2031/VBIAS pixel_2031/NB2 pixel_2031/AMP_IN pixel_2031/SF_IB
+ pixel_2031/PIX_OUT pixel_2031/CSA_VREF pixel
Xpixel_1341 pixel_1341/gring pixel_1341/VDD pixel_1341/GND pixel_1341/VREF pixel_1341/ROW_SEL
+ pixel_1341/NB1 pixel_1341/VBIAS pixel_1341/NB2 pixel_1341/AMP_IN pixel_1341/SF_IB
+ pixel_1341/PIX_OUT pixel_1341/CSA_VREF pixel
Xpixel_1330 pixel_1330/gring pixel_1330/VDD pixel_1330/GND pixel_1330/VREF pixel_1330/ROW_SEL
+ pixel_1330/NB1 pixel_1330/VBIAS pixel_1330/NB2 pixel_1330/AMP_IN pixel_1330/SF_IB
+ pixel_1330/PIX_OUT pixel_1330/CSA_VREF pixel
Xpixel_2086 pixel_2086/gring pixel_2086/VDD pixel_2086/GND pixel_2086/VREF pixel_2086/ROW_SEL
+ pixel_2086/NB1 pixel_2086/VBIAS pixel_2086/NB2 pixel_2086/AMP_IN pixel_2086/SF_IB
+ pixel_2086/PIX_OUT pixel_2086/CSA_VREF pixel
Xpixel_2075 pixel_2075/gring pixel_2075/VDD pixel_2075/GND pixel_2075/VREF pixel_2075/ROW_SEL
+ pixel_2075/NB1 pixel_2075/VBIAS pixel_2075/NB2 pixel_2075/AMP_IN pixel_2075/SF_IB
+ pixel_2075/PIX_OUT pixel_2075/CSA_VREF pixel
Xpixel_2064 pixel_2064/gring pixel_2064/VDD pixel_2064/GND pixel_2064/VREF pixel_2064/ROW_SEL
+ pixel_2064/NB1 pixel_2064/VBIAS pixel_2064/NB2 pixel_2064/AMP_IN pixel_2064/SF_IB
+ pixel_2064/PIX_OUT pixel_2064/CSA_VREF pixel
Xpixel_1385 pixel_1385/gring pixel_1385/VDD pixel_1385/GND pixel_1385/VREF pixel_1385/ROW_SEL
+ pixel_1385/NB1 pixel_1385/VBIAS pixel_1385/NB2 pixel_1385/AMP_IN pixel_1385/SF_IB
+ pixel_1385/PIX_OUT pixel_1385/CSA_VREF pixel
Xpixel_1374 pixel_1374/gring pixel_1374/VDD pixel_1374/GND pixel_1374/VREF pixel_1374/ROW_SEL
+ pixel_1374/NB1 pixel_1374/VBIAS pixel_1374/NB2 pixel_1374/AMP_IN pixel_1374/SF_IB
+ pixel_1374/PIX_OUT pixel_1374/CSA_VREF pixel
Xpixel_1363 pixel_1363/gring pixel_1363/VDD pixel_1363/GND pixel_1363/VREF pixel_1363/ROW_SEL
+ pixel_1363/NB1 pixel_1363/VBIAS pixel_1363/NB2 pixel_1363/AMP_IN pixel_1363/SF_IB
+ pixel_1363/PIX_OUT pixel_1363/CSA_VREF pixel
Xpixel_1352 pixel_1352/gring pixel_1352/VDD pixel_1352/GND pixel_1352/VREF pixel_1352/ROW_SEL
+ pixel_1352/NB1 pixel_1352/VBIAS pixel_1352/NB2 pixel_1352/AMP_IN pixel_1352/SF_IB
+ pixel_1352/PIX_OUT pixel_1352/CSA_VREF pixel
Xpixel_2097 pixel_2097/gring pixel_2097/VDD pixel_2097/GND pixel_2097/VREF pixel_2097/ROW_SEL
+ pixel_2097/NB1 pixel_2097/VBIAS pixel_2097/NB2 pixel_2097/AMP_IN pixel_2097/SF_IB
+ pixel_2097/PIX_OUT pixel_2097/CSA_VREF pixel
Xpixel_1396 pixel_1396/gring pixel_1396/VDD pixel_1396/GND pixel_1396/VREF pixel_1396/ROW_SEL
+ pixel_1396/NB1 pixel_1396/VBIAS pixel_1396/NB2 pixel_1396/AMP_IN pixel_1396/SF_IB
+ pixel_1396/PIX_OUT pixel_1396/CSA_VREF pixel
Xpixel_9693 pixel_9693/gring pixel_9693/VDD pixel_9693/GND pixel_9693/VREF pixel_9693/ROW_SEL
+ pixel_9693/NB1 pixel_9693/VBIAS pixel_9693/NB2 pixel_9693/AMP_IN pixel_9693/SF_IB
+ pixel_9693/PIX_OUT pixel_9693/CSA_VREF pixel
Xpixel_9660 pixel_9660/gring pixel_9660/VDD pixel_9660/GND pixel_9660/VREF pixel_9660/ROW_SEL
+ pixel_9660/NB1 pixel_9660/VBIAS pixel_9660/NB2 pixel_9660/AMP_IN pixel_9660/SF_IB
+ pixel_9660/PIX_OUT pixel_9660/CSA_VREF pixel
Xpixel_9671 pixel_9671/gring pixel_9671/VDD pixel_9671/GND pixel_9671/VREF pixel_9671/ROW_SEL
+ pixel_9671/NB1 pixel_9671/VBIAS pixel_9671/NB2 pixel_9671/AMP_IN pixel_9671/SF_IB
+ pixel_9671/PIX_OUT pixel_9671/CSA_VREF pixel
Xpixel_9682 pixel_9682/gring pixel_9682/VDD pixel_9682/GND pixel_9682/VREF pixel_9682/ROW_SEL
+ pixel_9682/NB1 pixel_9682/VBIAS pixel_9682/NB2 pixel_9682/AMP_IN pixel_9682/SF_IB
+ pixel_9682/PIX_OUT pixel_9682/CSA_VREF pixel
Xpixel_8981 pixel_8981/gring pixel_8981/VDD pixel_8981/GND pixel_8981/VREF pixel_8981/ROW_SEL
+ pixel_8981/NB1 pixel_8981/VBIAS pixel_8981/NB2 pixel_8981/AMP_IN pixel_8981/SF_IB
+ pixel_8981/PIX_OUT pixel_8981/CSA_VREF pixel
Xpixel_8970 pixel_8970/gring pixel_8970/VDD pixel_8970/GND pixel_8970/VREF pixel_8970/ROW_SEL
+ pixel_8970/NB1 pixel_8970/VBIAS pixel_8970/NB2 pixel_8970/AMP_IN pixel_8970/SF_IB
+ pixel_8970/PIX_OUT pixel_8970/CSA_VREF pixel
Xpixel_8992 pixel_8992/gring pixel_8992/VDD pixel_8992/GND pixel_8992/VREF pixel_8992/ROW_SEL
+ pixel_8992/NB1 pixel_8992/VBIAS pixel_8992/NB2 pixel_8992/AMP_IN pixel_8992/SF_IB
+ pixel_8992/PIX_OUT pixel_8992/CSA_VREF pixel
Xpixel_7009 pixel_7009/gring pixel_7009/VDD pixel_7009/GND pixel_7009/VREF pixel_7009/ROW_SEL
+ pixel_7009/NB1 pixel_7009/VBIAS pixel_7009/NB2 pixel_7009/AMP_IN pixel_7009/SF_IB
+ pixel_7009/PIX_OUT pixel_7009/CSA_VREF pixel
Xpixel_6308 pixel_6308/gring pixel_6308/VDD pixel_6308/GND pixel_6308/VREF pixel_6308/ROW_SEL
+ pixel_6308/NB1 pixel_6308/VBIAS pixel_6308/NB2 pixel_6308/AMP_IN pixel_6308/SF_IB
+ pixel_6308/PIX_OUT pixel_6308/CSA_VREF pixel
Xpixel_6319 pixel_6319/gring pixel_6319/VDD pixel_6319/GND pixel_6319/VREF pixel_6319/ROW_SEL
+ pixel_6319/NB1 pixel_6319/VBIAS pixel_6319/NB2 pixel_6319/AMP_IN pixel_6319/SF_IB
+ pixel_6319/PIX_OUT pixel_6319/CSA_VREF pixel
Xpixel_5607 pixel_5607/gring pixel_5607/VDD pixel_5607/GND pixel_5607/VREF pixel_5607/ROW_SEL
+ pixel_5607/NB1 pixel_5607/VBIAS pixel_5607/NB2 pixel_5607/AMP_IN pixel_5607/SF_IB
+ pixel_5607/PIX_OUT pixel_5607/CSA_VREF pixel
Xpixel_5618 pixel_5618/gring pixel_5618/VDD pixel_5618/GND pixel_5618/VREF pixel_5618/ROW_SEL
+ pixel_5618/NB1 pixel_5618/VBIAS pixel_5618/NB2 pixel_5618/AMP_IN pixel_5618/SF_IB
+ pixel_5618/PIX_OUT pixel_5618/CSA_VREF pixel
Xpixel_5629 pixel_5629/gring pixel_5629/VDD pixel_5629/GND pixel_5629/VREF pixel_5629/ROW_SEL
+ pixel_5629/NB1 pixel_5629/VBIAS pixel_5629/NB2 pixel_5629/AMP_IN pixel_5629/SF_IB
+ pixel_5629/PIX_OUT pixel_5629/CSA_VREF pixel
Xpixel_923 pixel_923/gring pixel_923/VDD pixel_923/GND pixel_923/VREF pixel_923/ROW_SEL
+ pixel_923/NB1 pixel_923/VBIAS pixel_923/NB2 pixel_923/AMP_IN pixel_923/SF_IB pixel_923/PIX_OUT
+ pixel_923/CSA_VREF pixel
Xpixel_912 pixel_912/gring pixel_912/VDD pixel_912/GND pixel_912/VREF pixel_912/ROW_SEL
+ pixel_912/NB1 pixel_912/VBIAS pixel_912/NB2 pixel_912/AMP_IN pixel_912/SF_IB pixel_912/PIX_OUT
+ pixel_912/CSA_VREF pixel
Xpixel_901 pixel_901/gring pixel_901/VDD pixel_901/GND pixel_901/VREF pixel_901/ROW_SEL
+ pixel_901/NB1 pixel_901/VBIAS pixel_901/NB2 pixel_901/AMP_IN pixel_901/SF_IB pixel_901/PIX_OUT
+ pixel_901/CSA_VREF pixel
Xpixel_4906 pixel_4906/gring pixel_4906/VDD pixel_4906/GND pixel_4906/VREF pixel_4906/ROW_SEL
+ pixel_4906/NB1 pixel_4906/VBIAS pixel_4906/NB2 pixel_4906/AMP_IN pixel_4906/SF_IB
+ pixel_4906/PIX_OUT pixel_4906/CSA_VREF pixel
Xpixel_4917 pixel_4917/gring pixel_4917/VDD pixel_4917/GND pixel_4917/VREF pixel_4917/ROW_SEL
+ pixel_4917/NB1 pixel_4917/VBIAS pixel_4917/NB2 pixel_4917/AMP_IN pixel_4917/SF_IB
+ pixel_4917/PIX_OUT pixel_4917/CSA_VREF pixel
Xpixel_4928 pixel_4928/gring pixel_4928/VDD pixel_4928/GND pixel_4928/VREF pixel_4928/ROW_SEL
+ pixel_4928/NB1 pixel_4928/VBIAS pixel_4928/NB2 pixel_4928/AMP_IN pixel_4928/SF_IB
+ pixel_4928/PIX_OUT pixel_4928/CSA_VREF pixel
Xpixel_967 pixel_967/gring pixel_967/VDD pixel_967/GND pixel_967/VREF pixel_967/ROW_SEL
+ pixel_967/NB1 pixel_967/VBIAS pixel_967/NB2 pixel_967/AMP_IN pixel_967/SF_IB pixel_967/PIX_OUT
+ pixel_967/CSA_VREF pixel
Xpixel_956 pixel_956/gring pixel_956/VDD pixel_956/GND pixel_956/VREF pixel_956/ROW_SEL
+ pixel_956/NB1 pixel_956/VBIAS pixel_956/NB2 pixel_956/AMP_IN pixel_956/SF_IB pixel_956/PIX_OUT
+ pixel_956/CSA_VREF pixel
Xpixel_945 pixel_945/gring pixel_945/VDD pixel_945/GND pixel_945/VREF pixel_945/ROW_SEL
+ pixel_945/NB1 pixel_945/VBIAS pixel_945/NB2 pixel_945/AMP_IN pixel_945/SF_IB pixel_945/PIX_OUT
+ pixel_945/CSA_VREF pixel
Xpixel_934 pixel_934/gring pixel_934/VDD pixel_934/GND pixel_934/VREF pixel_934/ROW_SEL
+ pixel_934/NB1 pixel_934/VBIAS pixel_934/NB2 pixel_934/AMP_IN pixel_934/SF_IB pixel_934/PIX_OUT
+ pixel_934/CSA_VREF pixel
Xpixel_4939 pixel_4939/gring pixel_4939/VDD pixel_4939/GND pixel_4939/VREF pixel_4939/ROW_SEL
+ pixel_4939/NB1 pixel_4939/VBIAS pixel_4939/NB2 pixel_4939/AMP_IN pixel_4939/SF_IB
+ pixel_4939/PIX_OUT pixel_4939/CSA_VREF pixel
Xpixel_989 pixel_989/gring pixel_989/VDD pixel_989/GND pixel_989/VREF pixel_989/ROW_SEL
+ pixel_989/NB1 pixel_989/VBIAS pixel_989/NB2 pixel_989/AMP_IN pixel_989/SF_IB pixel_989/PIX_OUT
+ pixel_989/CSA_VREF pixel
Xpixel_978 pixel_978/gring pixel_978/VDD pixel_978/GND pixel_978/VREF pixel_978/ROW_SEL
+ pixel_978/NB1 pixel_978/VBIAS pixel_978/NB2 pixel_978/AMP_IN pixel_978/SF_IB pixel_978/PIX_OUT
+ pixel_978/CSA_VREF pixel
Xpixel_8200 pixel_8200/gring pixel_8200/VDD pixel_8200/GND pixel_8200/VREF pixel_8200/ROW_SEL
+ pixel_8200/NB1 pixel_8200/VBIAS pixel_8200/NB2 pixel_8200/AMP_IN pixel_8200/SF_IB
+ pixel_8200/PIX_OUT pixel_8200/CSA_VREF pixel
Xpixel_8211 pixel_8211/gring pixel_8211/VDD pixel_8211/GND pixel_8211/VREF pixel_8211/ROW_SEL
+ pixel_8211/NB1 pixel_8211/VBIAS pixel_8211/NB2 pixel_8211/AMP_IN pixel_8211/SF_IB
+ pixel_8211/PIX_OUT pixel_8211/CSA_VREF pixel
Xpixel_8222 pixel_8222/gring pixel_8222/VDD pixel_8222/GND pixel_8222/VREF pixel_8222/ROW_SEL
+ pixel_8222/NB1 pixel_8222/VBIAS pixel_8222/NB2 pixel_8222/AMP_IN pixel_8222/SF_IB
+ pixel_8222/PIX_OUT pixel_8222/CSA_VREF pixel
Xpixel_8233 pixel_8233/gring pixel_8233/VDD pixel_8233/GND pixel_8233/VREF pixel_8233/ROW_SEL
+ pixel_8233/NB1 pixel_8233/VBIAS pixel_8233/NB2 pixel_8233/AMP_IN pixel_8233/SF_IB
+ pixel_8233/PIX_OUT pixel_8233/CSA_VREF pixel
Xpixel_8244 pixel_8244/gring pixel_8244/VDD pixel_8244/GND pixel_8244/VREF pixel_8244/ROW_SEL
+ pixel_8244/NB1 pixel_8244/VBIAS pixel_8244/NB2 pixel_8244/AMP_IN pixel_8244/SF_IB
+ pixel_8244/PIX_OUT pixel_8244/CSA_VREF pixel
Xpixel_8255 pixel_8255/gring pixel_8255/VDD pixel_8255/GND pixel_8255/VREF pixel_8255/ROW_SEL
+ pixel_8255/NB1 pixel_8255/VBIAS pixel_8255/NB2 pixel_8255/AMP_IN pixel_8255/SF_IB
+ pixel_8255/PIX_OUT pixel_8255/CSA_VREF pixel
Xpixel_8266 pixel_8266/gring pixel_8266/VDD pixel_8266/GND pixel_8266/VREF pixel_8266/ROW_SEL
+ pixel_8266/NB1 pixel_8266/VBIAS pixel_8266/NB2 pixel_8266/AMP_IN pixel_8266/SF_IB
+ pixel_8266/PIX_OUT pixel_8266/CSA_VREF pixel
Xpixel_8277 pixel_8277/gring pixel_8277/VDD pixel_8277/GND pixel_8277/VREF pixel_8277/ROW_SEL
+ pixel_8277/NB1 pixel_8277/VBIAS pixel_8277/NB2 pixel_8277/AMP_IN pixel_8277/SF_IB
+ pixel_8277/PIX_OUT pixel_8277/CSA_VREF pixel
Xpixel_7510 pixel_7510/gring pixel_7510/VDD pixel_7510/GND pixel_7510/VREF pixel_7510/ROW_SEL
+ pixel_7510/NB1 pixel_7510/VBIAS pixel_7510/NB2 pixel_7510/AMP_IN pixel_7510/SF_IB
+ pixel_7510/PIX_OUT pixel_7510/CSA_VREF pixel
Xpixel_7521 pixel_7521/gring pixel_7521/VDD pixel_7521/GND pixel_7521/VREF pixel_7521/ROW_SEL
+ pixel_7521/NB1 pixel_7521/VBIAS pixel_7521/NB2 pixel_7521/AMP_IN pixel_7521/SF_IB
+ pixel_7521/PIX_OUT pixel_7521/CSA_VREF pixel
Xpixel_7532 pixel_7532/gring pixel_7532/VDD pixel_7532/GND pixel_7532/VREF pixel_7532/ROW_SEL
+ pixel_7532/NB1 pixel_7532/VBIAS pixel_7532/NB2 pixel_7532/AMP_IN pixel_7532/SF_IB
+ pixel_7532/PIX_OUT pixel_7532/CSA_VREF pixel
Xpixel_8288 pixel_8288/gring pixel_8288/VDD pixel_8288/GND pixel_8288/VREF pixel_8288/ROW_SEL
+ pixel_8288/NB1 pixel_8288/VBIAS pixel_8288/NB2 pixel_8288/AMP_IN pixel_8288/SF_IB
+ pixel_8288/PIX_OUT pixel_8288/CSA_VREF pixel
Xpixel_8299 pixel_8299/gring pixel_8299/VDD pixel_8299/GND pixel_8299/VREF pixel_8299/ROW_SEL
+ pixel_8299/NB1 pixel_8299/VBIAS pixel_8299/NB2 pixel_8299/AMP_IN pixel_8299/SF_IB
+ pixel_8299/PIX_OUT pixel_8299/CSA_VREF pixel
Xpixel_7543 pixel_7543/gring pixel_7543/VDD pixel_7543/GND pixel_7543/VREF pixel_7543/ROW_SEL
+ pixel_7543/NB1 pixel_7543/VBIAS pixel_7543/NB2 pixel_7543/AMP_IN pixel_7543/SF_IB
+ pixel_7543/PIX_OUT pixel_7543/CSA_VREF pixel
Xpixel_7554 pixel_7554/gring pixel_7554/VDD pixel_7554/GND pixel_7554/VREF pixel_7554/ROW_SEL
+ pixel_7554/NB1 pixel_7554/VBIAS pixel_7554/NB2 pixel_7554/AMP_IN pixel_7554/SF_IB
+ pixel_7554/PIX_OUT pixel_7554/CSA_VREF pixel
Xpixel_7565 pixel_7565/gring pixel_7565/VDD pixel_7565/GND pixel_7565/VREF pixel_7565/ROW_SEL
+ pixel_7565/NB1 pixel_7565/VBIAS pixel_7565/NB2 pixel_7565/AMP_IN pixel_7565/SF_IB
+ pixel_7565/PIX_OUT pixel_7565/CSA_VREF pixel
Xpixel_6820 pixel_6820/gring pixel_6820/VDD pixel_6820/GND pixel_6820/VREF pixel_6820/ROW_SEL
+ pixel_6820/NB1 pixel_6820/VBIAS pixel_6820/NB2 pixel_6820/AMP_IN pixel_6820/SF_IB
+ pixel_6820/PIX_OUT pixel_6820/CSA_VREF pixel
Xpixel_7576 pixel_7576/gring pixel_7576/VDD pixel_7576/GND pixel_7576/VREF pixel_7576/ROW_SEL
+ pixel_7576/NB1 pixel_7576/VBIAS pixel_7576/NB2 pixel_7576/AMP_IN pixel_7576/SF_IB
+ pixel_7576/PIX_OUT pixel_7576/CSA_VREF pixel
Xpixel_7587 pixel_7587/gring pixel_7587/VDD pixel_7587/GND pixel_7587/VREF pixel_7587/ROW_SEL
+ pixel_7587/NB1 pixel_7587/VBIAS pixel_7587/NB2 pixel_7587/AMP_IN pixel_7587/SF_IB
+ pixel_7587/PIX_OUT pixel_7587/CSA_VREF pixel
Xpixel_7598 pixel_7598/gring pixel_7598/VDD pixel_7598/GND pixel_7598/VREF pixel_7598/ROW_SEL
+ pixel_7598/NB1 pixel_7598/VBIAS pixel_7598/NB2 pixel_7598/AMP_IN pixel_7598/SF_IB
+ pixel_7598/PIX_OUT pixel_7598/CSA_VREF pixel
Xpixel_6831 pixel_6831/gring pixel_6831/VDD pixel_6831/GND pixel_6831/VREF pixel_6831/ROW_SEL
+ pixel_6831/NB1 pixel_6831/VBIAS pixel_6831/NB2 pixel_6831/AMP_IN pixel_6831/SF_IB
+ pixel_6831/PIX_OUT pixel_6831/CSA_VREF pixel
Xpixel_6842 pixel_6842/gring pixel_6842/VDD pixel_6842/GND pixel_6842/VREF pixel_6842/ROW_SEL
+ pixel_6842/NB1 pixel_6842/VBIAS pixel_6842/NB2 pixel_6842/AMP_IN pixel_6842/SF_IB
+ pixel_6842/PIX_OUT pixel_6842/CSA_VREF pixel
Xpixel_6853 pixel_6853/gring pixel_6853/VDD pixel_6853/GND pixel_6853/VREF pixel_6853/ROW_SEL
+ pixel_6853/NB1 pixel_6853/VBIAS pixel_6853/NB2 pixel_6853/AMP_IN pixel_6853/SF_IB
+ pixel_6853/PIX_OUT pixel_6853/CSA_VREF pixel
Xpixel_6864 pixel_6864/gring pixel_6864/VDD pixel_6864/GND pixel_6864/VREF pixel_6864/ROW_SEL
+ pixel_6864/NB1 pixel_6864/VBIAS pixel_6864/NB2 pixel_6864/AMP_IN pixel_6864/SF_IB
+ pixel_6864/PIX_OUT pixel_6864/CSA_VREF pixel
Xpixel_6875 pixel_6875/gring pixel_6875/VDD pixel_6875/GND pixel_6875/VREF pixel_6875/ROW_SEL
+ pixel_6875/NB1 pixel_6875/VBIAS pixel_6875/NB2 pixel_6875/AMP_IN pixel_6875/SF_IB
+ pixel_6875/PIX_OUT pixel_6875/CSA_VREF pixel
Xpixel_6886 pixel_6886/gring pixel_6886/VDD pixel_6886/GND pixel_6886/VREF pixel_6886/ROW_SEL
+ pixel_6886/NB1 pixel_6886/VBIAS pixel_6886/NB2 pixel_6886/AMP_IN pixel_6886/SF_IB
+ pixel_6886/PIX_OUT pixel_6886/CSA_VREF pixel
Xpixel_6897 pixel_6897/gring pixel_6897/VDD pixel_6897/GND pixel_6897/VREF pixel_6897/ROW_SEL
+ pixel_6897/NB1 pixel_6897/VBIAS pixel_6897/NB2 pixel_6897/AMP_IN pixel_6897/SF_IB
+ pixel_6897/PIX_OUT pixel_6897/CSA_VREF pixel
Xpixel_1160 pixel_1160/gring pixel_1160/VDD pixel_1160/GND pixel_1160/VREF pixel_1160/ROW_SEL
+ pixel_1160/NB1 pixel_1160/VBIAS pixel_1160/NB2 pixel_1160/AMP_IN pixel_1160/SF_IB
+ pixel_1160/PIX_OUT pixel_1160/CSA_VREF pixel
Xpixel_1193 pixel_1193/gring pixel_1193/VDD pixel_1193/GND pixel_1193/VREF pixel_1193/ROW_SEL
+ pixel_1193/NB1 pixel_1193/VBIAS pixel_1193/NB2 pixel_1193/AMP_IN pixel_1193/SF_IB
+ pixel_1193/PIX_OUT pixel_1193/CSA_VREF pixel
Xpixel_1182 pixel_1182/gring pixel_1182/VDD pixel_1182/GND pixel_1182/VREF pixel_1182/ROW_SEL
+ pixel_1182/NB1 pixel_1182/VBIAS pixel_1182/NB2 pixel_1182/AMP_IN pixel_1182/SF_IB
+ pixel_1182/PIX_OUT pixel_1182/CSA_VREF pixel
Xpixel_1171 pixel_1171/gring pixel_1171/VDD pixel_1171/GND pixel_1171/VREF pixel_1171/ROW_SEL
+ pixel_1171/NB1 pixel_1171/VBIAS pixel_1171/NB2 pixel_1171/AMP_IN pixel_1171/SF_IB
+ pixel_1171/PIX_OUT pixel_1171/CSA_VREF pixel
Xpixel_9490 pixel_9490/gring pixel_9490/VDD pixel_9490/GND pixel_9490/VREF pixel_9490/ROW_SEL
+ pixel_9490/NB1 pixel_9490/VBIAS pixel_9490/NB2 pixel_9490/AMP_IN pixel_9490/SF_IB
+ pixel_9490/PIX_OUT pixel_9490/CSA_VREF pixel
Xpixel_219 pixel_219/gring pixel_219/VDD pixel_219/GND pixel_219/VREF pixel_219/ROW_SEL
+ pixel_219/NB1 pixel_219/VBIAS pixel_219/NB2 pixel_219/AMP_IN pixel_219/SF_IB pixel_219/PIX_OUT
+ pixel_219/CSA_VREF pixel
Xpixel_208 pixel_208/gring pixel_208/VDD pixel_208/GND pixel_208/VREF pixel_208/ROW_SEL
+ pixel_208/NB1 pixel_208/VBIAS pixel_208/NB2 pixel_208/AMP_IN pixel_208/SF_IB pixel_208/PIX_OUT
+ pixel_208/CSA_VREF pixel
Xpixel_6105 pixel_6105/gring pixel_6105/VDD pixel_6105/GND pixel_6105/VREF pixel_6105/ROW_SEL
+ pixel_6105/NB1 pixel_6105/VBIAS pixel_6105/NB2 pixel_6105/AMP_IN pixel_6105/SF_IB
+ pixel_6105/PIX_OUT pixel_6105/CSA_VREF pixel
Xpixel_6116 pixel_6116/gring pixel_6116/VDD pixel_6116/GND pixel_6116/VREF pixel_6116/ROW_SEL
+ pixel_6116/NB1 pixel_6116/VBIAS pixel_6116/NB2 pixel_6116/AMP_IN pixel_6116/SF_IB
+ pixel_6116/PIX_OUT pixel_6116/CSA_VREF pixel
Xpixel_6127 pixel_6127/gring pixel_6127/VDD pixel_6127/GND pixel_6127/VREF pixel_6127/ROW_SEL
+ pixel_6127/NB1 pixel_6127/VBIAS pixel_6127/NB2 pixel_6127/AMP_IN pixel_6127/SF_IB
+ pixel_6127/PIX_OUT pixel_6127/CSA_VREF pixel
Xpixel_6138 pixel_6138/gring pixel_6138/VDD pixel_6138/GND pixel_6138/VREF pixel_6138/ROW_SEL
+ pixel_6138/NB1 pixel_6138/VBIAS pixel_6138/NB2 pixel_6138/AMP_IN pixel_6138/SF_IB
+ pixel_6138/PIX_OUT pixel_6138/CSA_VREF pixel
Xpixel_6149 pixel_6149/gring pixel_6149/VDD pixel_6149/GND pixel_6149/VREF pixel_6149/ROW_SEL
+ pixel_6149/NB1 pixel_6149/VBIAS pixel_6149/NB2 pixel_6149/AMP_IN pixel_6149/SF_IB
+ pixel_6149/PIX_OUT pixel_6149/CSA_VREF pixel
Xpixel_5404 pixel_5404/gring pixel_5404/VDD pixel_5404/GND pixel_5404/VREF pixel_5404/ROW_SEL
+ pixel_5404/NB1 pixel_5404/VBIAS pixel_5404/NB2 pixel_5404/AMP_IN pixel_5404/SF_IB
+ pixel_5404/PIX_OUT pixel_5404/CSA_VREF pixel
Xpixel_5415 pixel_5415/gring pixel_5415/VDD pixel_5415/GND pixel_5415/VREF pixel_5415/ROW_SEL
+ pixel_5415/NB1 pixel_5415/VBIAS pixel_5415/NB2 pixel_5415/AMP_IN pixel_5415/SF_IB
+ pixel_5415/PIX_OUT pixel_5415/CSA_VREF pixel
Xpixel_5426 pixel_5426/gring pixel_5426/VDD pixel_5426/GND pixel_5426/VREF pixel_5426/ROW_SEL
+ pixel_5426/NB1 pixel_5426/VBIAS pixel_5426/NB2 pixel_5426/AMP_IN pixel_5426/SF_IB
+ pixel_5426/PIX_OUT pixel_5426/CSA_VREF pixel
Xpixel_5437 pixel_5437/gring pixel_5437/VDD pixel_5437/GND pixel_5437/VREF pixel_5437/ROW_SEL
+ pixel_5437/NB1 pixel_5437/VBIAS pixel_5437/NB2 pixel_5437/AMP_IN pixel_5437/SF_IB
+ pixel_5437/PIX_OUT pixel_5437/CSA_VREF pixel
Xpixel_5448 pixel_5448/gring pixel_5448/VDD pixel_5448/GND pixel_5448/VREF pixel_5448/ROW_SEL
+ pixel_5448/NB1 pixel_5448/VBIAS pixel_5448/NB2 pixel_5448/AMP_IN pixel_5448/SF_IB
+ pixel_5448/PIX_OUT pixel_5448/CSA_VREF pixel
Xpixel_4703 pixel_4703/gring pixel_4703/VDD pixel_4703/GND pixel_4703/VREF pixel_4703/ROW_SEL
+ pixel_4703/NB1 pixel_4703/VBIAS pixel_4703/NB2 pixel_4703/AMP_IN pixel_4703/SF_IB
+ pixel_4703/PIX_OUT pixel_4703/CSA_VREF pixel
Xpixel_742 pixel_742/gring pixel_742/VDD pixel_742/GND pixel_742/VREF pixel_742/ROW_SEL
+ pixel_742/NB1 pixel_742/VBIAS pixel_742/NB2 pixel_742/AMP_IN pixel_742/SF_IB pixel_742/PIX_OUT
+ pixel_742/CSA_VREF pixel
Xpixel_731 pixel_731/gring pixel_731/VDD pixel_731/GND pixel_731/VREF pixel_731/ROW_SEL
+ pixel_731/NB1 pixel_731/VBIAS pixel_731/NB2 pixel_731/AMP_IN pixel_731/SF_IB pixel_731/PIX_OUT
+ pixel_731/CSA_VREF pixel
Xpixel_720 pixel_720/gring pixel_720/VDD pixel_720/GND pixel_720/VREF pixel_720/ROW_SEL
+ pixel_720/NB1 pixel_720/VBIAS pixel_720/NB2 pixel_720/AMP_IN pixel_720/SF_IB pixel_720/PIX_OUT
+ pixel_720/CSA_VREF pixel
Xpixel_5459 pixel_5459/gring pixel_5459/VDD pixel_5459/GND pixel_5459/VREF pixel_5459/ROW_SEL
+ pixel_5459/NB1 pixel_5459/VBIAS pixel_5459/NB2 pixel_5459/AMP_IN pixel_5459/SF_IB
+ pixel_5459/PIX_OUT pixel_5459/CSA_VREF pixel
Xpixel_4714 pixel_4714/gring pixel_4714/VDD pixel_4714/GND pixel_4714/VREF pixel_4714/ROW_SEL
+ pixel_4714/NB1 pixel_4714/VBIAS pixel_4714/NB2 pixel_4714/AMP_IN pixel_4714/SF_IB
+ pixel_4714/PIX_OUT pixel_4714/CSA_VREF pixel
Xpixel_4725 pixel_4725/gring pixel_4725/VDD pixel_4725/GND pixel_4725/VREF pixel_4725/ROW_SEL
+ pixel_4725/NB1 pixel_4725/VBIAS pixel_4725/NB2 pixel_4725/AMP_IN pixel_4725/SF_IB
+ pixel_4725/PIX_OUT pixel_4725/CSA_VREF pixel
Xpixel_4736 pixel_4736/gring pixel_4736/VDD pixel_4736/GND pixel_4736/VREF pixel_4736/ROW_SEL
+ pixel_4736/NB1 pixel_4736/VBIAS pixel_4736/NB2 pixel_4736/AMP_IN pixel_4736/SF_IB
+ pixel_4736/PIX_OUT pixel_4736/CSA_VREF pixel
Xpixel_775 pixel_775/gring pixel_775/VDD pixel_775/GND pixel_775/VREF pixel_775/ROW_SEL
+ pixel_775/NB1 pixel_775/VBIAS pixel_775/NB2 pixel_775/AMP_IN pixel_775/SF_IB pixel_775/PIX_OUT
+ pixel_775/CSA_VREF pixel
Xpixel_764 pixel_764/gring pixel_764/VDD pixel_764/GND pixel_764/VREF pixel_764/ROW_SEL
+ pixel_764/NB1 pixel_764/VBIAS pixel_764/NB2 pixel_764/AMP_IN pixel_764/SF_IB pixel_764/PIX_OUT
+ pixel_764/CSA_VREF pixel
Xpixel_753 pixel_753/gring pixel_753/VDD pixel_753/GND pixel_753/VREF pixel_753/ROW_SEL
+ pixel_753/NB1 pixel_753/VBIAS pixel_753/NB2 pixel_753/AMP_IN pixel_753/SF_IB pixel_753/PIX_OUT
+ pixel_753/CSA_VREF pixel
Xpixel_4747 pixel_4747/gring pixel_4747/VDD pixel_4747/GND pixel_4747/VREF pixel_4747/ROW_SEL
+ pixel_4747/NB1 pixel_4747/VBIAS pixel_4747/NB2 pixel_4747/AMP_IN pixel_4747/SF_IB
+ pixel_4747/PIX_OUT pixel_4747/CSA_VREF pixel
Xpixel_4758 pixel_4758/gring pixel_4758/VDD pixel_4758/GND pixel_4758/VREF pixel_4758/ROW_SEL
+ pixel_4758/NB1 pixel_4758/VBIAS pixel_4758/NB2 pixel_4758/AMP_IN pixel_4758/SF_IB
+ pixel_4758/PIX_OUT pixel_4758/CSA_VREF pixel
Xpixel_4769 pixel_4769/gring pixel_4769/VDD pixel_4769/GND pixel_4769/VREF pixel_4769/ROW_SEL
+ pixel_4769/NB1 pixel_4769/VBIAS pixel_4769/NB2 pixel_4769/AMP_IN pixel_4769/SF_IB
+ pixel_4769/PIX_OUT pixel_4769/CSA_VREF pixel
Xpixel_797 pixel_797/gring pixel_797/VDD pixel_797/GND pixel_797/VREF pixel_797/ROW_SEL
+ pixel_797/NB1 pixel_797/VBIAS pixel_797/NB2 pixel_797/AMP_IN pixel_797/SF_IB pixel_797/PIX_OUT
+ pixel_797/CSA_VREF pixel
Xpixel_786 pixel_786/gring pixel_786/VDD pixel_786/GND pixel_786/VREF pixel_786/ROW_SEL
+ pixel_786/NB1 pixel_786/VBIAS pixel_786/NB2 pixel_786/AMP_IN pixel_786/SF_IB pixel_786/PIX_OUT
+ pixel_786/CSA_VREF pixel
Xpixel_8030 pixel_8030/gring pixel_8030/VDD pixel_8030/GND pixel_8030/VREF pixel_8030/ROW_SEL
+ pixel_8030/NB1 pixel_8030/VBIAS pixel_8030/NB2 pixel_8030/AMP_IN pixel_8030/SF_IB
+ pixel_8030/PIX_OUT pixel_8030/CSA_VREF pixel
Xpixel_8041 pixel_8041/gring pixel_8041/VDD pixel_8041/GND pixel_8041/VREF pixel_8041/ROW_SEL
+ pixel_8041/NB1 pixel_8041/VBIAS pixel_8041/NB2 pixel_8041/AMP_IN pixel_8041/SF_IB
+ pixel_8041/PIX_OUT pixel_8041/CSA_VREF pixel
Xpixel_8052 pixel_8052/gring pixel_8052/VDD pixel_8052/GND pixel_8052/VREF pixel_8052/ROW_SEL
+ pixel_8052/NB1 pixel_8052/VBIAS pixel_8052/NB2 pixel_8052/AMP_IN pixel_8052/SF_IB
+ pixel_8052/PIX_OUT pixel_8052/CSA_VREF pixel
Xpixel_8063 pixel_8063/gring pixel_8063/VDD pixel_8063/GND pixel_8063/VREF pixel_8063/ROW_SEL
+ pixel_8063/NB1 pixel_8063/VBIAS pixel_8063/NB2 pixel_8063/AMP_IN pixel_8063/SF_IB
+ pixel_8063/PIX_OUT pixel_8063/CSA_VREF pixel
Xpixel_8074 pixel_8074/gring pixel_8074/VDD pixel_8074/GND pixel_8074/VREF pixel_8074/ROW_SEL
+ pixel_8074/NB1 pixel_8074/VBIAS pixel_8074/NB2 pixel_8074/AMP_IN pixel_8074/SF_IB
+ pixel_8074/PIX_OUT pixel_8074/CSA_VREF pixel
Xpixel_8085 pixel_8085/gring pixel_8085/VDD pixel_8085/GND pixel_8085/VREF pixel_8085/ROW_SEL
+ pixel_8085/NB1 pixel_8085/VBIAS pixel_8085/NB2 pixel_8085/AMP_IN pixel_8085/SF_IB
+ pixel_8085/PIX_OUT pixel_8085/CSA_VREF pixel
Xpixel_7340 pixel_7340/gring pixel_7340/VDD pixel_7340/GND pixel_7340/VREF pixel_7340/ROW_SEL
+ pixel_7340/NB1 pixel_7340/VBIAS pixel_7340/NB2 pixel_7340/AMP_IN pixel_7340/SF_IB
+ pixel_7340/PIX_OUT pixel_7340/CSA_VREF pixel
Xpixel_8096 pixel_8096/gring pixel_8096/VDD pixel_8096/GND pixel_8096/VREF pixel_8096/ROW_SEL
+ pixel_8096/NB1 pixel_8096/VBIAS pixel_8096/NB2 pixel_8096/AMP_IN pixel_8096/SF_IB
+ pixel_8096/PIX_OUT pixel_8096/CSA_VREF pixel
Xpixel_7351 pixel_7351/gring pixel_7351/VDD pixel_7351/GND pixel_7351/VREF pixel_7351/ROW_SEL
+ pixel_7351/NB1 pixel_7351/VBIAS pixel_7351/NB2 pixel_7351/AMP_IN pixel_7351/SF_IB
+ pixel_7351/PIX_OUT pixel_7351/CSA_VREF pixel
Xpixel_7362 pixel_7362/gring pixel_7362/VDD pixel_7362/GND pixel_7362/VREF pixel_7362/ROW_SEL
+ pixel_7362/NB1 pixel_7362/VBIAS pixel_7362/NB2 pixel_7362/AMP_IN pixel_7362/SF_IB
+ pixel_7362/PIX_OUT pixel_7362/CSA_VREF pixel
Xpixel_7373 pixel_7373/gring pixel_7373/VDD pixel_7373/GND pixel_7373/VREF pixel_7373/ROW_SEL
+ pixel_7373/NB1 pixel_7373/VBIAS pixel_7373/NB2 pixel_7373/AMP_IN pixel_7373/SF_IB
+ pixel_7373/PIX_OUT pixel_7373/CSA_VREF pixel
Xpixel_7384 pixel_7384/gring pixel_7384/VDD pixel_7384/GND pixel_7384/VREF pixel_7384/ROW_SEL
+ pixel_7384/NB1 pixel_7384/VBIAS pixel_7384/NB2 pixel_7384/AMP_IN pixel_7384/SF_IB
+ pixel_7384/PIX_OUT pixel_7384/CSA_VREF pixel
Xpixel_7395 pixel_7395/gring pixel_7395/VDD pixel_7395/GND pixel_7395/VREF pixel_7395/ROW_SEL
+ pixel_7395/NB1 pixel_7395/VBIAS pixel_7395/NB2 pixel_7395/AMP_IN pixel_7395/SF_IB
+ pixel_7395/PIX_OUT pixel_7395/CSA_VREF pixel
Xpixel_6650 pixel_6650/gring pixel_6650/VDD pixel_6650/GND pixel_6650/VREF pixel_6650/ROW_SEL
+ pixel_6650/NB1 pixel_6650/VBIAS pixel_6650/NB2 pixel_6650/AMP_IN pixel_6650/SF_IB
+ pixel_6650/PIX_OUT pixel_6650/CSA_VREF pixel
Xpixel_6661 pixel_6661/gring pixel_6661/VDD pixel_6661/GND pixel_6661/VREF pixel_6661/ROW_SEL
+ pixel_6661/NB1 pixel_6661/VBIAS pixel_6661/NB2 pixel_6661/AMP_IN pixel_6661/SF_IB
+ pixel_6661/PIX_OUT pixel_6661/CSA_VREF pixel
Xpixel_6672 pixel_6672/gring pixel_6672/VDD pixel_6672/GND pixel_6672/VREF pixel_6672/ROW_SEL
+ pixel_6672/NB1 pixel_6672/VBIAS pixel_6672/NB2 pixel_6672/AMP_IN pixel_6672/SF_IB
+ pixel_6672/PIX_OUT pixel_6672/CSA_VREF pixel
Xpixel_6683 pixel_6683/gring pixel_6683/VDD pixel_6683/GND pixel_6683/VREF pixel_6683/ROW_SEL
+ pixel_6683/NB1 pixel_6683/VBIAS pixel_6683/NB2 pixel_6683/AMP_IN pixel_6683/SF_IB
+ pixel_6683/PIX_OUT pixel_6683/CSA_VREF pixel
Xpixel_6694 pixel_6694/gring pixel_6694/VDD pixel_6694/GND pixel_6694/VREF pixel_6694/ROW_SEL
+ pixel_6694/NB1 pixel_6694/VBIAS pixel_6694/NB2 pixel_6694/AMP_IN pixel_6694/SF_IB
+ pixel_6694/PIX_OUT pixel_6694/CSA_VREF pixel
Xpixel_5960 pixel_5960/gring pixel_5960/VDD pixel_5960/GND pixel_5960/VREF pixel_5960/ROW_SEL
+ pixel_5960/NB1 pixel_5960/VBIAS pixel_5960/NB2 pixel_5960/AMP_IN pixel_5960/SF_IB
+ pixel_5960/PIX_OUT pixel_5960/CSA_VREF pixel
Xpixel_5971 pixel_5971/gring pixel_5971/VDD pixel_5971/GND pixel_5971/VREF pixel_5971/ROW_SEL
+ pixel_5971/NB1 pixel_5971/VBIAS pixel_5971/NB2 pixel_5971/AMP_IN pixel_5971/SF_IB
+ pixel_5971/PIX_OUT pixel_5971/CSA_VREF pixel
Xpixel_5982 pixel_5982/gring pixel_5982/VDD pixel_5982/GND pixel_5982/VREF pixel_5982/ROW_SEL
+ pixel_5982/NB1 pixel_5982/VBIAS pixel_5982/NB2 pixel_5982/AMP_IN pixel_5982/SF_IB
+ pixel_5982/PIX_OUT pixel_5982/CSA_VREF pixel
Xpixel_5993 pixel_5993/gring pixel_5993/VDD pixel_5993/GND pixel_5993/VREF pixel_5993/ROW_SEL
+ pixel_5993/NB1 pixel_5993/VBIAS pixel_5993/NB2 pixel_5993/AMP_IN pixel_5993/SF_IB
+ pixel_5993/PIX_OUT pixel_5993/CSA_VREF pixel
Xpixel_3309 pixel_3309/gring pixel_3309/VDD pixel_3309/GND pixel_3309/VREF pixel_3309/ROW_SEL
+ pixel_3309/NB1 pixel_3309/VBIAS pixel_3309/NB2 pixel_3309/AMP_IN pixel_3309/SF_IB
+ pixel_3309/PIX_OUT pixel_3309/CSA_VREF pixel
Xpixel_2619 pixel_2619/gring pixel_2619/VDD pixel_2619/GND pixel_2619/VREF pixel_2619/ROW_SEL
+ pixel_2619/NB1 pixel_2619/VBIAS pixel_2619/NB2 pixel_2619/AMP_IN pixel_2619/SF_IB
+ pixel_2619/PIX_OUT pixel_2619/CSA_VREF pixel
Xpixel_2608 pixel_2608/gring pixel_2608/VDD pixel_2608/GND pixel_2608/VREF pixel_2608/ROW_SEL
+ pixel_2608/NB1 pixel_2608/VBIAS pixel_2608/NB2 pixel_2608/AMP_IN pixel_2608/SF_IB
+ pixel_2608/PIX_OUT pixel_2608/CSA_VREF pixel
Xpixel_1907 pixel_1907/gring pixel_1907/VDD pixel_1907/GND pixel_1907/VREF pixel_1907/ROW_SEL
+ pixel_1907/NB1 pixel_1907/VBIAS pixel_1907/NB2 pixel_1907/AMP_IN pixel_1907/SF_IB
+ pixel_1907/PIX_OUT pixel_1907/CSA_VREF pixel
Xpixel_1929 pixel_1929/gring pixel_1929/VDD pixel_1929/GND pixel_1929/VREF pixel_1929/ROW_SEL
+ pixel_1929/NB1 pixel_1929/VBIAS pixel_1929/NB2 pixel_1929/AMP_IN pixel_1929/SF_IB
+ pixel_1929/PIX_OUT pixel_1929/CSA_VREF pixel
Xpixel_1918 pixel_1918/gring pixel_1918/VDD pixel_1918/GND pixel_1918/VREF pixel_1918/ROW_SEL
+ pixel_1918/NB1 pixel_1918/VBIAS pixel_1918/NB2 pixel_1918/AMP_IN pixel_1918/SF_IB
+ pixel_1918/PIX_OUT pixel_1918/CSA_VREF pixel
Xpixel_5201 pixel_5201/gring pixel_5201/VDD pixel_5201/GND pixel_5201/VREF pixel_5201/ROW_SEL
+ pixel_5201/NB1 pixel_5201/VBIAS pixel_5201/NB2 pixel_5201/AMP_IN pixel_5201/SF_IB
+ pixel_5201/PIX_OUT pixel_5201/CSA_VREF pixel
Xpixel_5212 pixel_5212/gring pixel_5212/VDD pixel_5212/GND pixel_5212/VREF pixel_5212/ROW_SEL
+ pixel_5212/NB1 pixel_5212/VBIAS pixel_5212/NB2 pixel_5212/AMP_IN pixel_5212/SF_IB
+ pixel_5212/PIX_OUT pixel_5212/CSA_VREF pixel
Xpixel_5223 pixel_5223/gring pixel_5223/VDD pixel_5223/GND pixel_5223/VREF pixel_5223/ROW_SEL
+ pixel_5223/NB1 pixel_5223/VBIAS pixel_5223/NB2 pixel_5223/AMP_IN pixel_5223/SF_IB
+ pixel_5223/PIX_OUT pixel_5223/CSA_VREF pixel
Xpixel_5234 pixel_5234/gring pixel_5234/VDD pixel_5234/GND pixel_5234/VREF pixel_5234/ROW_SEL
+ pixel_5234/NB1 pixel_5234/VBIAS pixel_5234/NB2 pixel_5234/AMP_IN pixel_5234/SF_IB
+ pixel_5234/PIX_OUT pixel_5234/CSA_VREF pixel
Xpixel_5245 pixel_5245/gring pixel_5245/VDD pixel_5245/GND pixel_5245/VREF pixel_5245/ROW_SEL
+ pixel_5245/NB1 pixel_5245/VBIAS pixel_5245/NB2 pixel_5245/AMP_IN pixel_5245/SF_IB
+ pixel_5245/PIX_OUT pixel_5245/CSA_VREF pixel
Xpixel_5256 pixel_5256/gring pixel_5256/VDD pixel_5256/GND pixel_5256/VREF pixel_5256/ROW_SEL
+ pixel_5256/NB1 pixel_5256/VBIAS pixel_5256/NB2 pixel_5256/AMP_IN pixel_5256/SF_IB
+ pixel_5256/PIX_OUT pixel_5256/CSA_VREF pixel
Xpixel_4500 pixel_4500/gring pixel_4500/VDD pixel_4500/GND pixel_4500/VREF pixel_4500/ROW_SEL
+ pixel_4500/NB1 pixel_4500/VBIAS pixel_4500/NB2 pixel_4500/AMP_IN pixel_4500/SF_IB
+ pixel_4500/PIX_OUT pixel_4500/CSA_VREF pixel
Xpixel_4511 pixel_4511/gring pixel_4511/VDD pixel_4511/GND pixel_4511/VREF pixel_4511/ROW_SEL
+ pixel_4511/NB1 pixel_4511/VBIAS pixel_4511/NB2 pixel_4511/AMP_IN pixel_4511/SF_IB
+ pixel_4511/PIX_OUT pixel_4511/CSA_VREF pixel
Xpixel_550 pixel_550/gring pixel_550/VDD pixel_550/GND pixel_550/VREF pixel_550/ROW_SEL
+ pixel_550/NB1 pixel_550/VBIAS pixel_550/NB2 pixel_550/AMP_IN pixel_550/SF_IB pixel_550/PIX_OUT
+ pixel_550/CSA_VREF pixel
Xpixel_5267 pixel_5267/gring pixel_5267/VDD pixel_5267/GND pixel_5267/VREF pixel_5267/ROW_SEL
+ pixel_5267/NB1 pixel_5267/VBIAS pixel_5267/NB2 pixel_5267/AMP_IN pixel_5267/SF_IB
+ pixel_5267/PIX_OUT pixel_5267/CSA_VREF pixel
Xpixel_5278 pixel_5278/gring pixel_5278/VDD pixel_5278/GND pixel_5278/VREF pixel_5278/ROW_SEL
+ pixel_5278/NB1 pixel_5278/VBIAS pixel_5278/NB2 pixel_5278/AMP_IN pixel_5278/SF_IB
+ pixel_5278/PIX_OUT pixel_5278/CSA_VREF pixel
Xpixel_5289 pixel_5289/gring pixel_5289/VDD pixel_5289/GND pixel_5289/VREF pixel_5289/ROW_SEL
+ pixel_5289/NB1 pixel_5289/VBIAS pixel_5289/NB2 pixel_5289/AMP_IN pixel_5289/SF_IB
+ pixel_5289/PIX_OUT pixel_5289/CSA_VREF pixel
Xpixel_4522 pixel_4522/gring pixel_4522/VDD pixel_4522/GND pixel_4522/VREF pixel_4522/ROW_SEL
+ pixel_4522/NB1 pixel_4522/VBIAS pixel_4522/NB2 pixel_4522/AMP_IN pixel_4522/SF_IB
+ pixel_4522/PIX_OUT pixel_4522/CSA_VREF pixel
Xpixel_4533 pixel_4533/gring pixel_4533/VDD pixel_4533/GND pixel_4533/VREF pixel_4533/ROW_SEL
+ pixel_4533/NB1 pixel_4533/VBIAS pixel_4533/NB2 pixel_4533/AMP_IN pixel_4533/SF_IB
+ pixel_4533/PIX_OUT pixel_4533/CSA_VREF pixel
Xpixel_4544 pixel_4544/gring pixel_4544/VDD pixel_4544/GND pixel_4544/VREF pixel_4544/ROW_SEL
+ pixel_4544/NB1 pixel_4544/VBIAS pixel_4544/NB2 pixel_4544/AMP_IN pixel_4544/SF_IB
+ pixel_4544/PIX_OUT pixel_4544/CSA_VREF pixel
Xpixel_4555 pixel_4555/gring pixel_4555/VDD pixel_4555/GND pixel_4555/VREF pixel_4555/ROW_SEL
+ pixel_4555/NB1 pixel_4555/VBIAS pixel_4555/NB2 pixel_4555/AMP_IN pixel_4555/SF_IB
+ pixel_4555/PIX_OUT pixel_4555/CSA_VREF pixel
Xpixel_3810 pixel_3810/gring pixel_3810/VDD pixel_3810/GND pixel_3810/VREF pixel_3810/ROW_SEL
+ pixel_3810/NB1 pixel_3810/VBIAS pixel_3810/NB2 pixel_3810/AMP_IN pixel_3810/SF_IB
+ pixel_3810/PIX_OUT pixel_3810/CSA_VREF pixel
Xpixel_583 pixel_583/gring pixel_583/VDD pixel_583/GND pixel_583/VREF pixel_583/ROW_SEL
+ pixel_583/NB1 pixel_583/VBIAS pixel_583/NB2 pixel_583/AMP_IN pixel_583/SF_IB pixel_583/PIX_OUT
+ pixel_583/CSA_VREF pixel
Xpixel_572 pixel_572/gring pixel_572/VDD pixel_572/GND pixel_572/VREF pixel_572/ROW_SEL
+ pixel_572/NB1 pixel_572/VBIAS pixel_572/NB2 pixel_572/AMP_IN pixel_572/SF_IB pixel_572/PIX_OUT
+ pixel_572/CSA_VREF pixel
Xpixel_561 pixel_561/gring pixel_561/VDD pixel_561/GND pixel_561/VREF pixel_561/ROW_SEL
+ pixel_561/NB1 pixel_561/VBIAS pixel_561/NB2 pixel_561/AMP_IN pixel_561/SF_IB pixel_561/PIX_OUT
+ pixel_561/CSA_VREF pixel
Xpixel_4566 pixel_4566/gring pixel_4566/VDD pixel_4566/GND pixel_4566/VREF pixel_4566/ROW_SEL
+ pixel_4566/NB1 pixel_4566/VBIAS pixel_4566/NB2 pixel_4566/AMP_IN pixel_4566/SF_IB
+ pixel_4566/PIX_OUT pixel_4566/CSA_VREF pixel
Xpixel_4577 pixel_4577/gring pixel_4577/VDD pixel_4577/GND pixel_4577/VREF pixel_4577/ROW_SEL
+ pixel_4577/NB1 pixel_4577/VBIAS pixel_4577/NB2 pixel_4577/AMP_IN pixel_4577/SF_IB
+ pixel_4577/PIX_OUT pixel_4577/CSA_VREF pixel
Xpixel_4588 pixel_4588/gring pixel_4588/VDD pixel_4588/GND pixel_4588/VREF pixel_4588/ROW_SEL
+ pixel_4588/NB1 pixel_4588/VBIAS pixel_4588/NB2 pixel_4588/AMP_IN pixel_4588/SF_IB
+ pixel_4588/PIX_OUT pixel_4588/CSA_VREF pixel
Xpixel_3821 pixel_3821/gring pixel_3821/VDD pixel_3821/GND pixel_3821/VREF pixel_3821/ROW_SEL
+ pixel_3821/NB1 pixel_3821/VBIAS pixel_3821/NB2 pixel_3821/AMP_IN pixel_3821/SF_IB
+ pixel_3821/PIX_OUT pixel_3821/CSA_VREF pixel
Xpixel_3832 pixel_3832/gring pixel_3832/VDD pixel_3832/GND pixel_3832/VREF pixel_3832/ROW_SEL
+ pixel_3832/NB1 pixel_3832/VBIAS pixel_3832/NB2 pixel_3832/AMP_IN pixel_3832/SF_IB
+ pixel_3832/PIX_OUT pixel_3832/CSA_VREF pixel
Xpixel_3843 pixel_3843/gring pixel_3843/VDD pixel_3843/GND pixel_3843/VREF pixel_3843/ROW_SEL
+ pixel_3843/NB1 pixel_3843/VBIAS pixel_3843/NB2 pixel_3843/AMP_IN pixel_3843/SF_IB
+ pixel_3843/PIX_OUT pixel_3843/CSA_VREF pixel
Xpixel_594 pixel_594/gring pixel_594/VDD pixel_594/GND pixel_594/VREF pixel_594/ROW_SEL
+ pixel_594/NB1 pixel_594/VBIAS pixel_594/NB2 pixel_594/AMP_IN pixel_594/SF_IB pixel_594/PIX_OUT
+ pixel_594/CSA_VREF pixel
Xpixel_3876 pixel_3876/gring pixel_3876/VDD pixel_3876/GND pixel_3876/VREF pixel_3876/ROW_SEL
+ pixel_3876/NB1 pixel_3876/VBIAS pixel_3876/NB2 pixel_3876/AMP_IN pixel_3876/SF_IB
+ pixel_3876/PIX_OUT pixel_3876/CSA_VREF pixel
Xpixel_3865 pixel_3865/gring pixel_3865/VDD pixel_3865/GND pixel_3865/VREF pixel_3865/ROW_SEL
+ pixel_3865/NB1 pixel_3865/VBIAS pixel_3865/NB2 pixel_3865/AMP_IN pixel_3865/SF_IB
+ pixel_3865/PIX_OUT pixel_3865/CSA_VREF pixel
Xpixel_3854 pixel_3854/gring pixel_3854/VDD pixel_3854/GND pixel_3854/VREF pixel_3854/ROW_SEL
+ pixel_3854/NB1 pixel_3854/VBIAS pixel_3854/NB2 pixel_3854/AMP_IN pixel_3854/SF_IB
+ pixel_3854/PIX_OUT pixel_3854/CSA_VREF pixel
Xpixel_4599 pixel_4599/gring pixel_4599/VDD pixel_4599/GND pixel_4599/VREF pixel_4599/ROW_SEL
+ pixel_4599/NB1 pixel_4599/VBIAS pixel_4599/NB2 pixel_4599/AMP_IN pixel_4599/SF_IB
+ pixel_4599/PIX_OUT pixel_4599/CSA_VREF pixel
Xpixel_3898 pixel_3898/gring pixel_3898/VDD pixel_3898/GND pixel_3898/VREF pixel_3898/ROW_SEL
+ pixel_3898/NB1 pixel_3898/VBIAS pixel_3898/NB2 pixel_3898/AMP_IN pixel_3898/SF_IB
+ pixel_3898/PIX_OUT pixel_3898/CSA_VREF pixel
Xpixel_3887 pixel_3887/gring pixel_3887/VDD pixel_3887/GND pixel_3887/VREF pixel_3887/ROW_SEL
+ pixel_3887/NB1 pixel_3887/VBIAS pixel_3887/NB2 pixel_3887/AMP_IN pixel_3887/SF_IB
+ pixel_3887/PIX_OUT pixel_3887/CSA_VREF pixel
Xpixel_7170 pixel_7170/gring pixel_7170/VDD pixel_7170/GND pixel_7170/VREF pixel_7170/ROW_SEL
+ pixel_7170/NB1 pixel_7170/VBIAS pixel_7170/NB2 pixel_7170/AMP_IN pixel_7170/SF_IB
+ pixel_7170/PIX_OUT pixel_7170/CSA_VREF pixel
Xpixel_7181 pixel_7181/gring pixel_7181/VDD pixel_7181/GND pixel_7181/VREF pixel_7181/ROW_SEL
+ pixel_7181/NB1 pixel_7181/VBIAS pixel_7181/NB2 pixel_7181/AMP_IN pixel_7181/SF_IB
+ pixel_7181/PIX_OUT pixel_7181/CSA_VREF pixel
Xpixel_7192 pixel_7192/gring pixel_7192/VDD pixel_7192/GND pixel_7192/VREF pixel_7192/ROW_SEL
+ pixel_7192/NB1 pixel_7192/VBIAS pixel_7192/NB2 pixel_7192/AMP_IN pixel_7192/SF_IB
+ pixel_7192/PIX_OUT pixel_7192/CSA_VREF pixel
Xpixel_6480 pixel_6480/gring pixel_6480/VDD pixel_6480/GND pixel_6480/VREF pixel_6480/ROW_SEL
+ pixel_6480/NB1 pixel_6480/VBIAS pixel_6480/NB2 pixel_6480/AMP_IN pixel_6480/SF_IB
+ pixel_6480/PIX_OUT pixel_6480/CSA_VREF pixel
Xpixel_6491 pixel_6491/gring pixel_6491/VDD pixel_6491/GND pixel_6491/VREF pixel_6491/ROW_SEL
+ pixel_6491/NB1 pixel_6491/VBIAS pixel_6491/NB2 pixel_6491/AMP_IN pixel_6491/SF_IB
+ pixel_6491/PIX_OUT pixel_6491/CSA_VREF pixel
Xpixel_5790 pixel_5790/gring pixel_5790/VDD pixel_5790/GND pixel_5790/VREF pixel_5790/ROW_SEL
+ pixel_5790/NB1 pixel_5790/VBIAS pixel_5790/NB2 pixel_5790/AMP_IN pixel_5790/SF_IB
+ pixel_5790/PIX_OUT pixel_5790/CSA_VREF pixel
Xpixel_3139 pixel_3139/gring pixel_3139/VDD pixel_3139/GND pixel_3139/VREF pixel_3139/ROW_SEL
+ pixel_3139/NB1 pixel_3139/VBIAS pixel_3139/NB2 pixel_3139/AMP_IN pixel_3139/SF_IB
+ pixel_3139/PIX_OUT pixel_3139/CSA_VREF pixel
Xpixel_3128 pixel_3128/gring pixel_3128/VDD pixel_3128/GND pixel_3128/VREF pixel_3128/ROW_SEL
+ pixel_3128/NB1 pixel_3128/VBIAS pixel_3128/NB2 pixel_3128/AMP_IN pixel_3128/SF_IB
+ pixel_3128/PIX_OUT pixel_3128/CSA_VREF pixel
Xpixel_3117 pixel_3117/gring pixel_3117/VDD pixel_3117/GND pixel_3117/VREF pixel_3117/ROW_SEL
+ pixel_3117/NB1 pixel_3117/VBIAS pixel_3117/NB2 pixel_3117/AMP_IN pixel_3117/SF_IB
+ pixel_3117/PIX_OUT pixel_3117/CSA_VREF pixel
Xpixel_3106 pixel_3106/gring pixel_3106/VDD pixel_3106/GND pixel_3106/VREF pixel_3106/ROW_SEL
+ pixel_3106/NB1 pixel_3106/VBIAS pixel_3106/NB2 pixel_3106/AMP_IN pixel_3106/SF_IB
+ pixel_3106/PIX_OUT pixel_3106/CSA_VREF pixel
Xpixel_2427 pixel_2427/gring pixel_2427/VDD pixel_2427/GND pixel_2427/VREF pixel_2427/ROW_SEL
+ pixel_2427/NB1 pixel_2427/VBIAS pixel_2427/NB2 pixel_2427/AMP_IN pixel_2427/SF_IB
+ pixel_2427/PIX_OUT pixel_2427/CSA_VREF pixel
Xpixel_2416 pixel_2416/gring pixel_2416/VDD pixel_2416/GND pixel_2416/VREF pixel_2416/ROW_SEL
+ pixel_2416/NB1 pixel_2416/VBIAS pixel_2416/NB2 pixel_2416/AMP_IN pixel_2416/SF_IB
+ pixel_2416/PIX_OUT pixel_2416/CSA_VREF pixel
Xpixel_2405 pixel_2405/gring pixel_2405/VDD pixel_2405/GND pixel_2405/VREF pixel_2405/ROW_SEL
+ pixel_2405/NB1 pixel_2405/VBIAS pixel_2405/NB2 pixel_2405/AMP_IN pixel_2405/SF_IB
+ pixel_2405/PIX_OUT pixel_2405/CSA_VREF pixel
Xpixel_1726 pixel_1726/gring pixel_1726/VDD pixel_1726/GND pixel_1726/VREF pixel_1726/ROW_SEL
+ pixel_1726/NB1 pixel_1726/VBIAS pixel_1726/NB2 pixel_1726/AMP_IN pixel_1726/SF_IB
+ pixel_1726/PIX_OUT pixel_1726/CSA_VREF pixel
Xpixel_1715 pixel_1715/gring pixel_1715/VDD pixel_1715/GND pixel_1715/VREF pixel_1715/ROW_SEL
+ pixel_1715/NB1 pixel_1715/VBIAS pixel_1715/NB2 pixel_1715/AMP_IN pixel_1715/SF_IB
+ pixel_1715/PIX_OUT pixel_1715/CSA_VREF pixel
Xpixel_1704 pixel_1704/gring pixel_1704/VDD pixel_1704/GND pixel_1704/VREF pixel_1704/ROW_SEL
+ pixel_1704/NB1 pixel_1704/VBIAS pixel_1704/NB2 pixel_1704/AMP_IN pixel_1704/SF_IB
+ pixel_1704/PIX_OUT pixel_1704/CSA_VREF pixel
Xpixel_2449 pixel_2449/gring pixel_2449/VDD pixel_2449/GND pixel_2449/VREF pixel_2449/ROW_SEL
+ pixel_2449/NB1 pixel_2449/VBIAS pixel_2449/NB2 pixel_2449/AMP_IN pixel_2449/SF_IB
+ pixel_2449/PIX_OUT pixel_2449/CSA_VREF pixel
Xpixel_2438 pixel_2438/gring pixel_2438/VDD pixel_2438/GND pixel_2438/VREF pixel_2438/ROW_SEL
+ pixel_2438/NB1 pixel_2438/VBIAS pixel_2438/NB2 pixel_2438/AMP_IN pixel_2438/SF_IB
+ pixel_2438/PIX_OUT pixel_2438/CSA_VREF pixel
Xpixel_1759 pixel_1759/gring pixel_1759/VDD pixel_1759/GND pixel_1759/VREF pixel_1759/ROW_SEL
+ pixel_1759/NB1 pixel_1759/VBIAS pixel_1759/NB2 pixel_1759/AMP_IN pixel_1759/SF_IB
+ pixel_1759/PIX_OUT pixel_1759/CSA_VREF pixel
Xpixel_1748 pixel_1748/gring pixel_1748/VDD pixel_1748/GND pixel_1748/VREF pixel_1748/ROW_SEL
+ pixel_1748/NB1 pixel_1748/VBIAS pixel_1748/NB2 pixel_1748/AMP_IN pixel_1748/SF_IB
+ pixel_1748/PIX_OUT pixel_1748/CSA_VREF pixel
Xpixel_1737 pixel_1737/gring pixel_1737/VDD pixel_1737/GND pixel_1737/VREF pixel_1737/ROW_SEL
+ pixel_1737/NB1 pixel_1737/VBIAS pixel_1737/NB2 pixel_1737/AMP_IN pixel_1737/SF_IB
+ pixel_1737/PIX_OUT pixel_1737/CSA_VREF pixel
Xpixel_5020 pixel_5020/gring pixel_5020/VDD pixel_5020/GND pixel_5020/VREF pixel_5020/ROW_SEL
+ pixel_5020/NB1 pixel_5020/VBIAS pixel_5020/NB2 pixel_5020/AMP_IN pixel_5020/SF_IB
+ pixel_5020/PIX_OUT pixel_5020/CSA_VREF pixel
Xpixel_5031 pixel_5031/gring pixel_5031/VDD pixel_5031/GND pixel_5031/VREF pixel_5031/ROW_SEL
+ pixel_5031/NB1 pixel_5031/VBIAS pixel_5031/NB2 pixel_5031/AMP_IN pixel_5031/SF_IB
+ pixel_5031/PIX_OUT pixel_5031/CSA_VREF pixel
Xpixel_5042 pixel_5042/gring pixel_5042/VDD pixel_5042/GND pixel_5042/VREF pixel_5042/ROW_SEL
+ pixel_5042/NB1 pixel_5042/VBIAS pixel_5042/NB2 pixel_5042/AMP_IN pixel_5042/SF_IB
+ pixel_5042/PIX_OUT pixel_5042/CSA_VREF pixel
Xpixel_5053 pixel_5053/gring pixel_5053/VDD pixel_5053/GND pixel_5053/VREF pixel_5053/ROW_SEL
+ pixel_5053/NB1 pixel_5053/VBIAS pixel_5053/NB2 pixel_5053/AMP_IN pixel_5053/SF_IB
+ pixel_5053/PIX_OUT pixel_5053/CSA_VREF pixel
Xpixel_5064 pixel_5064/gring pixel_5064/VDD pixel_5064/GND pixel_5064/VREF pixel_5064/ROW_SEL
+ pixel_5064/NB1 pixel_5064/VBIAS pixel_5064/NB2 pixel_5064/AMP_IN pixel_5064/SF_IB
+ pixel_5064/PIX_OUT pixel_5064/CSA_VREF pixel
Xpixel_5075 pixel_5075/gring pixel_5075/VDD pixel_5075/GND pixel_5075/VREF pixel_5075/ROW_SEL
+ pixel_5075/NB1 pixel_5075/VBIAS pixel_5075/NB2 pixel_5075/AMP_IN pixel_5075/SF_IB
+ pixel_5075/PIX_OUT pixel_5075/CSA_VREF pixel
Xpixel_5086 pixel_5086/gring pixel_5086/VDD pixel_5086/GND pixel_5086/VREF pixel_5086/ROW_SEL
+ pixel_5086/NB1 pixel_5086/VBIAS pixel_5086/NB2 pixel_5086/AMP_IN pixel_5086/SF_IB
+ pixel_5086/PIX_OUT pixel_5086/CSA_VREF pixel
Xpixel_5097 pixel_5097/gring pixel_5097/VDD pixel_5097/GND pixel_5097/VREF pixel_5097/ROW_SEL
+ pixel_5097/NB1 pixel_5097/VBIAS pixel_5097/NB2 pixel_5097/AMP_IN pixel_5097/SF_IB
+ pixel_5097/PIX_OUT pixel_5097/CSA_VREF pixel
Xpixel_4330 pixel_4330/gring pixel_4330/VDD pixel_4330/GND pixel_4330/VREF pixel_4330/ROW_SEL
+ pixel_4330/NB1 pixel_4330/VBIAS pixel_4330/NB2 pixel_4330/AMP_IN pixel_4330/SF_IB
+ pixel_4330/PIX_OUT pixel_4330/CSA_VREF pixel
Xpixel_4341 pixel_4341/gring pixel_4341/VDD pixel_4341/GND pixel_4341/VREF pixel_4341/ROW_SEL
+ pixel_4341/NB1 pixel_4341/VBIAS pixel_4341/NB2 pixel_4341/AMP_IN pixel_4341/SF_IB
+ pixel_4341/PIX_OUT pixel_4341/CSA_VREF pixel
Xpixel_4352 pixel_4352/gring pixel_4352/VDD pixel_4352/GND pixel_4352/VREF pixel_4352/ROW_SEL
+ pixel_4352/NB1 pixel_4352/VBIAS pixel_4352/NB2 pixel_4352/AMP_IN pixel_4352/SF_IB
+ pixel_4352/PIX_OUT pixel_4352/CSA_VREF pixel
Xpixel_4363 pixel_4363/gring pixel_4363/VDD pixel_4363/GND pixel_4363/VREF pixel_4363/ROW_SEL
+ pixel_4363/NB1 pixel_4363/VBIAS pixel_4363/NB2 pixel_4363/AMP_IN pixel_4363/SF_IB
+ pixel_4363/PIX_OUT pixel_4363/CSA_VREF pixel
Xpixel_391 pixel_391/gring pixel_391/VDD pixel_391/GND pixel_391/VREF pixel_391/ROW_SEL
+ pixel_391/NB1 pixel_391/VBIAS pixel_391/NB2 pixel_391/AMP_IN pixel_391/SF_IB pixel_391/PIX_OUT
+ pixel_391/CSA_VREF pixel
Xpixel_380 pixel_380/gring pixel_380/VDD pixel_380/GND pixel_380/VREF pixel_380/ROW_SEL
+ pixel_380/NB1 pixel_380/VBIAS pixel_380/NB2 pixel_380/AMP_IN pixel_380/SF_IB pixel_380/PIX_OUT
+ pixel_380/CSA_VREF pixel
Xpixel_3651 pixel_3651/gring pixel_3651/VDD pixel_3651/GND pixel_3651/VREF pixel_3651/ROW_SEL
+ pixel_3651/NB1 pixel_3651/VBIAS pixel_3651/NB2 pixel_3651/AMP_IN pixel_3651/SF_IB
+ pixel_3651/PIX_OUT pixel_3651/CSA_VREF pixel
Xpixel_3640 pixel_3640/gring pixel_3640/VDD pixel_3640/GND pixel_3640/VREF pixel_3640/ROW_SEL
+ pixel_3640/NB1 pixel_3640/VBIAS pixel_3640/NB2 pixel_3640/AMP_IN pixel_3640/SF_IB
+ pixel_3640/PIX_OUT pixel_3640/CSA_VREF pixel
Xpixel_4374 pixel_4374/gring pixel_4374/VDD pixel_4374/GND pixel_4374/VREF pixel_4374/ROW_SEL
+ pixel_4374/NB1 pixel_4374/VBIAS pixel_4374/NB2 pixel_4374/AMP_IN pixel_4374/SF_IB
+ pixel_4374/PIX_OUT pixel_4374/CSA_VREF pixel
Xpixel_4385 pixel_4385/gring pixel_4385/VDD pixel_4385/GND pixel_4385/VREF pixel_4385/ROW_SEL
+ pixel_4385/NB1 pixel_4385/VBIAS pixel_4385/NB2 pixel_4385/AMP_IN pixel_4385/SF_IB
+ pixel_4385/PIX_OUT pixel_4385/CSA_VREF pixel
Xpixel_4396 pixel_4396/gring pixel_4396/VDD pixel_4396/GND pixel_4396/VREF pixel_4396/ROW_SEL
+ pixel_4396/NB1 pixel_4396/VBIAS pixel_4396/NB2 pixel_4396/AMP_IN pixel_4396/SF_IB
+ pixel_4396/PIX_OUT pixel_4396/CSA_VREF pixel
Xpixel_2950 pixel_2950/gring pixel_2950/VDD pixel_2950/GND pixel_2950/VREF pixel_2950/ROW_SEL
+ pixel_2950/NB1 pixel_2950/VBIAS pixel_2950/NB2 pixel_2950/AMP_IN pixel_2950/SF_IB
+ pixel_2950/PIX_OUT pixel_2950/CSA_VREF pixel
Xpixel_3695 pixel_3695/gring pixel_3695/VDD pixel_3695/GND pixel_3695/VREF pixel_3695/ROW_SEL
+ pixel_3695/NB1 pixel_3695/VBIAS pixel_3695/NB2 pixel_3695/AMP_IN pixel_3695/SF_IB
+ pixel_3695/PIX_OUT pixel_3695/CSA_VREF pixel
Xpixel_3684 pixel_3684/gring pixel_3684/VDD pixel_3684/GND pixel_3684/VREF pixel_3684/ROW_SEL
+ pixel_3684/NB1 pixel_3684/VBIAS pixel_3684/NB2 pixel_3684/AMP_IN pixel_3684/SF_IB
+ pixel_3684/PIX_OUT pixel_3684/CSA_VREF pixel
Xpixel_3673 pixel_3673/gring pixel_3673/VDD pixel_3673/GND pixel_3673/VREF pixel_3673/ROW_SEL
+ pixel_3673/NB1 pixel_3673/VBIAS pixel_3673/NB2 pixel_3673/AMP_IN pixel_3673/SF_IB
+ pixel_3673/PIX_OUT pixel_3673/CSA_VREF pixel
Xpixel_3662 pixel_3662/gring pixel_3662/VDD pixel_3662/GND pixel_3662/VREF pixel_3662/ROW_SEL
+ pixel_3662/NB1 pixel_3662/VBIAS pixel_3662/NB2 pixel_3662/AMP_IN pixel_3662/SF_IB
+ pixel_3662/PIX_OUT pixel_3662/CSA_VREF pixel
Xpixel_2983 pixel_2983/gring pixel_2983/VDD pixel_2983/GND pixel_2983/VREF pixel_2983/ROW_SEL
+ pixel_2983/NB1 pixel_2983/VBIAS pixel_2983/NB2 pixel_2983/AMP_IN pixel_2983/SF_IB
+ pixel_2983/PIX_OUT pixel_2983/CSA_VREF pixel
Xpixel_2972 pixel_2972/gring pixel_2972/VDD pixel_2972/GND pixel_2972/VREF pixel_2972/ROW_SEL
+ pixel_2972/NB1 pixel_2972/VBIAS pixel_2972/NB2 pixel_2972/AMP_IN pixel_2972/SF_IB
+ pixel_2972/PIX_OUT pixel_2972/CSA_VREF pixel
Xpixel_2961 pixel_2961/gring pixel_2961/VDD pixel_2961/GND pixel_2961/VREF pixel_2961/ROW_SEL
+ pixel_2961/NB1 pixel_2961/VBIAS pixel_2961/NB2 pixel_2961/AMP_IN pixel_2961/SF_IB
+ pixel_2961/PIX_OUT pixel_2961/CSA_VREF pixel
Xpixel_2994 pixel_2994/gring pixel_2994/VDD pixel_2994/GND pixel_2994/VREF pixel_2994/ROW_SEL
+ pixel_2994/NB1 pixel_2994/VBIAS pixel_2994/NB2 pixel_2994/AMP_IN pixel_2994/SF_IB
+ pixel_2994/PIX_OUT pixel_2994/CSA_VREF pixel
Xpixel_9319 pixel_9319/gring pixel_9319/VDD pixel_9319/GND pixel_9319/VREF pixel_9319/ROW_SEL
+ pixel_9319/NB1 pixel_9319/VBIAS pixel_9319/NB2 pixel_9319/AMP_IN pixel_9319/SF_IB
+ pixel_9319/PIX_OUT pixel_9319/CSA_VREF pixel
Xpixel_9308 pixel_9308/gring pixel_9308/VDD pixel_9308/GND pixel_9308/VREF pixel_9308/ROW_SEL
+ pixel_9308/NB1 pixel_9308/VBIAS pixel_9308/NB2 pixel_9308/AMP_IN pixel_9308/SF_IB
+ pixel_9308/PIX_OUT pixel_9308/CSA_VREF pixel
Xpixel_8618 pixel_8618/gring pixel_8618/VDD pixel_8618/GND pixel_8618/VREF pixel_8618/ROW_SEL
+ pixel_8618/NB1 pixel_8618/VBIAS pixel_8618/NB2 pixel_8618/AMP_IN pixel_8618/SF_IB
+ pixel_8618/PIX_OUT pixel_8618/CSA_VREF pixel
Xpixel_8607 pixel_8607/gring pixel_8607/VDD pixel_8607/GND pixel_8607/VREF pixel_8607/ROW_SEL
+ pixel_8607/NB1 pixel_8607/VBIAS pixel_8607/NB2 pixel_8607/AMP_IN pixel_8607/SF_IB
+ pixel_8607/PIX_OUT pixel_8607/CSA_VREF pixel
Xpixel_8629 pixel_8629/gring pixel_8629/VDD pixel_8629/GND pixel_8629/VREF pixel_8629/ROW_SEL
+ pixel_8629/NB1 pixel_8629/VBIAS pixel_8629/NB2 pixel_8629/AMP_IN pixel_8629/SF_IB
+ pixel_8629/PIX_OUT pixel_8629/CSA_VREF pixel
Xpixel_7906 pixel_7906/gring pixel_7906/VDD pixel_7906/GND pixel_7906/VREF pixel_7906/ROW_SEL
+ pixel_7906/NB1 pixel_7906/VBIAS pixel_7906/NB2 pixel_7906/AMP_IN pixel_7906/SF_IB
+ pixel_7906/PIX_OUT pixel_7906/CSA_VREF pixel
Xpixel_7917 pixel_7917/gring pixel_7917/VDD pixel_7917/GND pixel_7917/VREF pixel_7917/ROW_SEL
+ pixel_7917/NB1 pixel_7917/VBIAS pixel_7917/NB2 pixel_7917/AMP_IN pixel_7917/SF_IB
+ pixel_7917/PIX_OUT pixel_7917/CSA_VREF pixel
Xpixel_7928 pixel_7928/gring pixel_7928/VDD pixel_7928/GND pixel_7928/VREF pixel_7928/ROW_SEL
+ pixel_7928/NB1 pixel_7928/VBIAS pixel_7928/NB2 pixel_7928/AMP_IN pixel_7928/SF_IB
+ pixel_7928/PIX_OUT pixel_7928/CSA_VREF pixel
Xpixel_7939 pixel_7939/gring pixel_7939/VDD pixel_7939/GND pixel_7939/VREF pixel_7939/ROW_SEL
+ pixel_7939/NB1 pixel_7939/VBIAS pixel_7939/NB2 pixel_7939/AMP_IN pixel_7939/SF_IB
+ pixel_7939/PIX_OUT pixel_7939/CSA_VREF pixel
Xpixel_2202 pixel_2202/gring pixel_2202/VDD pixel_2202/GND pixel_2202/VREF pixel_2202/ROW_SEL
+ pixel_2202/NB1 pixel_2202/VBIAS pixel_2202/NB2 pixel_2202/AMP_IN pixel_2202/SF_IB
+ pixel_2202/PIX_OUT pixel_2202/CSA_VREF pixel
Xpixel_2235 pixel_2235/gring pixel_2235/VDD pixel_2235/GND pixel_2235/VREF pixel_2235/ROW_SEL
+ pixel_2235/NB1 pixel_2235/VBIAS pixel_2235/NB2 pixel_2235/AMP_IN pixel_2235/SF_IB
+ pixel_2235/PIX_OUT pixel_2235/CSA_VREF pixel
Xpixel_2224 pixel_2224/gring pixel_2224/VDD pixel_2224/GND pixel_2224/VREF pixel_2224/ROW_SEL
+ pixel_2224/NB1 pixel_2224/VBIAS pixel_2224/NB2 pixel_2224/AMP_IN pixel_2224/SF_IB
+ pixel_2224/PIX_OUT pixel_2224/CSA_VREF pixel
Xpixel_2213 pixel_2213/gring pixel_2213/VDD pixel_2213/GND pixel_2213/VREF pixel_2213/ROW_SEL
+ pixel_2213/NB1 pixel_2213/VBIAS pixel_2213/NB2 pixel_2213/AMP_IN pixel_2213/SF_IB
+ pixel_2213/PIX_OUT pixel_2213/CSA_VREF pixel
Xpixel_1534 pixel_1534/gring pixel_1534/VDD pixel_1534/GND pixel_1534/VREF pixel_1534/ROW_SEL
+ pixel_1534/NB1 pixel_1534/VBIAS pixel_1534/NB2 pixel_1534/AMP_IN pixel_1534/SF_IB
+ pixel_1534/PIX_OUT pixel_1534/CSA_VREF pixel
Xpixel_1523 pixel_1523/gring pixel_1523/VDD pixel_1523/GND pixel_1523/VREF pixel_1523/ROW_SEL
+ pixel_1523/NB1 pixel_1523/VBIAS pixel_1523/NB2 pixel_1523/AMP_IN pixel_1523/SF_IB
+ pixel_1523/PIX_OUT pixel_1523/CSA_VREF pixel
Xpixel_1512 pixel_1512/gring pixel_1512/VDD pixel_1512/GND pixel_1512/VREF pixel_1512/ROW_SEL
+ pixel_1512/NB1 pixel_1512/VBIAS pixel_1512/NB2 pixel_1512/AMP_IN pixel_1512/SF_IB
+ pixel_1512/PIX_OUT pixel_1512/CSA_VREF pixel
Xpixel_1501 pixel_1501/gring pixel_1501/VDD pixel_1501/GND pixel_1501/VREF pixel_1501/ROW_SEL
+ pixel_1501/NB1 pixel_1501/VBIAS pixel_1501/NB2 pixel_1501/AMP_IN pixel_1501/SF_IB
+ pixel_1501/PIX_OUT pixel_1501/CSA_VREF pixel
Xpixel_2279 pixel_2279/gring pixel_2279/VDD pixel_2279/GND pixel_2279/VREF pixel_2279/ROW_SEL
+ pixel_2279/NB1 pixel_2279/VBIAS pixel_2279/NB2 pixel_2279/AMP_IN pixel_2279/SF_IB
+ pixel_2279/PIX_OUT pixel_2279/CSA_VREF pixel
Xpixel_2268 pixel_2268/gring pixel_2268/VDD pixel_2268/GND pixel_2268/VREF pixel_2268/ROW_SEL
+ pixel_2268/NB1 pixel_2268/VBIAS pixel_2268/NB2 pixel_2268/AMP_IN pixel_2268/SF_IB
+ pixel_2268/PIX_OUT pixel_2268/CSA_VREF pixel
Xpixel_2257 pixel_2257/gring pixel_2257/VDD pixel_2257/GND pixel_2257/VREF pixel_2257/ROW_SEL
+ pixel_2257/NB1 pixel_2257/VBIAS pixel_2257/NB2 pixel_2257/AMP_IN pixel_2257/SF_IB
+ pixel_2257/PIX_OUT pixel_2257/CSA_VREF pixel
Xpixel_2246 pixel_2246/gring pixel_2246/VDD pixel_2246/GND pixel_2246/VREF pixel_2246/ROW_SEL
+ pixel_2246/NB1 pixel_2246/VBIAS pixel_2246/NB2 pixel_2246/AMP_IN pixel_2246/SF_IB
+ pixel_2246/PIX_OUT pixel_2246/CSA_VREF pixel
Xpixel_1567 pixel_1567/gring pixel_1567/VDD pixel_1567/GND pixel_1567/VREF pixel_1567/ROW_SEL
+ pixel_1567/NB1 pixel_1567/VBIAS pixel_1567/NB2 pixel_1567/AMP_IN pixel_1567/SF_IB
+ pixel_1567/PIX_OUT pixel_1567/CSA_VREF pixel
Xpixel_1556 pixel_1556/gring pixel_1556/VDD pixel_1556/GND pixel_1556/VREF pixel_1556/ROW_SEL
+ pixel_1556/NB1 pixel_1556/VBIAS pixel_1556/NB2 pixel_1556/AMP_IN pixel_1556/SF_IB
+ pixel_1556/PIX_OUT pixel_1556/CSA_VREF pixel
Xpixel_1545 pixel_1545/gring pixel_1545/VDD pixel_1545/GND pixel_1545/VREF pixel_1545/ROW_SEL
+ pixel_1545/NB1 pixel_1545/VBIAS pixel_1545/NB2 pixel_1545/AMP_IN pixel_1545/SF_IB
+ pixel_1545/PIX_OUT pixel_1545/CSA_VREF pixel
Xpixel_1589 pixel_1589/gring pixel_1589/VDD pixel_1589/GND pixel_1589/VREF pixel_1589/ROW_SEL
+ pixel_1589/NB1 pixel_1589/VBIAS pixel_1589/NB2 pixel_1589/AMP_IN pixel_1589/SF_IB
+ pixel_1589/PIX_OUT pixel_1589/CSA_VREF pixel
Xpixel_1578 pixel_1578/gring pixel_1578/VDD pixel_1578/GND pixel_1578/VREF pixel_1578/ROW_SEL
+ pixel_1578/NB1 pixel_1578/VBIAS pixel_1578/NB2 pixel_1578/AMP_IN pixel_1578/SF_IB
+ pixel_1578/PIX_OUT pixel_1578/CSA_VREF pixel
Xpixel_9842 pixel_9842/gring pixel_9842/VDD pixel_9842/GND pixel_9842/VREF pixel_9842/ROW_SEL
+ pixel_9842/NB1 pixel_9842/VBIAS pixel_9842/NB2 pixel_9842/AMP_IN pixel_9842/SF_IB
+ pixel_9842/PIX_OUT pixel_9842/CSA_VREF pixel
Xpixel_9831 pixel_9831/gring pixel_9831/VDD pixel_9831/GND pixel_9831/VREF pixel_9831/ROW_SEL
+ pixel_9831/NB1 pixel_9831/VBIAS pixel_9831/NB2 pixel_9831/AMP_IN pixel_9831/SF_IB
+ pixel_9831/PIX_OUT pixel_9831/CSA_VREF pixel
Xpixel_9820 pixel_9820/gring pixel_9820/VDD pixel_9820/GND pixel_9820/VREF pixel_9820/ROW_SEL
+ pixel_9820/NB1 pixel_9820/VBIAS pixel_9820/NB2 pixel_9820/AMP_IN pixel_9820/SF_IB
+ pixel_9820/PIX_OUT pixel_9820/CSA_VREF pixel
Xpixel_9853 pixel_9853/gring pixel_9853/VDD pixel_9853/GND pixel_9853/VREF pixel_9853/ROW_SEL
+ pixel_9853/NB1 pixel_9853/VBIAS pixel_9853/NB2 pixel_9853/AMP_IN pixel_9853/SF_IB
+ pixel_9853/PIX_OUT pixel_9853/CSA_VREF pixel
Xpixel_9864 pixel_9864/gring pixel_9864/VDD pixel_9864/GND pixel_9864/VREF pixel_9864/ROW_SEL
+ pixel_9864/NB1 pixel_9864/VBIAS pixel_9864/NB2 pixel_9864/AMP_IN pixel_9864/SF_IB
+ pixel_9864/PIX_OUT pixel_9864/CSA_VREF pixel
Xpixel_9875 pixel_9875/gring pixel_9875/VDD pixel_9875/GND pixel_9875/VREF pixel_9875/ROW_SEL
+ pixel_9875/NB1 pixel_9875/VBIAS pixel_9875/NB2 pixel_9875/AMP_IN pixel_9875/SF_IB
+ pixel_9875/PIX_OUT pixel_9875/CSA_VREF pixel
Xpixel_9886 pixel_9886/gring pixel_9886/VDD pixel_9886/GND pixel_9886/VREF pixel_9886/ROW_SEL
+ pixel_9886/NB1 pixel_9886/VBIAS pixel_9886/NB2 pixel_9886/AMP_IN pixel_9886/SF_IB
+ pixel_9886/PIX_OUT pixel_9886/CSA_VREF pixel
Xpixel_9897 pixel_9897/gring pixel_9897/VDD pixel_9897/GND pixel_9897/VREF pixel_9897/ROW_SEL
+ pixel_9897/NB1 pixel_9897/VBIAS pixel_9897/NB2 pixel_9897/AMP_IN pixel_9897/SF_IB
+ pixel_9897/PIX_OUT pixel_9897/CSA_VREF pixel
Xpixel_4160 pixel_4160/gring pixel_4160/VDD pixel_4160/GND pixel_4160/VREF pixel_4160/ROW_SEL
+ pixel_4160/NB1 pixel_4160/VBIAS pixel_4160/NB2 pixel_4160/AMP_IN pixel_4160/SF_IB
+ pixel_4160/PIX_OUT pixel_4160/CSA_VREF pixel
Xpixel_4171 pixel_4171/gring pixel_4171/VDD pixel_4171/GND pixel_4171/VREF pixel_4171/ROW_SEL
+ pixel_4171/NB1 pixel_4171/VBIAS pixel_4171/NB2 pixel_4171/AMP_IN pixel_4171/SF_IB
+ pixel_4171/PIX_OUT pixel_4171/CSA_VREF pixel
Xpixel_4182 pixel_4182/gring pixel_4182/VDD pixel_4182/GND pixel_4182/VREF pixel_4182/ROW_SEL
+ pixel_4182/NB1 pixel_4182/VBIAS pixel_4182/NB2 pixel_4182/AMP_IN pixel_4182/SF_IB
+ pixel_4182/PIX_OUT pixel_4182/CSA_VREF pixel
Xpixel_4193 pixel_4193/gring pixel_4193/VDD pixel_4193/GND pixel_4193/VREF pixel_4193/ROW_SEL
+ pixel_4193/NB1 pixel_4193/VBIAS pixel_4193/NB2 pixel_4193/AMP_IN pixel_4193/SF_IB
+ pixel_4193/PIX_OUT pixel_4193/CSA_VREF pixel
Xpixel_3492 pixel_3492/gring pixel_3492/VDD pixel_3492/GND pixel_3492/VREF pixel_3492/ROW_SEL
+ pixel_3492/NB1 pixel_3492/VBIAS pixel_3492/NB2 pixel_3492/AMP_IN pixel_3492/SF_IB
+ pixel_3492/PIX_OUT pixel_3492/CSA_VREF pixel
Xpixel_3481 pixel_3481/gring pixel_3481/VDD pixel_3481/GND pixel_3481/VREF pixel_3481/ROW_SEL
+ pixel_3481/NB1 pixel_3481/VBIAS pixel_3481/NB2 pixel_3481/AMP_IN pixel_3481/SF_IB
+ pixel_3481/PIX_OUT pixel_3481/CSA_VREF pixel
Xpixel_3470 pixel_3470/gring pixel_3470/VDD pixel_3470/GND pixel_3470/VREF pixel_3470/ROW_SEL
+ pixel_3470/NB1 pixel_3470/VBIAS pixel_3470/NB2 pixel_3470/AMP_IN pixel_3470/SF_IB
+ pixel_3470/PIX_OUT pixel_3470/CSA_VREF pixel
Xpixel_2791 pixel_2791/gring pixel_2791/VDD pixel_2791/GND pixel_2791/VREF pixel_2791/ROW_SEL
+ pixel_2791/NB1 pixel_2791/VBIAS pixel_2791/NB2 pixel_2791/AMP_IN pixel_2791/SF_IB
+ pixel_2791/PIX_OUT pixel_2791/CSA_VREF pixel
Xpixel_2780 pixel_2780/gring pixel_2780/VDD pixel_2780/GND pixel_2780/VREF pixel_2780/ROW_SEL
+ pixel_2780/NB1 pixel_2780/VBIAS pixel_2780/NB2 pixel_2780/AMP_IN pixel_2780/SF_IB
+ pixel_2780/PIX_OUT pixel_2780/CSA_VREF pixel
Xpixel_9127 pixel_9127/gring pixel_9127/VDD pixel_9127/GND pixel_9127/VREF pixel_9127/ROW_SEL
+ pixel_9127/NB1 pixel_9127/VBIAS pixel_9127/NB2 pixel_9127/AMP_IN pixel_9127/SF_IB
+ pixel_9127/PIX_OUT pixel_9127/CSA_VREF pixel
Xpixel_9116 pixel_9116/gring pixel_9116/VDD pixel_9116/GND pixel_9116/VREF pixel_9116/ROW_SEL
+ pixel_9116/NB1 pixel_9116/VBIAS pixel_9116/NB2 pixel_9116/AMP_IN pixel_9116/SF_IB
+ pixel_9116/PIX_OUT pixel_9116/CSA_VREF pixel
Xpixel_9105 pixel_9105/gring pixel_9105/VDD pixel_9105/GND pixel_9105/VREF pixel_9105/ROW_SEL
+ pixel_9105/NB1 pixel_9105/VBIAS pixel_9105/NB2 pixel_9105/AMP_IN pixel_9105/SF_IB
+ pixel_9105/PIX_OUT pixel_9105/CSA_VREF pixel
Xpixel_8426 pixel_8426/gring pixel_8426/VDD pixel_8426/GND pixel_8426/VREF pixel_8426/ROW_SEL
+ pixel_8426/NB1 pixel_8426/VBIAS pixel_8426/NB2 pixel_8426/AMP_IN pixel_8426/SF_IB
+ pixel_8426/PIX_OUT pixel_8426/CSA_VREF pixel
Xpixel_8415 pixel_8415/gring pixel_8415/VDD pixel_8415/GND pixel_8415/VREF pixel_8415/ROW_SEL
+ pixel_8415/NB1 pixel_8415/VBIAS pixel_8415/NB2 pixel_8415/AMP_IN pixel_8415/SF_IB
+ pixel_8415/PIX_OUT pixel_8415/CSA_VREF pixel
Xpixel_8404 pixel_8404/gring pixel_8404/VDD pixel_8404/GND pixel_8404/VREF pixel_8404/ROW_SEL
+ pixel_8404/NB1 pixel_8404/VBIAS pixel_8404/NB2 pixel_8404/AMP_IN pixel_8404/SF_IB
+ pixel_8404/PIX_OUT pixel_8404/CSA_VREF pixel
Xpixel_9149 pixel_9149/gring pixel_9149/VDD pixel_9149/GND pixel_9149/VREF pixel_9149/ROW_SEL
+ pixel_9149/NB1 pixel_9149/VBIAS pixel_9149/NB2 pixel_9149/AMP_IN pixel_9149/SF_IB
+ pixel_9149/PIX_OUT pixel_9149/CSA_VREF pixel
Xpixel_9138 pixel_9138/gring pixel_9138/VDD pixel_9138/GND pixel_9138/VREF pixel_9138/ROW_SEL
+ pixel_9138/NB1 pixel_9138/VBIAS pixel_9138/NB2 pixel_9138/AMP_IN pixel_9138/SF_IB
+ pixel_9138/PIX_OUT pixel_9138/CSA_VREF pixel
Xpixel_8437 pixel_8437/gring pixel_8437/VDD pixel_8437/GND pixel_8437/VREF pixel_8437/ROW_SEL
+ pixel_8437/NB1 pixel_8437/VBIAS pixel_8437/NB2 pixel_8437/AMP_IN pixel_8437/SF_IB
+ pixel_8437/PIX_OUT pixel_8437/CSA_VREF pixel
Xpixel_8448 pixel_8448/gring pixel_8448/VDD pixel_8448/GND pixel_8448/VREF pixel_8448/ROW_SEL
+ pixel_8448/NB1 pixel_8448/VBIAS pixel_8448/NB2 pixel_8448/AMP_IN pixel_8448/SF_IB
+ pixel_8448/PIX_OUT pixel_8448/CSA_VREF pixel
Xpixel_8459 pixel_8459/gring pixel_8459/VDD pixel_8459/GND pixel_8459/VREF pixel_8459/ROW_SEL
+ pixel_8459/NB1 pixel_8459/VBIAS pixel_8459/NB2 pixel_8459/AMP_IN pixel_8459/SF_IB
+ pixel_8459/PIX_OUT pixel_8459/CSA_VREF pixel
Xpixel_7703 pixel_7703/gring pixel_7703/VDD pixel_7703/GND pixel_7703/VREF pixel_7703/ROW_SEL
+ pixel_7703/NB1 pixel_7703/VBIAS pixel_7703/NB2 pixel_7703/AMP_IN pixel_7703/SF_IB
+ pixel_7703/PIX_OUT pixel_7703/CSA_VREF pixel
Xpixel_7714 pixel_7714/gring pixel_7714/VDD pixel_7714/GND pixel_7714/VREF pixel_7714/ROW_SEL
+ pixel_7714/NB1 pixel_7714/VBIAS pixel_7714/NB2 pixel_7714/AMP_IN pixel_7714/SF_IB
+ pixel_7714/PIX_OUT pixel_7714/CSA_VREF pixel
Xpixel_7725 pixel_7725/gring pixel_7725/VDD pixel_7725/GND pixel_7725/VREF pixel_7725/ROW_SEL
+ pixel_7725/NB1 pixel_7725/VBIAS pixel_7725/NB2 pixel_7725/AMP_IN pixel_7725/SF_IB
+ pixel_7725/PIX_OUT pixel_7725/CSA_VREF pixel
Xpixel_7736 pixel_7736/gring pixel_7736/VDD pixel_7736/GND pixel_7736/VREF pixel_7736/ROW_SEL
+ pixel_7736/NB1 pixel_7736/VBIAS pixel_7736/NB2 pixel_7736/AMP_IN pixel_7736/SF_IB
+ pixel_7736/PIX_OUT pixel_7736/CSA_VREF pixel
Xpixel_7747 pixel_7747/gring pixel_7747/VDD pixel_7747/GND pixel_7747/VREF pixel_7747/ROW_SEL
+ pixel_7747/NB1 pixel_7747/VBIAS pixel_7747/NB2 pixel_7747/AMP_IN pixel_7747/SF_IB
+ pixel_7747/PIX_OUT pixel_7747/CSA_VREF pixel
Xpixel_7758 pixel_7758/gring pixel_7758/VDD pixel_7758/GND pixel_7758/VREF pixel_7758/ROW_SEL
+ pixel_7758/NB1 pixel_7758/VBIAS pixel_7758/NB2 pixel_7758/AMP_IN pixel_7758/SF_IB
+ pixel_7758/PIX_OUT pixel_7758/CSA_VREF pixel
Xpixel_7769 pixel_7769/gring pixel_7769/VDD pixel_7769/GND pixel_7769/VREF pixel_7769/ROW_SEL
+ pixel_7769/NB1 pixel_7769/VBIAS pixel_7769/NB2 pixel_7769/AMP_IN pixel_7769/SF_IB
+ pixel_7769/PIX_OUT pixel_7769/CSA_VREF pixel
Xpixel_2010 pixel_2010/gring pixel_2010/VDD pixel_2010/GND pixel_2010/VREF pixel_2010/ROW_SEL
+ pixel_2010/NB1 pixel_2010/VBIAS pixel_2010/NB2 pixel_2010/AMP_IN pixel_2010/SF_IB
+ pixel_2010/PIX_OUT pixel_2010/CSA_VREF pixel
Xpixel_2054 pixel_2054/gring pixel_2054/VDD pixel_2054/GND pixel_2054/VREF pixel_2054/ROW_SEL
+ pixel_2054/NB1 pixel_2054/VBIAS pixel_2054/NB2 pixel_2054/AMP_IN pixel_2054/SF_IB
+ pixel_2054/PIX_OUT pixel_2054/CSA_VREF pixel
Xpixel_2043 pixel_2043/gring pixel_2043/VDD pixel_2043/GND pixel_2043/VREF pixel_2043/ROW_SEL
+ pixel_2043/NB1 pixel_2043/VBIAS pixel_2043/NB2 pixel_2043/AMP_IN pixel_2043/SF_IB
+ pixel_2043/PIX_OUT pixel_2043/CSA_VREF pixel
Xpixel_2032 pixel_2032/gring pixel_2032/VDD pixel_2032/GND pixel_2032/VREF pixel_2032/ROW_SEL
+ pixel_2032/NB1 pixel_2032/VBIAS pixel_2032/NB2 pixel_2032/AMP_IN pixel_2032/SF_IB
+ pixel_2032/PIX_OUT pixel_2032/CSA_VREF pixel
Xpixel_2021 pixel_2021/gring pixel_2021/VDD pixel_2021/GND pixel_2021/VREF pixel_2021/ROW_SEL
+ pixel_2021/NB1 pixel_2021/VBIAS pixel_2021/NB2 pixel_2021/AMP_IN pixel_2021/SF_IB
+ pixel_2021/PIX_OUT pixel_2021/CSA_VREF pixel
Xpixel_1342 pixel_1342/gring pixel_1342/VDD pixel_1342/GND pixel_1342/VREF pixel_1342/ROW_SEL
+ pixel_1342/NB1 pixel_1342/VBIAS pixel_1342/NB2 pixel_1342/AMP_IN pixel_1342/SF_IB
+ pixel_1342/PIX_OUT pixel_1342/CSA_VREF pixel
Xpixel_1331 pixel_1331/gring pixel_1331/VDD pixel_1331/GND pixel_1331/VREF pixel_1331/ROW_SEL
+ pixel_1331/NB1 pixel_1331/VBIAS pixel_1331/NB2 pixel_1331/AMP_IN pixel_1331/SF_IB
+ pixel_1331/PIX_OUT pixel_1331/CSA_VREF pixel
Xpixel_1320 pixel_1320/gring pixel_1320/VDD pixel_1320/GND pixel_1320/VREF pixel_1320/ROW_SEL
+ pixel_1320/NB1 pixel_1320/VBIAS pixel_1320/NB2 pixel_1320/AMP_IN pixel_1320/SF_IB
+ pixel_1320/PIX_OUT pixel_1320/CSA_VREF pixel
Xpixel_2087 pixel_2087/gring pixel_2087/VDD pixel_2087/GND pixel_2087/VREF pixel_2087/ROW_SEL
+ pixel_2087/NB1 pixel_2087/VBIAS pixel_2087/NB2 pixel_2087/AMP_IN pixel_2087/SF_IB
+ pixel_2087/PIX_OUT pixel_2087/CSA_VREF pixel
Xpixel_2076 pixel_2076/gring pixel_2076/VDD pixel_2076/GND pixel_2076/VREF pixel_2076/ROW_SEL
+ pixel_2076/NB1 pixel_2076/VBIAS pixel_2076/NB2 pixel_2076/AMP_IN pixel_2076/SF_IB
+ pixel_2076/PIX_OUT pixel_2076/CSA_VREF pixel
Xpixel_2065 pixel_2065/gring pixel_2065/VDD pixel_2065/GND pixel_2065/VREF pixel_2065/ROW_SEL
+ pixel_2065/NB1 pixel_2065/VBIAS pixel_2065/NB2 pixel_2065/AMP_IN pixel_2065/SF_IB
+ pixel_2065/PIX_OUT pixel_2065/CSA_VREF pixel
Xpixel_1375 pixel_1375/gring pixel_1375/VDD pixel_1375/GND pixel_1375/VREF pixel_1375/ROW_SEL
+ pixel_1375/NB1 pixel_1375/VBIAS pixel_1375/NB2 pixel_1375/AMP_IN pixel_1375/SF_IB
+ pixel_1375/PIX_OUT pixel_1375/CSA_VREF pixel
Xpixel_1364 pixel_1364/gring pixel_1364/VDD pixel_1364/GND pixel_1364/VREF pixel_1364/ROW_SEL
+ pixel_1364/NB1 pixel_1364/VBIAS pixel_1364/NB2 pixel_1364/AMP_IN pixel_1364/SF_IB
+ pixel_1364/PIX_OUT pixel_1364/CSA_VREF pixel
Xpixel_1353 pixel_1353/gring pixel_1353/VDD pixel_1353/GND pixel_1353/VREF pixel_1353/ROW_SEL
+ pixel_1353/NB1 pixel_1353/VBIAS pixel_1353/NB2 pixel_1353/AMP_IN pixel_1353/SF_IB
+ pixel_1353/PIX_OUT pixel_1353/CSA_VREF pixel
Xpixel_2098 pixel_2098/gring pixel_2098/VDD pixel_2098/GND pixel_2098/VREF pixel_2098/ROW_SEL
+ pixel_2098/NB1 pixel_2098/VBIAS pixel_2098/NB2 pixel_2098/AMP_IN pixel_2098/SF_IB
+ pixel_2098/PIX_OUT pixel_2098/CSA_VREF pixel
Xpixel_1397 pixel_1397/gring pixel_1397/VDD pixel_1397/GND pixel_1397/VREF pixel_1397/ROW_SEL
+ pixel_1397/NB1 pixel_1397/VBIAS pixel_1397/NB2 pixel_1397/AMP_IN pixel_1397/SF_IB
+ pixel_1397/PIX_OUT pixel_1397/CSA_VREF pixel
Xpixel_1386 pixel_1386/gring pixel_1386/VDD pixel_1386/GND pixel_1386/VREF pixel_1386/ROW_SEL
+ pixel_1386/NB1 pixel_1386/VBIAS pixel_1386/NB2 pixel_1386/AMP_IN pixel_1386/SF_IB
+ pixel_1386/PIX_OUT pixel_1386/CSA_VREF pixel
Xpixel_9650 pixel_9650/gring pixel_9650/VDD pixel_9650/GND pixel_9650/VREF pixel_9650/ROW_SEL
+ pixel_9650/NB1 pixel_9650/VBIAS pixel_9650/NB2 pixel_9650/AMP_IN pixel_9650/SF_IB
+ pixel_9650/PIX_OUT pixel_9650/CSA_VREF pixel
Xpixel_9661 pixel_9661/gring pixel_9661/VDD pixel_9661/GND pixel_9661/VREF pixel_9661/ROW_SEL
+ pixel_9661/NB1 pixel_9661/VBIAS pixel_9661/NB2 pixel_9661/AMP_IN pixel_9661/SF_IB
+ pixel_9661/PIX_OUT pixel_9661/CSA_VREF pixel
Xpixel_9672 pixel_9672/gring pixel_9672/VDD pixel_9672/GND pixel_9672/VREF pixel_9672/ROW_SEL
+ pixel_9672/NB1 pixel_9672/VBIAS pixel_9672/NB2 pixel_9672/AMP_IN pixel_9672/SF_IB
+ pixel_9672/PIX_OUT pixel_9672/CSA_VREF pixel
Xpixel_9683 pixel_9683/gring pixel_9683/VDD pixel_9683/GND pixel_9683/VREF pixel_9683/ROW_SEL
+ pixel_9683/NB1 pixel_9683/VBIAS pixel_9683/NB2 pixel_9683/AMP_IN pixel_9683/SF_IB
+ pixel_9683/PIX_OUT pixel_9683/CSA_VREF pixel
Xpixel_8982 pixel_8982/gring pixel_8982/VDD pixel_8982/GND pixel_8982/VREF pixel_8982/ROW_SEL
+ pixel_8982/NB1 pixel_8982/VBIAS pixel_8982/NB2 pixel_8982/AMP_IN pixel_8982/SF_IB
+ pixel_8982/PIX_OUT pixel_8982/CSA_VREF pixel
Xpixel_8971 pixel_8971/gring pixel_8971/VDD pixel_8971/GND pixel_8971/VREF pixel_8971/ROW_SEL
+ pixel_8971/NB1 pixel_8971/VBIAS pixel_8971/NB2 pixel_8971/AMP_IN pixel_8971/SF_IB
+ pixel_8971/PIX_OUT pixel_8971/CSA_VREF pixel
Xpixel_8960 pixel_8960/gring pixel_8960/VDD pixel_8960/GND pixel_8960/VREF pixel_8960/ROW_SEL
+ pixel_8960/NB1 pixel_8960/VBIAS pixel_8960/NB2 pixel_8960/AMP_IN pixel_8960/SF_IB
+ pixel_8960/PIX_OUT pixel_8960/CSA_VREF pixel
Xpixel_9694 pixel_9694/gring pixel_9694/VDD pixel_9694/GND pixel_9694/VREF pixel_9694/ROW_SEL
+ pixel_9694/NB1 pixel_9694/VBIAS pixel_9694/NB2 pixel_9694/AMP_IN pixel_9694/SF_IB
+ pixel_9694/PIX_OUT pixel_9694/CSA_VREF pixel
Xpixel_8993 pixel_8993/gring pixel_8993/VDD pixel_8993/GND pixel_8993/VREF pixel_8993/ROW_SEL
+ pixel_8993/NB1 pixel_8993/VBIAS pixel_8993/NB2 pixel_8993/AMP_IN pixel_8993/SF_IB
+ pixel_8993/PIX_OUT pixel_8993/CSA_VREF pixel
Xpixel_6309 pixel_6309/gring pixel_6309/VDD pixel_6309/GND pixel_6309/VREF pixel_6309/ROW_SEL
+ pixel_6309/NB1 pixel_6309/VBIAS pixel_6309/NB2 pixel_6309/AMP_IN pixel_6309/SF_IB
+ pixel_6309/PIX_OUT pixel_6309/CSA_VREF pixel
Xpixel_5608 pixel_5608/gring pixel_5608/VDD pixel_5608/GND pixel_5608/VREF pixel_5608/ROW_SEL
+ pixel_5608/NB1 pixel_5608/VBIAS pixel_5608/NB2 pixel_5608/AMP_IN pixel_5608/SF_IB
+ pixel_5608/PIX_OUT pixel_5608/CSA_VREF pixel
Xpixel_5619 pixel_5619/gring pixel_5619/VDD pixel_5619/GND pixel_5619/VREF pixel_5619/ROW_SEL
+ pixel_5619/NB1 pixel_5619/VBIAS pixel_5619/NB2 pixel_5619/AMP_IN pixel_5619/SF_IB
+ pixel_5619/PIX_OUT pixel_5619/CSA_VREF pixel
Xpixel_924 pixel_924/gring pixel_924/VDD pixel_924/GND pixel_924/VREF pixel_924/ROW_SEL
+ pixel_924/NB1 pixel_924/VBIAS pixel_924/NB2 pixel_924/AMP_IN pixel_924/SF_IB pixel_924/PIX_OUT
+ pixel_924/CSA_VREF pixel
Xpixel_913 pixel_913/gring pixel_913/VDD pixel_913/GND pixel_913/VREF pixel_913/ROW_SEL
+ pixel_913/NB1 pixel_913/VBIAS pixel_913/NB2 pixel_913/AMP_IN pixel_913/SF_IB pixel_913/PIX_OUT
+ pixel_913/CSA_VREF pixel
Xpixel_902 pixel_902/gring pixel_902/VDD pixel_902/GND pixel_902/VREF pixel_902/ROW_SEL
+ pixel_902/NB1 pixel_902/VBIAS pixel_902/NB2 pixel_902/AMP_IN pixel_902/SF_IB pixel_902/PIX_OUT
+ pixel_902/CSA_VREF pixel
Xpixel_4907 pixel_4907/gring pixel_4907/VDD pixel_4907/GND pixel_4907/VREF pixel_4907/ROW_SEL
+ pixel_4907/NB1 pixel_4907/VBIAS pixel_4907/NB2 pixel_4907/AMP_IN pixel_4907/SF_IB
+ pixel_4907/PIX_OUT pixel_4907/CSA_VREF pixel
Xpixel_4918 pixel_4918/gring pixel_4918/VDD pixel_4918/GND pixel_4918/VREF pixel_4918/ROW_SEL
+ pixel_4918/NB1 pixel_4918/VBIAS pixel_4918/NB2 pixel_4918/AMP_IN pixel_4918/SF_IB
+ pixel_4918/PIX_OUT pixel_4918/CSA_VREF pixel
Xpixel_4929 pixel_4929/gring pixel_4929/VDD pixel_4929/GND pixel_4929/VREF pixel_4929/ROW_SEL
+ pixel_4929/NB1 pixel_4929/VBIAS pixel_4929/NB2 pixel_4929/AMP_IN pixel_4929/SF_IB
+ pixel_4929/PIX_OUT pixel_4929/CSA_VREF pixel
Xpixel_957 pixel_957/gring pixel_957/VDD pixel_957/GND pixel_957/VREF pixel_957/ROW_SEL
+ pixel_957/NB1 pixel_957/VBIAS pixel_957/NB2 pixel_957/AMP_IN pixel_957/SF_IB pixel_957/PIX_OUT
+ pixel_957/CSA_VREF pixel
Xpixel_946 pixel_946/gring pixel_946/VDD pixel_946/GND pixel_946/VREF pixel_946/ROW_SEL
+ pixel_946/NB1 pixel_946/VBIAS pixel_946/NB2 pixel_946/AMP_IN pixel_946/SF_IB pixel_946/PIX_OUT
+ pixel_946/CSA_VREF pixel
Xpixel_935 pixel_935/gring pixel_935/VDD pixel_935/GND pixel_935/VREF pixel_935/ROW_SEL
+ pixel_935/NB1 pixel_935/VBIAS pixel_935/NB2 pixel_935/AMP_IN pixel_935/SF_IB pixel_935/PIX_OUT
+ pixel_935/CSA_VREF pixel
Xpixel_979 pixel_979/gring pixel_979/VDD pixel_979/GND pixel_979/VREF pixel_979/ROW_SEL
+ pixel_979/NB1 pixel_979/VBIAS pixel_979/NB2 pixel_979/AMP_IN pixel_979/SF_IB pixel_979/PIX_OUT
+ pixel_979/CSA_VREF pixel
Xpixel_968 pixel_968/gring pixel_968/VDD pixel_968/GND pixel_968/VREF pixel_968/ROW_SEL
+ pixel_968/NB1 pixel_968/VBIAS pixel_968/NB2 pixel_968/AMP_IN pixel_968/SF_IB pixel_968/PIX_OUT
+ pixel_968/CSA_VREF pixel
Xpixel_8201 pixel_8201/gring pixel_8201/VDD pixel_8201/GND pixel_8201/VREF pixel_8201/ROW_SEL
+ pixel_8201/NB1 pixel_8201/VBIAS pixel_8201/NB2 pixel_8201/AMP_IN pixel_8201/SF_IB
+ pixel_8201/PIX_OUT pixel_8201/CSA_VREF pixel
Xpixel_8212 pixel_8212/gring pixel_8212/VDD pixel_8212/GND pixel_8212/VREF pixel_8212/ROW_SEL
+ pixel_8212/NB1 pixel_8212/VBIAS pixel_8212/NB2 pixel_8212/AMP_IN pixel_8212/SF_IB
+ pixel_8212/PIX_OUT pixel_8212/CSA_VREF pixel
Xpixel_8223 pixel_8223/gring pixel_8223/VDD pixel_8223/GND pixel_8223/VREF pixel_8223/ROW_SEL
+ pixel_8223/NB1 pixel_8223/VBIAS pixel_8223/NB2 pixel_8223/AMP_IN pixel_8223/SF_IB
+ pixel_8223/PIX_OUT pixel_8223/CSA_VREF pixel
Xpixel_8234 pixel_8234/gring pixel_8234/VDD pixel_8234/GND pixel_8234/VREF pixel_8234/ROW_SEL
+ pixel_8234/NB1 pixel_8234/VBIAS pixel_8234/NB2 pixel_8234/AMP_IN pixel_8234/SF_IB
+ pixel_8234/PIX_OUT pixel_8234/CSA_VREF pixel
Xpixel_8245 pixel_8245/gring pixel_8245/VDD pixel_8245/GND pixel_8245/VREF pixel_8245/ROW_SEL
+ pixel_8245/NB1 pixel_8245/VBIAS pixel_8245/NB2 pixel_8245/AMP_IN pixel_8245/SF_IB
+ pixel_8245/PIX_OUT pixel_8245/CSA_VREF pixel
Xpixel_8256 pixel_8256/gring pixel_8256/VDD pixel_8256/GND pixel_8256/VREF pixel_8256/ROW_SEL
+ pixel_8256/NB1 pixel_8256/VBIAS pixel_8256/NB2 pixel_8256/AMP_IN pixel_8256/SF_IB
+ pixel_8256/PIX_OUT pixel_8256/CSA_VREF pixel
Xpixel_8267 pixel_8267/gring pixel_8267/VDD pixel_8267/GND pixel_8267/VREF pixel_8267/ROW_SEL
+ pixel_8267/NB1 pixel_8267/VBIAS pixel_8267/NB2 pixel_8267/AMP_IN pixel_8267/SF_IB
+ pixel_8267/PIX_OUT pixel_8267/CSA_VREF pixel
Xpixel_7500 pixel_7500/gring pixel_7500/VDD pixel_7500/GND pixel_7500/VREF pixel_7500/ROW_SEL
+ pixel_7500/NB1 pixel_7500/VBIAS pixel_7500/NB2 pixel_7500/AMP_IN pixel_7500/SF_IB
+ pixel_7500/PIX_OUT pixel_7500/CSA_VREF pixel
Xpixel_7511 pixel_7511/gring pixel_7511/VDD pixel_7511/GND pixel_7511/VREF pixel_7511/ROW_SEL
+ pixel_7511/NB1 pixel_7511/VBIAS pixel_7511/NB2 pixel_7511/AMP_IN pixel_7511/SF_IB
+ pixel_7511/PIX_OUT pixel_7511/CSA_VREF pixel
Xpixel_7522 pixel_7522/gring pixel_7522/VDD pixel_7522/GND pixel_7522/VREF pixel_7522/ROW_SEL
+ pixel_7522/NB1 pixel_7522/VBIAS pixel_7522/NB2 pixel_7522/AMP_IN pixel_7522/SF_IB
+ pixel_7522/PIX_OUT pixel_7522/CSA_VREF pixel
Xpixel_7533 pixel_7533/gring pixel_7533/VDD pixel_7533/GND pixel_7533/VREF pixel_7533/ROW_SEL
+ pixel_7533/NB1 pixel_7533/VBIAS pixel_7533/NB2 pixel_7533/AMP_IN pixel_7533/SF_IB
+ pixel_7533/PIX_OUT pixel_7533/CSA_VREF pixel
Xpixel_8278 pixel_8278/gring pixel_8278/VDD pixel_8278/GND pixel_8278/VREF pixel_8278/ROW_SEL
+ pixel_8278/NB1 pixel_8278/VBIAS pixel_8278/NB2 pixel_8278/AMP_IN pixel_8278/SF_IB
+ pixel_8278/PIX_OUT pixel_8278/CSA_VREF pixel
Xpixel_8289 pixel_8289/gring pixel_8289/VDD pixel_8289/GND pixel_8289/VREF pixel_8289/ROW_SEL
+ pixel_8289/NB1 pixel_8289/VBIAS pixel_8289/NB2 pixel_8289/AMP_IN pixel_8289/SF_IB
+ pixel_8289/PIX_OUT pixel_8289/CSA_VREF pixel
Xpixel_7544 pixel_7544/gring pixel_7544/VDD pixel_7544/GND pixel_7544/VREF pixel_7544/ROW_SEL
+ pixel_7544/NB1 pixel_7544/VBIAS pixel_7544/NB2 pixel_7544/AMP_IN pixel_7544/SF_IB
+ pixel_7544/PIX_OUT pixel_7544/CSA_VREF pixel
Xpixel_7555 pixel_7555/gring pixel_7555/VDD pixel_7555/GND pixel_7555/VREF pixel_7555/ROW_SEL
+ pixel_7555/NB1 pixel_7555/VBIAS pixel_7555/NB2 pixel_7555/AMP_IN pixel_7555/SF_IB
+ pixel_7555/PIX_OUT pixel_7555/CSA_VREF pixel
Xpixel_7566 pixel_7566/gring pixel_7566/VDD pixel_7566/GND pixel_7566/VREF pixel_7566/ROW_SEL
+ pixel_7566/NB1 pixel_7566/VBIAS pixel_7566/NB2 pixel_7566/AMP_IN pixel_7566/SF_IB
+ pixel_7566/PIX_OUT pixel_7566/CSA_VREF pixel
Xpixel_6810 pixel_6810/gring pixel_6810/VDD pixel_6810/GND pixel_6810/VREF pixel_6810/ROW_SEL
+ pixel_6810/NB1 pixel_6810/VBIAS pixel_6810/NB2 pixel_6810/AMP_IN pixel_6810/SF_IB
+ pixel_6810/PIX_OUT pixel_6810/CSA_VREF pixel
Xpixel_6821 pixel_6821/gring pixel_6821/VDD pixel_6821/GND pixel_6821/VREF pixel_6821/ROW_SEL
+ pixel_6821/NB1 pixel_6821/VBIAS pixel_6821/NB2 pixel_6821/AMP_IN pixel_6821/SF_IB
+ pixel_6821/PIX_OUT pixel_6821/CSA_VREF pixel
Xpixel_7577 pixel_7577/gring pixel_7577/VDD pixel_7577/GND pixel_7577/VREF pixel_7577/ROW_SEL
+ pixel_7577/NB1 pixel_7577/VBIAS pixel_7577/NB2 pixel_7577/AMP_IN pixel_7577/SF_IB
+ pixel_7577/PIX_OUT pixel_7577/CSA_VREF pixel
Xpixel_7588 pixel_7588/gring pixel_7588/VDD pixel_7588/GND pixel_7588/VREF pixel_7588/ROW_SEL
+ pixel_7588/NB1 pixel_7588/VBIAS pixel_7588/NB2 pixel_7588/AMP_IN pixel_7588/SF_IB
+ pixel_7588/PIX_OUT pixel_7588/CSA_VREF pixel
Xpixel_7599 pixel_7599/gring pixel_7599/VDD pixel_7599/GND pixel_7599/VREF pixel_7599/ROW_SEL
+ pixel_7599/NB1 pixel_7599/VBIAS pixel_7599/NB2 pixel_7599/AMP_IN pixel_7599/SF_IB
+ pixel_7599/PIX_OUT pixel_7599/CSA_VREF pixel
Xpixel_6832 pixel_6832/gring pixel_6832/VDD pixel_6832/GND pixel_6832/VREF pixel_6832/ROW_SEL
+ pixel_6832/NB1 pixel_6832/VBIAS pixel_6832/NB2 pixel_6832/AMP_IN pixel_6832/SF_IB
+ pixel_6832/PIX_OUT pixel_6832/CSA_VREF pixel
Xpixel_6843 pixel_6843/gring pixel_6843/VDD pixel_6843/GND pixel_6843/VREF pixel_6843/ROW_SEL
+ pixel_6843/NB1 pixel_6843/VBIAS pixel_6843/NB2 pixel_6843/AMP_IN pixel_6843/SF_IB
+ pixel_6843/PIX_OUT pixel_6843/CSA_VREF pixel
Xpixel_6854 pixel_6854/gring pixel_6854/VDD pixel_6854/GND pixel_6854/VREF pixel_6854/ROW_SEL
+ pixel_6854/NB1 pixel_6854/VBIAS pixel_6854/NB2 pixel_6854/AMP_IN pixel_6854/SF_IB
+ pixel_6854/PIX_OUT pixel_6854/CSA_VREF pixel
Xpixel_6865 pixel_6865/gring pixel_6865/VDD pixel_6865/GND pixel_6865/VREF pixel_6865/ROW_SEL
+ pixel_6865/NB1 pixel_6865/VBIAS pixel_6865/NB2 pixel_6865/AMP_IN pixel_6865/SF_IB
+ pixel_6865/PIX_OUT pixel_6865/CSA_VREF pixel
Xpixel_6876 pixel_6876/gring pixel_6876/VDD pixel_6876/GND pixel_6876/VREF pixel_6876/ROW_SEL
+ pixel_6876/NB1 pixel_6876/VBIAS pixel_6876/NB2 pixel_6876/AMP_IN pixel_6876/SF_IB
+ pixel_6876/PIX_OUT pixel_6876/CSA_VREF pixel
Xpixel_6887 pixel_6887/gring pixel_6887/VDD pixel_6887/GND pixel_6887/VREF pixel_6887/ROW_SEL
+ pixel_6887/NB1 pixel_6887/VBIAS pixel_6887/NB2 pixel_6887/AMP_IN pixel_6887/SF_IB
+ pixel_6887/PIX_OUT pixel_6887/CSA_VREF pixel
Xpixel_6898 pixel_6898/gring pixel_6898/VDD pixel_6898/GND pixel_6898/VREF pixel_6898/ROW_SEL
+ pixel_6898/NB1 pixel_6898/VBIAS pixel_6898/NB2 pixel_6898/AMP_IN pixel_6898/SF_IB
+ pixel_6898/PIX_OUT pixel_6898/CSA_VREF pixel
Xpixel_1150 pixel_1150/gring pixel_1150/VDD pixel_1150/GND pixel_1150/VREF pixel_1150/ROW_SEL
+ pixel_1150/NB1 pixel_1150/VBIAS pixel_1150/NB2 pixel_1150/AMP_IN pixel_1150/SF_IB
+ pixel_1150/PIX_OUT pixel_1150/CSA_VREF pixel
Xpixel_1183 pixel_1183/gring pixel_1183/VDD pixel_1183/GND pixel_1183/VREF pixel_1183/ROW_SEL
+ pixel_1183/NB1 pixel_1183/VBIAS pixel_1183/NB2 pixel_1183/AMP_IN pixel_1183/SF_IB
+ pixel_1183/PIX_OUT pixel_1183/CSA_VREF pixel
Xpixel_1172 pixel_1172/gring pixel_1172/VDD pixel_1172/GND pixel_1172/VREF pixel_1172/ROW_SEL
+ pixel_1172/NB1 pixel_1172/VBIAS pixel_1172/NB2 pixel_1172/AMP_IN pixel_1172/SF_IB
+ pixel_1172/PIX_OUT pixel_1172/CSA_VREF pixel
Xpixel_1161 pixel_1161/gring pixel_1161/VDD pixel_1161/GND pixel_1161/VREF pixel_1161/ROW_SEL
+ pixel_1161/NB1 pixel_1161/VBIAS pixel_1161/NB2 pixel_1161/AMP_IN pixel_1161/SF_IB
+ pixel_1161/PIX_OUT pixel_1161/CSA_VREF pixel
Xpixel_1194 pixel_1194/gring pixel_1194/VDD pixel_1194/GND pixel_1194/VREF pixel_1194/ROW_SEL
+ pixel_1194/NB1 pixel_1194/VBIAS pixel_1194/NB2 pixel_1194/AMP_IN pixel_1194/SF_IB
+ pixel_1194/PIX_OUT pixel_1194/CSA_VREF pixel
Xpixel_9491 pixel_9491/gring pixel_9491/VDD pixel_9491/GND pixel_9491/VREF pixel_9491/ROW_SEL
+ pixel_9491/NB1 pixel_9491/VBIAS pixel_9491/NB2 pixel_9491/AMP_IN pixel_9491/SF_IB
+ pixel_9491/PIX_OUT pixel_9491/CSA_VREF pixel
Xpixel_9480 pixel_9480/gring pixel_9480/VDD pixel_9480/GND pixel_9480/VREF pixel_9480/ROW_SEL
+ pixel_9480/NB1 pixel_9480/VBIAS pixel_9480/NB2 pixel_9480/AMP_IN pixel_9480/SF_IB
+ pixel_9480/PIX_OUT pixel_9480/CSA_VREF pixel
Xpixel_8790 pixel_8790/gring pixel_8790/VDD pixel_8790/GND pixel_8790/VREF pixel_8790/ROW_SEL
+ pixel_8790/NB1 pixel_8790/VBIAS pixel_8790/NB2 pixel_8790/AMP_IN pixel_8790/SF_IB
+ pixel_8790/PIX_OUT pixel_8790/CSA_VREF pixel
Xpixel_209 pixel_209/gring pixel_209/VDD pixel_209/GND pixel_209/VREF pixel_209/ROW_SEL
+ pixel_209/NB1 pixel_209/VBIAS pixel_209/NB2 pixel_209/AMP_IN pixel_209/SF_IB pixel_209/PIX_OUT
+ pixel_209/CSA_VREF pixel
Xpixel_6106 pixel_6106/gring pixel_6106/VDD pixel_6106/GND pixel_6106/VREF pixel_6106/ROW_SEL
+ pixel_6106/NB1 pixel_6106/VBIAS pixel_6106/NB2 pixel_6106/AMP_IN pixel_6106/SF_IB
+ pixel_6106/PIX_OUT pixel_6106/CSA_VREF pixel
Xpixel_6117 pixel_6117/gring pixel_6117/VDD pixel_6117/GND pixel_6117/VREF pixel_6117/ROW_SEL
+ pixel_6117/NB1 pixel_6117/VBIAS pixel_6117/NB2 pixel_6117/AMP_IN pixel_6117/SF_IB
+ pixel_6117/PIX_OUT pixel_6117/CSA_VREF pixel
Xpixel_6128 pixel_6128/gring pixel_6128/VDD pixel_6128/GND pixel_6128/VREF pixel_6128/ROW_SEL
+ pixel_6128/NB1 pixel_6128/VBIAS pixel_6128/NB2 pixel_6128/AMP_IN pixel_6128/SF_IB
+ pixel_6128/PIX_OUT pixel_6128/CSA_VREF pixel
Xpixel_6139 pixel_6139/gring pixel_6139/VDD pixel_6139/GND pixel_6139/VREF pixel_6139/ROW_SEL
+ pixel_6139/NB1 pixel_6139/VBIAS pixel_6139/NB2 pixel_6139/AMP_IN pixel_6139/SF_IB
+ pixel_6139/PIX_OUT pixel_6139/CSA_VREF pixel
Xpixel_5405 pixel_5405/gring pixel_5405/VDD pixel_5405/GND pixel_5405/VREF pixel_5405/ROW_SEL
+ pixel_5405/NB1 pixel_5405/VBIAS pixel_5405/NB2 pixel_5405/AMP_IN pixel_5405/SF_IB
+ pixel_5405/PIX_OUT pixel_5405/CSA_VREF pixel
Xpixel_5416 pixel_5416/gring pixel_5416/VDD pixel_5416/GND pixel_5416/VREF pixel_5416/ROW_SEL
+ pixel_5416/NB1 pixel_5416/VBIAS pixel_5416/NB2 pixel_5416/AMP_IN pixel_5416/SF_IB
+ pixel_5416/PIX_OUT pixel_5416/CSA_VREF pixel
Xpixel_5427 pixel_5427/gring pixel_5427/VDD pixel_5427/GND pixel_5427/VREF pixel_5427/ROW_SEL
+ pixel_5427/NB1 pixel_5427/VBIAS pixel_5427/NB2 pixel_5427/AMP_IN pixel_5427/SF_IB
+ pixel_5427/PIX_OUT pixel_5427/CSA_VREF pixel
Xpixel_5438 pixel_5438/gring pixel_5438/VDD pixel_5438/GND pixel_5438/VREF pixel_5438/ROW_SEL
+ pixel_5438/NB1 pixel_5438/VBIAS pixel_5438/NB2 pixel_5438/AMP_IN pixel_5438/SF_IB
+ pixel_5438/PIX_OUT pixel_5438/CSA_VREF pixel
Xpixel_4704 pixel_4704/gring pixel_4704/VDD pixel_4704/GND pixel_4704/VREF pixel_4704/ROW_SEL
+ pixel_4704/NB1 pixel_4704/VBIAS pixel_4704/NB2 pixel_4704/AMP_IN pixel_4704/SF_IB
+ pixel_4704/PIX_OUT pixel_4704/CSA_VREF pixel
Xpixel_732 pixel_732/gring pixel_732/VDD pixel_732/GND pixel_732/VREF pixel_732/ROW_SEL
+ pixel_732/NB1 pixel_732/VBIAS pixel_732/NB2 pixel_732/AMP_IN pixel_732/SF_IB pixel_732/PIX_OUT
+ pixel_732/CSA_VREF pixel
Xpixel_721 pixel_721/gring pixel_721/VDD pixel_721/GND pixel_721/VREF pixel_721/ROW_SEL
+ pixel_721/NB1 pixel_721/VBIAS pixel_721/NB2 pixel_721/AMP_IN pixel_721/SF_IB pixel_721/PIX_OUT
+ pixel_721/CSA_VREF pixel
Xpixel_710 pixel_710/gring pixel_710/VDD pixel_710/GND pixel_710/VREF pixel_710/ROW_SEL
+ pixel_710/NB1 pixel_710/VBIAS pixel_710/NB2 pixel_710/AMP_IN pixel_710/SF_IB pixel_710/PIX_OUT
+ pixel_710/CSA_VREF pixel
Xpixel_5449 pixel_5449/gring pixel_5449/VDD pixel_5449/GND pixel_5449/VREF pixel_5449/ROW_SEL
+ pixel_5449/NB1 pixel_5449/VBIAS pixel_5449/NB2 pixel_5449/AMP_IN pixel_5449/SF_IB
+ pixel_5449/PIX_OUT pixel_5449/CSA_VREF pixel
Xpixel_4715 pixel_4715/gring pixel_4715/VDD pixel_4715/GND pixel_4715/VREF pixel_4715/ROW_SEL
+ pixel_4715/NB1 pixel_4715/VBIAS pixel_4715/NB2 pixel_4715/AMP_IN pixel_4715/SF_IB
+ pixel_4715/PIX_OUT pixel_4715/CSA_VREF pixel
Xpixel_4726 pixel_4726/gring pixel_4726/VDD pixel_4726/GND pixel_4726/VREF pixel_4726/ROW_SEL
+ pixel_4726/NB1 pixel_4726/VBIAS pixel_4726/NB2 pixel_4726/AMP_IN pixel_4726/SF_IB
+ pixel_4726/PIX_OUT pixel_4726/CSA_VREF pixel
Xpixel_4737 pixel_4737/gring pixel_4737/VDD pixel_4737/GND pixel_4737/VREF pixel_4737/ROW_SEL
+ pixel_4737/NB1 pixel_4737/VBIAS pixel_4737/NB2 pixel_4737/AMP_IN pixel_4737/SF_IB
+ pixel_4737/PIX_OUT pixel_4737/CSA_VREF pixel
Xpixel_765 pixel_765/gring pixel_765/VDD pixel_765/GND pixel_765/VREF pixel_765/ROW_SEL
+ pixel_765/NB1 pixel_765/VBIAS pixel_765/NB2 pixel_765/AMP_IN pixel_765/SF_IB pixel_765/PIX_OUT
+ pixel_765/CSA_VREF pixel
Xpixel_754 pixel_754/gring pixel_754/VDD pixel_754/GND pixel_754/VREF pixel_754/ROW_SEL
+ pixel_754/NB1 pixel_754/VBIAS pixel_754/NB2 pixel_754/AMP_IN pixel_754/SF_IB pixel_754/PIX_OUT
+ pixel_754/CSA_VREF pixel
Xpixel_743 pixel_743/gring pixel_743/VDD pixel_743/GND pixel_743/VREF pixel_743/ROW_SEL
+ pixel_743/NB1 pixel_743/VBIAS pixel_743/NB2 pixel_743/AMP_IN pixel_743/SF_IB pixel_743/PIX_OUT
+ pixel_743/CSA_VREF pixel
Xpixel_4748 pixel_4748/gring pixel_4748/VDD pixel_4748/GND pixel_4748/VREF pixel_4748/ROW_SEL
+ pixel_4748/NB1 pixel_4748/VBIAS pixel_4748/NB2 pixel_4748/AMP_IN pixel_4748/SF_IB
+ pixel_4748/PIX_OUT pixel_4748/CSA_VREF pixel
Xpixel_4759 pixel_4759/gring pixel_4759/VDD pixel_4759/GND pixel_4759/VREF pixel_4759/ROW_SEL
+ pixel_4759/NB1 pixel_4759/VBIAS pixel_4759/NB2 pixel_4759/AMP_IN pixel_4759/SF_IB
+ pixel_4759/PIX_OUT pixel_4759/CSA_VREF pixel
Xpixel_798 pixel_798/gring pixel_798/VDD pixel_798/GND pixel_798/VREF pixel_798/ROW_SEL
+ pixel_798/NB1 pixel_798/VBIAS pixel_798/NB2 pixel_798/AMP_IN pixel_798/SF_IB pixel_798/PIX_OUT
+ pixel_798/CSA_VREF pixel
Xpixel_787 pixel_787/gring pixel_787/VDD pixel_787/GND pixel_787/VREF pixel_787/ROW_SEL
+ pixel_787/NB1 pixel_787/VBIAS pixel_787/NB2 pixel_787/AMP_IN pixel_787/SF_IB pixel_787/PIX_OUT
+ pixel_787/CSA_VREF pixel
Xpixel_776 pixel_776/gring pixel_776/VDD pixel_776/GND pixel_776/VREF pixel_776/ROW_SEL
+ pixel_776/NB1 pixel_776/VBIAS pixel_776/NB2 pixel_776/AMP_IN pixel_776/SF_IB pixel_776/PIX_OUT
+ pixel_776/CSA_VREF pixel
Xpixel_8020 pixel_8020/gring pixel_8020/VDD pixel_8020/GND pixel_8020/VREF pixel_8020/ROW_SEL
+ pixel_8020/NB1 pixel_8020/VBIAS pixel_8020/NB2 pixel_8020/AMP_IN pixel_8020/SF_IB
+ pixel_8020/PIX_OUT pixel_8020/CSA_VREF pixel
Xpixel_8031 pixel_8031/gring pixel_8031/VDD pixel_8031/GND pixel_8031/VREF pixel_8031/ROW_SEL
+ pixel_8031/NB1 pixel_8031/VBIAS pixel_8031/NB2 pixel_8031/AMP_IN pixel_8031/SF_IB
+ pixel_8031/PIX_OUT pixel_8031/CSA_VREF pixel
Xpixel_8042 pixel_8042/gring pixel_8042/VDD pixel_8042/GND pixel_8042/VREF pixel_8042/ROW_SEL
+ pixel_8042/NB1 pixel_8042/VBIAS pixel_8042/NB2 pixel_8042/AMP_IN pixel_8042/SF_IB
+ pixel_8042/PIX_OUT pixel_8042/CSA_VREF pixel
Xpixel_8053 pixel_8053/gring pixel_8053/VDD pixel_8053/GND pixel_8053/VREF pixel_8053/ROW_SEL
+ pixel_8053/NB1 pixel_8053/VBIAS pixel_8053/NB2 pixel_8053/AMP_IN pixel_8053/SF_IB
+ pixel_8053/PIX_OUT pixel_8053/CSA_VREF pixel
Xpixel_8064 pixel_8064/gring pixel_8064/VDD pixel_8064/GND pixel_8064/VREF pixel_8064/ROW_SEL
+ pixel_8064/NB1 pixel_8064/VBIAS pixel_8064/NB2 pixel_8064/AMP_IN pixel_8064/SF_IB
+ pixel_8064/PIX_OUT pixel_8064/CSA_VREF pixel
Xpixel_8075 pixel_8075/gring pixel_8075/VDD pixel_8075/GND pixel_8075/VREF pixel_8075/ROW_SEL
+ pixel_8075/NB1 pixel_8075/VBIAS pixel_8075/NB2 pixel_8075/AMP_IN pixel_8075/SF_IB
+ pixel_8075/PIX_OUT pixel_8075/CSA_VREF pixel
Xpixel_8086 pixel_8086/gring pixel_8086/VDD pixel_8086/GND pixel_8086/VREF pixel_8086/ROW_SEL
+ pixel_8086/NB1 pixel_8086/VBIAS pixel_8086/NB2 pixel_8086/AMP_IN pixel_8086/SF_IB
+ pixel_8086/PIX_OUT pixel_8086/CSA_VREF pixel
Xpixel_7330 pixel_7330/gring pixel_7330/VDD pixel_7330/GND pixel_7330/VREF pixel_7330/ROW_SEL
+ pixel_7330/NB1 pixel_7330/VBIAS pixel_7330/NB2 pixel_7330/AMP_IN pixel_7330/SF_IB
+ pixel_7330/PIX_OUT pixel_7330/CSA_VREF pixel
Xpixel_7341 pixel_7341/gring pixel_7341/VDD pixel_7341/GND pixel_7341/VREF pixel_7341/ROW_SEL
+ pixel_7341/NB1 pixel_7341/VBIAS pixel_7341/NB2 pixel_7341/AMP_IN pixel_7341/SF_IB
+ pixel_7341/PIX_OUT pixel_7341/CSA_VREF pixel
Xpixel_8097 pixel_8097/gring pixel_8097/VDD pixel_8097/GND pixel_8097/VREF pixel_8097/ROW_SEL
+ pixel_8097/NB1 pixel_8097/VBIAS pixel_8097/NB2 pixel_8097/AMP_IN pixel_8097/SF_IB
+ pixel_8097/PIX_OUT pixel_8097/CSA_VREF pixel
Xpixel_7352 pixel_7352/gring pixel_7352/VDD pixel_7352/GND pixel_7352/VREF pixel_7352/ROW_SEL
+ pixel_7352/NB1 pixel_7352/VBIAS pixel_7352/NB2 pixel_7352/AMP_IN pixel_7352/SF_IB
+ pixel_7352/PIX_OUT pixel_7352/CSA_VREF pixel
Xpixel_7363 pixel_7363/gring pixel_7363/VDD pixel_7363/GND pixel_7363/VREF pixel_7363/ROW_SEL
+ pixel_7363/NB1 pixel_7363/VBIAS pixel_7363/NB2 pixel_7363/AMP_IN pixel_7363/SF_IB
+ pixel_7363/PIX_OUT pixel_7363/CSA_VREF pixel
Xpixel_7374 pixel_7374/gring pixel_7374/VDD pixel_7374/GND pixel_7374/VREF pixel_7374/ROW_SEL
+ pixel_7374/NB1 pixel_7374/VBIAS pixel_7374/NB2 pixel_7374/AMP_IN pixel_7374/SF_IB
+ pixel_7374/PIX_OUT pixel_7374/CSA_VREF pixel
Xpixel_7385 pixel_7385/gring pixel_7385/VDD pixel_7385/GND pixel_7385/VREF pixel_7385/ROW_SEL
+ pixel_7385/NB1 pixel_7385/VBIAS pixel_7385/NB2 pixel_7385/AMP_IN pixel_7385/SF_IB
+ pixel_7385/PIX_OUT pixel_7385/CSA_VREF pixel
Xpixel_7396 pixel_7396/gring pixel_7396/VDD pixel_7396/GND pixel_7396/VREF pixel_7396/ROW_SEL
+ pixel_7396/NB1 pixel_7396/VBIAS pixel_7396/NB2 pixel_7396/AMP_IN pixel_7396/SF_IB
+ pixel_7396/PIX_OUT pixel_7396/CSA_VREF pixel
Xpixel_6640 pixel_6640/gring pixel_6640/VDD pixel_6640/GND pixel_6640/VREF pixel_6640/ROW_SEL
+ pixel_6640/NB1 pixel_6640/VBIAS pixel_6640/NB2 pixel_6640/AMP_IN pixel_6640/SF_IB
+ pixel_6640/PIX_OUT pixel_6640/CSA_VREF pixel
Xpixel_6651 pixel_6651/gring pixel_6651/VDD pixel_6651/GND pixel_6651/VREF pixel_6651/ROW_SEL
+ pixel_6651/NB1 pixel_6651/VBIAS pixel_6651/NB2 pixel_6651/AMP_IN pixel_6651/SF_IB
+ pixel_6651/PIX_OUT pixel_6651/CSA_VREF pixel
Xpixel_6662 pixel_6662/gring pixel_6662/VDD pixel_6662/GND pixel_6662/VREF pixel_6662/ROW_SEL
+ pixel_6662/NB1 pixel_6662/VBIAS pixel_6662/NB2 pixel_6662/AMP_IN pixel_6662/SF_IB
+ pixel_6662/PIX_OUT pixel_6662/CSA_VREF pixel
Xpixel_6673 pixel_6673/gring pixel_6673/VDD pixel_6673/GND pixel_6673/VREF pixel_6673/ROW_SEL
+ pixel_6673/NB1 pixel_6673/VBIAS pixel_6673/NB2 pixel_6673/AMP_IN pixel_6673/SF_IB
+ pixel_6673/PIX_OUT pixel_6673/CSA_VREF pixel
Xpixel_6684 pixel_6684/gring pixel_6684/VDD pixel_6684/GND pixel_6684/VREF pixel_6684/ROW_SEL
+ pixel_6684/NB1 pixel_6684/VBIAS pixel_6684/NB2 pixel_6684/AMP_IN pixel_6684/SF_IB
+ pixel_6684/PIX_OUT pixel_6684/CSA_VREF pixel
Xpixel_6695 pixel_6695/gring pixel_6695/VDD pixel_6695/GND pixel_6695/VREF pixel_6695/ROW_SEL
+ pixel_6695/NB1 pixel_6695/VBIAS pixel_6695/NB2 pixel_6695/AMP_IN pixel_6695/SF_IB
+ pixel_6695/PIX_OUT pixel_6695/CSA_VREF pixel
Xpixel_5950 pixel_5950/gring pixel_5950/VDD pixel_5950/GND pixel_5950/VREF pixel_5950/ROW_SEL
+ pixel_5950/NB1 pixel_5950/VBIAS pixel_5950/NB2 pixel_5950/AMP_IN pixel_5950/SF_IB
+ pixel_5950/PIX_OUT pixel_5950/CSA_VREF pixel
Xpixel_5961 pixel_5961/gring pixel_5961/VDD pixel_5961/GND pixel_5961/VREF pixel_5961/ROW_SEL
+ pixel_5961/NB1 pixel_5961/VBIAS pixel_5961/NB2 pixel_5961/AMP_IN pixel_5961/SF_IB
+ pixel_5961/PIX_OUT pixel_5961/CSA_VREF pixel
Xpixel_5972 pixel_5972/gring pixel_5972/VDD pixel_5972/GND pixel_5972/VREF pixel_5972/ROW_SEL
+ pixel_5972/NB1 pixel_5972/VBIAS pixel_5972/NB2 pixel_5972/AMP_IN pixel_5972/SF_IB
+ pixel_5972/PIX_OUT pixel_5972/CSA_VREF pixel
Xpixel_5983 pixel_5983/gring pixel_5983/VDD pixel_5983/GND pixel_5983/VREF pixel_5983/ROW_SEL
+ pixel_5983/NB1 pixel_5983/VBIAS pixel_5983/NB2 pixel_5983/AMP_IN pixel_5983/SF_IB
+ pixel_5983/PIX_OUT pixel_5983/CSA_VREF pixel
Xpixel_5994 pixel_5994/gring pixel_5994/VDD pixel_5994/GND pixel_5994/VREF pixel_5994/ROW_SEL
+ pixel_5994/NB1 pixel_5994/VBIAS pixel_5994/NB2 pixel_5994/AMP_IN pixel_5994/SF_IB
+ pixel_5994/PIX_OUT pixel_5994/CSA_VREF pixel
Xpixel_2609 pixel_2609/gring pixel_2609/VDD pixel_2609/GND pixel_2609/VREF pixel_2609/ROW_SEL
+ pixel_2609/NB1 pixel_2609/VBIAS pixel_2609/NB2 pixel_2609/AMP_IN pixel_2609/SF_IB
+ pixel_2609/PIX_OUT pixel_2609/CSA_VREF pixel
Xpixel_1908 pixel_1908/gring pixel_1908/VDD pixel_1908/GND pixel_1908/VREF pixel_1908/ROW_SEL
+ pixel_1908/NB1 pixel_1908/VBIAS pixel_1908/NB2 pixel_1908/AMP_IN pixel_1908/SF_IB
+ pixel_1908/PIX_OUT pixel_1908/CSA_VREF pixel
Xpixel_1919 pixel_1919/gring pixel_1919/VDD pixel_1919/GND pixel_1919/VREF pixel_1919/ROW_SEL
+ pixel_1919/NB1 pixel_1919/VBIAS pixel_1919/NB2 pixel_1919/AMP_IN pixel_1919/SF_IB
+ pixel_1919/PIX_OUT pixel_1919/CSA_VREF pixel
Xpixel_5202 pixel_5202/gring pixel_5202/VDD pixel_5202/GND pixel_5202/VREF pixel_5202/ROW_SEL
+ pixel_5202/NB1 pixel_5202/VBIAS pixel_5202/NB2 pixel_5202/AMP_IN pixel_5202/SF_IB
+ pixel_5202/PIX_OUT pixel_5202/CSA_VREF pixel
Xpixel_5213 pixel_5213/gring pixel_5213/VDD pixel_5213/GND pixel_5213/VREF pixel_5213/ROW_SEL
+ pixel_5213/NB1 pixel_5213/VBIAS pixel_5213/NB2 pixel_5213/AMP_IN pixel_5213/SF_IB
+ pixel_5213/PIX_OUT pixel_5213/CSA_VREF pixel
Xpixel_5224 pixel_5224/gring pixel_5224/VDD pixel_5224/GND pixel_5224/VREF pixel_5224/ROW_SEL
+ pixel_5224/NB1 pixel_5224/VBIAS pixel_5224/NB2 pixel_5224/AMP_IN pixel_5224/SF_IB
+ pixel_5224/PIX_OUT pixel_5224/CSA_VREF pixel
Xpixel_5235 pixel_5235/gring pixel_5235/VDD pixel_5235/GND pixel_5235/VREF pixel_5235/ROW_SEL
+ pixel_5235/NB1 pixel_5235/VBIAS pixel_5235/NB2 pixel_5235/AMP_IN pixel_5235/SF_IB
+ pixel_5235/PIX_OUT pixel_5235/CSA_VREF pixel
Xpixel_5246 pixel_5246/gring pixel_5246/VDD pixel_5246/GND pixel_5246/VREF pixel_5246/ROW_SEL
+ pixel_5246/NB1 pixel_5246/VBIAS pixel_5246/NB2 pixel_5246/AMP_IN pixel_5246/SF_IB
+ pixel_5246/PIX_OUT pixel_5246/CSA_VREF pixel
Xpixel_5257 pixel_5257/gring pixel_5257/VDD pixel_5257/GND pixel_5257/VREF pixel_5257/ROW_SEL
+ pixel_5257/NB1 pixel_5257/VBIAS pixel_5257/NB2 pixel_5257/AMP_IN pixel_5257/SF_IB
+ pixel_5257/PIX_OUT pixel_5257/CSA_VREF pixel
Xpixel_4501 pixel_4501/gring pixel_4501/VDD pixel_4501/GND pixel_4501/VREF pixel_4501/ROW_SEL
+ pixel_4501/NB1 pixel_4501/VBIAS pixel_4501/NB2 pixel_4501/AMP_IN pixel_4501/SF_IB
+ pixel_4501/PIX_OUT pixel_4501/CSA_VREF pixel
Xpixel_4512 pixel_4512/gring pixel_4512/VDD pixel_4512/GND pixel_4512/VREF pixel_4512/ROW_SEL
+ pixel_4512/NB1 pixel_4512/VBIAS pixel_4512/NB2 pixel_4512/AMP_IN pixel_4512/SF_IB
+ pixel_4512/PIX_OUT pixel_4512/CSA_VREF pixel
Xpixel_540 pixel_540/gring pixel_540/VDD pixel_540/GND pixel_540/VREF pixel_540/ROW_SEL
+ pixel_540/NB1 pixel_540/VBIAS pixel_540/NB2 pixel_540/AMP_IN pixel_540/SF_IB pixel_540/PIX_OUT
+ pixel_540/CSA_VREF pixel
Xpixel_5268 pixel_5268/gring pixel_5268/VDD pixel_5268/GND pixel_5268/VREF pixel_5268/ROW_SEL
+ pixel_5268/NB1 pixel_5268/VBIAS pixel_5268/NB2 pixel_5268/AMP_IN pixel_5268/SF_IB
+ pixel_5268/PIX_OUT pixel_5268/CSA_VREF pixel
Xpixel_5279 pixel_5279/gring pixel_5279/VDD pixel_5279/GND pixel_5279/VREF pixel_5279/ROW_SEL
+ pixel_5279/NB1 pixel_5279/VBIAS pixel_5279/NB2 pixel_5279/AMP_IN pixel_5279/SF_IB
+ pixel_5279/PIX_OUT pixel_5279/CSA_VREF pixel
Xpixel_4523 pixel_4523/gring pixel_4523/VDD pixel_4523/GND pixel_4523/VREF pixel_4523/ROW_SEL
+ pixel_4523/NB1 pixel_4523/VBIAS pixel_4523/NB2 pixel_4523/AMP_IN pixel_4523/SF_IB
+ pixel_4523/PIX_OUT pixel_4523/CSA_VREF pixel
Xpixel_4534 pixel_4534/gring pixel_4534/VDD pixel_4534/GND pixel_4534/VREF pixel_4534/ROW_SEL
+ pixel_4534/NB1 pixel_4534/VBIAS pixel_4534/NB2 pixel_4534/AMP_IN pixel_4534/SF_IB
+ pixel_4534/PIX_OUT pixel_4534/CSA_VREF pixel
Xpixel_4545 pixel_4545/gring pixel_4545/VDD pixel_4545/GND pixel_4545/VREF pixel_4545/ROW_SEL
+ pixel_4545/NB1 pixel_4545/VBIAS pixel_4545/NB2 pixel_4545/AMP_IN pixel_4545/SF_IB
+ pixel_4545/PIX_OUT pixel_4545/CSA_VREF pixel
Xpixel_3800 pixel_3800/gring pixel_3800/VDD pixel_3800/GND pixel_3800/VREF pixel_3800/ROW_SEL
+ pixel_3800/NB1 pixel_3800/VBIAS pixel_3800/NB2 pixel_3800/AMP_IN pixel_3800/SF_IB
+ pixel_3800/PIX_OUT pixel_3800/CSA_VREF pixel
Xpixel_584 pixel_584/gring pixel_584/VDD pixel_584/GND pixel_584/VREF pixel_584/ROW_SEL
+ pixel_584/NB1 pixel_584/VBIAS pixel_584/NB2 pixel_584/AMP_IN pixel_584/SF_IB pixel_584/PIX_OUT
+ pixel_584/CSA_VREF pixel
Xpixel_573 pixel_573/gring pixel_573/VDD pixel_573/GND pixel_573/VREF pixel_573/ROW_SEL
+ pixel_573/NB1 pixel_573/VBIAS pixel_573/NB2 pixel_573/AMP_IN pixel_573/SF_IB pixel_573/PIX_OUT
+ pixel_573/CSA_VREF pixel
Xpixel_562 pixel_562/gring pixel_562/VDD pixel_562/GND pixel_562/VREF pixel_562/ROW_SEL
+ pixel_562/NB1 pixel_562/VBIAS pixel_562/NB2 pixel_562/AMP_IN pixel_562/SF_IB pixel_562/PIX_OUT
+ pixel_562/CSA_VREF pixel
Xpixel_551 pixel_551/gring pixel_551/VDD pixel_551/GND pixel_551/VREF pixel_551/ROW_SEL
+ pixel_551/NB1 pixel_551/VBIAS pixel_551/NB2 pixel_551/AMP_IN pixel_551/SF_IB pixel_551/PIX_OUT
+ pixel_551/CSA_VREF pixel
Xpixel_3844 pixel_3844/gring pixel_3844/VDD pixel_3844/GND pixel_3844/VREF pixel_3844/ROW_SEL
+ pixel_3844/NB1 pixel_3844/VBIAS pixel_3844/NB2 pixel_3844/AMP_IN pixel_3844/SF_IB
+ pixel_3844/PIX_OUT pixel_3844/CSA_VREF pixel
Xpixel_4556 pixel_4556/gring pixel_4556/VDD pixel_4556/GND pixel_4556/VREF pixel_4556/ROW_SEL
+ pixel_4556/NB1 pixel_4556/VBIAS pixel_4556/NB2 pixel_4556/AMP_IN pixel_4556/SF_IB
+ pixel_4556/PIX_OUT pixel_4556/CSA_VREF pixel
Xpixel_4567 pixel_4567/gring pixel_4567/VDD pixel_4567/GND pixel_4567/VREF pixel_4567/ROW_SEL
+ pixel_4567/NB1 pixel_4567/VBIAS pixel_4567/NB2 pixel_4567/AMP_IN pixel_4567/SF_IB
+ pixel_4567/PIX_OUT pixel_4567/CSA_VREF pixel
Xpixel_4578 pixel_4578/gring pixel_4578/VDD pixel_4578/GND pixel_4578/VREF pixel_4578/ROW_SEL
+ pixel_4578/NB1 pixel_4578/VBIAS pixel_4578/NB2 pixel_4578/AMP_IN pixel_4578/SF_IB
+ pixel_4578/PIX_OUT pixel_4578/CSA_VREF pixel
Xpixel_3811 pixel_3811/gring pixel_3811/VDD pixel_3811/GND pixel_3811/VREF pixel_3811/ROW_SEL
+ pixel_3811/NB1 pixel_3811/VBIAS pixel_3811/NB2 pixel_3811/AMP_IN pixel_3811/SF_IB
+ pixel_3811/PIX_OUT pixel_3811/CSA_VREF pixel
Xpixel_3822 pixel_3822/gring pixel_3822/VDD pixel_3822/GND pixel_3822/VREF pixel_3822/ROW_SEL
+ pixel_3822/NB1 pixel_3822/VBIAS pixel_3822/NB2 pixel_3822/AMP_IN pixel_3822/SF_IB
+ pixel_3822/PIX_OUT pixel_3822/CSA_VREF pixel
Xpixel_3833 pixel_3833/gring pixel_3833/VDD pixel_3833/GND pixel_3833/VREF pixel_3833/ROW_SEL
+ pixel_3833/NB1 pixel_3833/VBIAS pixel_3833/NB2 pixel_3833/AMP_IN pixel_3833/SF_IB
+ pixel_3833/PIX_OUT pixel_3833/CSA_VREF pixel
Xpixel_595 pixel_595/gring pixel_595/VDD pixel_595/GND pixel_595/VREF pixel_595/ROW_SEL
+ pixel_595/NB1 pixel_595/VBIAS pixel_595/NB2 pixel_595/AMP_IN pixel_595/SF_IB pixel_595/PIX_OUT
+ pixel_595/CSA_VREF pixel
Xpixel_3877 pixel_3877/gring pixel_3877/VDD pixel_3877/GND pixel_3877/VREF pixel_3877/ROW_SEL
+ pixel_3877/NB1 pixel_3877/VBIAS pixel_3877/NB2 pixel_3877/AMP_IN pixel_3877/SF_IB
+ pixel_3877/PIX_OUT pixel_3877/CSA_VREF pixel
Xpixel_3866 pixel_3866/gring pixel_3866/VDD pixel_3866/GND pixel_3866/VREF pixel_3866/ROW_SEL
+ pixel_3866/NB1 pixel_3866/VBIAS pixel_3866/NB2 pixel_3866/AMP_IN pixel_3866/SF_IB
+ pixel_3866/PIX_OUT pixel_3866/CSA_VREF pixel
Xpixel_3855 pixel_3855/gring pixel_3855/VDD pixel_3855/GND pixel_3855/VREF pixel_3855/ROW_SEL
+ pixel_3855/NB1 pixel_3855/VBIAS pixel_3855/NB2 pixel_3855/AMP_IN pixel_3855/SF_IB
+ pixel_3855/PIX_OUT pixel_3855/CSA_VREF pixel
Xpixel_4589 pixel_4589/gring pixel_4589/VDD pixel_4589/GND pixel_4589/VREF pixel_4589/ROW_SEL
+ pixel_4589/NB1 pixel_4589/VBIAS pixel_4589/NB2 pixel_4589/AMP_IN pixel_4589/SF_IB
+ pixel_4589/PIX_OUT pixel_4589/CSA_VREF pixel
Xpixel_3899 pixel_3899/gring pixel_3899/VDD pixel_3899/GND pixel_3899/VREF pixel_3899/ROW_SEL
+ pixel_3899/NB1 pixel_3899/VBIAS pixel_3899/NB2 pixel_3899/AMP_IN pixel_3899/SF_IB
+ pixel_3899/PIX_OUT pixel_3899/CSA_VREF pixel
Xpixel_3888 pixel_3888/gring pixel_3888/VDD pixel_3888/GND pixel_3888/VREF pixel_3888/ROW_SEL
+ pixel_3888/NB1 pixel_3888/VBIAS pixel_3888/NB2 pixel_3888/AMP_IN pixel_3888/SF_IB
+ pixel_3888/PIX_OUT pixel_3888/CSA_VREF pixel
Xpixel_7160 pixel_7160/gring pixel_7160/VDD pixel_7160/GND pixel_7160/VREF pixel_7160/ROW_SEL
+ pixel_7160/NB1 pixel_7160/VBIAS pixel_7160/NB2 pixel_7160/AMP_IN pixel_7160/SF_IB
+ pixel_7160/PIX_OUT pixel_7160/CSA_VREF pixel
Xpixel_7171 pixel_7171/gring pixel_7171/VDD pixel_7171/GND pixel_7171/VREF pixel_7171/ROW_SEL
+ pixel_7171/NB1 pixel_7171/VBIAS pixel_7171/NB2 pixel_7171/AMP_IN pixel_7171/SF_IB
+ pixel_7171/PIX_OUT pixel_7171/CSA_VREF pixel
Xpixel_7182 pixel_7182/gring pixel_7182/VDD pixel_7182/GND pixel_7182/VREF pixel_7182/ROW_SEL
+ pixel_7182/NB1 pixel_7182/VBIAS pixel_7182/NB2 pixel_7182/AMP_IN pixel_7182/SF_IB
+ pixel_7182/PIX_OUT pixel_7182/CSA_VREF pixel
Xpixel_7193 pixel_7193/gring pixel_7193/VDD pixel_7193/GND pixel_7193/VREF pixel_7193/ROW_SEL
+ pixel_7193/NB1 pixel_7193/VBIAS pixel_7193/NB2 pixel_7193/AMP_IN pixel_7193/SF_IB
+ pixel_7193/PIX_OUT pixel_7193/CSA_VREF pixel
Xpixel_6470 pixel_6470/gring pixel_6470/VDD pixel_6470/GND pixel_6470/VREF pixel_6470/ROW_SEL
+ pixel_6470/NB1 pixel_6470/VBIAS pixel_6470/NB2 pixel_6470/AMP_IN pixel_6470/SF_IB
+ pixel_6470/PIX_OUT pixel_6470/CSA_VREF pixel
Xpixel_6481 pixel_6481/gring pixel_6481/VDD pixel_6481/GND pixel_6481/VREF pixel_6481/ROW_SEL
+ pixel_6481/NB1 pixel_6481/VBIAS pixel_6481/NB2 pixel_6481/AMP_IN pixel_6481/SF_IB
+ pixel_6481/PIX_OUT pixel_6481/CSA_VREF pixel
Xpixel_6492 pixel_6492/gring pixel_6492/VDD pixel_6492/GND pixel_6492/VREF pixel_6492/ROW_SEL
+ pixel_6492/NB1 pixel_6492/VBIAS pixel_6492/NB2 pixel_6492/AMP_IN pixel_6492/SF_IB
+ pixel_6492/PIX_OUT pixel_6492/CSA_VREF pixel
Xpixel_5780 pixel_5780/gring pixel_5780/VDD pixel_5780/GND pixel_5780/VREF pixel_5780/ROW_SEL
+ pixel_5780/NB1 pixel_5780/VBIAS pixel_5780/NB2 pixel_5780/AMP_IN pixel_5780/SF_IB
+ pixel_5780/PIX_OUT pixel_5780/CSA_VREF pixel
Xpixel_5791 pixel_5791/gring pixel_5791/VDD pixel_5791/GND pixel_5791/VREF pixel_5791/ROW_SEL
+ pixel_5791/NB1 pixel_5791/VBIAS pixel_5791/NB2 pixel_5791/AMP_IN pixel_5791/SF_IB
+ pixel_5791/PIX_OUT pixel_5791/CSA_VREF pixel
Xpixel_3129 pixel_3129/gring pixel_3129/VDD pixel_3129/GND pixel_3129/VREF pixel_3129/ROW_SEL
+ pixel_3129/NB1 pixel_3129/VBIAS pixel_3129/NB2 pixel_3129/AMP_IN pixel_3129/SF_IB
+ pixel_3129/PIX_OUT pixel_3129/CSA_VREF pixel
Xpixel_3118 pixel_3118/gring pixel_3118/VDD pixel_3118/GND pixel_3118/VREF pixel_3118/ROW_SEL
+ pixel_3118/NB1 pixel_3118/VBIAS pixel_3118/NB2 pixel_3118/AMP_IN pixel_3118/SF_IB
+ pixel_3118/PIX_OUT pixel_3118/CSA_VREF pixel
Xpixel_3107 pixel_3107/gring pixel_3107/VDD pixel_3107/GND pixel_3107/VREF pixel_3107/ROW_SEL
+ pixel_3107/NB1 pixel_3107/VBIAS pixel_3107/NB2 pixel_3107/AMP_IN pixel_3107/SF_IB
+ pixel_3107/PIX_OUT pixel_3107/CSA_VREF pixel
Xpixel_2428 pixel_2428/gring pixel_2428/VDD pixel_2428/GND pixel_2428/VREF pixel_2428/ROW_SEL
+ pixel_2428/NB1 pixel_2428/VBIAS pixel_2428/NB2 pixel_2428/AMP_IN pixel_2428/SF_IB
+ pixel_2428/PIX_OUT pixel_2428/CSA_VREF pixel
Xpixel_2417 pixel_2417/gring pixel_2417/VDD pixel_2417/GND pixel_2417/VREF pixel_2417/ROW_SEL
+ pixel_2417/NB1 pixel_2417/VBIAS pixel_2417/NB2 pixel_2417/AMP_IN pixel_2417/SF_IB
+ pixel_2417/PIX_OUT pixel_2417/CSA_VREF pixel
Xpixel_2406 pixel_2406/gring pixel_2406/VDD pixel_2406/GND pixel_2406/VREF pixel_2406/ROW_SEL
+ pixel_2406/NB1 pixel_2406/VBIAS pixel_2406/NB2 pixel_2406/AMP_IN pixel_2406/SF_IB
+ pixel_2406/PIX_OUT pixel_2406/CSA_VREF pixel
Xpixel_1716 pixel_1716/gring pixel_1716/VDD pixel_1716/GND pixel_1716/VREF pixel_1716/ROW_SEL
+ pixel_1716/NB1 pixel_1716/VBIAS pixel_1716/NB2 pixel_1716/AMP_IN pixel_1716/SF_IB
+ pixel_1716/PIX_OUT pixel_1716/CSA_VREF pixel
Xpixel_1705 pixel_1705/gring pixel_1705/VDD pixel_1705/GND pixel_1705/VREF pixel_1705/ROW_SEL
+ pixel_1705/NB1 pixel_1705/VBIAS pixel_1705/NB2 pixel_1705/AMP_IN pixel_1705/SF_IB
+ pixel_1705/PIX_OUT pixel_1705/CSA_VREF pixel
Xpixel_2439 pixel_2439/gring pixel_2439/VDD pixel_2439/GND pixel_2439/VREF pixel_2439/ROW_SEL
+ pixel_2439/NB1 pixel_2439/VBIAS pixel_2439/NB2 pixel_2439/AMP_IN pixel_2439/SF_IB
+ pixel_2439/PIX_OUT pixel_2439/CSA_VREF pixel
Xpixel_1749 pixel_1749/gring pixel_1749/VDD pixel_1749/GND pixel_1749/VREF pixel_1749/ROW_SEL
+ pixel_1749/NB1 pixel_1749/VBIAS pixel_1749/NB2 pixel_1749/AMP_IN pixel_1749/SF_IB
+ pixel_1749/PIX_OUT pixel_1749/CSA_VREF pixel
Xpixel_1738 pixel_1738/gring pixel_1738/VDD pixel_1738/GND pixel_1738/VREF pixel_1738/ROW_SEL
+ pixel_1738/NB1 pixel_1738/VBIAS pixel_1738/NB2 pixel_1738/AMP_IN pixel_1738/SF_IB
+ pixel_1738/PIX_OUT pixel_1738/CSA_VREF pixel
Xpixel_1727 pixel_1727/gring pixel_1727/VDD pixel_1727/GND pixel_1727/VREF pixel_1727/ROW_SEL
+ pixel_1727/NB1 pixel_1727/VBIAS pixel_1727/NB2 pixel_1727/AMP_IN pixel_1727/SF_IB
+ pixel_1727/PIX_OUT pixel_1727/CSA_VREF pixel
Xpixel_5010 pixel_5010/gring pixel_5010/VDD pixel_5010/GND pixel_5010/VREF pixel_5010/ROW_SEL
+ pixel_5010/NB1 pixel_5010/VBIAS pixel_5010/NB2 pixel_5010/AMP_IN pixel_5010/SF_IB
+ pixel_5010/PIX_OUT pixel_5010/CSA_VREF pixel
Xpixel_5021 pixel_5021/gring pixel_5021/VDD pixel_5021/GND pixel_5021/VREF pixel_5021/ROW_SEL
+ pixel_5021/NB1 pixel_5021/VBIAS pixel_5021/NB2 pixel_5021/AMP_IN pixel_5021/SF_IB
+ pixel_5021/PIX_OUT pixel_5021/CSA_VREF pixel
Xpixel_5032 pixel_5032/gring pixel_5032/VDD pixel_5032/GND pixel_5032/VREF pixel_5032/ROW_SEL
+ pixel_5032/NB1 pixel_5032/VBIAS pixel_5032/NB2 pixel_5032/AMP_IN pixel_5032/SF_IB
+ pixel_5032/PIX_OUT pixel_5032/CSA_VREF pixel
Xpixel_5043 pixel_5043/gring pixel_5043/VDD pixel_5043/GND pixel_5043/VREF pixel_5043/ROW_SEL
+ pixel_5043/NB1 pixel_5043/VBIAS pixel_5043/NB2 pixel_5043/AMP_IN pixel_5043/SF_IB
+ pixel_5043/PIX_OUT pixel_5043/CSA_VREF pixel
Xpixel_5054 pixel_5054/gring pixel_5054/VDD pixel_5054/GND pixel_5054/VREF pixel_5054/ROW_SEL
+ pixel_5054/NB1 pixel_5054/VBIAS pixel_5054/NB2 pixel_5054/AMP_IN pixel_5054/SF_IB
+ pixel_5054/PIX_OUT pixel_5054/CSA_VREF pixel
Xpixel_5065 pixel_5065/gring pixel_5065/VDD pixel_5065/GND pixel_5065/VREF pixel_5065/ROW_SEL
+ pixel_5065/NB1 pixel_5065/VBIAS pixel_5065/NB2 pixel_5065/AMP_IN pixel_5065/SF_IB
+ pixel_5065/PIX_OUT pixel_5065/CSA_VREF pixel
Xpixel_4320 pixel_4320/gring pixel_4320/VDD pixel_4320/GND pixel_4320/VREF pixel_4320/ROW_SEL
+ pixel_4320/NB1 pixel_4320/VBIAS pixel_4320/NB2 pixel_4320/AMP_IN pixel_4320/SF_IB
+ pixel_4320/PIX_OUT pixel_4320/CSA_VREF pixel
Xpixel_5076 pixel_5076/gring pixel_5076/VDD pixel_5076/GND pixel_5076/VREF pixel_5076/ROW_SEL
+ pixel_5076/NB1 pixel_5076/VBIAS pixel_5076/NB2 pixel_5076/AMP_IN pixel_5076/SF_IB
+ pixel_5076/PIX_OUT pixel_5076/CSA_VREF pixel
Xpixel_5087 pixel_5087/gring pixel_5087/VDD pixel_5087/GND pixel_5087/VREF pixel_5087/ROW_SEL
+ pixel_5087/NB1 pixel_5087/VBIAS pixel_5087/NB2 pixel_5087/AMP_IN pixel_5087/SF_IB
+ pixel_5087/PIX_OUT pixel_5087/CSA_VREF pixel
Xpixel_5098 pixel_5098/gring pixel_5098/VDD pixel_5098/GND pixel_5098/VREF pixel_5098/ROW_SEL
+ pixel_5098/NB1 pixel_5098/VBIAS pixel_5098/NB2 pixel_5098/AMP_IN pixel_5098/SF_IB
+ pixel_5098/PIX_OUT pixel_5098/CSA_VREF pixel
Xpixel_4331 pixel_4331/gring pixel_4331/VDD pixel_4331/GND pixel_4331/VREF pixel_4331/ROW_SEL
+ pixel_4331/NB1 pixel_4331/VBIAS pixel_4331/NB2 pixel_4331/AMP_IN pixel_4331/SF_IB
+ pixel_4331/PIX_OUT pixel_4331/CSA_VREF pixel
Xpixel_4342 pixel_4342/gring pixel_4342/VDD pixel_4342/GND pixel_4342/VREF pixel_4342/ROW_SEL
+ pixel_4342/NB1 pixel_4342/VBIAS pixel_4342/NB2 pixel_4342/AMP_IN pixel_4342/SF_IB
+ pixel_4342/PIX_OUT pixel_4342/CSA_VREF pixel
Xpixel_4353 pixel_4353/gring pixel_4353/VDD pixel_4353/GND pixel_4353/VREF pixel_4353/ROW_SEL
+ pixel_4353/NB1 pixel_4353/VBIAS pixel_4353/NB2 pixel_4353/AMP_IN pixel_4353/SF_IB
+ pixel_4353/PIX_OUT pixel_4353/CSA_VREF pixel
Xpixel_392 pixel_392/gring pixel_392/VDD pixel_392/GND pixel_392/VREF pixel_392/ROW_SEL
+ pixel_392/NB1 pixel_392/VBIAS pixel_392/NB2 pixel_392/AMP_IN pixel_392/SF_IB pixel_392/PIX_OUT
+ pixel_392/CSA_VREF pixel
Xpixel_381 pixel_381/gring pixel_381/VDD pixel_381/GND pixel_381/VREF pixel_381/ROW_SEL
+ pixel_381/NB1 pixel_381/VBIAS pixel_381/NB2 pixel_381/AMP_IN pixel_381/SF_IB pixel_381/PIX_OUT
+ pixel_381/CSA_VREF pixel
Xpixel_370 pixel_370/gring pixel_370/VDD pixel_370/GND pixel_370/VREF pixel_370/ROW_SEL
+ pixel_370/NB1 pixel_370/VBIAS pixel_370/NB2 pixel_370/AMP_IN pixel_370/SF_IB pixel_370/PIX_OUT
+ pixel_370/CSA_VREF pixel
Xpixel_3652 pixel_3652/gring pixel_3652/VDD pixel_3652/GND pixel_3652/VREF pixel_3652/ROW_SEL
+ pixel_3652/NB1 pixel_3652/VBIAS pixel_3652/NB2 pixel_3652/AMP_IN pixel_3652/SF_IB
+ pixel_3652/PIX_OUT pixel_3652/CSA_VREF pixel
Xpixel_3641 pixel_3641/gring pixel_3641/VDD pixel_3641/GND pixel_3641/VREF pixel_3641/ROW_SEL
+ pixel_3641/NB1 pixel_3641/VBIAS pixel_3641/NB2 pixel_3641/AMP_IN pixel_3641/SF_IB
+ pixel_3641/PIX_OUT pixel_3641/CSA_VREF pixel
Xpixel_3630 pixel_3630/gring pixel_3630/VDD pixel_3630/GND pixel_3630/VREF pixel_3630/ROW_SEL
+ pixel_3630/NB1 pixel_3630/VBIAS pixel_3630/NB2 pixel_3630/AMP_IN pixel_3630/SF_IB
+ pixel_3630/PIX_OUT pixel_3630/CSA_VREF pixel
Xpixel_4364 pixel_4364/gring pixel_4364/VDD pixel_4364/GND pixel_4364/VREF pixel_4364/ROW_SEL
+ pixel_4364/NB1 pixel_4364/VBIAS pixel_4364/NB2 pixel_4364/AMP_IN pixel_4364/SF_IB
+ pixel_4364/PIX_OUT pixel_4364/CSA_VREF pixel
Xpixel_4375 pixel_4375/gring pixel_4375/VDD pixel_4375/GND pixel_4375/VREF pixel_4375/ROW_SEL
+ pixel_4375/NB1 pixel_4375/VBIAS pixel_4375/NB2 pixel_4375/AMP_IN pixel_4375/SF_IB
+ pixel_4375/PIX_OUT pixel_4375/CSA_VREF pixel
Xpixel_4386 pixel_4386/gring pixel_4386/VDD pixel_4386/GND pixel_4386/VREF pixel_4386/ROW_SEL
+ pixel_4386/NB1 pixel_4386/VBIAS pixel_4386/NB2 pixel_4386/AMP_IN pixel_4386/SF_IB
+ pixel_4386/PIX_OUT pixel_4386/CSA_VREF pixel
Xpixel_4397 pixel_4397/gring pixel_4397/VDD pixel_4397/GND pixel_4397/VREF pixel_4397/ROW_SEL
+ pixel_4397/NB1 pixel_4397/VBIAS pixel_4397/NB2 pixel_4397/AMP_IN pixel_4397/SF_IB
+ pixel_4397/PIX_OUT pixel_4397/CSA_VREF pixel
Xpixel_2940 pixel_2940/gring pixel_2940/VDD pixel_2940/GND pixel_2940/VREF pixel_2940/ROW_SEL
+ pixel_2940/NB1 pixel_2940/VBIAS pixel_2940/NB2 pixel_2940/AMP_IN pixel_2940/SF_IB
+ pixel_2940/PIX_OUT pixel_2940/CSA_VREF pixel
Xpixel_3685 pixel_3685/gring pixel_3685/VDD pixel_3685/GND pixel_3685/VREF pixel_3685/ROW_SEL
+ pixel_3685/NB1 pixel_3685/VBIAS pixel_3685/NB2 pixel_3685/AMP_IN pixel_3685/SF_IB
+ pixel_3685/PIX_OUT pixel_3685/CSA_VREF pixel
Xpixel_3674 pixel_3674/gring pixel_3674/VDD pixel_3674/GND pixel_3674/VREF pixel_3674/ROW_SEL
+ pixel_3674/NB1 pixel_3674/VBIAS pixel_3674/NB2 pixel_3674/AMP_IN pixel_3674/SF_IB
+ pixel_3674/PIX_OUT pixel_3674/CSA_VREF pixel
Xpixel_3663 pixel_3663/gring pixel_3663/VDD pixel_3663/GND pixel_3663/VREF pixel_3663/ROW_SEL
+ pixel_3663/NB1 pixel_3663/VBIAS pixel_3663/NB2 pixel_3663/AMP_IN pixel_3663/SF_IB
+ pixel_3663/PIX_OUT pixel_3663/CSA_VREF pixel
Xpixel_2973 pixel_2973/gring pixel_2973/VDD pixel_2973/GND pixel_2973/VREF pixel_2973/ROW_SEL
+ pixel_2973/NB1 pixel_2973/VBIAS pixel_2973/NB2 pixel_2973/AMP_IN pixel_2973/SF_IB
+ pixel_2973/PIX_OUT pixel_2973/CSA_VREF pixel
Xpixel_2962 pixel_2962/gring pixel_2962/VDD pixel_2962/GND pixel_2962/VREF pixel_2962/ROW_SEL
+ pixel_2962/NB1 pixel_2962/VBIAS pixel_2962/NB2 pixel_2962/AMP_IN pixel_2962/SF_IB
+ pixel_2962/PIX_OUT pixel_2962/CSA_VREF pixel
Xpixel_2951 pixel_2951/gring pixel_2951/VDD pixel_2951/GND pixel_2951/VREF pixel_2951/ROW_SEL
+ pixel_2951/NB1 pixel_2951/VBIAS pixel_2951/NB2 pixel_2951/AMP_IN pixel_2951/SF_IB
+ pixel_2951/PIX_OUT pixel_2951/CSA_VREF pixel
Xpixel_3696 pixel_3696/gring pixel_3696/VDD pixel_3696/GND pixel_3696/VREF pixel_3696/ROW_SEL
+ pixel_3696/NB1 pixel_3696/VBIAS pixel_3696/NB2 pixel_3696/AMP_IN pixel_3696/SF_IB
+ pixel_3696/PIX_OUT pixel_3696/CSA_VREF pixel
Xpixel_2995 pixel_2995/gring pixel_2995/VDD pixel_2995/GND pixel_2995/VREF pixel_2995/ROW_SEL
+ pixel_2995/NB1 pixel_2995/VBIAS pixel_2995/NB2 pixel_2995/AMP_IN pixel_2995/SF_IB
+ pixel_2995/PIX_OUT pixel_2995/CSA_VREF pixel
Xpixel_2984 pixel_2984/gring pixel_2984/VDD pixel_2984/GND pixel_2984/VREF pixel_2984/ROW_SEL
+ pixel_2984/NB1 pixel_2984/VBIAS pixel_2984/NB2 pixel_2984/AMP_IN pixel_2984/SF_IB
+ pixel_2984/PIX_OUT pixel_2984/CSA_VREF pixel
Xpixel_9309 pixel_9309/gring pixel_9309/VDD pixel_9309/GND pixel_9309/VREF pixel_9309/ROW_SEL
+ pixel_9309/NB1 pixel_9309/VBIAS pixel_9309/NB2 pixel_9309/AMP_IN pixel_9309/SF_IB
+ pixel_9309/PIX_OUT pixel_9309/CSA_VREF pixel
Xpixel_8608 pixel_8608/gring pixel_8608/VDD pixel_8608/GND pixel_8608/VREF pixel_8608/ROW_SEL
+ pixel_8608/NB1 pixel_8608/VBIAS pixel_8608/NB2 pixel_8608/AMP_IN pixel_8608/SF_IB
+ pixel_8608/PIX_OUT pixel_8608/CSA_VREF pixel
Xpixel_8619 pixel_8619/gring pixel_8619/VDD pixel_8619/GND pixel_8619/VREF pixel_8619/ROW_SEL
+ pixel_8619/NB1 pixel_8619/VBIAS pixel_8619/NB2 pixel_8619/AMP_IN pixel_8619/SF_IB
+ pixel_8619/PIX_OUT pixel_8619/CSA_VREF pixel
Xpixel_7907 pixel_7907/gring pixel_7907/VDD pixel_7907/GND pixel_7907/VREF pixel_7907/ROW_SEL
+ pixel_7907/NB1 pixel_7907/VBIAS pixel_7907/NB2 pixel_7907/AMP_IN pixel_7907/SF_IB
+ pixel_7907/PIX_OUT pixel_7907/CSA_VREF pixel
Xpixel_7918 pixel_7918/gring pixel_7918/VDD pixel_7918/GND pixel_7918/VREF pixel_7918/ROW_SEL
+ pixel_7918/NB1 pixel_7918/VBIAS pixel_7918/NB2 pixel_7918/AMP_IN pixel_7918/SF_IB
+ pixel_7918/PIX_OUT pixel_7918/CSA_VREF pixel
Xpixel_7929 pixel_7929/gring pixel_7929/VDD pixel_7929/GND pixel_7929/VREF pixel_7929/ROW_SEL
+ pixel_7929/NB1 pixel_7929/VBIAS pixel_7929/NB2 pixel_7929/AMP_IN pixel_7929/SF_IB
+ pixel_7929/PIX_OUT pixel_7929/CSA_VREF pixel
Xpixel_2203 pixel_2203/gring pixel_2203/VDD pixel_2203/GND pixel_2203/VREF pixel_2203/ROW_SEL
+ pixel_2203/NB1 pixel_2203/VBIAS pixel_2203/NB2 pixel_2203/AMP_IN pixel_2203/SF_IB
+ pixel_2203/PIX_OUT pixel_2203/CSA_VREF pixel
Xpixel_2236 pixel_2236/gring pixel_2236/VDD pixel_2236/GND pixel_2236/VREF pixel_2236/ROW_SEL
+ pixel_2236/NB1 pixel_2236/VBIAS pixel_2236/NB2 pixel_2236/AMP_IN pixel_2236/SF_IB
+ pixel_2236/PIX_OUT pixel_2236/CSA_VREF pixel
Xpixel_2225 pixel_2225/gring pixel_2225/VDD pixel_2225/GND pixel_2225/VREF pixel_2225/ROW_SEL
+ pixel_2225/NB1 pixel_2225/VBIAS pixel_2225/NB2 pixel_2225/AMP_IN pixel_2225/SF_IB
+ pixel_2225/PIX_OUT pixel_2225/CSA_VREF pixel
Xpixel_2214 pixel_2214/gring pixel_2214/VDD pixel_2214/GND pixel_2214/VREF pixel_2214/ROW_SEL
+ pixel_2214/NB1 pixel_2214/VBIAS pixel_2214/NB2 pixel_2214/AMP_IN pixel_2214/SF_IB
+ pixel_2214/PIX_OUT pixel_2214/CSA_VREF pixel
Xpixel_1524 pixel_1524/gring pixel_1524/VDD pixel_1524/GND pixel_1524/VREF pixel_1524/ROW_SEL
+ pixel_1524/NB1 pixel_1524/VBIAS pixel_1524/NB2 pixel_1524/AMP_IN pixel_1524/SF_IB
+ pixel_1524/PIX_OUT pixel_1524/CSA_VREF pixel
Xpixel_1513 pixel_1513/gring pixel_1513/VDD pixel_1513/GND pixel_1513/VREF pixel_1513/ROW_SEL
+ pixel_1513/NB1 pixel_1513/VBIAS pixel_1513/NB2 pixel_1513/AMP_IN pixel_1513/SF_IB
+ pixel_1513/PIX_OUT pixel_1513/CSA_VREF pixel
Xpixel_1502 pixel_1502/gring pixel_1502/VDD pixel_1502/GND pixel_1502/VREF pixel_1502/ROW_SEL
+ pixel_1502/NB1 pixel_1502/VBIAS pixel_1502/NB2 pixel_1502/AMP_IN pixel_1502/SF_IB
+ pixel_1502/PIX_OUT pixel_1502/CSA_VREF pixel
Xpixel_2269 pixel_2269/gring pixel_2269/VDD pixel_2269/GND pixel_2269/VREF pixel_2269/ROW_SEL
+ pixel_2269/NB1 pixel_2269/VBIAS pixel_2269/NB2 pixel_2269/AMP_IN pixel_2269/SF_IB
+ pixel_2269/PIX_OUT pixel_2269/CSA_VREF pixel
Xpixel_2258 pixel_2258/gring pixel_2258/VDD pixel_2258/GND pixel_2258/VREF pixel_2258/ROW_SEL
+ pixel_2258/NB1 pixel_2258/VBIAS pixel_2258/NB2 pixel_2258/AMP_IN pixel_2258/SF_IB
+ pixel_2258/PIX_OUT pixel_2258/CSA_VREF pixel
Xpixel_2247 pixel_2247/gring pixel_2247/VDD pixel_2247/GND pixel_2247/VREF pixel_2247/ROW_SEL
+ pixel_2247/NB1 pixel_2247/VBIAS pixel_2247/NB2 pixel_2247/AMP_IN pixel_2247/SF_IB
+ pixel_2247/PIX_OUT pixel_2247/CSA_VREF pixel
Xpixel_1568 pixel_1568/gring pixel_1568/VDD pixel_1568/GND pixel_1568/VREF pixel_1568/ROW_SEL
+ pixel_1568/NB1 pixel_1568/VBIAS pixel_1568/NB2 pixel_1568/AMP_IN pixel_1568/SF_IB
+ pixel_1568/PIX_OUT pixel_1568/CSA_VREF pixel
Xpixel_1557 pixel_1557/gring pixel_1557/VDD pixel_1557/GND pixel_1557/VREF pixel_1557/ROW_SEL
+ pixel_1557/NB1 pixel_1557/VBIAS pixel_1557/NB2 pixel_1557/AMP_IN pixel_1557/SF_IB
+ pixel_1557/PIX_OUT pixel_1557/CSA_VREF pixel
Xpixel_1546 pixel_1546/gring pixel_1546/VDD pixel_1546/GND pixel_1546/VREF pixel_1546/ROW_SEL
+ pixel_1546/NB1 pixel_1546/VBIAS pixel_1546/NB2 pixel_1546/AMP_IN pixel_1546/SF_IB
+ pixel_1546/PIX_OUT pixel_1546/CSA_VREF pixel
Xpixel_1535 pixel_1535/gring pixel_1535/VDD pixel_1535/GND pixel_1535/VREF pixel_1535/ROW_SEL
+ pixel_1535/NB1 pixel_1535/VBIAS pixel_1535/NB2 pixel_1535/AMP_IN pixel_1535/SF_IB
+ pixel_1535/PIX_OUT pixel_1535/CSA_VREF pixel
Xpixel_1579 pixel_1579/gring pixel_1579/VDD pixel_1579/GND pixel_1579/VREF pixel_1579/ROW_SEL
+ pixel_1579/NB1 pixel_1579/VBIAS pixel_1579/NB2 pixel_1579/AMP_IN pixel_1579/SF_IB
+ pixel_1579/PIX_OUT pixel_1579/CSA_VREF pixel
Xpixel_9832 pixel_9832/gring pixel_9832/VDD pixel_9832/GND pixel_9832/VREF pixel_9832/ROW_SEL
+ pixel_9832/NB1 pixel_9832/VBIAS pixel_9832/NB2 pixel_9832/AMP_IN pixel_9832/SF_IB
+ pixel_9832/PIX_OUT pixel_9832/CSA_VREF pixel
Xpixel_9821 pixel_9821/gring pixel_9821/VDD pixel_9821/GND pixel_9821/VREF pixel_9821/ROW_SEL
+ pixel_9821/NB1 pixel_9821/VBIAS pixel_9821/NB2 pixel_9821/AMP_IN pixel_9821/SF_IB
+ pixel_9821/PIX_OUT pixel_9821/CSA_VREF pixel
Xpixel_9810 pixel_9810/gring pixel_9810/VDD pixel_9810/GND pixel_9810/VREF pixel_9810/ROW_SEL
+ pixel_9810/NB1 pixel_9810/VBIAS pixel_9810/NB2 pixel_9810/AMP_IN pixel_9810/SF_IB
+ pixel_9810/PIX_OUT pixel_9810/CSA_VREF pixel
Xpixel_9843 pixel_9843/gring pixel_9843/VDD pixel_9843/GND pixel_9843/VREF pixel_9843/ROW_SEL
+ pixel_9843/NB1 pixel_9843/VBIAS pixel_9843/NB2 pixel_9843/AMP_IN pixel_9843/SF_IB
+ pixel_9843/PIX_OUT pixel_9843/CSA_VREF pixel
Xpixel_9854 pixel_9854/gring pixel_9854/VDD pixel_9854/GND pixel_9854/VREF pixel_9854/ROW_SEL
+ pixel_9854/NB1 pixel_9854/VBIAS pixel_9854/NB2 pixel_9854/AMP_IN pixel_9854/SF_IB
+ pixel_9854/PIX_OUT pixel_9854/CSA_VREF pixel
Xpixel_9865 pixel_9865/gring pixel_9865/VDD pixel_9865/GND pixel_9865/VREF pixel_9865/ROW_SEL
+ pixel_9865/NB1 pixel_9865/VBIAS pixel_9865/NB2 pixel_9865/AMP_IN pixel_9865/SF_IB
+ pixel_9865/PIX_OUT pixel_9865/CSA_VREF pixel
Xpixel_9876 pixel_9876/gring pixel_9876/VDD pixel_9876/GND pixel_9876/VREF pixel_9876/ROW_SEL
+ pixel_9876/NB1 pixel_9876/VBIAS pixel_9876/NB2 pixel_9876/AMP_IN pixel_9876/SF_IB
+ pixel_9876/PIX_OUT pixel_9876/CSA_VREF pixel
Xpixel_9887 pixel_9887/gring pixel_9887/VDD pixel_9887/GND pixel_9887/VREF pixel_9887/ROW_SEL
+ pixel_9887/NB1 pixel_9887/VBIAS pixel_9887/NB2 pixel_9887/AMP_IN pixel_9887/SF_IB
+ pixel_9887/PIX_OUT pixel_9887/CSA_VREF pixel
Xpixel_9898 pixel_9898/gring pixel_9898/VDD pixel_9898/GND pixel_9898/VREF pixel_9898/ROW_SEL
+ pixel_9898/NB1 pixel_9898/VBIAS pixel_9898/NB2 pixel_9898/AMP_IN pixel_9898/SF_IB
+ pixel_9898/PIX_OUT pixel_9898/CSA_VREF pixel
Xpixel_4150 pixel_4150/gring pixel_4150/VDD pixel_4150/GND pixel_4150/VREF pixel_4150/ROW_SEL
+ pixel_4150/NB1 pixel_4150/VBIAS pixel_4150/NB2 pixel_4150/AMP_IN pixel_4150/SF_IB
+ pixel_4150/PIX_OUT pixel_4150/CSA_VREF pixel
Xpixel_4161 pixel_4161/gring pixel_4161/VDD pixel_4161/GND pixel_4161/VREF pixel_4161/ROW_SEL
+ pixel_4161/NB1 pixel_4161/VBIAS pixel_4161/NB2 pixel_4161/AMP_IN pixel_4161/SF_IB
+ pixel_4161/PIX_OUT pixel_4161/CSA_VREF pixel
Xpixel_3460 pixel_3460/gring pixel_3460/VDD pixel_3460/GND pixel_3460/VREF pixel_3460/ROW_SEL
+ pixel_3460/NB1 pixel_3460/VBIAS pixel_3460/NB2 pixel_3460/AMP_IN pixel_3460/SF_IB
+ pixel_3460/PIX_OUT pixel_3460/CSA_VREF pixel
Xpixel_4172 pixel_4172/gring pixel_4172/VDD pixel_4172/GND pixel_4172/VREF pixel_4172/ROW_SEL
+ pixel_4172/NB1 pixel_4172/VBIAS pixel_4172/NB2 pixel_4172/AMP_IN pixel_4172/SF_IB
+ pixel_4172/PIX_OUT pixel_4172/CSA_VREF pixel
Xpixel_4183 pixel_4183/gring pixel_4183/VDD pixel_4183/GND pixel_4183/VREF pixel_4183/ROW_SEL
+ pixel_4183/NB1 pixel_4183/VBIAS pixel_4183/NB2 pixel_4183/AMP_IN pixel_4183/SF_IB
+ pixel_4183/PIX_OUT pixel_4183/CSA_VREF pixel
Xpixel_4194 pixel_4194/gring pixel_4194/VDD pixel_4194/GND pixel_4194/VREF pixel_4194/ROW_SEL
+ pixel_4194/NB1 pixel_4194/VBIAS pixel_4194/NB2 pixel_4194/AMP_IN pixel_4194/SF_IB
+ pixel_4194/PIX_OUT pixel_4194/CSA_VREF pixel
Xpixel_3493 pixel_3493/gring pixel_3493/VDD pixel_3493/GND pixel_3493/VREF pixel_3493/ROW_SEL
+ pixel_3493/NB1 pixel_3493/VBIAS pixel_3493/NB2 pixel_3493/AMP_IN pixel_3493/SF_IB
+ pixel_3493/PIX_OUT pixel_3493/CSA_VREF pixel
Xpixel_3482 pixel_3482/gring pixel_3482/VDD pixel_3482/GND pixel_3482/VREF pixel_3482/ROW_SEL
+ pixel_3482/NB1 pixel_3482/VBIAS pixel_3482/NB2 pixel_3482/AMP_IN pixel_3482/SF_IB
+ pixel_3482/PIX_OUT pixel_3482/CSA_VREF pixel
Xpixel_3471 pixel_3471/gring pixel_3471/VDD pixel_3471/GND pixel_3471/VREF pixel_3471/ROW_SEL
+ pixel_3471/NB1 pixel_3471/VBIAS pixel_3471/NB2 pixel_3471/AMP_IN pixel_3471/SF_IB
+ pixel_3471/PIX_OUT pixel_3471/CSA_VREF pixel
Xpixel_2792 pixel_2792/gring pixel_2792/VDD pixel_2792/GND pixel_2792/VREF pixel_2792/ROW_SEL
+ pixel_2792/NB1 pixel_2792/VBIAS pixel_2792/NB2 pixel_2792/AMP_IN pixel_2792/SF_IB
+ pixel_2792/PIX_OUT pixel_2792/CSA_VREF pixel
Xpixel_2781 pixel_2781/gring pixel_2781/VDD pixel_2781/GND pixel_2781/VREF pixel_2781/ROW_SEL
+ pixel_2781/NB1 pixel_2781/VBIAS pixel_2781/NB2 pixel_2781/AMP_IN pixel_2781/SF_IB
+ pixel_2781/PIX_OUT pixel_2781/CSA_VREF pixel
Xpixel_2770 pixel_2770/gring pixel_2770/VDD pixel_2770/GND pixel_2770/VREF pixel_2770/ROW_SEL
+ pixel_2770/NB1 pixel_2770/VBIAS pixel_2770/NB2 pixel_2770/AMP_IN pixel_2770/SF_IB
+ pixel_2770/PIX_OUT pixel_2770/CSA_VREF pixel
Xpixel_9128 pixel_9128/gring pixel_9128/VDD pixel_9128/GND pixel_9128/VREF pixel_9128/ROW_SEL
+ pixel_9128/NB1 pixel_9128/VBIAS pixel_9128/NB2 pixel_9128/AMP_IN pixel_9128/SF_IB
+ pixel_9128/PIX_OUT pixel_9128/CSA_VREF pixel
Xpixel_9117 pixel_9117/gring pixel_9117/VDD pixel_9117/GND pixel_9117/VREF pixel_9117/ROW_SEL
+ pixel_9117/NB1 pixel_9117/VBIAS pixel_9117/NB2 pixel_9117/AMP_IN pixel_9117/SF_IB
+ pixel_9117/PIX_OUT pixel_9117/CSA_VREF pixel
Xpixel_9106 pixel_9106/gring pixel_9106/VDD pixel_9106/GND pixel_9106/VREF pixel_9106/ROW_SEL
+ pixel_9106/NB1 pixel_9106/VBIAS pixel_9106/NB2 pixel_9106/AMP_IN pixel_9106/SF_IB
+ pixel_9106/PIX_OUT pixel_9106/CSA_VREF pixel
Xpixel_8416 pixel_8416/gring pixel_8416/VDD pixel_8416/GND pixel_8416/VREF pixel_8416/ROW_SEL
+ pixel_8416/NB1 pixel_8416/VBIAS pixel_8416/NB2 pixel_8416/AMP_IN pixel_8416/SF_IB
+ pixel_8416/PIX_OUT pixel_8416/CSA_VREF pixel
Xpixel_8405 pixel_8405/gring pixel_8405/VDD pixel_8405/GND pixel_8405/VREF pixel_8405/ROW_SEL
+ pixel_8405/NB1 pixel_8405/VBIAS pixel_8405/NB2 pixel_8405/AMP_IN pixel_8405/SF_IB
+ pixel_8405/PIX_OUT pixel_8405/CSA_VREF pixel
Xpixel_9139 pixel_9139/gring pixel_9139/VDD pixel_9139/GND pixel_9139/VREF pixel_9139/ROW_SEL
+ pixel_9139/NB1 pixel_9139/VBIAS pixel_9139/NB2 pixel_9139/AMP_IN pixel_9139/SF_IB
+ pixel_9139/PIX_OUT pixel_9139/CSA_VREF pixel
Xpixel_8427 pixel_8427/gring pixel_8427/VDD pixel_8427/GND pixel_8427/VREF pixel_8427/ROW_SEL
+ pixel_8427/NB1 pixel_8427/VBIAS pixel_8427/NB2 pixel_8427/AMP_IN pixel_8427/SF_IB
+ pixel_8427/PIX_OUT pixel_8427/CSA_VREF pixel
Xpixel_8438 pixel_8438/gring pixel_8438/VDD pixel_8438/GND pixel_8438/VREF pixel_8438/ROW_SEL
+ pixel_8438/NB1 pixel_8438/VBIAS pixel_8438/NB2 pixel_8438/AMP_IN pixel_8438/SF_IB
+ pixel_8438/PIX_OUT pixel_8438/CSA_VREF pixel
Xpixel_8449 pixel_8449/gring pixel_8449/VDD pixel_8449/GND pixel_8449/VREF pixel_8449/ROW_SEL
+ pixel_8449/NB1 pixel_8449/VBIAS pixel_8449/NB2 pixel_8449/AMP_IN pixel_8449/SF_IB
+ pixel_8449/PIX_OUT pixel_8449/CSA_VREF pixel
Xpixel_7704 pixel_7704/gring pixel_7704/VDD pixel_7704/GND pixel_7704/VREF pixel_7704/ROW_SEL
+ pixel_7704/NB1 pixel_7704/VBIAS pixel_7704/NB2 pixel_7704/AMP_IN pixel_7704/SF_IB
+ pixel_7704/PIX_OUT pixel_7704/CSA_VREF pixel
Xpixel_7715 pixel_7715/gring pixel_7715/VDD pixel_7715/GND pixel_7715/VREF pixel_7715/ROW_SEL
+ pixel_7715/NB1 pixel_7715/VBIAS pixel_7715/NB2 pixel_7715/AMP_IN pixel_7715/SF_IB
+ pixel_7715/PIX_OUT pixel_7715/CSA_VREF pixel
Xpixel_7726 pixel_7726/gring pixel_7726/VDD pixel_7726/GND pixel_7726/VREF pixel_7726/ROW_SEL
+ pixel_7726/NB1 pixel_7726/VBIAS pixel_7726/NB2 pixel_7726/AMP_IN pixel_7726/SF_IB
+ pixel_7726/PIX_OUT pixel_7726/CSA_VREF pixel
Xpixel_7737 pixel_7737/gring pixel_7737/VDD pixel_7737/GND pixel_7737/VREF pixel_7737/ROW_SEL
+ pixel_7737/NB1 pixel_7737/VBIAS pixel_7737/NB2 pixel_7737/AMP_IN pixel_7737/SF_IB
+ pixel_7737/PIX_OUT pixel_7737/CSA_VREF pixel
Xpixel_7748 pixel_7748/gring pixel_7748/VDD pixel_7748/GND pixel_7748/VREF pixel_7748/ROW_SEL
+ pixel_7748/NB1 pixel_7748/VBIAS pixel_7748/NB2 pixel_7748/AMP_IN pixel_7748/SF_IB
+ pixel_7748/PIX_OUT pixel_7748/CSA_VREF pixel
Xpixel_7759 pixel_7759/gring pixel_7759/VDD pixel_7759/GND pixel_7759/VREF pixel_7759/ROW_SEL
+ pixel_7759/NB1 pixel_7759/VBIAS pixel_7759/NB2 pixel_7759/AMP_IN pixel_7759/SF_IB
+ pixel_7759/PIX_OUT pixel_7759/CSA_VREF pixel
Xpixel_2011 pixel_2011/gring pixel_2011/VDD pixel_2011/GND pixel_2011/VREF pixel_2011/ROW_SEL
+ pixel_2011/NB1 pixel_2011/VBIAS pixel_2011/NB2 pixel_2011/AMP_IN pixel_2011/SF_IB
+ pixel_2011/PIX_OUT pixel_2011/CSA_VREF pixel
Xpixel_2000 pixel_2000/gring pixel_2000/VDD pixel_2000/GND pixel_2000/VREF pixel_2000/ROW_SEL
+ pixel_2000/NB1 pixel_2000/VBIAS pixel_2000/NB2 pixel_2000/AMP_IN pixel_2000/SF_IB
+ pixel_2000/PIX_OUT pixel_2000/CSA_VREF pixel
Xpixel_2044 pixel_2044/gring pixel_2044/VDD pixel_2044/GND pixel_2044/VREF pixel_2044/ROW_SEL
+ pixel_2044/NB1 pixel_2044/VBIAS pixel_2044/NB2 pixel_2044/AMP_IN pixel_2044/SF_IB
+ pixel_2044/PIX_OUT pixel_2044/CSA_VREF pixel
Xpixel_2033 pixel_2033/gring pixel_2033/VDD pixel_2033/GND pixel_2033/VREF pixel_2033/ROW_SEL
+ pixel_2033/NB1 pixel_2033/VBIAS pixel_2033/NB2 pixel_2033/AMP_IN pixel_2033/SF_IB
+ pixel_2033/PIX_OUT pixel_2033/CSA_VREF pixel
Xpixel_2022 pixel_2022/gring pixel_2022/VDD pixel_2022/GND pixel_2022/VREF pixel_2022/ROW_SEL
+ pixel_2022/NB1 pixel_2022/VBIAS pixel_2022/NB2 pixel_2022/AMP_IN pixel_2022/SF_IB
+ pixel_2022/PIX_OUT pixel_2022/CSA_VREF pixel
Xpixel_1332 pixel_1332/gring pixel_1332/VDD pixel_1332/GND pixel_1332/VREF pixel_1332/ROW_SEL
+ pixel_1332/NB1 pixel_1332/VBIAS pixel_1332/NB2 pixel_1332/AMP_IN pixel_1332/SF_IB
+ pixel_1332/PIX_OUT pixel_1332/CSA_VREF pixel
Xpixel_1321 pixel_1321/gring pixel_1321/VDD pixel_1321/GND pixel_1321/VREF pixel_1321/ROW_SEL
+ pixel_1321/NB1 pixel_1321/VBIAS pixel_1321/NB2 pixel_1321/AMP_IN pixel_1321/SF_IB
+ pixel_1321/PIX_OUT pixel_1321/CSA_VREF pixel
Xpixel_1310 pixel_1310/gring pixel_1310/VDD pixel_1310/GND pixel_1310/VREF pixel_1310/ROW_SEL
+ pixel_1310/NB1 pixel_1310/VBIAS pixel_1310/NB2 pixel_1310/AMP_IN pixel_1310/SF_IB
+ pixel_1310/PIX_OUT pixel_1310/CSA_VREF pixel
Xpixel_2077 pixel_2077/gring pixel_2077/VDD pixel_2077/GND pixel_2077/VREF pixel_2077/ROW_SEL
+ pixel_2077/NB1 pixel_2077/VBIAS pixel_2077/NB2 pixel_2077/AMP_IN pixel_2077/SF_IB
+ pixel_2077/PIX_OUT pixel_2077/CSA_VREF pixel
Xpixel_2066 pixel_2066/gring pixel_2066/VDD pixel_2066/GND pixel_2066/VREF pixel_2066/ROW_SEL
+ pixel_2066/NB1 pixel_2066/VBIAS pixel_2066/NB2 pixel_2066/AMP_IN pixel_2066/SF_IB
+ pixel_2066/PIX_OUT pixel_2066/CSA_VREF pixel
Xpixel_2055 pixel_2055/gring pixel_2055/VDD pixel_2055/GND pixel_2055/VREF pixel_2055/ROW_SEL
+ pixel_2055/NB1 pixel_2055/VBIAS pixel_2055/NB2 pixel_2055/AMP_IN pixel_2055/SF_IB
+ pixel_2055/PIX_OUT pixel_2055/CSA_VREF pixel
Xpixel_1376 pixel_1376/gring pixel_1376/VDD pixel_1376/GND pixel_1376/VREF pixel_1376/ROW_SEL
+ pixel_1376/NB1 pixel_1376/VBIAS pixel_1376/NB2 pixel_1376/AMP_IN pixel_1376/SF_IB
+ pixel_1376/PIX_OUT pixel_1376/CSA_VREF pixel
Xpixel_1365 pixel_1365/gring pixel_1365/VDD pixel_1365/GND pixel_1365/VREF pixel_1365/ROW_SEL
+ pixel_1365/NB1 pixel_1365/VBIAS pixel_1365/NB2 pixel_1365/AMP_IN pixel_1365/SF_IB
+ pixel_1365/PIX_OUT pixel_1365/CSA_VREF pixel
Xpixel_1354 pixel_1354/gring pixel_1354/VDD pixel_1354/GND pixel_1354/VREF pixel_1354/ROW_SEL
+ pixel_1354/NB1 pixel_1354/VBIAS pixel_1354/NB2 pixel_1354/AMP_IN pixel_1354/SF_IB
+ pixel_1354/PIX_OUT pixel_1354/CSA_VREF pixel
Xpixel_1343 pixel_1343/gring pixel_1343/VDD pixel_1343/GND pixel_1343/VREF pixel_1343/ROW_SEL
+ pixel_1343/NB1 pixel_1343/VBIAS pixel_1343/NB2 pixel_1343/AMP_IN pixel_1343/SF_IB
+ pixel_1343/PIX_OUT pixel_1343/CSA_VREF pixel
Xpixel_2099 pixel_2099/gring pixel_2099/VDD pixel_2099/GND pixel_2099/VREF pixel_2099/ROW_SEL
+ pixel_2099/NB1 pixel_2099/VBIAS pixel_2099/NB2 pixel_2099/AMP_IN pixel_2099/SF_IB
+ pixel_2099/PIX_OUT pixel_2099/CSA_VREF pixel
Xpixel_2088 pixel_2088/gring pixel_2088/VDD pixel_2088/GND pixel_2088/VREF pixel_2088/ROW_SEL
+ pixel_2088/NB1 pixel_2088/VBIAS pixel_2088/NB2 pixel_2088/AMP_IN pixel_2088/SF_IB
+ pixel_2088/PIX_OUT pixel_2088/CSA_VREF pixel
Xpixel_1398 pixel_1398/gring pixel_1398/VDD pixel_1398/GND pixel_1398/VREF pixel_1398/ROW_SEL
+ pixel_1398/NB1 pixel_1398/VBIAS pixel_1398/NB2 pixel_1398/AMP_IN pixel_1398/SF_IB
+ pixel_1398/PIX_OUT pixel_1398/CSA_VREF pixel
Xpixel_1387 pixel_1387/gring pixel_1387/VDD pixel_1387/GND pixel_1387/VREF pixel_1387/ROW_SEL
+ pixel_1387/NB1 pixel_1387/VBIAS pixel_1387/NB2 pixel_1387/AMP_IN pixel_1387/SF_IB
+ pixel_1387/PIX_OUT pixel_1387/CSA_VREF pixel
Xpixel_9640 pixel_9640/gring pixel_9640/VDD pixel_9640/GND pixel_9640/VREF pixel_9640/ROW_SEL
+ pixel_9640/NB1 pixel_9640/VBIAS pixel_9640/NB2 pixel_9640/AMP_IN pixel_9640/SF_IB
+ pixel_9640/PIX_OUT pixel_9640/CSA_VREF pixel
Xpixel_9684 pixel_9684/gring pixel_9684/VDD pixel_9684/GND pixel_9684/VREF pixel_9684/ROW_SEL
+ pixel_9684/NB1 pixel_9684/VBIAS pixel_9684/NB2 pixel_9684/AMP_IN pixel_9684/SF_IB
+ pixel_9684/PIX_OUT pixel_9684/CSA_VREF pixel
Xpixel_9651 pixel_9651/gring pixel_9651/VDD pixel_9651/GND pixel_9651/VREF pixel_9651/ROW_SEL
+ pixel_9651/NB1 pixel_9651/VBIAS pixel_9651/NB2 pixel_9651/AMP_IN pixel_9651/SF_IB
+ pixel_9651/PIX_OUT pixel_9651/CSA_VREF pixel
Xpixel_9662 pixel_9662/gring pixel_9662/VDD pixel_9662/GND pixel_9662/VREF pixel_9662/ROW_SEL
+ pixel_9662/NB1 pixel_9662/VBIAS pixel_9662/NB2 pixel_9662/AMP_IN pixel_9662/SF_IB
+ pixel_9662/PIX_OUT pixel_9662/CSA_VREF pixel
Xpixel_9673 pixel_9673/gring pixel_9673/VDD pixel_9673/GND pixel_9673/VREF pixel_9673/ROW_SEL
+ pixel_9673/NB1 pixel_9673/VBIAS pixel_9673/NB2 pixel_9673/AMP_IN pixel_9673/SF_IB
+ pixel_9673/PIX_OUT pixel_9673/CSA_VREF pixel
Xpixel_8972 pixel_8972/gring pixel_8972/VDD pixel_8972/GND pixel_8972/VREF pixel_8972/ROW_SEL
+ pixel_8972/NB1 pixel_8972/VBIAS pixel_8972/NB2 pixel_8972/AMP_IN pixel_8972/SF_IB
+ pixel_8972/PIX_OUT pixel_8972/CSA_VREF pixel
Xpixel_8961 pixel_8961/gring pixel_8961/VDD pixel_8961/GND pixel_8961/VREF pixel_8961/ROW_SEL
+ pixel_8961/NB1 pixel_8961/VBIAS pixel_8961/NB2 pixel_8961/AMP_IN pixel_8961/SF_IB
+ pixel_8961/PIX_OUT pixel_8961/CSA_VREF pixel
Xpixel_8950 pixel_8950/gring pixel_8950/VDD pixel_8950/GND pixel_8950/VREF pixel_8950/ROW_SEL
+ pixel_8950/NB1 pixel_8950/VBIAS pixel_8950/NB2 pixel_8950/AMP_IN pixel_8950/SF_IB
+ pixel_8950/PIX_OUT pixel_8950/CSA_VREF pixel
Xpixel_9695 pixel_9695/gring pixel_9695/VDD pixel_9695/GND pixel_9695/VREF pixel_9695/ROW_SEL
+ pixel_9695/NB1 pixel_9695/VBIAS pixel_9695/NB2 pixel_9695/AMP_IN pixel_9695/SF_IB
+ pixel_9695/PIX_OUT pixel_9695/CSA_VREF pixel
Xpixel_8994 pixel_8994/gring pixel_8994/VDD pixel_8994/GND pixel_8994/VREF pixel_8994/ROW_SEL
+ pixel_8994/NB1 pixel_8994/VBIAS pixel_8994/NB2 pixel_8994/AMP_IN pixel_8994/SF_IB
+ pixel_8994/PIX_OUT pixel_8994/CSA_VREF pixel
Xpixel_8983 pixel_8983/gring pixel_8983/VDD pixel_8983/GND pixel_8983/VREF pixel_8983/ROW_SEL
+ pixel_8983/NB1 pixel_8983/VBIAS pixel_8983/NB2 pixel_8983/AMP_IN pixel_8983/SF_IB
+ pixel_8983/PIX_OUT pixel_8983/CSA_VREF pixel
Xpixel_3290 pixel_3290/gring pixel_3290/VDD pixel_3290/GND pixel_3290/VREF pixel_3290/ROW_SEL
+ pixel_3290/NB1 pixel_3290/VBIAS pixel_3290/NB2 pixel_3290/AMP_IN pixel_3290/SF_IB
+ pixel_3290/PIX_OUT pixel_3290/CSA_VREF pixel
Xpixel_5609 pixel_5609/gring pixel_5609/VDD pixel_5609/GND pixel_5609/VREF pixel_5609/ROW_SEL
+ pixel_5609/NB1 pixel_5609/VBIAS pixel_5609/NB2 pixel_5609/AMP_IN pixel_5609/SF_IB
+ pixel_5609/PIX_OUT pixel_5609/CSA_VREF pixel
Xpixel_914 pixel_914/gring pixel_914/VDD pixel_914/GND pixel_914/VREF pixel_914/ROW_SEL
+ pixel_914/NB1 pixel_914/VBIAS pixel_914/NB2 pixel_914/AMP_IN pixel_914/SF_IB pixel_914/PIX_OUT
+ pixel_914/CSA_VREF pixel
Xpixel_903 pixel_903/gring pixel_903/VDD pixel_903/GND pixel_903/VREF pixel_903/ROW_SEL
+ pixel_903/NB1 pixel_903/VBIAS pixel_903/NB2 pixel_903/AMP_IN pixel_903/SF_IB pixel_903/PIX_OUT
+ pixel_903/CSA_VREF pixel
Xpixel_4908 pixel_4908/gring pixel_4908/VDD pixel_4908/GND pixel_4908/VREF pixel_4908/ROW_SEL
+ pixel_4908/NB1 pixel_4908/VBIAS pixel_4908/NB2 pixel_4908/AMP_IN pixel_4908/SF_IB
+ pixel_4908/PIX_OUT pixel_4908/CSA_VREF pixel
Xpixel_4919 pixel_4919/gring pixel_4919/VDD pixel_4919/GND pixel_4919/VREF pixel_4919/ROW_SEL
+ pixel_4919/NB1 pixel_4919/VBIAS pixel_4919/NB2 pixel_4919/AMP_IN pixel_4919/SF_IB
+ pixel_4919/PIX_OUT pixel_4919/CSA_VREF pixel
Xpixel_958 pixel_958/gring pixel_958/VDD pixel_958/GND pixel_958/VREF pixel_958/ROW_SEL
+ pixel_958/NB1 pixel_958/VBIAS pixel_958/NB2 pixel_958/AMP_IN pixel_958/SF_IB pixel_958/PIX_OUT
+ pixel_958/CSA_VREF pixel
Xpixel_947 pixel_947/gring pixel_947/VDD pixel_947/GND pixel_947/VREF pixel_947/ROW_SEL
+ pixel_947/NB1 pixel_947/VBIAS pixel_947/NB2 pixel_947/AMP_IN pixel_947/SF_IB pixel_947/PIX_OUT
+ pixel_947/CSA_VREF pixel
Xpixel_936 pixel_936/gring pixel_936/VDD pixel_936/GND pixel_936/VREF pixel_936/ROW_SEL
+ pixel_936/NB1 pixel_936/VBIAS pixel_936/NB2 pixel_936/AMP_IN pixel_936/SF_IB pixel_936/PIX_OUT
+ pixel_936/CSA_VREF pixel
Xpixel_925 pixel_925/gring pixel_925/VDD pixel_925/GND pixel_925/VREF pixel_925/ROW_SEL
+ pixel_925/NB1 pixel_925/VBIAS pixel_925/NB2 pixel_925/AMP_IN pixel_925/SF_IB pixel_925/PIX_OUT
+ pixel_925/CSA_VREF pixel
Xpixel_969 pixel_969/gring pixel_969/VDD pixel_969/GND pixel_969/VREF pixel_969/ROW_SEL
+ pixel_969/NB1 pixel_969/VBIAS pixel_969/NB2 pixel_969/AMP_IN pixel_969/SF_IB pixel_969/PIX_OUT
+ pixel_969/CSA_VREF pixel
Xpixel_8202 pixel_8202/gring pixel_8202/VDD pixel_8202/GND pixel_8202/VREF pixel_8202/ROW_SEL
+ pixel_8202/NB1 pixel_8202/VBIAS pixel_8202/NB2 pixel_8202/AMP_IN pixel_8202/SF_IB
+ pixel_8202/PIX_OUT pixel_8202/CSA_VREF pixel
Xpixel_8213 pixel_8213/gring pixel_8213/VDD pixel_8213/GND pixel_8213/VREF pixel_8213/ROW_SEL
+ pixel_8213/NB1 pixel_8213/VBIAS pixel_8213/NB2 pixel_8213/AMP_IN pixel_8213/SF_IB
+ pixel_8213/PIX_OUT pixel_8213/CSA_VREF pixel
Xpixel_8224 pixel_8224/gring pixel_8224/VDD pixel_8224/GND pixel_8224/VREF pixel_8224/ROW_SEL
+ pixel_8224/NB1 pixel_8224/VBIAS pixel_8224/NB2 pixel_8224/AMP_IN pixel_8224/SF_IB
+ pixel_8224/PIX_OUT pixel_8224/CSA_VREF pixel
Xpixel_8235 pixel_8235/gring pixel_8235/VDD pixel_8235/GND pixel_8235/VREF pixel_8235/ROW_SEL
+ pixel_8235/NB1 pixel_8235/VBIAS pixel_8235/NB2 pixel_8235/AMP_IN pixel_8235/SF_IB
+ pixel_8235/PIX_OUT pixel_8235/CSA_VREF pixel
Xpixel_8246 pixel_8246/gring pixel_8246/VDD pixel_8246/GND pixel_8246/VREF pixel_8246/ROW_SEL
+ pixel_8246/NB1 pixel_8246/VBIAS pixel_8246/NB2 pixel_8246/AMP_IN pixel_8246/SF_IB
+ pixel_8246/PIX_OUT pixel_8246/CSA_VREF pixel
Xpixel_8257 pixel_8257/gring pixel_8257/VDD pixel_8257/GND pixel_8257/VREF pixel_8257/ROW_SEL
+ pixel_8257/NB1 pixel_8257/VBIAS pixel_8257/NB2 pixel_8257/AMP_IN pixel_8257/SF_IB
+ pixel_8257/PIX_OUT pixel_8257/CSA_VREF pixel
Xpixel_8268 pixel_8268/gring pixel_8268/VDD pixel_8268/GND pixel_8268/VREF pixel_8268/ROW_SEL
+ pixel_8268/NB1 pixel_8268/VBIAS pixel_8268/NB2 pixel_8268/AMP_IN pixel_8268/SF_IB
+ pixel_8268/PIX_OUT pixel_8268/CSA_VREF pixel
Xpixel_7501 pixel_7501/gring pixel_7501/VDD pixel_7501/GND pixel_7501/VREF pixel_7501/ROW_SEL
+ pixel_7501/NB1 pixel_7501/VBIAS pixel_7501/NB2 pixel_7501/AMP_IN pixel_7501/SF_IB
+ pixel_7501/PIX_OUT pixel_7501/CSA_VREF pixel
Xpixel_7512 pixel_7512/gring pixel_7512/VDD pixel_7512/GND pixel_7512/VREF pixel_7512/ROW_SEL
+ pixel_7512/NB1 pixel_7512/VBIAS pixel_7512/NB2 pixel_7512/AMP_IN pixel_7512/SF_IB
+ pixel_7512/PIX_OUT pixel_7512/CSA_VREF pixel
Xpixel_7523 pixel_7523/gring pixel_7523/VDD pixel_7523/GND pixel_7523/VREF pixel_7523/ROW_SEL
+ pixel_7523/NB1 pixel_7523/VBIAS pixel_7523/NB2 pixel_7523/AMP_IN pixel_7523/SF_IB
+ pixel_7523/PIX_OUT pixel_7523/CSA_VREF pixel
Xpixel_8279 pixel_8279/gring pixel_8279/VDD pixel_8279/GND pixel_8279/VREF pixel_8279/ROW_SEL
+ pixel_8279/NB1 pixel_8279/VBIAS pixel_8279/NB2 pixel_8279/AMP_IN pixel_8279/SF_IB
+ pixel_8279/PIX_OUT pixel_8279/CSA_VREF pixel
Xpixel_7534 pixel_7534/gring pixel_7534/VDD pixel_7534/GND pixel_7534/VREF pixel_7534/ROW_SEL
+ pixel_7534/NB1 pixel_7534/VBIAS pixel_7534/NB2 pixel_7534/AMP_IN pixel_7534/SF_IB
+ pixel_7534/PIX_OUT pixel_7534/CSA_VREF pixel
Xpixel_7545 pixel_7545/gring pixel_7545/VDD pixel_7545/GND pixel_7545/VREF pixel_7545/ROW_SEL
+ pixel_7545/NB1 pixel_7545/VBIAS pixel_7545/NB2 pixel_7545/AMP_IN pixel_7545/SF_IB
+ pixel_7545/PIX_OUT pixel_7545/CSA_VREF pixel
Xpixel_7556 pixel_7556/gring pixel_7556/VDD pixel_7556/GND pixel_7556/VREF pixel_7556/ROW_SEL
+ pixel_7556/NB1 pixel_7556/VBIAS pixel_7556/NB2 pixel_7556/AMP_IN pixel_7556/SF_IB
+ pixel_7556/PIX_OUT pixel_7556/CSA_VREF pixel
Xpixel_6800 pixel_6800/gring pixel_6800/VDD pixel_6800/GND pixel_6800/VREF pixel_6800/ROW_SEL
+ pixel_6800/NB1 pixel_6800/VBIAS pixel_6800/NB2 pixel_6800/AMP_IN pixel_6800/SF_IB
+ pixel_6800/PIX_OUT pixel_6800/CSA_VREF pixel
Xpixel_6811 pixel_6811/gring pixel_6811/VDD pixel_6811/GND pixel_6811/VREF pixel_6811/ROW_SEL
+ pixel_6811/NB1 pixel_6811/VBIAS pixel_6811/NB2 pixel_6811/AMP_IN pixel_6811/SF_IB
+ pixel_6811/PIX_OUT pixel_6811/CSA_VREF pixel
Xpixel_7567 pixel_7567/gring pixel_7567/VDD pixel_7567/GND pixel_7567/VREF pixel_7567/ROW_SEL
+ pixel_7567/NB1 pixel_7567/VBIAS pixel_7567/NB2 pixel_7567/AMP_IN pixel_7567/SF_IB
+ pixel_7567/PIX_OUT pixel_7567/CSA_VREF pixel
Xpixel_7578 pixel_7578/gring pixel_7578/VDD pixel_7578/GND pixel_7578/VREF pixel_7578/ROW_SEL
+ pixel_7578/NB1 pixel_7578/VBIAS pixel_7578/NB2 pixel_7578/AMP_IN pixel_7578/SF_IB
+ pixel_7578/PIX_OUT pixel_7578/CSA_VREF pixel
Xpixel_7589 pixel_7589/gring pixel_7589/VDD pixel_7589/GND pixel_7589/VREF pixel_7589/ROW_SEL
+ pixel_7589/NB1 pixel_7589/VBIAS pixel_7589/NB2 pixel_7589/AMP_IN pixel_7589/SF_IB
+ pixel_7589/PIX_OUT pixel_7589/CSA_VREF pixel
Xpixel_6822 pixel_6822/gring pixel_6822/VDD pixel_6822/GND pixel_6822/VREF pixel_6822/ROW_SEL
+ pixel_6822/NB1 pixel_6822/VBIAS pixel_6822/NB2 pixel_6822/AMP_IN pixel_6822/SF_IB
+ pixel_6822/PIX_OUT pixel_6822/CSA_VREF pixel
Xpixel_6833 pixel_6833/gring pixel_6833/VDD pixel_6833/GND pixel_6833/VREF pixel_6833/ROW_SEL
+ pixel_6833/NB1 pixel_6833/VBIAS pixel_6833/NB2 pixel_6833/AMP_IN pixel_6833/SF_IB
+ pixel_6833/PIX_OUT pixel_6833/CSA_VREF pixel
Xpixel_6844 pixel_6844/gring pixel_6844/VDD pixel_6844/GND pixel_6844/VREF pixel_6844/ROW_SEL
+ pixel_6844/NB1 pixel_6844/VBIAS pixel_6844/NB2 pixel_6844/AMP_IN pixel_6844/SF_IB
+ pixel_6844/PIX_OUT pixel_6844/CSA_VREF pixel
Xpixel_6855 pixel_6855/gring pixel_6855/VDD pixel_6855/GND pixel_6855/VREF pixel_6855/ROW_SEL
+ pixel_6855/NB1 pixel_6855/VBIAS pixel_6855/NB2 pixel_6855/AMP_IN pixel_6855/SF_IB
+ pixel_6855/PIX_OUT pixel_6855/CSA_VREF pixel
Xpixel_6866 pixel_6866/gring pixel_6866/VDD pixel_6866/GND pixel_6866/VREF pixel_6866/ROW_SEL
+ pixel_6866/NB1 pixel_6866/VBIAS pixel_6866/NB2 pixel_6866/AMP_IN pixel_6866/SF_IB
+ pixel_6866/PIX_OUT pixel_6866/CSA_VREF pixel
Xpixel_6877 pixel_6877/gring pixel_6877/VDD pixel_6877/GND pixel_6877/VREF pixel_6877/ROW_SEL
+ pixel_6877/NB1 pixel_6877/VBIAS pixel_6877/NB2 pixel_6877/AMP_IN pixel_6877/SF_IB
+ pixel_6877/PIX_OUT pixel_6877/CSA_VREF pixel
Xpixel_6888 pixel_6888/gring pixel_6888/VDD pixel_6888/GND pixel_6888/VREF pixel_6888/ROW_SEL
+ pixel_6888/NB1 pixel_6888/VBIAS pixel_6888/NB2 pixel_6888/AMP_IN pixel_6888/SF_IB
+ pixel_6888/PIX_OUT pixel_6888/CSA_VREF pixel
Xpixel_6899 pixel_6899/gring pixel_6899/VDD pixel_6899/GND pixel_6899/VREF pixel_6899/ROW_SEL
+ pixel_6899/NB1 pixel_6899/VBIAS pixel_6899/NB2 pixel_6899/AMP_IN pixel_6899/SF_IB
+ pixel_6899/PIX_OUT pixel_6899/CSA_VREF pixel
Xpixel_1151 pixel_1151/gring pixel_1151/VDD pixel_1151/GND pixel_1151/VREF pixel_1151/ROW_SEL
+ pixel_1151/NB1 pixel_1151/VBIAS pixel_1151/NB2 pixel_1151/AMP_IN pixel_1151/SF_IB
+ pixel_1151/PIX_OUT pixel_1151/CSA_VREF pixel
Xpixel_1140 pixel_1140/gring pixel_1140/VDD pixel_1140/GND pixel_1140/VREF pixel_1140/ROW_SEL
+ pixel_1140/NB1 pixel_1140/VBIAS pixel_1140/NB2 pixel_1140/AMP_IN pixel_1140/SF_IB
+ pixel_1140/PIX_OUT pixel_1140/CSA_VREF pixel
Xpixel_1184 pixel_1184/gring pixel_1184/VDD pixel_1184/GND pixel_1184/VREF pixel_1184/ROW_SEL
+ pixel_1184/NB1 pixel_1184/VBIAS pixel_1184/NB2 pixel_1184/AMP_IN pixel_1184/SF_IB
+ pixel_1184/PIX_OUT pixel_1184/CSA_VREF pixel
Xpixel_1173 pixel_1173/gring pixel_1173/VDD pixel_1173/GND pixel_1173/VREF pixel_1173/ROW_SEL
+ pixel_1173/NB1 pixel_1173/VBIAS pixel_1173/NB2 pixel_1173/AMP_IN pixel_1173/SF_IB
+ pixel_1173/PIX_OUT pixel_1173/CSA_VREF pixel
Xpixel_1162 pixel_1162/gring pixel_1162/VDD pixel_1162/GND pixel_1162/VREF pixel_1162/ROW_SEL
+ pixel_1162/NB1 pixel_1162/VBIAS pixel_1162/NB2 pixel_1162/AMP_IN pixel_1162/SF_IB
+ pixel_1162/PIX_OUT pixel_1162/CSA_VREF pixel
Xpixel_1195 pixel_1195/gring pixel_1195/VDD pixel_1195/GND pixel_1195/VREF pixel_1195/ROW_SEL
+ pixel_1195/NB1 pixel_1195/VBIAS pixel_1195/NB2 pixel_1195/AMP_IN pixel_1195/SF_IB
+ pixel_1195/PIX_OUT pixel_1195/CSA_VREF pixel
Xpixel_9492 pixel_9492/gring pixel_9492/VDD pixel_9492/GND pixel_9492/VREF pixel_9492/ROW_SEL
+ pixel_9492/NB1 pixel_9492/VBIAS pixel_9492/NB2 pixel_9492/AMP_IN pixel_9492/SF_IB
+ pixel_9492/PIX_OUT pixel_9492/CSA_VREF pixel
Xpixel_9481 pixel_9481/gring pixel_9481/VDD pixel_9481/GND pixel_9481/VREF pixel_9481/ROW_SEL
+ pixel_9481/NB1 pixel_9481/VBIAS pixel_9481/NB2 pixel_9481/AMP_IN pixel_9481/SF_IB
+ pixel_9481/PIX_OUT pixel_9481/CSA_VREF pixel
Xpixel_9470 pixel_9470/gring pixel_9470/VDD pixel_9470/GND pixel_9470/VREF pixel_9470/ROW_SEL
+ pixel_9470/NB1 pixel_9470/VBIAS pixel_9470/NB2 pixel_9470/AMP_IN pixel_9470/SF_IB
+ pixel_9470/PIX_OUT pixel_9470/CSA_VREF pixel
Xpixel_8780 pixel_8780/gring pixel_8780/VDD pixel_8780/GND pixel_8780/VREF pixel_8780/ROW_SEL
+ pixel_8780/NB1 pixel_8780/VBIAS pixel_8780/NB2 pixel_8780/AMP_IN pixel_8780/SF_IB
+ pixel_8780/PIX_OUT pixel_8780/CSA_VREF pixel
Xpixel_8791 pixel_8791/gring pixel_8791/VDD pixel_8791/GND pixel_8791/VREF pixel_8791/ROW_SEL
+ pixel_8791/NB1 pixel_8791/VBIAS pixel_8791/NB2 pixel_8791/AMP_IN pixel_8791/SF_IB
+ pixel_8791/PIX_OUT pixel_8791/CSA_VREF pixel
Xpixel_6107 pixel_6107/gring pixel_6107/VDD pixel_6107/GND pixel_6107/VREF pixel_6107/ROW_SEL
+ pixel_6107/NB1 pixel_6107/VBIAS pixel_6107/NB2 pixel_6107/AMP_IN pixel_6107/SF_IB
+ pixel_6107/PIX_OUT pixel_6107/CSA_VREF pixel
Xpixel_6118 pixel_6118/gring pixel_6118/VDD pixel_6118/GND pixel_6118/VREF pixel_6118/ROW_SEL
+ pixel_6118/NB1 pixel_6118/VBIAS pixel_6118/NB2 pixel_6118/AMP_IN pixel_6118/SF_IB
+ pixel_6118/PIX_OUT pixel_6118/CSA_VREF pixel
Xpixel_6129 pixel_6129/gring pixel_6129/VDD pixel_6129/GND pixel_6129/VREF pixel_6129/ROW_SEL
+ pixel_6129/NB1 pixel_6129/VBIAS pixel_6129/NB2 pixel_6129/AMP_IN pixel_6129/SF_IB
+ pixel_6129/PIX_OUT pixel_6129/CSA_VREF pixel
Xpixel_5406 pixel_5406/gring pixel_5406/VDD pixel_5406/GND pixel_5406/VREF pixel_5406/ROW_SEL
+ pixel_5406/NB1 pixel_5406/VBIAS pixel_5406/NB2 pixel_5406/AMP_IN pixel_5406/SF_IB
+ pixel_5406/PIX_OUT pixel_5406/CSA_VREF pixel
Xpixel_5417 pixel_5417/gring pixel_5417/VDD pixel_5417/GND pixel_5417/VREF pixel_5417/ROW_SEL
+ pixel_5417/NB1 pixel_5417/VBIAS pixel_5417/NB2 pixel_5417/AMP_IN pixel_5417/SF_IB
+ pixel_5417/PIX_OUT pixel_5417/CSA_VREF pixel
Xpixel_5428 pixel_5428/gring pixel_5428/VDD pixel_5428/GND pixel_5428/VREF pixel_5428/ROW_SEL
+ pixel_5428/NB1 pixel_5428/VBIAS pixel_5428/NB2 pixel_5428/AMP_IN pixel_5428/SF_IB
+ pixel_5428/PIX_OUT pixel_5428/CSA_VREF pixel
Xpixel_5439 pixel_5439/gring pixel_5439/VDD pixel_5439/GND pixel_5439/VREF pixel_5439/ROW_SEL
+ pixel_5439/NB1 pixel_5439/VBIAS pixel_5439/NB2 pixel_5439/AMP_IN pixel_5439/SF_IB
+ pixel_5439/PIX_OUT pixel_5439/CSA_VREF pixel
Xpixel_733 pixel_733/gring pixel_733/VDD pixel_733/GND pixel_733/VREF pixel_733/ROW_SEL
+ pixel_733/NB1 pixel_733/VBIAS pixel_733/NB2 pixel_733/AMP_IN pixel_733/SF_IB pixel_733/PIX_OUT
+ pixel_733/CSA_VREF pixel
Xpixel_722 pixel_722/gring pixel_722/VDD pixel_722/GND pixel_722/VREF pixel_722/ROW_SEL
+ pixel_722/NB1 pixel_722/VBIAS pixel_722/NB2 pixel_722/AMP_IN pixel_722/SF_IB pixel_722/PIX_OUT
+ pixel_722/CSA_VREF pixel
Xpixel_711 pixel_711/gring pixel_711/VDD pixel_711/GND pixel_711/VREF pixel_711/ROW_SEL
+ pixel_711/NB1 pixel_711/VBIAS pixel_711/NB2 pixel_711/AMP_IN pixel_711/SF_IB pixel_711/PIX_OUT
+ pixel_711/CSA_VREF pixel
Xpixel_700 pixel_700/gring pixel_700/VDD pixel_700/GND pixel_700/VREF pixel_700/ROW_SEL
+ pixel_700/NB1 pixel_700/VBIAS pixel_700/NB2 pixel_700/AMP_IN pixel_700/SF_IB pixel_700/PIX_OUT
+ pixel_700/CSA_VREF pixel
Xpixel_4705 pixel_4705/gring pixel_4705/VDD pixel_4705/GND pixel_4705/VREF pixel_4705/ROW_SEL
+ pixel_4705/NB1 pixel_4705/VBIAS pixel_4705/NB2 pixel_4705/AMP_IN pixel_4705/SF_IB
+ pixel_4705/PIX_OUT pixel_4705/CSA_VREF pixel
Xpixel_4716 pixel_4716/gring pixel_4716/VDD pixel_4716/GND pixel_4716/VREF pixel_4716/ROW_SEL
+ pixel_4716/NB1 pixel_4716/VBIAS pixel_4716/NB2 pixel_4716/AMP_IN pixel_4716/SF_IB
+ pixel_4716/PIX_OUT pixel_4716/CSA_VREF pixel
Xpixel_4727 pixel_4727/gring pixel_4727/VDD pixel_4727/GND pixel_4727/VREF pixel_4727/ROW_SEL
+ pixel_4727/NB1 pixel_4727/VBIAS pixel_4727/NB2 pixel_4727/AMP_IN pixel_4727/SF_IB
+ pixel_4727/PIX_OUT pixel_4727/CSA_VREF pixel
Xpixel_766 pixel_766/gring pixel_766/VDD pixel_766/GND pixel_766/VREF pixel_766/ROW_SEL
+ pixel_766/NB1 pixel_766/VBIAS pixel_766/NB2 pixel_766/AMP_IN pixel_766/SF_IB pixel_766/PIX_OUT
+ pixel_766/CSA_VREF pixel
Xpixel_755 pixel_755/gring pixel_755/VDD pixel_755/GND pixel_755/VREF pixel_755/ROW_SEL
+ pixel_755/NB1 pixel_755/VBIAS pixel_755/NB2 pixel_755/AMP_IN pixel_755/SF_IB pixel_755/PIX_OUT
+ pixel_755/CSA_VREF pixel
Xpixel_744 pixel_744/gring pixel_744/VDD pixel_744/GND pixel_744/VREF pixel_744/ROW_SEL
+ pixel_744/NB1 pixel_744/VBIAS pixel_744/NB2 pixel_744/AMP_IN pixel_744/SF_IB pixel_744/PIX_OUT
+ pixel_744/CSA_VREF pixel
Xpixel_4738 pixel_4738/gring pixel_4738/VDD pixel_4738/GND pixel_4738/VREF pixel_4738/ROW_SEL
+ pixel_4738/NB1 pixel_4738/VBIAS pixel_4738/NB2 pixel_4738/AMP_IN pixel_4738/SF_IB
+ pixel_4738/PIX_OUT pixel_4738/CSA_VREF pixel
Xpixel_4749 pixel_4749/gring pixel_4749/VDD pixel_4749/GND pixel_4749/VREF pixel_4749/ROW_SEL
+ pixel_4749/NB1 pixel_4749/VBIAS pixel_4749/NB2 pixel_4749/AMP_IN pixel_4749/SF_IB
+ pixel_4749/PIX_OUT pixel_4749/CSA_VREF pixel
Xpixel_799 pixel_799/gring pixel_799/VDD pixel_799/GND pixel_799/VREF pixel_799/ROW_SEL
+ pixel_799/NB1 pixel_799/VBIAS pixel_799/NB2 pixel_799/AMP_IN pixel_799/SF_IB pixel_799/PIX_OUT
+ pixel_799/CSA_VREF pixel
Xpixel_788 pixel_788/gring pixel_788/VDD pixel_788/GND pixel_788/VREF pixel_788/ROW_SEL
+ pixel_788/NB1 pixel_788/VBIAS pixel_788/NB2 pixel_788/AMP_IN pixel_788/SF_IB pixel_788/PIX_OUT
+ pixel_788/CSA_VREF pixel
Xpixel_777 pixel_777/gring pixel_777/VDD pixel_777/GND pixel_777/VREF pixel_777/ROW_SEL
+ pixel_777/NB1 pixel_777/VBIAS pixel_777/NB2 pixel_777/AMP_IN pixel_777/SF_IB pixel_777/PIX_OUT
+ pixel_777/CSA_VREF pixel
Xpixel_8010 pixel_8010/gring pixel_8010/VDD pixel_8010/GND pixel_8010/VREF pixel_8010/ROW_SEL
+ pixel_8010/NB1 pixel_8010/VBIAS pixel_8010/NB2 pixel_8010/AMP_IN pixel_8010/SF_IB
+ pixel_8010/PIX_OUT pixel_8010/CSA_VREF pixel
Xpixel_8021 pixel_8021/gring pixel_8021/VDD pixel_8021/GND pixel_8021/VREF pixel_8021/ROW_SEL
+ pixel_8021/NB1 pixel_8021/VBIAS pixel_8021/NB2 pixel_8021/AMP_IN pixel_8021/SF_IB
+ pixel_8021/PIX_OUT pixel_8021/CSA_VREF pixel
Xpixel_8032 pixel_8032/gring pixel_8032/VDD pixel_8032/GND pixel_8032/VREF pixel_8032/ROW_SEL
+ pixel_8032/NB1 pixel_8032/VBIAS pixel_8032/NB2 pixel_8032/AMP_IN pixel_8032/SF_IB
+ pixel_8032/PIX_OUT pixel_8032/CSA_VREF pixel
Xpixel_8043 pixel_8043/gring pixel_8043/VDD pixel_8043/GND pixel_8043/VREF pixel_8043/ROW_SEL
+ pixel_8043/NB1 pixel_8043/VBIAS pixel_8043/NB2 pixel_8043/AMP_IN pixel_8043/SF_IB
+ pixel_8043/PIX_OUT pixel_8043/CSA_VREF pixel
Xpixel_8054 pixel_8054/gring pixel_8054/VDD pixel_8054/GND pixel_8054/VREF pixel_8054/ROW_SEL
+ pixel_8054/NB1 pixel_8054/VBIAS pixel_8054/NB2 pixel_8054/AMP_IN pixel_8054/SF_IB
+ pixel_8054/PIX_OUT pixel_8054/CSA_VREF pixel
Xpixel_8065 pixel_8065/gring pixel_8065/VDD pixel_8065/GND pixel_8065/VREF pixel_8065/ROW_SEL
+ pixel_8065/NB1 pixel_8065/VBIAS pixel_8065/NB2 pixel_8065/AMP_IN pixel_8065/SF_IB
+ pixel_8065/PIX_OUT pixel_8065/CSA_VREF pixel
Xpixel_8076 pixel_8076/gring pixel_8076/VDD pixel_8076/GND pixel_8076/VREF pixel_8076/ROW_SEL
+ pixel_8076/NB1 pixel_8076/VBIAS pixel_8076/NB2 pixel_8076/AMP_IN pixel_8076/SF_IB
+ pixel_8076/PIX_OUT pixel_8076/CSA_VREF pixel
Xpixel_7320 pixel_7320/gring pixel_7320/VDD pixel_7320/GND pixel_7320/VREF pixel_7320/ROW_SEL
+ pixel_7320/NB1 pixel_7320/VBIAS pixel_7320/NB2 pixel_7320/AMP_IN pixel_7320/SF_IB
+ pixel_7320/PIX_OUT pixel_7320/CSA_VREF pixel
Xpixel_7331 pixel_7331/gring pixel_7331/VDD pixel_7331/GND pixel_7331/VREF pixel_7331/ROW_SEL
+ pixel_7331/NB1 pixel_7331/VBIAS pixel_7331/NB2 pixel_7331/AMP_IN pixel_7331/SF_IB
+ pixel_7331/PIX_OUT pixel_7331/CSA_VREF pixel
Xpixel_8087 pixel_8087/gring pixel_8087/VDD pixel_8087/GND pixel_8087/VREF pixel_8087/ROW_SEL
+ pixel_8087/NB1 pixel_8087/VBIAS pixel_8087/NB2 pixel_8087/AMP_IN pixel_8087/SF_IB
+ pixel_8087/PIX_OUT pixel_8087/CSA_VREF pixel
Xpixel_8098 pixel_8098/gring pixel_8098/VDD pixel_8098/GND pixel_8098/VREF pixel_8098/ROW_SEL
+ pixel_8098/NB1 pixel_8098/VBIAS pixel_8098/NB2 pixel_8098/AMP_IN pixel_8098/SF_IB
+ pixel_8098/PIX_OUT pixel_8098/CSA_VREF pixel
Xpixel_7342 pixel_7342/gring pixel_7342/VDD pixel_7342/GND pixel_7342/VREF pixel_7342/ROW_SEL
+ pixel_7342/NB1 pixel_7342/VBIAS pixel_7342/NB2 pixel_7342/AMP_IN pixel_7342/SF_IB
+ pixel_7342/PIX_OUT pixel_7342/CSA_VREF pixel
Xpixel_7353 pixel_7353/gring pixel_7353/VDD pixel_7353/GND pixel_7353/VREF pixel_7353/ROW_SEL
+ pixel_7353/NB1 pixel_7353/VBIAS pixel_7353/NB2 pixel_7353/AMP_IN pixel_7353/SF_IB
+ pixel_7353/PIX_OUT pixel_7353/CSA_VREF pixel
Xpixel_7364 pixel_7364/gring pixel_7364/VDD pixel_7364/GND pixel_7364/VREF pixel_7364/ROW_SEL
+ pixel_7364/NB1 pixel_7364/VBIAS pixel_7364/NB2 pixel_7364/AMP_IN pixel_7364/SF_IB
+ pixel_7364/PIX_OUT pixel_7364/CSA_VREF pixel
Xpixel_7375 pixel_7375/gring pixel_7375/VDD pixel_7375/GND pixel_7375/VREF pixel_7375/ROW_SEL
+ pixel_7375/NB1 pixel_7375/VBIAS pixel_7375/NB2 pixel_7375/AMP_IN pixel_7375/SF_IB
+ pixel_7375/PIX_OUT pixel_7375/CSA_VREF pixel
Xpixel_6630 pixel_6630/gring pixel_6630/VDD pixel_6630/GND pixel_6630/VREF pixel_6630/ROW_SEL
+ pixel_6630/NB1 pixel_6630/VBIAS pixel_6630/NB2 pixel_6630/AMP_IN pixel_6630/SF_IB
+ pixel_6630/PIX_OUT pixel_6630/CSA_VREF pixel
Xpixel_7386 pixel_7386/gring pixel_7386/VDD pixel_7386/GND pixel_7386/VREF pixel_7386/ROW_SEL
+ pixel_7386/NB1 pixel_7386/VBIAS pixel_7386/NB2 pixel_7386/AMP_IN pixel_7386/SF_IB
+ pixel_7386/PIX_OUT pixel_7386/CSA_VREF pixel
Xpixel_7397 pixel_7397/gring pixel_7397/VDD pixel_7397/GND pixel_7397/VREF pixel_7397/ROW_SEL
+ pixel_7397/NB1 pixel_7397/VBIAS pixel_7397/NB2 pixel_7397/AMP_IN pixel_7397/SF_IB
+ pixel_7397/PIX_OUT pixel_7397/CSA_VREF pixel
Xpixel_6641 pixel_6641/gring pixel_6641/VDD pixel_6641/GND pixel_6641/VREF pixel_6641/ROW_SEL
+ pixel_6641/NB1 pixel_6641/VBIAS pixel_6641/NB2 pixel_6641/AMP_IN pixel_6641/SF_IB
+ pixel_6641/PIX_OUT pixel_6641/CSA_VREF pixel
Xpixel_6652 pixel_6652/gring pixel_6652/VDD pixel_6652/GND pixel_6652/VREF pixel_6652/ROW_SEL
+ pixel_6652/NB1 pixel_6652/VBIAS pixel_6652/NB2 pixel_6652/AMP_IN pixel_6652/SF_IB
+ pixel_6652/PIX_OUT pixel_6652/CSA_VREF pixel
Xpixel_6663 pixel_6663/gring pixel_6663/VDD pixel_6663/GND pixel_6663/VREF pixel_6663/ROW_SEL
+ pixel_6663/NB1 pixel_6663/VBIAS pixel_6663/NB2 pixel_6663/AMP_IN pixel_6663/SF_IB
+ pixel_6663/PIX_OUT pixel_6663/CSA_VREF pixel
Xpixel_6674 pixel_6674/gring pixel_6674/VDD pixel_6674/GND pixel_6674/VREF pixel_6674/ROW_SEL
+ pixel_6674/NB1 pixel_6674/VBIAS pixel_6674/NB2 pixel_6674/AMP_IN pixel_6674/SF_IB
+ pixel_6674/PIX_OUT pixel_6674/CSA_VREF pixel
Xpixel_6685 pixel_6685/gring pixel_6685/VDD pixel_6685/GND pixel_6685/VREF pixel_6685/ROW_SEL
+ pixel_6685/NB1 pixel_6685/VBIAS pixel_6685/NB2 pixel_6685/AMP_IN pixel_6685/SF_IB
+ pixel_6685/PIX_OUT pixel_6685/CSA_VREF pixel
Xpixel_6696 pixel_6696/gring pixel_6696/VDD pixel_6696/GND pixel_6696/VREF pixel_6696/ROW_SEL
+ pixel_6696/NB1 pixel_6696/VBIAS pixel_6696/NB2 pixel_6696/AMP_IN pixel_6696/SF_IB
+ pixel_6696/PIX_OUT pixel_6696/CSA_VREF pixel
Xpixel_5940 pixel_5940/gring pixel_5940/VDD pixel_5940/GND pixel_5940/VREF pixel_5940/ROW_SEL
+ pixel_5940/NB1 pixel_5940/VBIAS pixel_5940/NB2 pixel_5940/AMP_IN pixel_5940/SF_IB
+ pixel_5940/PIX_OUT pixel_5940/CSA_VREF pixel
Xpixel_5951 pixel_5951/gring pixel_5951/VDD pixel_5951/GND pixel_5951/VREF pixel_5951/ROW_SEL
+ pixel_5951/NB1 pixel_5951/VBIAS pixel_5951/NB2 pixel_5951/AMP_IN pixel_5951/SF_IB
+ pixel_5951/PIX_OUT pixel_5951/CSA_VREF pixel
Xpixel_5962 pixel_5962/gring pixel_5962/VDD pixel_5962/GND pixel_5962/VREF pixel_5962/ROW_SEL
+ pixel_5962/NB1 pixel_5962/VBIAS pixel_5962/NB2 pixel_5962/AMP_IN pixel_5962/SF_IB
+ pixel_5962/PIX_OUT pixel_5962/CSA_VREF pixel
Xpixel_5973 pixel_5973/gring pixel_5973/VDD pixel_5973/GND pixel_5973/VREF pixel_5973/ROW_SEL
+ pixel_5973/NB1 pixel_5973/VBIAS pixel_5973/NB2 pixel_5973/AMP_IN pixel_5973/SF_IB
+ pixel_5973/PIX_OUT pixel_5973/CSA_VREF pixel
Xpixel_5984 pixel_5984/gring pixel_5984/VDD pixel_5984/GND pixel_5984/VREF pixel_5984/ROW_SEL
+ pixel_5984/NB1 pixel_5984/VBIAS pixel_5984/NB2 pixel_5984/AMP_IN pixel_5984/SF_IB
+ pixel_5984/PIX_OUT pixel_5984/CSA_VREF pixel
Xpixel_5995 pixel_5995/gring pixel_5995/VDD pixel_5995/GND pixel_5995/VREF pixel_5995/ROW_SEL
+ pixel_5995/NB1 pixel_5995/VBIAS pixel_5995/NB2 pixel_5995/AMP_IN pixel_5995/SF_IB
+ pixel_5995/PIX_OUT pixel_5995/CSA_VREF pixel
Xpixel_1909 pixel_1909/gring pixel_1909/VDD pixel_1909/GND pixel_1909/VREF pixel_1909/ROW_SEL
+ pixel_1909/NB1 pixel_1909/VBIAS pixel_1909/NB2 pixel_1909/AMP_IN pixel_1909/SF_IB
+ pixel_1909/PIX_OUT pixel_1909/CSA_VREF pixel
Xpixel_5203 pixel_5203/gring pixel_5203/VDD pixel_5203/GND pixel_5203/VREF pixel_5203/ROW_SEL
+ pixel_5203/NB1 pixel_5203/VBIAS pixel_5203/NB2 pixel_5203/AMP_IN pixel_5203/SF_IB
+ pixel_5203/PIX_OUT pixel_5203/CSA_VREF pixel
Xpixel_5214 pixel_5214/gring pixel_5214/VDD pixel_5214/GND pixel_5214/VREF pixel_5214/ROW_SEL
+ pixel_5214/NB1 pixel_5214/VBIAS pixel_5214/NB2 pixel_5214/AMP_IN pixel_5214/SF_IB
+ pixel_5214/PIX_OUT pixel_5214/CSA_VREF pixel
Xpixel_5225 pixel_5225/gring pixel_5225/VDD pixel_5225/GND pixel_5225/VREF pixel_5225/ROW_SEL
+ pixel_5225/NB1 pixel_5225/VBIAS pixel_5225/NB2 pixel_5225/AMP_IN pixel_5225/SF_IB
+ pixel_5225/PIX_OUT pixel_5225/CSA_VREF pixel
Xpixel_5236 pixel_5236/gring pixel_5236/VDD pixel_5236/GND pixel_5236/VREF pixel_5236/ROW_SEL
+ pixel_5236/NB1 pixel_5236/VBIAS pixel_5236/NB2 pixel_5236/AMP_IN pixel_5236/SF_IB
+ pixel_5236/PIX_OUT pixel_5236/CSA_VREF pixel
Xpixel_5247 pixel_5247/gring pixel_5247/VDD pixel_5247/GND pixel_5247/VREF pixel_5247/ROW_SEL
+ pixel_5247/NB1 pixel_5247/VBIAS pixel_5247/NB2 pixel_5247/AMP_IN pixel_5247/SF_IB
+ pixel_5247/PIX_OUT pixel_5247/CSA_VREF pixel
Xpixel_4502 pixel_4502/gring pixel_4502/VDD pixel_4502/GND pixel_4502/VREF pixel_4502/ROW_SEL
+ pixel_4502/NB1 pixel_4502/VBIAS pixel_4502/NB2 pixel_4502/AMP_IN pixel_4502/SF_IB
+ pixel_4502/PIX_OUT pixel_4502/CSA_VREF pixel
Xpixel_541 pixel_541/gring pixel_541/VDD pixel_541/GND pixel_541/VREF pixel_541/ROW_SEL
+ pixel_541/NB1 pixel_541/VBIAS pixel_541/NB2 pixel_541/AMP_IN pixel_541/SF_IB pixel_541/PIX_OUT
+ pixel_541/CSA_VREF pixel
Xpixel_530 pixel_530/gring pixel_530/VDD pixel_530/GND pixel_530/VREF pixel_530/ROW_SEL
+ pixel_530/NB1 pixel_530/VBIAS pixel_530/NB2 pixel_530/AMP_IN pixel_530/SF_IB pixel_530/PIX_OUT
+ pixel_530/CSA_VREF pixel
Xpixel_5258 pixel_5258/gring pixel_5258/VDD pixel_5258/GND pixel_5258/VREF pixel_5258/ROW_SEL
+ pixel_5258/NB1 pixel_5258/VBIAS pixel_5258/NB2 pixel_5258/AMP_IN pixel_5258/SF_IB
+ pixel_5258/PIX_OUT pixel_5258/CSA_VREF pixel
Xpixel_5269 pixel_5269/gring pixel_5269/VDD pixel_5269/GND pixel_5269/VREF pixel_5269/ROW_SEL
+ pixel_5269/NB1 pixel_5269/VBIAS pixel_5269/NB2 pixel_5269/AMP_IN pixel_5269/SF_IB
+ pixel_5269/PIX_OUT pixel_5269/CSA_VREF pixel
Xpixel_4513 pixel_4513/gring pixel_4513/VDD pixel_4513/GND pixel_4513/VREF pixel_4513/ROW_SEL
+ pixel_4513/NB1 pixel_4513/VBIAS pixel_4513/NB2 pixel_4513/AMP_IN pixel_4513/SF_IB
+ pixel_4513/PIX_OUT pixel_4513/CSA_VREF pixel
Xpixel_4524 pixel_4524/gring pixel_4524/VDD pixel_4524/GND pixel_4524/VREF pixel_4524/ROW_SEL
+ pixel_4524/NB1 pixel_4524/VBIAS pixel_4524/NB2 pixel_4524/AMP_IN pixel_4524/SF_IB
+ pixel_4524/PIX_OUT pixel_4524/CSA_VREF pixel
Xpixel_4535 pixel_4535/gring pixel_4535/VDD pixel_4535/GND pixel_4535/VREF pixel_4535/ROW_SEL
+ pixel_4535/NB1 pixel_4535/VBIAS pixel_4535/NB2 pixel_4535/AMP_IN pixel_4535/SF_IB
+ pixel_4535/PIX_OUT pixel_4535/CSA_VREF pixel
Xpixel_4546 pixel_4546/gring pixel_4546/VDD pixel_4546/GND pixel_4546/VREF pixel_4546/ROW_SEL
+ pixel_4546/NB1 pixel_4546/VBIAS pixel_4546/NB2 pixel_4546/AMP_IN pixel_4546/SF_IB
+ pixel_4546/PIX_OUT pixel_4546/CSA_VREF pixel
Xpixel_3801 pixel_3801/gring pixel_3801/VDD pixel_3801/GND pixel_3801/VREF pixel_3801/ROW_SEL
+ pixel_3801/NB1 pixel_3801/VBIAS pixel_3801/NB2 pixel_3801/AMP_IN pixel_3801/SF_IB
+ pixel_3801/PIX_OUT pixel_3801/CSA_VREF pixel
Xpixel_574 pixel_574/gring pixel_574/VDD pixel_574/GND pixel_574/VREF pixel_574/ROW_SEL
+ pixel_574/NB1 pixel_574/VBIAS pixel_574/NB2 pixel_574/AMP_IN pixel_574/SF_IB pixel_574/PIX_OUT
+ pixel_574/CSA_VREF pixel
Xpixel_563 pixel_563/gring pixel_563/VDD pixel_563/GND pixel_563/VREF pixel_563/ROW_SEL
+ pixel_563/NB1 pixel_563/VBIAS pixel_563/NB2 pixel_563/AMP_IN pixel_563/SF_IB pixel_563/PIX_OUT
+ pixel_563/CSA_VREF pixel
Xpixel_552 pixel_552/gring pixel_552/VDD pixel_552/GND pixel_552/VREF pixel_552/ROW_SEL
+ pixel_552/NB1 pixel_552/VBIAS pixel_552/NB2 pixel_552/AMP_IN pixel_552/SF_IB pixel_552/PIX_OUT
+ pixel_552/CSA_VREF pixel
Xpixel_4557 pixel_4557/gring pixel_4557/VDD pixel_4557/GND pixel_4557/VREF pixel_4557/ROW_SEL
+ pixel_4557/NB1 pixel_4557/VBIAS pixel_4557/NB2 pixel_4557/AMP_IN pixel_4557/SF_IB
+ pixel_4557/PIX_OUT pixel_4557/CSA_VREF pixel
Xpixel_4568 pixel_4568/gring pixel_4568/VDD pixel_4568/GND pixel_4568/VREF pixel_4568/ROW_SEL
+ pixel_4568/NB1 pixel_4568/VBIAS pixel_4568/NB2 pixel_4568/AMP_IN pixel_4568/SF_IB
+ pixel_4568/PIX_OUT pixel_4568/CSA_VREF pixel
Xpixel_4579 pixel_4579/gring pixel_4579/VDD pixel_4579/GND pixel_4579/VREF pixel_4579/ROW_SEL
+ pixel_4579/NB1 pixel_4579/VBIAS pixel_4579/NB2 pixel_4579/AMP_IN pixel_4579/SF_IB
+ pixel_4579/PIX_OUT pixel_4579/CSA_VREF pixel
Xpixel_3812 pixel_3812/gring pixel_3812/VDD pixel_3812/GND pixel_3812/VREF pixel_3812/ROW_SEL
+ pixel_3812/NB1 pixel_3812/VBIAS pixel_3812/NB2 pixel_3812/AMP_IN pixel_3812/SF_IB
+ pixel_3812/PIX_OUT pixel_3812/CSA_VREF pixel
Xpixel_3823 pixel_3823/gring pixel_3823/VDD pixel_3823/GND pixel_3823/VREF pixel_3823/ROW_SEL
+ pixel_3823/NB1 pixel_3823/VBIAS pixel_3823/NB2 pixel_3823/AMP_IN pixel_3823/SF_IB
+ pixel_3823/PIX_OUT pixel_3823/CSA_VREF pixel
Xpixel_3834 pixel_3834/gring pixel_3834/VDD pixel_3834/GND pixel_3834/VREF pixel_3834/ROW_SEL
+ pixel_3834/NB1 pixel_3834/VBIAS pixel_3834/NB2 pixel_3834/AMP_IN pixel_3834/SF_IB
+ pixel_3834/PIX_OUT pixel_3834/CSA_VREF pixel
Xpixel_596 pixel_596/gring pixel_596/VDD pixel_596/GND pixel_596/VREF pixel_596/ROW_SEL
+ pixel_596/NB1 pixel_596/VBIAS pixel_596/NB2 pixel_596/AMP_IN pixel_596/SF_IB pixel_596/PIX_OUT
+ pixel_596/CSA_VREF pixel
Xpixel_585 pixel_585/gring pixel_585/VDD pixel_585/GND pixel_585/VREF pixel_585/ROW_SEL
+ pixel_585/NB1 pixel_585/VBIAS pixel_585/NB2 pixel_585/AMP_IN pixel_585/SF_IB pixel_585/PIX_OUT
+ pixel_585/CSA_VREF pixel
Xpixel_3867 pixel_3867/gring pixel_3867/VDD pixel_3867/GND pixel_3867/VREF pixel_3867/ROW_SEL
+ pixel_3867/NB1 pixel_3867/VBIAS pixel_3867/NB2 pixel_3867/AMP_IN pixel_3867/SF_IB
+ pixel_3867/PIX_OUT pixel_3867/CSA_VREF pixel
Xpixel_3856 pixel_3856/gring pixel_3856/VDD pixel_3856/GND pixel_3856/VREF pixel_3856/ROW_SEL
+ pixel_3856/NB1 pixel_3856/VBIAS pixel_3856/NB2 pixel_3856/AMP_IN pixel_3856/SF_IB
+ pixel_3856/PIX_OUT pixel_3856/CSA_VREF pixel
Xpixel_3845 pixel_3845/gring pixel_3845/VDD pixel_3845/GND pixel_3845/VREF pixel_3845/ROW_SEL
+ pixel_3845/NB1 pixel_3845/VBIAS pixel_3845/NB2 pixel_3845/AMP_IN pixel_3845/SF_IB
+ pixel_3845/PIX_OUT pixel_3845/CSA_VREF pixel
Xpixel_3889 pixel_3889/gring pixel_3889/VDD pixel_3889/GND pixel_3889/VREF pixel_3889/ROW_SEL
+ pixel_3889/NB1 pixel_3889/VBIAS pixel_3889/NB2 pixel_3889/AMP_IN pixel_3889/SF_IB
+ pixel_3889/PIX_OUT pixel_3889/CSA_VREF pixel
Xpixel_3878 pixel_3878/gring pixel_3878/VDD pixel_3878/GND pixel_3878/VREF pixel_3878/ROW_SEL
+ pixel_3878/NB1 pixel_3878/VBIAS pixel_3878/NB2 pixel_3878/AMP_IN pixel_3878/SF_IB
+ pixel_3878/PIX_OUT pixel_3878/CSA_VREF pixel
Xpixel_7150 pixel_7150/gring pixel_7150/VDD pixel_7150/GND pixel_7150/VREF pixel_7150/ROW_SEL
+ pixel_7150/NB1 pixel_7150/VBIAS pixel_7150/NB2 pixel_7150/AMP_IN pixel_7150/SF_IB
+ pixel_7150/PIX_OUT pixel_7150/CSA_VREF pixel
Xpixel_7161 pixel_7161/gring pixel_7161/VDD pixel_7161/GND pixel_7161/VREF pixel_7161/ROW_SEL
+ pixel_7161/NB1 pixel_7161/VBIAS pixel_7161/NB2 pixel_7161/AMP_IN pixel_7161/SF_IB
+ pixel_7161/PIX_OUT pixel_7161/CSA_VREF pixel
Xpixel_7172 pixel_7172/gring pixel_7172/VDD pixel_7172/GND pixel_7172/VREF pixel_7172/ROW_SEL
+ pixel_7172/NB1 pixel_7172/VBIAS pixel_7172/NB2 pixel_7172/AMP_IN pixel_7172/SF_IB
+ pixel_7172/PIX_OUT pixel_7172/CSA_VREF pixel
Xpixel_7183 pixel_7183/gring pixel_7183/VDD pixel_7183/GND pixel_7183/VREF pixel_7183/ROW_SEL
+ pixel_7183/NB1 pixel_7183/VBIAS pixel_7183/NB2 pixel_7183/AMP_IN pixel_7183/SF_IB
+ pixel_7183/PIX_OUT pixel_7183/CSA_VREF pixel
Xpixel_7194 pixel_7194/gring pixel_7194/VDD pixel_7194/GND pixel_7194/VREF pixel_7194/ROW_SEL
+ pixel_7194/NB1 pixel_7194/VBIAS pixel_7194/NB2 pixel_7194/AMP_IN pixel_7194/SF_IB
+ pixel_7194/PIX_OUT pixel_7194/CSA_VREF pixel
Xpixel_6460 pixel_6460/gring pixel_6460/VDD pixel_6460/GND pixel_6460/VREF pixel_6460/ROW_SEL
+ pixel_6460/NB1 pixel_6460/VBIAS pixel_6460/NB2 pixel_6460/AMP_IN pixel_6460/SF_IB
+ pixel_6460/PIX_OUT pixel_6460/CSA_VREF pixel
Xpixel_6471 pixel_6471/gring pixel_6471/VDD pixel_6471/GND pixel_6471/VREF pixel_6471/ROW_SEL
+ pixel_6471/NB1 pixel_6471/VBIAS pixel_6471/NB2 pixel_6471/AMP_IN pixel_6471/SF_IB
+ pixel_6471/PIX_OUT pixel_6471/CSA_VREF pixel
Xpixel_6482 pixel_6482/gring pixel_6482/VDD pixel_6482/GND pixel_6482/VREF pixel_6482/ROW_SEL
+ pixel_6482/NB1 pixel_6482/VBIAS pixel_6482/NB2 pixel_6482/AMP_IN pixel_6482/SF_IB
+ pixel_6482/PIX_OUT pixel_6482/CSA_VREF pixel
Xpixel_6493 pixel_6493/gring pixel_6493/VDD pixel_6493/GND pixel_6493/VREF pixel_6493/ROW_SEL
+ pixel_6493/NB1 pixel_6493/VBIAS pixel_6493/NB2 pixel_6493/AMP_IN pixel_6493/SF_IB
+ pixel_6493/PIX_OUT pixel_6493/CSA_VREF pixel
Xpixel_5770 pixel_5770/gring pixel_5770/VDD pixel_5770/GND pixel_5770/VREF pixel_5770/ROW_SEL
+ pixel_5770/NB1 pixel_5770/VBIAS pixel_5770/NB2 pixel_5770/AMP_IN pixel_5770/SF_IB
+ pixel_5770/PIX_OUT pixel_5770/CSA_VREF pixel
Xpixel_5781 pixel_5781/gring pixel_5781/VDD pixel_5781/GND pixel_5781/VREF pixel_5781/ROW_SEL
+ pixel_5781/NB1 pixel_5781/VBIAS pixel_5781/NB2 pixel_5781/AMP_IN pixel_5781/SF_IB
+ pixel_5781/PIX_OUT pixel_5781/CSA_VREF pixel
Xpixel_5792 pixel_5792/gring pixel_5792/VDD pixel_5792/GND pixel_5792/VREF pixel_5792/ROW_SEL
+ pixel_5792/NB1 pixel_5792/VBIAS pixel_5792/NB2 pixel_5792/AMP_IN pixel_5792/SF_IB
+ pixel_5792/PIX_OUT pixel_5792/CSA_VREF pixel
Xpixel_3119 pixel_3119/gring pixel_3119/VDD pixel_3119/GND pixel_3119/VREF pixel_3119/ROW_SEL
+ pixel_3119/NB1 pixel_3119/VBIAS pixel_3119/NB2 pixel_3119/AMP_IN pixel_3119/SF_IB
+ pixel_3119/PIX_OUT pixel_3119/CSA_VREF pixel
Xpixel_3108 pixel_3108/gring pixel_3108/VDD pixel_3108/GND pixel_3108/VREF pixel_3108/ROW_SEL
+ pixel_3108/NB1 pixel_3108/VBIAS pixel_3108/NB2 pixel_3108/AMP_IN pixel_3108/SF_IB
+ pixel_3108/PIX_OUT pixel_3108/CSA_VREF pixel
Xpixel_2418 pixel_2418/gring pixel_2418/VDD pixel_2418/GND pixel_2418/VREF pixel_2418/ROW_SEL
+ pixel_2418/NB1 pixel_2418/VBIAS pixel_2418/NB2 pixel_2418/AMP_IN pixel_2418/SF_IB
+ pixel_2418/PIX_OUT pixel_2418/CSA_VREF pixel
Xpixel_2407 pixel_2407/gring pixel_2407/VDD pixel_2407/GND pixel_2407/VREF pixel_2407/ROW_SEL
+ pixel_2407/NB1 pixel_2407/VBIAS pixel_2407/NB2 pixel_2407/AMP_IN pixel_2407/SF_IB
+ pixel_2407/PIX_OUT pixel_2407/CSA_VREF pixel
Xpixel_1717 pixel_1717/gring pixel_1717/VDD pixel_1717/GND pixel_1717/VREF pixel_1717/ROW_SEL
+ pixel_1717/NB1 pixel_1717/VBIAS pixel_1717/NB2 pixel_1717/AMP_IN pixel_1717/SF_IB
+ pixel_1717/PIX_OUT pixel_1717/CSA_VREF pixel
Xpixel_1706 pixel_1706/gring pixel_1706/VDD pixel_1706/GND pixel_1706/VREF pixel_1706/ROW_SEL
+ pixel_1706/NB1 pixel_1706/VBIAS pixel_1706/NB2 pixel_1706/AMP_IN pixel_1706/SF_IB
+ pixel_1706/PIX_OUT pixel_1706/CSA_VREF pixel
Xpixel_2429 pixel_2429/gring pixel_2429/VDD pixel_2429/GND pixel_2429/VREF pixel_2429/ROW_SEL
+ pixel_2429/NB1 pixel_2429/VBIAS pixel_2429/NB2 pixel_2429/AMP_IN pixel_2429/SF_IB
+ pixel_2429/PIX_OUT pixel_2429/CSA_VREF pixel
Xpixel_1739 pixel_1739/gring pixel_1739/VDD pixel_1739/GND pixel_1739/VREF pixel_1739/ROW_SEL
+ pixel_1739/NB1 pixel_1739/VBIAS pixel_1739/NB2 pixel_1739/AMP_IN pixel_1739/SF_IB
+ pixel_1739/PIX_OUT pixel_1739/CSA_VREF pixel
Xpixel_1728 pixel_1728/gring pixel_1728/VDD pixel_1728/GND pixel_1728/VREF pixel_1728/ROW_SEL
+ pixel_1728/NB1 pixel_1728/VBIAS pixel_1728/NB2 pixel_1728/AMP_IN pixel_1728/SF_IB
+ pixel_1728/PIX_OUT pixel_1728/CSA_VREF pixel
Xpixel_5000 pixel_5000/gring pixel_5000/VDD pixel_5000/GND pixel_5000/VREF pixel_5000/ROW_SEL
+ pixel_5000/NB1 pixel_5000/VBIAS pixel_5000/NB2 pixel_5000/AMP_IN pixel_5000/SF_IB
+ pixel_5000/PIX_OUT pixel_5000/CSA_VREF pixel
Xpixel_5011 pixel_5011/gring pixel_5011/VDD pixel_5011/GND pixel_5011/VREF pixel_5011/ROW_SEL
+ pixel_5011/NB1 pixel_5011/VBIAS pixel_5011/NB2 pixel_5011/AMP_IN pixel_5011/SF_IB
+ pixel_5011/PIX_OUT pixel_5011/CSA_VREF pixel
Xpixel_5022 pixel_5022/gring pixel_5022/VDD pixel_5022/GND pixel_5022/VREF pixel_5022/ROW_SEL
+ pixel_5022/NB1 pixel_5022/VBIAS pixel_5022/NB2 pixel_5022/AMP_IN pixel_5022/SF_IB
+ pixel_5022/PIX_OUT pixel_5022/CSA_VREF pixel
Xpixel_5033 pixel_5033/gring pixel_5033/VDD pixel_5033/GND pixel_5033/VREF pixel_5033/ROW_SEL
+ pixel_5033/NB1 pixel_5033/VBIAS pixel_5033/NB2 pixel_5033/AMP_IN pixel_5033/SF_IB
+ pixel_5033/PIX_OUT pixel_5033/CSA_VREF pixel
Xpixel_5044 pixel_5044/gring pixel_5044/VDD pixel_5044/GND pixel_5044/VREF pixel_5044/ROW_SEL
+ pixel_5044/NB1 pixel_5044/VBIAS pixel_5044/NB2 pixel_5044/AMP_IN pixel_5044/SF_IB
+ pixel_5044/PIX_OUT pixel_5044/CSA_VREF pixel
Xpixel_5055 pixel_5055/gring pixel_5055/VDD pixel_5055/GND pixel_5055/VREF pixel_5055/ROW_SEL
+ pixel_5055/NB1 pixel_5055/VBIAS pixel_5055/NB2 pixel_5055/AMP_IN pixel_5055/SF_IB
+ pixel_5055/PIX_OUT pixel_5055/CSA_VREF pixel
Xpixel_4310 pixel_4310/gring pixel_4310/VDD pixel_4310/GND pixel_4310/VREF pixel_4310/ROW_SEL
+ pixel_4310/NB1 pixel_4310/VBIAS pixel_4310/NB2 pixel_4310/AMP_IN pixel_4310/SF_IB
+ pixel_4310/PIX_OUT pixel_4310/CSA_VREF pixel
Xpixel_5066 pixel_5066/gring pixel_5066/VDD pixel_5066/GND pixel_5066/VREF pixel_5066/ROW_SEL
+ pixel_5066/NB1 pixel_5066/VBIAS pixel_5066/NB2 pixel_5066/AMP_IN pixel_5066/SF_IB
+ pixel_5066/PIX_OUT pixel_5066/CSA_VREF pixel
Xpixel_5077 pixel_5077/gring pixel_5077/VDD pixel_5077/GND pixel_5077/VREF pixel_5077/ROW_SEL
+ pixel_5077/NB1 pixel_5077/VBIAS pixel_5077/NB2 pixel_5077/AMP_IN pixel_5077/SF_IB
+ pixel_5077/PIX_OUT pixel_5077/CSA_VREF pixel
Xpixel_5088 pixel_5088/gring pixel_5088/VDD pixel_5088/GND pixel_5088/VREF pixel_5088/ROW_SEL
+ pixel_5088/NB1 pixel_5088/VBIAS pixel_5088/NB2 pixel_5088/AMP_IN pixel_5088/SF_IB
+ pixel_5088/PIX_OUT pixel_5088/CSA_VREF pixel
Xpixel_5099 pixel_5099/gring pixel_5099/VDD pixel_5099/GND pixel_5099/VREF pixel_5099/ROW_SEL
+ pixel_5099/NB1 pixel_5099/VBIAS pixel_5099/NB2 pixel_5099/AMP_IN pixel_5099/SF_IB
+ pixel_5099/PIX_OUT pixel_5099/CSA_VREF pixel
Xpixel_4321 pixel_4321/gring pixel_4321/VDD pixel_4321/GND pixel_4321/VREF pixel_4321/ROW_SEL
+ pixel_4321/NB1 pixel_4321/VBIAS pixel_4321/NB2 pixel_4321/AMP_IN pixel_4321/SF_IB
+ pixel_4321/PIX_OUT pixel_4321/CSA_VREF pixel
Xpixel_4332 pixel_4332/gring pixel_4332/VDD pixel_4332/GND pixel_4332/VREF pixel_4332/ROW_SEL
+ pixel_4332/NB1 pixel_4332/VBIAS pixel_4332/NB2 pixel_4332/AMP_IN pixel_4332/SF_IB
+ pixel_4332/PIX_OUT pixel_4332/CSA_VREF pixel
Xpixel_4343 pixel_4343/gring pixel_4343/VDD pixel_4343/GND pixel_4343/VREF pixel_4343/ROW_SEL
+ pixel_4343/NB1 pixel_4343/VBIAS pixel_4343/NB2 pixel_4343/AMP_IN pixel_4343/SF_IB
+ pixel_4343/PIX_OUT pixel_4343/CSA_VREF pixel
Xpixel_4354 pixel_4354/gring pixel_4354/VDD pixel_4354/GND pixel_4354/VREF pixel_4354/ROW_SEL
+ pixel_4354/NB1 pixel_4354/VBIAS pixel_4354/NB2 pixel_4354/AMP_IN pixel_4354/SF_IB
+ pixel_4354/PIX_OUT pixel_4354/CSA_VREF pixel
Xpixel_382 pixel_382/gring pixel_382/VDD pixel_382/GND pixel_382/VREF pixel_382/ROW_SEL
+ pixel_382/NB1 pixel_382/VBIAS pixel_382/NB2 pixel_382/AMP_IN pixel_382/SF_IB pixel_382/PIX_OUT
+ pixel_382/CSA_VREF pixel
Xpixel_371 pixel_371/gring pixel_371/VDD pixel_371/GND pixel_371/VREF pixel_371/ROW_SEL
+ pixel_371/NB1 pixel_371/VBIAS pixel_371/NB2 pixel_371/AMP_IN pixel_371/SF_IB pixel_371/PIX_OUT
+ pixel_371/CSA_VREF pixel
Xpixel_360 pixel_360/gring pixel_360/VDD pixel_360/GND pixel_360/VREF pixel_360/ROW_SEL
+ pixel_360/NB1 pixel_360/VBIAS pixel_360/NB2 pixel_360/AMP_IN pixel_360/SF_IB pixel_360/PIX_OUT
+ pixel_360/CSA_VREF pixel
Xpixel_3642 pixel_3642/gring pixel_3642/VDD pixel_3642/GND pixel_3642/VREF pixel_3642/ROW_SEL
+ pixel_3642/NB1 pixel_3642/VBIAS pixel_3642/NB2 pixel_3642/AMP_IN pixel_3642/SF_IB
+ pixel_3642/PIX_OUT pixel_3642/CSA_VREF pixel
Xpixel_3631 pixel_3631/gring pixel_3631/VDD pixel_3631/GND pixel_3631/VREF pixel_3631/ROW_SEL
+ pixel_3631/NB1 pixel_3631/VBIAS pixel_3631/NB2 pixel_3631/AMP_IN pixel_3631/SF_IB
+ pixel_3631/PIX_OUT pixel_3631/CSA_VREF pixel
Xpixel_3620 pixel_3620/gring pixel_3620/VDD pixel_3620/GND pixel_3620/VREF pixel_3620/ROW_SEL
+ pixel_3620/NB1 pixel_3620/VBIAS pixel_3620/NB2 pixel_3620/AMP_IN pixel_3620/SF_IB
+ pixel_3620/PIX_OUT pixel_3620/CSA_VREF pixel
Xpixel_4365 pixel_4365/gring pixel_4365/VDD pixel_4365/GND pixel_4365/VREF pixel_4365/ROW_SEL
+ pixel_4365/NB1 pixel_4365/VBIAS pixel_4365/NB2 pixel_4365/AMP_IN pixel_4365/SF_IB
+ pixel_4365/PIX_OUT pixel_4365/CSA_VREF pixel
Xpixel_4376 pixel_4376/gring pixel_4376/VDD pixel_4376/GND pixel_4376/VREF pixel_4376/ROW_SEL
+ pixel_4376/NB1 pixel_4376/VBIAS pixel_4376/NB2 pixel_4376/AMP_IN pixel_4376/SF_IB
+ pixel_4376/PIX_OUT pixel_4376/CSA_VREF pixel
Xpixel_4387 pixel_4387/gring pixel_4387/VDD pixel_4387/GND pixel_4387/VREF pixel_4387/ROW_SEL
+ pixel_4387/NB1 pixel_4387/VBIAS pixel_4387/NB2 pixel_4387/AMP_IN pixel_4387/SF_IB
+ pixel_4387/PIX_OUT pixel_4387/CSA_VREF pixel
Xpixel_393 pixel_393/gring pixel_393/VDD pixel_393/GND pixel_393/VREF pixel_393/ROW_SEL
+ pixel_393/NB1 pixel_393/VBIAS pixel_393/NB2 pixel_393/AMP_IN pixel_393/SF_IB pixel_393/PIX_OUT
+ pixel_393/CSA_VREF pixel
Xpixel_2941 pixel_2941/gring pixel_2941/VDD pixel_2941/GND pixel_2941/VREF pixel_2941/ROW_SEL
+ pixel_2941/NB1 pixel_2941/VBIAS pixel_2941/NB2 pixel_2941/AMP_IN pixel_2941/SF_IB
+ pixel_2941/PIX_OUT pixel_2941/CSA_VREF pixel
Xpixel_2930 pixel_2930/gring pixel_2930/VDD pixel_2930/GND pixel_2930/VREF pixel_2930/ROW_SEL
+ pixel_2930/NB1 pixel_2930/VBIAS pixel_2930/NB2 pixel_2930/AMP_IN pixel_2930/SF_IB
+ pixel_2930/PIX_OUT pixel_2930/CSA_VREF pixel
Xpixel_3686 pixel_3686/gring pixel_3686/VDD pixel_3686/GND pixel_3686/VREF pixel_3686/ROW_SEL
+ pixel_3686/NB1 pixel_3686/VBIAS pixel_3686/NB2 pixel_3686/AMP_IN pixel_3686/SF_IB
+ pixel_3686/PIX_OUT pixel_3686/CSA_VREF pixel
Xpixel_3675 pixel_3675/gring pixel_3675/VDD pixel_3675/GND pixel_3675/VREF pixel_3675/ROW_SEL
+ pixel_3675/NB1 pixel_3675/VBIAS pixel_3675/NB2 pixel_3675/AMP_IN pixel_3675/SF_IB
+ pixel_3675/PIX_OUT pixel_3675/CSA_VREF pixel
Xpixel_3664 pixel_3664/gring pixel_3664/VDD pixel_3664/GND pixel_3664/VREF pixel_3664/ROW_SEL
+ pixel_3664/NB1 pixel_3664/VBIAS pixel_3664/NB2 pixel_3664/AMP_IN pixel_3664/SF_IB
+ pixel_3664/PIX_OUT pixel_3664/CSA_VREF pixel
Xpixel_3653 pixel_3653/gring pixel_3653/VDD pixel_3653/GND pixel_3653/VREF pixel_3653/ROW_SEL
+ pixel_3653/NB1 pixel_3653/VBIAS pixel_3653/NB2 pixel_3653/AMP_IN pixel_3653/SF_IB
+ pixel_3653/PIX_OUT pixel_3653/CSA_VREF pixel
Xpixel_4398 pixel_4398/gring pixel_4398/VDD pixel_4398/GND pixel_4398/VREF pixel_4398/ROW_SEL
+ pixel_4398/NB1 pixel_4398/VBIAS pixel_4398/NB2 pixel_4398/AMP_IN pixel_4398/SF_IB
+ pixel_4398/PIX_OUT pixel_4398/CSA_VREF pixel
Xpixel_2974 pixel_2974/gring pixel_2974/VDD pixel_2974/GND pixel_2974/VREF pixel_2974/ROW_SEL
+ pixel_2974/NB1 pixel_2974/VBIAS pixel_2974/NB2 pixel_2974/AMP_IN pixel_2974/SF_IB
+ pixel_2974/PIX_OUT pixel_2974/CSA_VREF pixel
Xpixel_2963 pixel_2963/gring pixel_2963/VDD pixel_2963/GND pixel_2963/VREF pixel_2963/ROW_SEL
+ pixel_2963/NB1 pixel_2963/VBIAS pixel_2963/NB2 pixel_2963/AMP_IN pixel_2963/SF_IB
+ pixel_2963/PIX_OUT pixel_2963/CSA_VREF pixel
Xpixel_2952 pixel_2952/gring pixel_2952/VDD pixel_2952/GND pixel_2952/VREF pixel_2952/ROW_SEL
+ pixel_2952/NB1 pixel_2952/VBIAS pixel_2952/NB2 pixel_2952/AMP_IN pixel_2952/SF_IB
+ pixel_2952/PIX_OUT pixel_2952/CSA_VREF pixel
Xpixel_3697 pixel_3697/gring pixel_3697/VDD pixel_3697/GND pixel_3697/VREF pixel_3697/ROW_SEL
+ pixel_3697/NB1 pixel_3697/VBIAS pixel_3697/NB2 pixel_3697/AMP_IN pixel_3697/SF_IB
+ pixel_3697/PIX_OUT pixel_3697/CSA_VREF pixel
Xpixel_2996 pixel_2996/gring pixel_2996/VDD pixel_2996/GND pixel_2996/VREF pixel_2996/ROW_SEL
+ pixel_2996/NB1 pixel_2996/VBIAS pixel_2996/NB2 pixel_2996/AMP_IN pixel_2996/SF_IB
+ pixel_2996/PIX_OUT pixel_2996/CSA_VREF pixel
Xpixel_2985 pixel_2985/gring pixel_2985/VDD pixel_2985/GND pixel_2985/VREF pixel_2985/ROW_SEL
+ pixel_2985/NB1 pixel_2985/VBIAS pixel_2985/NB2 pixel_2985/AMP_IN pixel_2985/SF_IB
+ pixel_2985/PIX_OUT pixel_2985/CSA_VREF pixel
Xpixel_6290 pixel_6290/gring pixel_6290/VDD pixel_6290/GND pixel_6290/VREF pixel_6290/ROW_SEL
+ pixel_6290/NB1 pixel_6290/VBIAS pixel_6290/NB2 pixel_6290/AMP_IN pixel_6290/SF_IB
+ pixel_6290/PIX_OUT pixel_6290/CSA_VREF pixel
Xpixel_8609 pixel_8609/gring pixel_8609/VDD pixel_8609/GND pixel_8609/VREF pixel_8609/ROW_SEL
+ pixel_8609/NB1 pixel_8609/VBIAS pixel_8609/NB2 pixel_8609/AMP_IN pixel_8609/SF_IB
+ pixel_8609/PIX_OUT pixel_8609/CSA_VREF pixel
Xpixel_7908 pixel_7908/gring pixel_7908/VDD pixel_7908/GND pixel_7908/VREF pixel_7908/ROW_SEL
+ pixel_7908/NB1 pixel_7908/VBIAS pixel_7908/NB2 pixel_7908/AMP_IN pixel_7908/SF_IB
+ pixel_7908/PIX_OUT pixel_7908/CSA_VREF pixel
Xpixel_7919 pixel_7919/gring pixel_7919/VDD pixel_7919/GND pixel_7919/VREF pixel_7919/ROW_SEL
+ pixel_7919/NB1 pixel_7919/VBIAS pixel_7919/NB2 pixel_7919/AMP_IN pixel_7919/SF_IB
+ pixel_7919/PIX_OUT pixel_7919/CSA_VREF pixel
Xpixel_2226 pixel_2226/gring pixel_2226/VDD pixel_2226/GND pixel_2226/VREF pixel_2226/ROW_SEL
+ pixel_2226/NB1 pixel_2226/VBIAS pixel_2226/NB2 pixel_2226/AMP_IN pixel_2226/SF_IB
+ pixel_2226/PIX_OUT pixel_2226/CSA_VREF pixel
Xpixel_2215 pixel_2215/gring pixel_2215/VDD pixel_2215/GND pixel_2215/VREF pixel_2215/ROW_SEL
+ pixel_2215/NB1 pixel_2215/VBIAS pixel_2215/NB2 pixel_2215/AMP_IN pixel_2215/SF_IB
+ pixel_2215/PIX_OUT pixel_2215/CSA_VREF pixel
Xpixel_2204 pixel_2204/gring pixel_2204/VDD pixel_2204/GND pixel_2204/VREF pixel_2204/ROW_SEL
+ pixel_2204/NB1 pixel_2204/VBIAS pixel_2204/NB2 pixel_2204/AMP_IN pixel_2204/SF_IB
+ pixel_2204/PIX_OUT pixel_2204/CSA_VREF pixel
Xpixel_1525 pixel_1525/gring pixel_1525/VDD pixel_1525/GND pixel_1525/VREF pixel_1525/ROW_SEL
+ pixel_1525/NB1 pixel_1525/VBIAS pixel_1525/NB2 pixel_1525/AMP_IN pixel_1525/SF_IB
+ pixel_1525/PIX_OUT pixel_1525/CSA_VREF pixel
Xpixel_1514 pixel_1514/gring pixel_1514/VDD pixel_1514/GND pixel_1514/VREF pixel_1514/ROW_SEL
+ pixel_1514/NB1 pixel_1514/VBIAS pixel_1514/NB2 pixel_1514/AMP_IN pixel_1514/SF_IB
+ pixel_1514/PIX_OUT pixel_1514/CSA_VREF pixel
Xpixel_1503 pixel_1503/gring pixel_1503/VDD pixel_1503/GND pixel_1503/VREF pixel_1503/ROW_SEL
+ pixel_1503/NB1 pixel_1503/VBIAS pixel_1503/NB2 pixel_1503/AMP_IN pixel_1503/SF_IB
+ pixel_1503/PIX_OUT pixel_1503/CSA_VREF pixel
Xpixel_2259 pixel_2259/gring pixel_2259/VDD pixel_2259/GND pixel_2259/VREF pixel_2259/ROW_SEL
+ pixel_2259/NB1 pixel_2259/VBIAS pixel_2259/NB2 pixel_2259/AMP_IN pixel_2259/SF_IB
+ pixel_2259/PIX_OUT pixel_2259/CSA_VREF pixel
Xpixel_2248 pixel_2248/gring pixel_2248/VDD pixel_2248/GND pixel_2248/VREF pixel_2248/ROW_SEL
+ pixel_2248/NB1 pixel_2248/VBIAS pixel_2248/NB2 pixel_2248/AMP_IN pixel_2248/SF_IB
+ pixel_2248/PIX_OUT pixel_2248/CSA_VREF pixel
Xpixel_2237 pixel_2237/gring pixel_2237/VDD pixel_2237/GND pixel_2237/VREF pixel_2237/ROW_SEL
+ pixel_2237/NB1 pixel_2237/VBIAS pixel_2237/NB2 pixel_2237/AMP_IN pixel_2237/SF_IB
+ pixel_2237/PIX_OUT pixel_2237/CSA_VREF pixel
Xpixel_1558 pixel_1558/gring pixel_1558/VDD pixel_1558/GND pixel_1558/VREF pixel_1558/ROW_SEL
+ pixel_1558/NB1 pixel_1558/VBIAS pixel_1558/NB2 pixel_1558/AMP_IN pixel_1558/SF_IB
+ pixel_1558/PIX_OUT pixel_1558/CSA_VREF pixel
Xpixel_1547 pixel_1547/gring pixel_1547/VDD pixel_1547/GND pixel_1547/VREF pixel_1547/ROW_SEL
+ pixel_1547/NB1 pixel_1547/VBIAS pixel_1547/NB2 pixel_1547/AMP_IN pixel_1547/SF_IB
+ pixel_1547/PIX_OUT pixel_1547/CSA_VREF pixel
Xpixel_1536 pixel_1536/gring pixel_1536/VDD pixel_1536/GND pixel_1536/VREF pixel_1536/ROW_SEL
+ pixel_1536/NB1 pixel_1536/VBIAS pixel_1536/NB2 pixel_1536/AMP_IN pixel_1536/SF_IB
+ pixel_1536/PIX_OUT pixel_1536/CSA_VREF pixel
Xpixel_1569 pixel_1569/gring pixel_1569/VDD pixel_1569/GND pixel_1569/VREF pixel_1569/ROW_SEL
+ pixel_1569/NB1 pixel_1569/VBIAS pixel_1569/NB2 pixel_1569/AMP_IN pixel_1569/SF_IB
+ pixel_1569/PIX_OUT pixel_1569/CSA_VREF pixel
Xpixel_9833 pixel_9833/gring pixel_9833/VDD pixel_9833/GND pixel_9833/VREF pixel_9833/ROW_SEL
+ pixel_9833/NB1 pixel_9833/VBIAS pixel_9833/NB2 pixel_9833/AMP_IN pixel_9833/SF_IB
+ pixel_9833/PIX_OUT pixel_9833/CSA_VREF pixel
Xpixel_9822 pixel_9822/gring pixel_9822/VDD pixel_9822/GND pixel_9822/VREF pixel_9822/ROW_SEL
+ pixel_9822/NB1 pixel_9822/VBIAS pixel_9822/NB2 pixel_9822/AMP_IN pixel_9822/SF_IB
+ pixel_9822/PIX_OUT pixel_9822/CSA_VREF pixel
Xpixel_9811 pixel_9811/gring pixel_9811/VDD pixel_9811/GND pixel_9811/VREF pixel_9811/ROW_SEL
+ pixel_9811/NB1 pixel_9811/VBIAS pixel_9811/NB2 pixel_9811/AMP_IN pixel_9811/SF_IB
+ pixel_9811/PIX_OUT pixel_9811/CSA_VREF pixel
Xpixel_9800 pixel_9800/gring pixel_9800/VDD pixel_9800/GND pixel_9800/VREF pixel_9800/ROW_SEL
+ pixel_9800/NB1 pixel_9800/VBIAS pixel_9800/NB2 pixel_9800/AMP_IN pixel_9800/SF_IB
+ pixel_9800/PIX_OUT pixel_9800/CSA_VREF pixel
Xpixel_9844 pixel_9844/gring pixel_9844/VDD pixel_9844/GND pixel_9844/VREF pixel_9844/ROW_SEL
+ pixel_9844/NB1 pixel_9844/VBIAS pixel_9844/NB2 pixel_9844/AMP_IN pixel_9844/SF_IB
+ pixel_9844/PIX_OUT pixel_9844/CSA_VREF pixel
Xpixel_9855 pixel_9855/gring pixel_9855/VDD pixel_9855/GND pixel_9855/VREF pixel_9855/ROW_SEL
+ pixel_9855/NB1 pixel_9855/VBIAS pixel_9855/NB2 pixel_9855/AMP_IN pixel_9855/SF_IB
+ pixel_9855/PIX_OUT pixel_9855/CSA_VREF pixel
Xpixel_9866 pixel_9866/gring pixel_9866/VDD pixel_9866/GND pixel_9866/VREF pixel_9866/ROW_SEL
+ pixel_9866/NB1 pixel_9866/VBIAS pixel_9866/NB2 pixel_9866/AMP_IN pixel_9866/SF_IB
+ pixel_9866/PIX_OUT pixel_9866/CSA_VREF pixel
Xpixel_9877 pixel_9877/gring pixel_9877/VDD pixel_9877/GND pixel_9877/VREF pixel_9877/ROW_SEL
+ pixel_9877/NB1 pixel_9877/VBIAS pixel_9877/NB2 pixel_9877/AMP_IN pixel_9877/SF_IB
+ pixel_9877/PIX_OUT pixel_9877/CSA_VREF pixel
Xpixel_9888 pixel_9888/gring pixel_9888/VDD pixel_9888/GND pixel_9888/VREF pixel_9888/ROW_SEL
+ pixel_9888/NB1 pixel_9888/VBIAS pixel_9888/NB2 pixel_9888/AMP_IN pixel_9888/SF_IB
+ pixel_9888/PIX_OUT pixel_9888/CSA_VREF pixel
Xpixel_9899 pixel_9899/gring pixel_9899/VDD pixel_9899/GND pixel_9899/VREF pixel_9899/ROW_SEL
+ pixel_9899/NB1 pixel_9899/VBIAS pixel_9899/NB2 pixel_9899/AMP_IN pixel_9899/SF_IB
+ pixel_9899/PIX_OUT pixel_9899/CSA_VREF pixel
Xpixel_4140 pixel_4140/gring pixel_4140/VDD pixel_4140/GND pixel_4140/VREF pixel_4140/ROW_SEL
+ pixel_4140/NB1 pixel_4140/VBIAS pixel_4140/NB2 pixel_4140/AMP_IN pixel_4140/SF_IB
+ pixel_4140/PIX_OUT pixel_4140/CSA_VREF pixel
Xpixel_4151 pixel_4151/gring pixel_4151/VDD pixel_4151/GND pixel_4151/VREF pixel_4151/ROW_SEL
+ pixel_4151/NB1 pixel_4151/VBIAS pixel_4151/NB2 pixel_4151/AMP_IN pixel_4151/SF_IB
+ pixel_4151/PIX_OUT pixel_4151/CSA_VREF pixel
Xpixel_4162 pixel_4162/gring pixel_4162/VDD pixel_4162/GND pixel_4162/VREF pixel_4162/ROW_SEL
+ pixel_4162/NB1 pixel_4162/VBIAS pixel_4162/NB2 pixel_4162/AMP_IN pixel_4162/SF_IB
+ pixel_4162/PIX_OUT pixel_4162/CSA_VREF pixel
Xpixel_190 pixel_190/gring pixel_190/VDD pixel_190/GND pixel_190/VREF pixel_190/ROW_SEL
+ pixel_190/NB1 pixel_190/VBIAS pixel_190/NB2 pixel_190/AMP_IN pixel_190/SF_IB pixel_190/PIX_OUT
+ pixel_190/CSA_VREF pixel
Xpixel_3450 pixel_3450/gring pixel_3450/VDD pixel_3450/GND pixel_3450/VREF pixel_3450/ROW_SEL
+ pixel_3450/NB1 pixel_3450/VBIAS pixel_3450/NB2 pixel_3450/AMP_IN pixel_3450/SF_IB
+ pixel_3450/PIX_OUT pixel_3450/CSA_VREF pixel
Xpixel_4173 pixel_4173/gring pixel_4173/VDD pixel_4173/GND pixel_4173/VREF pixel_4173/ROW_SEL
+ pixel_4173/NB1 pixel_4173/VBIAS pixel_4173/NB2 pixel_4173/AMP_IN pixel_4173/SF_IB
+ pixel_4173/PIX_OUT pixel_4173/CSA_VREF pixel
Xpixel_4184 pixel_4184/gring pixel_4184/VDD pixel_4184/GND pixel_4184/VREF pixel_4184/ROW_SEL
+ pixel_4184/NB1 pixel_4184/VBIAS pixel_4184/NB2 pixel_4184/AMP_IN pixel_4184/SF_IB
+ pixel_4184/PIX_OUT pixel_4184/CSA_VREF pixel
Xpixel_4195 pixel_4195/gring pixel_4195/VDD pixel_4195/GND pixel_4195/VREF pixel_4195/ROW_SEL
+ pixel_4195/NB1 pixel_4195/VBIAS pixel_4195/NB2 pixel_4195/AMP_IN pixel_4195/SF_IB
+ pixel_4195/PIX_OUT pixel_4195/CSA_VREF pixel
Xpixel_3494 pixel_3494/gring pixel_3494/VDD pixel_3494/GND pixel_3494/VREF pixel_3494/ROW_SEL
+ pixel_3494/NB1 pixel_3494/VBIAS pixel_3494/NB2 pixel_3494/AMP_IN pixel_3494/SF_IB
+ pixel_3494/PIX_OUT pixel_3494/CSA_VREF pixel
Xpixel_3483 pixel_3483/gring pixel_3483/VDD pixel_3483/GND pixel_3483/VREF pixel_3483/ROW_SEL
+ pixel_3483/NB1 pixel_3483/VBIAS pixel_3483/NB2 pixel_3483/AMP_IN pixel_3483/SF_IB
+ pixel_3483/PIX_OUT pixel_3483/CSA_VREF pixel
Xpixel_3472 pixel_3472/gring pixel_3472/VDD pixel_3472/GND pixel_3472/VREF pixel_3472/ROW_SEL
+ pixel_3472/NB1 pixel_3472/VBIAS pixel_3472/NB2 pixel_3472/AMP_IN pixel_3472/SF_IB
+ pixel_3472/PIX_OUT pixel_3472/CSA_VREF pixel
Xpixel_3461 pixel_3461/gring pixel_3461/VDD pixel_3461/GND pixel_3461/VREF pixel_3461/ROW_SEL
+ pixel_3461/NB1 pixel_3461/VBIAS pixel_3461/NB2 pixel_3461/AMP_IN pixel_3461/SF_IB
+ pixel_3461/PIX_OUT pixel_3461/CSA_VREF pixel
Xpixel_2782 pixel_2782/gring pixel_2782/VDD pixel_2782/GND pixel_2782/VREF pixel_2782/ROW_SEL
+ pixel_2782/NB1 pixel_2782/VBIAS pixel_2782/NB2 pixel_2782/AMP_IN pixel_2782/SF_IB
+ pixel_2782/PIX_OUT pixel_2782/CSA_VREF pixel
Xpixel_2771 pixel_2771/gring pixel_2771/VDD pixel_2771/GND pixel_2771/VREF pixel_2771/ROW_SEL
+ pixel_2771/NB1 pixel_2771/VBIAS pixel_2771/NB2 pixel_2771/AMP_IN pixel_2771/SF_IB
+ pixel_2771/PIX_OUT pixel_2771/CSA_VREF pixel
Xpixel_2760 pixel_2760/gring pixel_2760/VDD pixel_2760/GND pixel_2760/VREF pixel_2760/ROW_SEL
+ pixel_2760/NB1 pixel_2760/VBIAS pixel_2760/NB2 pixel_2760/AMP_IN pixel_2760/SF_IB
+ pixel_2760/PIX_OUT pixel_2760/CSA_VREF pixel
Xpixel_2793 pixel_2793/gring pixel_2793/VDD pixel_2793/GND pixel_2793/VREF pixel_2793/ROW_SEL
+ pixel_2793/NB1 pixel_2793/VBIAS pixel_2793/NB2 pixel_2793/AMP_IN pixel_2793/SF_IB
+ pixel_2793/PIX_OUT pixel_2793/CSA_VREF pixel
Xpixel_9118 pixel_9118/gring pixel_9118/VDD pixel_9118/GND pixel_9118/VREF pixel_9118/ROW_SEL
+ pixel_9118/NB1 pixel_9118/VBIAS pixel_9118/NB2 pixel_9118/AMP_IN pixel_9118/SF_IB
+ pixel_9118/PIX_OUT pixel_9118/CSA_VREF pixel
Xpixel_9107 pixel_9107/gring pixel_9107/VDD pixel_9107/GND pixel_9107/VREF pixel_9107/ROW_SEL
+ pixel_9107/NB1 pixel_9107/VBIAS pixel_9107/NB2 pixel_9107/AMP_IN pixel_9107/SF_IB
+ pixel_9107/PIX_OUT pixel_9107/CSA_VREF pixel
Xpixel_8417 pixel_8417/gring pixel_8417/VDD pixel_8417/GND pixel_8417/VREF pixel_8417/ROW_SEL
+ pixel_8417/NB1 pixel_8417/VBIAS pixel_8417/NB2 pixel_8417/AMP_IN pixel_8417/SF_IB
+ pixel_8417/PIX_OUT pixel_8417/CSA_VREF pixel
Xpixel_8406 pixel_8406/gring pixel_8406/VDD pixel_8406/GND pixel_8406/VREF pixel_8406/ROW_SEL
+ pixel_8406/NB1 pixel_8406/VBIAS pixel_8406/NB2 pixel_8406/AMP_IN pixel_8406/SF_IB
+ pixel_8406/PIX_OUT pixel_8406/CSA_VREF pixel
Xpixel_9129 pixel_9129/gring pixel_9129/VDD pixel_9129/GND pixel_9129/VREF pixel_9129/ROW_SEL
+ pixel_9129/NB1 pixel_9129/VBIAS pixel_9129/NB2 pixel_9129/AMP_IN pixel_9129/SF_IB
+ pixel_9129/PIX_OUT pixel_9129/CSA_VREF pixel
Xpixel_8428 pixel_8428/gring pixel_8428/VDD pixel_8428/GND pixel_8428/VREF pixel_8428/ROW_SEL
+ pixel_8428/NB1 pixel_8428/VBIAS pixel_8428/NB2 pixel_8428/AMP_IN pixel_8428/SF_IB
+ pixel_8428/PIX_OUT pixel_8428/CSA_VREF pixel
Xpixel_8439 pixel_8439/gring pixel_8439/VDD pixel_8439/GND pixel_8439/VREF pixel_8439/ROW_SEL
+ pixel_8439/NB1 pixel_8439/VBIAS pixel_8439/NB2 pixel_8439/AMP_IN pixel_8439/SF_IB
+ pixel_8439/PIX_OUT pixel_8439/CSA_VREF pixel
Xpixel_7705 pixel_7705/gring pixel_7705/VDD pixel_7705/GND pixel_7705/VREF pixel_7705/ROW_SEL
+ pixel_7705/NB1 pixel_7705/VBIAS pixel_7705/NB2 pixel_7705/AMP_IN pixel_7705/SF_IB
+ pixel_7705/PIX_OUT pixel_7705/CSA_VREF pixel
Xpixel_7716 pixel_7716/gring pixel_7716/VDD pixel_7716/GND pixel_7716/VREF pixel_7716/ROW_SEL
+ pixel_7716/NB1 pixel_7716/VBIAS pixel_7716/NB2 pixel_7716/AMP_IN pixel_7716/SF_IB
+ pixel_7716/PIX_OUT pixel_7716/CSA_VREF pixel
Xpixel_7727 pixel_7727/gring pixel_7727/VDD pixel_7727/GND pixel_7727/VREF pixel_7727/ROW_SEL
+ pixel_7727/NB1 pixel_7727/VBIAS pixel_7727/NB2 pixel_7727/AMP_IN pixel_7727/SF_IB
+ pixel_7727/PIX_OUT pixel_7727/CSA_VREF pixel
Xpixel_7738 pixel_7738/gring pixel_7738/VDD pixel_7738/GND pixel_7738/VREF pixel_7738/ROW_SEL
+ pixel_7738/NB1 pixel_7738/VBIAS pixel_7738/NB2 pixel_7738/AMP_IN pixel_7738/SF_IB
+ pixel_7738/PIX_OUT pixel_7738/CSA_VREF pixel
Xpixel_7749 pixel_7749/gring pixel_7749/VDD pixel_7749/GND pixel_7749/VREF pixel_7749/ROW_SEL
+ pixel_7749/NB1 pixel_7749/VBIAS pixel_7749/NB2 pixel_7749/AMP_IN pixel_7749/SF_IB
+ pixel_7749/PIX_OUT pixel_7749/CSA_VREF pixel
Xpixel_2001 pixel_2001/gring pixel_2001/VDD pixel_2001/GND pixel_2001/VREF pixel_2001/ROW_SEL
+ pixel_2001/NB1 pixel_2001/VBIAS pixel_2001/NB2 pixel_2001/AMP_IN pixel_2001/SF_IB
+ pixel_2001/PIX_OUT pixel_2001/CSA_VREF pixel
Xpixel_1300 pixel_1300/gring pixel_1300/VDD pixel_1300/GND pixel_1300/VREF pixel_1300/ROW_SEL
+ pixel_1300/NB1 pixel_1300/VBIAS pixel_1300/NB2 pixel_1300/AMP_IN pixel_1300/SF_IB
+ pixel_1300/PIX_OUT pixel_1300/CSA_VREF pixel
Xpixel_2045 pixel_2045/gring pixel_2045/VDD pixel_2045/GND pixel_2045/VREF pixel_2045/ROW_SEL
+ pixel_2045/NB1 pixel_2045/VBIAS pixel_2045/NB2 pixel_2045/AMP_IN pixel_2045/SF_IB
+ pixel_2045/PIX_OUT pixel_2045/CSA_VREF pixel
Xpixel_2034 pixel_2034/gring pixel_2034/VDD pixel_2034/GND pixel_2034/VREF pixel_2034/ROW_SEL
+ pixel_2034/NB1 pixel_2034/VBIAS pixel_2034/NB2 pixel_2034/AMP_IN pixel_2034/SF_IB
+ pixel_2034/PIX_OUT pixel_2034/CSA_VREF pixel
Xpixel_2023 pixel_2023/gring pixel_2023/VDD pixel_2023/GND pixel_2023/VREF pixel_2023/ROW_SEL
+ pixel_2023/NB1 pixel_2023/VBIAS pixel_2023/NB2 pixel_2023/AMP_IN pixel_2023/SF_IB
+ pixel_2023/PIX_OUT pixel_2023/CSA_VREF pixel
Xpixel_2012 pixel_2012/gring pixel_2012/VDD pixel_2012/GND pixel_2012/VREF pixel_2012/ROW_SEL
+ pixel_2012/NB1 pixel_2012/VBIAS pixel_2012/NB2 pixel_2012/AMP_IN pixel_2012/SF_IB
+ pixel_2012/PIX_OUT pixel_2012/CSA_VREF pixel
Xpixel_1333 pixel_1333/gring pixel_1333/VDD pixel_1333/GND pixel_1333/VREF pixel_1333/ROW_SEL
+ pixel_1333/NB1 pixel_1333/VBIAS pixel_1333/NB2 pixel_1333/AMP_IN pixel_1333/SF_IB
+ pixel_1333/PIX_OUT pixel_1333/CSA_VREF pixel
Xpixel_1322 pixel_1322/gring pixel_1322/VDD pixel_1322/GND pixel_1322/VREF pixel_1322/ROW_SEL
+ pixel_1322/NB1 pixel_1322/VBIAS pixel_1322/NB2 pixel_1322/AMP_IN pixel_1322/SF_IB
+ pixel_1322/PIX_OUT pixel_1322/CSA_VREF pixel
Xpixel_1311 pixel_1311/gring pixel_1311/VDD pixel_1311/GND pixel_1311/VREF pixel_1311/ROW_SEL
+ pixel_1311/NB1 pixel_1311/VBIAS pixel_1311/NB2 pixel_1311/AMP_IN pixel_1311/SF_IB
+ pixel_1311/PIX_OUT pixel_1311/CSA_VREF pixel
Xpixel_2078 pixel_2078/gring pixel_2078/VDD pixel_2078/GND pixel_2078/VREF pixel_2078/ROW_SEL
+ pixel_2078/NB1 pixel_2078/VBIAS pixel_2078/NB2 pixel_2078/AMP_IN pixel_2078/SF_IB
+ pixel_2078/PIX_OUT pixel_2078/CSA_VREF pixel
Xpixel_2067 pixel_2067/gring pixel_2067/VDD pixel_2067/GND pixel_2067/VREF pixel_2067/ROW_SEL
+ pixel_2067/NB1 pixel_2067/VBIAS pixel_2067/NB2 pixel_2067/AMP_IN pixel_2067/SF_IB
+ pixel_2067/PIX_OUT pixel_2067/CSA_VREF pixel
Xpixel_2056 pixel_2056/gring pixel_2056/VDD pixel_2056/GND pixel_2056/VREF pixel_2056/ROW_SEL
+ pixel_2056/NB1 pixel_2056/VBIAS pixel_2056/NB2 pixel_2056/AMP_IN pixel_2056/SF_IB
+ pixel_2056/PIX_OUT pixel_2056/CSA_VREF pixel
Xpixel_1366 pixel_1366/gring pixel_1366/VDD pixel_1366/GND pixel_1366/VREF pixel_1366/ROW_SEL
+ pixel_1366/NB1 pixel_1366/VBIAS pixel_1366/NB2 pixel_1366/AMP_IN pixel_1366/SF_IB
+ pixel_1366/PIX_OUT pixel_1366/CSA_VREF pixel
Xpixel_1355 pixel_1355/gring pixel_1355/VDD pixel_1355/GND pixel_1355/VREF pixel_1355/ROW_SEL
+ pixel_1355/NB1 pixel_1355/VBIAS pixel_1355/NB2 pixel_1355/AMP_IN pixel_1355/SF_IB
+ pixel_1355/PIX_OUT pixel_1355/CSA_VREF pixel
Xpixel_1344 pixel_1344/gring pixel_1344/VDD pixel_1344/GND pixel_1344/VREF pixel_1344/ROW_SEL
+ pixel_1344/NB1 pixel_1344/VBIAS pixel_1344/NB2 pixel_1344/AMP_IN pixel_1344/SF_IB
+ pixel_1344/PIX_OUT pixel_1344/CSA_VREF pixel
Xpixel_2089 pixel_2089/gring pixel_2089/VDD pixel_2089/GND pixel_2089/VREF pixel_2089/ROW_SEL
+ pixel_2089/NB1 pixel_2089/VBIAS pixel_2089/NB2 pixel_2089/AMP_IN pixel_2089/SF_IB
+ pixel_2089/PIX_OUT pixel_2089/CSA_VREF pixel
Xpixel_1399 pixel_1399/gring pixel_1399/VDD pixel_1399/GND pixel_1399/VREF pixel_1399/ROW_SEL
+ pixel_1399/NB1 pixel_1399/VBIAS pixel_1399/NB2 pixel_1399/AMP_IN pixel_1399/SF_IB
+ pixel_1399/PIX_OUT pixel_1399/CSA_VREF pixel
Xpixel_1388 pixel_1388/gring pixel_1388/VDD pixel_1388/GND pixel_1388/VREF pixel_1388/ROW_SEL
+ pixel_1388/NB1 pixel_1388/VBIAS pixel_1388/NB2 pixel_1388/AMP_IN pixel_1388/SF_IB
+ pixel_1388/PIX_OUT pixel_1388/CSA_VREF pixel
Xpixel_1377 pixel_1377/gring pixel_1377/VDD pixel_1377/GND pixel_1377/VREF pixel_1377/ROW_SEL
+ pixel_1377/NB1 pixel_1377/VBIAS pixel_1377/NB2 pixel_1377/AMP_IN pixel_1377/SF_IB
+ pixel_1377/PIX_OUT pixel_1377/CSA_VREF pixel
Xpixel_9630 pixel_9630/gring pixel_9630/VDD pixel_9630/GND pixel_9630/VREF pixel_9630/ROW_SEL
+ pixel_9630/NB1 pixel_9630/VBIAS pixel_9630/NB2 pixel_9630/AMP_IN pixel_9630/SF_IB
+ pixel_9630/PIX_OUT pixel_9630/CSA_VREF pixel
Xpixel_9641 pixel_9641/gring pixel_9641/VDD pixel_9641/GND pixel_9641/VREF pixel_9641/ROW_SEL
+ pixel_9641/NB1 pixel_9641/VBIAS pixel_9641/NB2 pixel_9641/AMP_IN pixel_9641/SF_IB
+ pixel_9641/PIX_OUT pixel_9641/CSA_VREF pixel
Xpixel_9652 pixel_9652/gring pixel_9652/VDD pixel_9652/GND pixel_9652/VREF pixel_9652/ROW_SEL
+ pixel_9652/NB1 pixel_9652/VBIAS pixel_9652/NB2 pixel_9652/AMP_IN pixel_9652/SF_IB
+ pixel_9652/PIX_OUT pixel_9652/CSA_VREF pixel
Xpixel_9663 pixel_9663/gring pixel_9663/VDD pixel_9663/GND pixel_9663/VREF pixel_9663/ROW_SEL
+ pixel_9663/NB1 pixel_9663/VBIAS pixel_9663/NB2 pixel_9663/AMP_IN pixel_9663/SF_IB
+ pixel_9663/PIX_OUT pixel_9663/CSA_VREF pixel
Xpixel_9674 pixel_9674/gring pixel_9674/VDD pixel_9674/GND pixel_9674/VREF pixel_9674/ROW_SEL
+ pixel_9674/NB1 pixel_9674/VBIAS pixel_9674/NB2 pixel_9674/AMP_IN pixel_9674/SF_IB
+ pixel_9674/PIX_OUT pixel_9674/CSA_VREF pixel
Xpixel_8973 pixel_8973/gring pixel_8973/VDD pixel_8973/GND pixel_8973/VREF pixel_8973/ROW_SEL
+ pixel_8973/NB1 pixel_8973/VBIAS pixel_8973/NB2 pixel_8973/AMP_IN pixel_8973/SF_IB
+ pixel_8973/PIX_OUT pixel_8973/CSA_VREF pixel
Xpixel_8962 pixel_8962/gring pixel_8962/VDD pixel_8962/GND pixel_8962/VREF pixel_8962/ROW_SEL
+ pixel_8962/NB1 pixel_8962/VBIAS pixel_8962/NB2 pixel_8962/AMP_IN pixel_8962/SF_IB
+ pixel_8962/PIX_OUT pixel_8962/CSA_VREF pixel
Xpixel_8951 pixel_8951/gring pixel_8951/VDD pixel_8951/GND pixel_8951/VREF pixel_8951/ROW_SEL
+ pixel_8951/NB1 pixel_8951/VBIAS pixel_8951/NB2 pixel_8951/AMP_IN pixel_8951/SF_IB
+ pixel_8951/PIX_OUT pixel_8951/CSA_VREF pixel
Xpixel_8940 pixel_8940/gring pixel_8940/VDD pixel_8940/GND pixel_8940/VREF pixel_8940/ROW_SEL
+ pixel_8940/NB1 pixel_8940/VBIAS pixel_8940/NB2 pixel_8940/AMP_IN pixel_8940/SF_IB
+ pixel_8940/PIX_OUT pixel_8940/CSA_VREF pixel
Xpixel_9696 pixel_9696/gring pixel_9696/VDD pixel_9696/GND pixel_9696/VREF pixel_9696/ROW_SEL
+ pixel_9696/NB1 pixel_9696/VBIAS pixel_9696/NB2 pixel_9696/AMP_IN pixel_9696/SF_IB
+ pixel_9696/PIX_OUT pixel_9696/CSA_VREF pixel
Xpixel_9685 pixel_9685/gring pixel_9685/VDD pixel_9685/GND pixel_9685/VREF pixel_9685/ROW_SEL
+ pixel_9685/NB1 pixel_9685/VBIAS pixel_9685/NB2 pixel_9685/AMP_IN pixel_9685/SF_IB
+ pixel_9685/PIX_OUT pixel_9685/CSA_VREF pixel
Xpixel_8995 pixel_8995/gring pixel_8995/VDD pixel_8995/GND pixel_8995/VREF pixel_8995/ROW_SEL
+ pixel_8995/NB1 pixel_8995/VBIAS pixel_8995/NB2 pixel_8995/AMP_IN pixel_8995/SF_IB
+ pixel_8995/PIX_OUT pixel_8995/CSA_VREF pixel
Xpixel_8984 pixel_8984/gring pixel_8984/VDD pixel_8984/GND pixel_8984/VREF pixel_8984/ROW_SEL
+ pixel_8984/NB1 pixel_8984/VBIAS pixel_8984/NB2 pixel_8984/AMP_IN pixel_8984/SF_IB
+ pixel_8984/PIX_OUT pixel_8984/CSA_VREF pixel
Xpixel_3291 pixel_3291/gring pixel_3291/VDD pixel_3291/GND pixel_3291/VREF pixel_3291/ROW_SEL
+ pixel_3291/NB1 pixel_3291/VBIAS pixel_3291/NB2 pixel_3291/AMP_IN pixel_3291/SF_IB
+ pixel_3291/PIX_OUT pixel_3291/CSA_VREF pixel
Xpixel_3280 pixel_3280/gring pixel_3280/VDD pixel_3280/GND pixel_3280/VREF pixel_3280/ROW_SEL
+ pixel_3280/NB1 pixel_3280/VBIAS pixel_3280/NB2 pixel_3280/AMP_IN pixel_3280/SF_IB
+ pixel_3280/PIX_OUT pixel_3280/CSA_VREF pixel
Xpixel_2590 pixel_2590/gring pixel_2590/VDD pixel_2590/GND pixel_2590/VREF pixel_2590/ROW_SEL
+ pixel_2590/NB1 pixel_2590/VBIAS pixel_2590/NB2 pixel_2590/AMP_IN pixel_2590/SF_IB
+ pixel_2590/PIX_OUT pixel_2590/CSA_VREF pixel
Xpixel_915 pixel_915/gring pixel_915/VDD pixel_915/GND pixel_915/VREF pixel_915/ROW_SEL
+ pixel_915/NB1 pixel_915/VBIAS pixel_915/NB2 pixel_915/AMP_IN pixel_915/SF_IB pixel_915/PIX_OUT
+ pixel_915/CSA_VREF pixel
Xpixel_904 pixel_904/gring pixel_904/VDD pixel_904/GND pixel_904/VREF pixel_904/ROW_SEL
+ pixel_904/NB1 pixel_904/VBIAS pixel_904/NB2 pixel_904/AMP_IN pixel_904/SF_IB pixel_904/PIX_OUT
+ pixel_904/CSA_VREF pixel
Xpixel_4909 pixel_4909/gring pixel_4909/VDD pixel_4909/GND pixel_4909/VREF pixel_4909/ROW_SEL
+ pixel_4909/NB1 pixel_4909/VBIAS pixel_4909/NB2 pixel_4909/AMP_IN pixel_4909/SF_IB
+ pixel_4909/PIX_OUT pixel_4909/CSA_VREF pixel
Xpixel_948 pixel_948/gring pixel_948/VDD pixel_948/GND pixel_948/VREF pixel_948/ROW_SEL
+ pixel_948/NB1 pixel_948/VBIAS pixel_948/NB2 pixel_948/AMP_IN pixel_948/SF_IB pixel_948/PIX_OUT
+ pixel_948/CSA_VREF pixel
Xpixel_937 pixel_937/gring pixel_937/VDD pixel_937/GND pixel_937/VREF pixel_937/ROW_SEL
+ pixel_937/NB1 pixel_937/VBIAS pixel_937/NB2 pixel_937/AMP_IN pixel_937/SF_IB pixel_937/PIX_OUT
+ pixel_937/CSA_VREF pixel
Xpixel_926 pixel_926/gring pixel_926/VDD pixel_926/GND pixel_926/VREF pixel_926/ROW_SEL
+ pixel_926/NB1 pixel_926/VBIAS pixel_926/NB2 pixel_926/AMP_IN pixel_926/SF_IB pixel_926/PIX_OUT
+ pixel_926/CSA_VREF pixel
Xpixel_959 pixel_959/gring pixel_959/VDD pixel_959/GND pixel_959/VREF pixel_959/ROW_SEL
+ pixel_959/NB1 pixel_959/VBIAS pixel_959/NB2 pixel_959/AMP_IN pixel_959/SF_IB pixel_959/PIX_OUT
+ pixel_959/CSA_VREF pixel
Xpixel_8203 pixel_8203/gring pixel_8203/VDD pixel_8203/GND pixel_8203/VREF pixel_8203/ROW_SEL
+ pixel_8203/NB1 pixel_8203/VBIAS pixel_8203/NB2 pixel_8203/AMP_IN pixel_8203/SF_IB
+ pixel_8203/PIX_OUT pixel_8203/CSA_VREF pixel
Xpixel_8214 pixel_8214/gring pixel_8214/VDD pixel_8214/GND pixel_8214/VREF pixel_8214/ROW_SEL
+ pixel_8214/NB1 pixel_8214/VBIAS pixel_8214/NB2 pixel_8214/AMP_IN pixel_8214/SF_IB
+ pixel_8214/PIX_OUT pixel_8214/CSA_VREF pixel
Xpixel_8225 pixel_8225/gring pixel_8225/VDD pixel_8225/GND pixel_8225/VREF pixel_8225/ROW_SEL
+ pixel_8225/NB1 pixel_8225/VBIAS pixel_8225/NB2 pixel_8225/AMP_IN pixel_8225/SF_IB
+ pixel_8225/PIX_OUT pixel_8225/CSA_VREF pixel
Xpixel_8236 pixel_8236/gring pixel_8236/VDD pixel_8236/GND pixel_8236/VREF pixel_8236/ROW_SEL
+ pixel_8236/NB1 pixel_8236/VBIAS pixel_8236/NB2 pixel_8236/AMP_IN pixel_8236/SF_IB
+ pixel_8236/PIX_OUT pixel_8236/CSA_VREF pixel
Xpixel_8247 pixel_8247/gring pixel_8247/VDD pixel_8247/GND pixel_8247/VREF pixel_8247/ROW_SEL
+ pixel_8247/NB1 pixel_8247/VBIAS pixel_8247/NB2 pixel_8247/AMP_IN pixel_8247/SF_IB
+ pixel_8247/PIX_OUT pixel_8247/CSA_VREF pixel
Xpixel_8258 pixel_8258/gring pixel_8258/VDD pixel_8258/GND pixel_8258/VREF pixel_8258/ROW_SEL
+ pixel_8258/NB1 pixel_8258/VBIAS pixel_8258/NB2 pixel_8258/AMP_IN pixel_8258/SF_IB
+ pixel_8258/PIX_OUT pixel_8258/CSA_VREF pixel
Xpixel_7502 pixel_7502/gring pixel_7502/VDD pixel_7502/GND pixel_7502/VREF pixel_7502/ROW_SEL
+ pixel_7502/NB1 pixel_7502/VBIAS pixel_7502/NB2 pixel_7502/AMP_IN pixel_7502/SF_IB
+ pixel_7502/PIX_OUT pixel_7502/CSA_VREF pixel
Xpixel_7513 pixel_7513/gring pixel_7513/VDD pixel_7513/GND pixel_7513/VREF pixel_7513/ROW_SEL
+ pixel_7513/NB1 pixel_7513/VBIAS pixel_7513/NB2 pixel_7513/AMP_IN pixel_7513/SF_IB
+ pixel_7513/PIX_OUT pixel_7513/CSA_VREF pixel
Xpixel_7524 pixel_7524/gring pixel_7524/VDD pixel_7524/GND pixel_7524/VREF pixel_7524/ROW_SEL
+ pixel_7524/NB1 pixel_7524/VBIAS pixel_7524/NB2 pixel_7524/AMP_IN pixel_7524/SF_IB
+ pixel_7524/PIX_OUT pixel_7524/CSA_VREF pixel
Xpixel_8269 pixel_8269/gring pixel_8269/VDD pixel_8269/GND pixel_8269/VREF pixel_8269/ROW_SEL
+ pixel_8269/NB1 pixel_8269/VBIAS pixel_8269/NB2 pixel_8269/AMP_IN pixel_8269/SF_IB
+ pixel_8269/PIX_OUT pixel_8269/CSA_VREF pixel
Xpixel_7535 pixel_7535/gring pixel_7535/VDD pixel_7535/GND pixel_7535/VREF pixel_7535/ROW_SEL
+ pixel_7535/NB1 pixel_7535/VBIAS pixel_7535/NB2 pixel_7535/AMP_IN pixel_7535/SF_IB
+ pixel_7535/PIX_OUT pixel_7535/CSA_VREF pixel
Xpixel_7546 pixel_7546/gring pixel_7546/VDD pixel_7546/GND pixel_7546/VREF pixel_7546/ROW_SEL
+ pixel_7546/NB1 pixel_7546/VBIAS pixel_7546/NB2 pixel_7546/AMP_IN pixel_7546/SF_IB
+ pixel_7546/PIX_OUT pixel_7546/CSA_VREF pixel
Xpixel_7557 pixel_7557/gring pixel_7557/VDD pixel_7557/GND pixel_7557/VREF pixel_7557/ROW_SEL
+ pixel_7557/NB1 pixel_7557/VBIAS pixel_7557/NB2 pixel_7557/AMP_IN pixel_7557/SF_IB
+ pixel_7557/PIX_OUT pixel_7557/CSA_VREF pixel
Xpixel_6801 pixel_6801/gring pixel_6801/VDD pixel_6801/GND pixel_6801/VREF pixel_6801/ROW_SEL
+ pixel_6801/NB1 pixel_6801/VBIAS pixel_6801/NB2 pixel_6801/AMP_IN pixel_6801/SF_IB
+ pixel_6801/PIX_OUT pixel_6801/CSA_VREF pixel
Xpixel_6812 pixel_6812/gring pixel_6812/VDD pixel_6812/GND pixel_6812/VREF pixel_6812/ROW_SEL
+ pixel_6812/NB1 pixel_6812/VBIAS pixel_6812/NB2 pixel_6812/AMP_IN pixel_6812/SF_IB
+ pixel_6812/PIX_OUT pixel_6812/CSA_VREF pixel
Xpixel_7568 pixel_7568/gring pixel_7568/VDD pixel_7568/GND pixel_7568/VREF pixel_7568/ROW_SEL
+ pixel_7568/NB1 pixel_7568/VBIAS pixel_7568/NB2 pixel_7568/AMP_IN pixel_7568/SF_IB
+ pixel_7568/PIX_OUT pixel_7568/CSA_VREF pixel
Xpixel_7579 pixel_7579/gring pixel_7579/VDD pixel_7579/GND pixel_7579/VREF pixel_7579/ROW_SEL
+ pixel_7579/NB1 pixel_7579/VBIAS pixel_7579/NB2 pixel_7579/AMP_IN pixel_7579/SF_IB
+ pixel_7579/PIX_OUT pixel_7579/CSA_VREF pixel
Xpixel_6823 pixel_6823/gring pixel_6823/VDD pixel_6823/GND pixel_6823/VREF pixel_6823/ROW_SEL
+ pixel_6823/NB1 pixel_6823/VBIAS pixel_6823/NB2 pixel_6823/AMP_IN pixel_6823/SF_IB
+ pixel_6823/PIX_OUT pixel_6823/CSA_VREF pixel
Xpixel_6834 pixel_6834/gring pixel_6834/VDD pixel_6834/GND pixel_6834/VREF pixel_6834/ROW_SEL
+ pixel_6834/NB1 pixel_6834/VBIAS pixel_6834/NB2 pixel_6834/AMP_IN pixel_6834/SF_IB
+ pixel_6834/PIX_OUT pixel_6834/CSA_VREF pixel
Xpixel_6845 pixel_6845/gring pixel_6845/VDD pixel_6845/GND pixel_6845/VREF pixel_6845/ROW_SEL
+ pixel_6845/NB1 pixel_6845/VBIAS pixel_6845/NB2 pixel_6845/AMP_IN pixel_6845/SF_IB
+ pixel_6845/PIX_OUT pixel_6845/CSA_VREF pixel
Xpixel_6856 pixel_6856/gring pixel_6856/VDD pixel_6856/GND pixel_6856/VREF pixel_6856/ROW_SEL
+ pixel_6856/NB1 pixel_6856/VBIAS pixel_6856/NB2 pixel_6856/AMP_IN pixel_6856/SF_IB
+ pixel_6856/PIX_OUT pixel_6856/CSA_VREF pixel
Xpixel_6867 pixel_6867/gring pixel_6867/VDD pixel_6867/GND pixel_6867/VREF pixel_6867/ROW_SEL
+ pixel_6867/NB1 pixel_6867/VBIAS pixel_6867/NB2 pixel_6867/AMP_IN pixel_6867/SF_IB
+ pixel_6867/PIX_OUT pixel_6867/CSA_VREF pixel
Xpixel_6878 pixel_6878/gring pixel_6878/VDD pixel_6878/GND pixel_6878/VREF pixel_6878/ROW_SEL
+ pixel_6878/NB1 pixel_6878/VBIAS pixel_6878/NB2 pixel_6878/AMP_IN pixel_6878/SF_IB
+ pixel_6878/PIX_OUT pixel_6878/CSA_VREF pixel
Xpixel_6889 pixel_6889/gring pixel_6889/VDD pixel_6889/GND pixel_6889/VREF pixel_6889/ROW_SEL
+ pixel_6889/NB1 pixel_6889/VBIAS pixel_6889/NB2 pixel_6889/AMP_IN pixel_6889/SF_IB
+ pixel_6889/PIX_OUT pixel_6889/CSA_VREF pixel
Xpixel_1141 pixel_1141/gring pixel_1141/VDD pixel_1141/GND pixel_1141/VREF pixel_1141/ROW_SEL
+ pixel_1141/NB1 pixel_1141/VBIAS pixel_1141/NB2 pixel_1141/AMP_IN pixel_1141/SF_IB
+ pixel_1141/PIX_OUT pixel_1141/CSA_VREF pixel
Xpixel_1130 pixel_1130/gring pixel_1130/VDD pixel_1130/GND pixel_1130/VREF pixel_1130/ROW_SEL
+ pixel_1130/NB1 pixel_1130/VBIAS pixel_1130/NB2 pixel_1130/AMP_IN pixel_1130/SF_IB
+ pixel_1130/PIX_OUT pixel_1130/CSA_VREF pixel
Xpixel_1174 pixel_1174/gring pixel_1174/VDD pixel_1174/GND pixel_1174/VREF pixel_1174/ROW_SEL
+ pixel_1174/NB1 pixel_1174/VBIAS pixel_1174/NB2 pixel_1174/AMP_IN pixel_1174/SF_IB
+ pixel_1174/PIX_OUT pixel_1174/CSA_VREF pixel
Xpixel_1163 pixel_1163/gring pixel_1163/VDD pixel_1163/GND pixel_1163/VREF pixel_1163/ROW_SEL
+ pixel_1163/NB1 pixel_1163/VBIAS pixel_1163/NB2 pixel_1163/AMP_IN pixel_1163/SF_IB
+ pixel_1163/PIX_OUT pixel_1163/CSA_VREF pixel
Xpixel_1152 pixel_1152/gring pixel_1152/VDD pixel_1152/GND pixel_1152/VREF pixel_1152/ROW_SEL
+ pixel_1152/NB1 pixel_1152/VBIAS pixel_1152/NB2 pixel_1152/AMP_IN pixel_1152/SF_IB
+ pixel_1152/PIX_OUT pixel_1152/CSA_VREF pixel
Xpixel_1196 pixel_1196/gring pixel_1196/VDD pixel_1196/GND pixel_1196/VREF pixel_1196/ROW_SEL
+ pixel_1196/NB1 pixel_1196/VBIAS pixel_1196/NB2 pixel_1196/AMP_IN pixel_1196/SF_IB
+ pixel_1196/PIX_OUT pixel_1196/CSA_VREF pixel
Xpixel_1185 pixel_1185/gring pixel_1185/VDD pixel_1185/GND pixel_1185/VREF pixel_1185/ROW_SEL
+ pixel_1185/NB1 pixel_1185/VBIAS pixel_1185/NB2 pixel_1185/AMP_IN pixel_1185/SF_IB
+ pixel_1185/PIX_OUT pixel_1185/CSA_VREF pixel
Xpixel_9482 pixel_9482/gring pixel_9482/VDD pixel_9482/GND pixel_9482/VREF pixel_9482/ROW_SEL
+ pixel_9482/NB1 pixel_9482/VBIAS pixel_9482/NB2 pixel_9482/AMP_IN pixel_9482/SF_IB
+ pixel_9482/PIX_OUT pixel_9482/CSA_VREF pixel
Xpixel_9471 pixel_9471/gring pixel_9471/VDD pixel_9471/GND pixel_9471/VREF pixel_9471/ROW_SEL
+ pixel_9471/NB1 pixel_9471/VBIAS pixel_9471/NB2 pixel_9471/AMP_IN pixel_9471/SF_IB
+ pixel_9471/PIX_OUT pixel_9471/CSA_VREF pixel
Xpixel_9460 pixel_9460/gring pixel_9460/VDD pixel_9460/GND pixel_9460/VREF pixel_9460/ROW_SEL
+ pixel_9460/NB1 pixel_9460/VBIAS pixel_9460/NB2 pixel_9460/AMP_IN pixel_9460/SF_IB
+ pixel_9460/PIX_OUT pixel_9460/CSA_VREF pixel
Xpixel_8781 pixel_8781/gring pixel_8781/VDD pixel_8781/GND pixel_8781/VREF pixel_8781/ROW_SEL
+ pixel_8781/NB1 pixel_8781/VBIAS pixel_8781/NB2 pixel_8781/AMP_IN pixel_8781/SF_IB
+ pixel_8781/PIX_OUT pixel_8781/CSA_VREF pixel
Xpixel_8770 pixel_8770/gring pixel_8770/VDD pixel_8770/GND pixel_8770/VREF pixel_8770/ROW_SEL
+ pixel_8770/NB1 pixel_8770/VBIAS pixel_8770/NB2 pixel_8770/AMP_IN pixel_8770/SF_IB
+ pixel_8770/PIX_OUT pixel_8770/CSA_VREF pixel
Xpixel_9493 pixel_9493/gring pixel_9493/VDD pixel_9493/GND pixel_9493/VREF pixel_9493/ROW_SEL
+ pixel_9493/NB1 pixel_9493/VBIAS pixel_9493/NB2 pixel_9493/AMP_IN pixel_9493/SF_IB
+ pixel_9493/PIX_OUT pixel_9493/CSA_VREF pixel
Xpixel_8792 pixel_8792/gring pixel_8792/VDD pixel_8792/GND pixel_8792/VREF pixel_8792/ROW_SEL
+ pixel_8792/NB1 pixel_8792/VBIAS pixel_8792/NB2 pixel_8792/AMP_IN pixel_8792/SF_IB
+ pixel_8792/PIX_OUT pixel_8792/CSA_VREF pixel
Xpixel_6108 pixel_6108/gring pixel_6108/VDD pixel_6108/GND pixel_6108/VREF pixel_6108/ROW_SEL
+ pixel_6108/NB1 pixel_6108/VBIAS pixel_6108/NB2 pixel_6108/AMP_IN pixel_6108/SF_IB
+ pixel_6108/PIX_OUT pixel_6108/CSA_VREF pixel
Xpixel_6119 pixel_6119/gring pixel_6119/VDD pixel_6119/GND pixel_6119/VREF pixel_6119/ROW_SEL
+ pixel_6119/NB1 pixel_6119/VBIAS pixel_6119/NB2 pixel_6119/AMP_IN pixel_6119/SF_IB
+ pixel_6119/PIX_OUT pixel_6119/CSA_VREF pixel
Xpixel_5407 pixel_5407/gring pixel_5407/VDD pixel_5407/GND pixel_5407/VREF pixel_5407/ROW_SEL
+ pixel_5407/NB1 pixel_5407/VBIAS pixel_5407/NB2 pixel_5407/AMP_IN pixel_5407/SF_IB
+ pixel_5407/PIX_OUT pixel_5407/CSA_VREF pixel
Xpixel_5418 pixel_5418/gring pixel_5418/VDD pixel_5418/GND pixel_5418/VREF pixel_5418/ROW_SEL
+ pixel_5418/NB1 pixel_5418/VBIAS pixel_5418/NB2 pixel_5418/AMP_IN pixel_5418/SF_IB
+ pixel_5418/PIX_OUT pixel_5418/CSA_VREF pixel
Xpixel_5429 pixel_5429/gring pixel_5429/VDD pixel_5429/GND pixel_5429/VREF pixel_5429/ROW_SEL
+ pixel_5429/NB1 pixel_5429/VBIAS pixel_5429/NB2 pixel_5429/AMP_IN pixel_5429/SF_IB
+ pixel_5429/PIX_OUT pixel_5429/CSA_VREF pixel
Xpixel_723 pixel_723/gring pixel_723/VDD pixel_723/GND pixel_723/VREF pixel_723/ROW_SEL
+ pixel_723/NB1 pixel_723/VBIAS pixel_723/NB2 pixel_723/AMP_IN pixel_723/SF_IB pixel_723/PIX_OUT
+ pixel_723/CSA_VREF pixel
Xpixel_712 pixel_712/gring pixel_712/VDD pixel_712/GND pixel_712/VREF pixel_712/ROW_SEL
+ pixel_712/NB1 pixel_712/VBIAS pixel_712/NB2 pixel_712/AMP_IN pixel_712/SF_IB pixel_712/PIX_OUT
+ pixel_712/CSA_VREF pixel
Xpixel_701 pixel_701/gring pixel_701/VDD pixel_701/GND pixel_701/VREF pixel_701/ROW_SEL
+ pixel_701/NB1 pixel_701/VBIAS pixel_701/NB2 pixel_701/AMP_IN pixel_701/SF_IB pixel_701/PIX_OUT
+ pixel_701/CSA_VREF pixel
Xpixel_4706 pixel_4706/gring pixel_4706/VDD pixel_4706/GND pixel_4706/VREF pixel_4706/ROW_SEL
+ pixel_4706/NB1 pixel_4706/VBIAS pixel_4706/NB2 pixel_4706/AMP_IN pixel_4706/SF_IB
+ pixel_4706/PIX_OUT pixel_4706/CSA_VREF pixel
Xpixel_4717 pixel_4717/gring pixel_4717/VDD pixel_4717/GND pixel_4717/VREF pixel_4717/ROW_SEL
+ pixel_4717/NB1 pixel_4717/VBIAS pixel_4717/NB2 pixel_4717/AMP_IN pixel_4717/SF_IB
+ pixel_4717/PIX_OUT pixel_4717/CSA_VREF pixel
Xpixel_4728 pixel_4728/gring pixel_4728/VDD pixel_4728/GND pixel_4728/VREF pixel_4728/ROW_SEL
+ pixel_4728/NB1 pixel_4728/VBIAS pixel_4728/NB2 pixel_4728/AMP_IN pixel_4728/SF_IB
+ pixel_4728/PIX_OUT pixel_4728/CSA_VREF pixel
Xpixel_756 pixel_756/gring pixel_756/VDD pixel_756/GND pixel_756/VREF pixel_756/ROW_SEL
+ pixel_756/NB1 pixel_756/VBIAS pixel_756/NB2 pixel_756/AMP_IN pixel_756/SF_IB pixel_756/PIX_OUT
+ pixel_756/CSA_VREF pixel
Xpixel_745 pixel_745/gring pixel_745/VDD pixel_745/GND pixel_745/VREF pixel_745/ROW_SEL
+ pixel_745/NB1 pixel_745/VBIAS pixel_745/NB2 pixel_745/AMP_IN pixel_745/SF_IB pixel_745/PIX_OUT
+ pixel_745/CSA_VREF pixel
Xpixel_734 pixel_734/gring pixel_734/VDD pixel_734/GND pixel_734/VREF pixel_734/ROW_SEL
+ pixel_734/NB1 pixel_734/VBIAS pixel_734/NB2 pixel_734/AMP_IN pixel_734/SF_IB pixel_734/PIX_OUT
+ pixel_734/CSA_VREF pixel
Xpixel_4739 pixel_4739/gring pixel_4739/VDD pixel_4739/GND pixel_4739/VREF pixel_4739/ROW_SEL
+ pixel_4739/NB1 pixel_4739/VBIAS pixel_4739/NB2 pixel_4739/AMP_IN pixel_4739/SF_IB
+ pixel_4739/PIX_OUT pixel_4739/CSA_VREF pixel
Xpixel_789 pixel_789/gring pixel_789/VDD pixel_789/GND pixel_789/VREF pixel_789/ROW_SEL
+ pixel_789/NB1 pixel_789/VBIAS pixel_789/NB2 pixel_789/AMP_IN pixel_789/SF_IB pixel_789/PIX_OUT
+ pixel_789/CSA_VREF pixel
Xpixel_778 pixel_778/gring pixel_778/VDD pixel_778/GND pixel_778/VREF pixel_778/ROW_SEL
+ pixel_778/NB1 pixel_778/VBIAS pixel_778/NB2 pixel_778/AMP_IN pixel_778/SF_IB pixel_778/PIX_OUT
+ pixel_778/CSA_VREF pixel
Xpixel_767 pixel_767/gring pixel_767/VDD pixel_767/GND pixel_767/VREF pixel_767/ROW_SEL
+ pixel_767/NB1 pixel_767/VBIAS pixel_767/NB2 pixel_767/AMP_IN pixel_767/SF_IB pixel_767/PIX_OUT
+ pixel_767/CSA_VREF pixel
Xpixel_8000 pixel_8000/gring pixel_8000/VDD pixel_8000/GND pixel_8000/VREF pixel_8000/ROW_SEL
+ pixel_8000/NB1 pixel_8000/VBIAS pixel_8000/NB2 pixel_8000/AMP_IN pixel_8000/SF_IB
+ pixel_8000/PIX_OUT pixel_8000/CSA_VREF pixel
Xpixel_8011 pixel_8011/gring pixel_8011/VDD pixel_8011/GND pixel_8011/VREF pixel_8011/ROW_SEL
+ pixel_8011/NB1 pixel_8011/VBIAS pixel_8011/NB2 pixel_8011/AMP_IN pixel_8011/SF_IB
+ pixel_8011/PIX_OUT pixel_8011/CSA_VREF pixel
Xpixel_8022 pixel_8022/gring pixel_8022/VDD pixel_8022/GND pixel_8022/VREF pixel_8022/ROW_SEL
+ pixel_8022/NB1 pixel_8022/VBIAS pixel_8022/NB2 pixel_8022/AMP_IN pixel_8022/SF_IB
+ pixel_8022/PIX_OUT pixel_8022/CSA_VREF pixel
Xpixel_8033 pixel_8033/gring pixel_8033/VDD pixel_8033/GND pixel_8033/VREF pixel_8033/ROW_SEL
+ pixel_8033/NB1 pixel_8033/VBIAS pixel_8033/NB2 pixel_8033/AMP_IN pixel_8033/SF_IB
+ pixel_8033/PIX_OUT pixel_8033/CSA_VREF pixel
Xpixel_8044 pixel_8044/gring pixel_8044/VDD pixel_8044/GND pixel_8044/VREF pixel_8044/ROW_SEL
+ pixel_8044/NB1 pixel_8044/VBIAS pixel_8044/NB2 pixel_8044/AMP_IN pixel_8044/SF_IB
+ pixel_8044/PIX_OUT pixel_8044/CSA_VREF pixel
Xpixel_8055 pixel_8055/gring pixel_8055/VDD pixel_8055/GND pixel_8055/VREF pixel_8055/ROW_SEL
+ pixel_8055/NB1 pixel_8055/VBIAS pixel_8055/NB2 pixel_8055/AMP_IN pixel_8055/SF_IB
+ pixel_8055/PIX_OUT pixel_8055/CSA_VREF pixel
Xpixel_8066 pixel_8066/gring pixel_8066/VDD pixel_8066/GND pixel_8066/VREF pixel_8066/ROW_SEL
+ pixel_8066/NB1 pixel_8066/VBIAS pixel_8066/NB2 pixel_8066/AMP_IN pixel_8066/SF_IB
+ pixel_8066/PIX_OUT pixel_8066/CSA_VREF pixel
Xpixel_8077 pixel_8077/gring pixel_8077/VDD pixel_8077/GND pixel_8077/VREF pixel_8077/ROW_SEL
+ pixel_8077/NB1 pixel_8077/VBIAS pixel_8077/NB2 pixel_8077/AMP_IN pixel_8077/SF_IB
+ pixel_8077/PIX_OUT pixel_8077/CSA_VREF pixel
Xpixel_7310 pixel_7310/gring pixel_7310/VDD pixel_7310/GND pixel_7310/VREF pixel_7310/ROW_SEL
+ pixel_7310/NB1 pixel_7310/VBIAS pixel_7310/NB2 pixel_7310/AMP_IN pixel_7310/SF_IB
+ pixel_7310/PIX_OUT pixel_7310/CSA_VREF pixel
Xpixel_7321 pixel_7321/gring pixel_7321/VDD pixel_7321/GND pixel_7321/VREF pixel_7321/ROW_SEL
+ pixel_7321/NB1 pixel_7321/VBIAS pixel_7321/NB2 pixel_7321/AMP_IN pixel_7321/SF_IB
+ pixel_7321/PIX_OUT pixel_7321/CSA_VREF pixel
Xpixel_7332 pixel_7332/gring pixel_7332/VDD pixel_7332/GND pixel_7332/VREF pixel_7332/ROW_SEL
+ pixel_7332/NB1 pixel_7332/VBIAS pixel_7332/NB2 pixel_7332/AMP_IN pixel_7332/SF_IB
+ pixel_7332/PIX_OUT pixel_7332/CSA_VREF pixel
Xpixel_8088 pixel_8088/gring pixel_8088/VDD pixel_8088/GND pixel_8088/VREF pixel_8088/ROW_SEL
+ pixel_8088/NB1 pixel_8088/VBIAS pixel_8088/NB2 pixel_8088/AMP_IN pixel_8088/SF_IB
+ pixel_8088/PIX_OUT pixel_8088/CSA_VREF pixel
Xpixel_8099 pixel_8099/gring pixel_8099/VDD pixel_8099/GND pixel_8099/VREF pixel_8099/ROW_SEL
+ pixel_8099/NB1 pixel_8099/VBIAS pixel_8099/NB2 pixel_8099/AMP_IN pixel_8099/SF_IB
+ pixel_8099/PIX_OUT pixel_8099/CSA_VREF pixel
Xpixel_7343 pixel_7343/gring pixel_7343/VDD pixel_7343/GND pixel_7343/VREF pixel_7343/ROW_SEL
+ pixel_7343/NB1 pixel_7343/VBIAS pixel_7343/NB2 pixel_7343/AMP_IN pixel_7343/SF_IB
+ pixel_7343/PIX_OUT pixel_7343/CSA_VREF pixel
Xpixel_7354 pixel_7354/gring pixel_7354/VDD pixel_7354/GND pixel_7354/VREF pixel_7354/ROW_SEL
+ pixel_7354/NB1 pixel_7354/VBIAS pixel_7354/NB2 pixel_7354/AMP_IN pixel_7354/SF_IB
+ pixel_7354/PIX_OUT pixel_7354/CSA_VREF pixel
Xpixel_7365 pixel_7365/gring pixel_7365/VDD pixel_7365/GND pixel_7365/VREF pixel_7365/ROW_SEL
+ pixel_7365/NB1 pixel_7365/VBIAS pixel_7365/NB2 pixel_7365/AMP_IN pixel_7365/SF_IB
+ pixel_7365/PIX_OUT pixel_7365/CSA_VREF pixel
Xpixel_6620 pixel_6620/gring pixel_6620/VDD pixel_6620/GND pixel_6620/VREF pixel_6620/ROW_SEL
+ pixel_6620/NB1 pixel_6620/VBIAS pixel_6620/NB2 pixel_6620/AMP_IN pixel_6620/SF_IB
+ pixel_6620/PIX_OUT pixel_6620/CSA_VREF pixel
Xpixel_7376 pixel_7376/gring pixel_7376/VDD pixel_7376/GND pixel_7376/VREF pixel_7376/ROW_SEL
+ pixel_7376/NB1 pixel_7376/VBIAS pixel_7376/NB2 pixel_7376/AMP_IN pixel_7376/SF_IB
+ pixel_7376/PIX_OUT pixel_7376/CSA_VREF pixel
Xpixel_7387 pixel_7387/gring pixel_7387/VDD pixel_7387/GND pixel_7387/VREF pixel_7387/ROW_SEL
+ pixel_7387/NB1 pixel_7387/VBIAS pixel_7387/NB2 pixel_7387/AMP_IN pixel_7387/SF_IB
+ pixel_7387/PIX_OUT pixel_7387/CSA_VREF pixel
Xpixel_7398 pixel_7398/gring pixel_7398/VDD pixel_7398/GND pixel_7398/VREF pixel_7398/ROW_SEL
+ pixel_7398/NB1 pixel_7398/VBIAS pixel_7398/NB2 pixel_7398/AMP_IN pixel_7398/SF_IB
+ pixel_7398/PIX_OUT pixel_7398/CSA_VREF pixel
Xpixel_6631 pixel_6631/gring pixel_6631/VDD pixel_6631/GND pixel_6631/VREF pixel_6631/ROW_SEL
+ pixel_6631/NB1 pixel_6631/VBIAS pixel_6631/NB2 pixel_6631/AMP_IN pixel_6631/SF_IB
+ pixel_6631/PIX_OUT pixel_6631/CSA_VREF pixel
Xpixel_6642 pixel_6642/gring pixel_6642/VDD pixel_6642/GND pixel_6642/VREF pixel_6642/ROW_SEL
+ pixel_6642/NB1 pixel_6642/VBIAS pixel_6642/NB2 pixel_6642/AMP_IN pixel_6642/SF_IB
+ pixel_6642/PIX_OUT pixel_6642/CSA_VREF pixel
Xpixel_6653 pixel_6653/gring pixel_6653/VDD pixel_6653/GND pixel_6653/VREF pixel_6653/ROW_SEL
+ pixel_6653/NB1 pixel_6653/VBIAS pixel_6653/NB2 pixel_6653/AMP_IN pixel_6653/SF_IB
+ pixel_6653/PIX_OUT pixel_6653/CSA_VREF pixel
Xpixel_6664 pixel_6664/gring pixel_6664/VDD pixel_6664/GND pixel_6664/VREF pixel_6664/ROW_SEL
+ pixel_6664/NB1 pixel_6664/VBIAS pixel_6664/NB2 pixel_6664/AMP_IN pixel_6664/SF_IB
+ pixel_6664/PIX_OUT pixel_6664/CSA_VREF pixel
Xpixel_6675 pixel_6675/gring pixel_6675/VDD pixel_6675/GND pixel_6675/VREF pixel_6675/ROW_SEL
+ pixel_6675/NB1 pixel_6675/VBIAS pixel_6675/NB2 pixel_6675/AMP_IN pixel_6675/SF_IB
+ pixel_6675/PIX_OUT pixel_6675/CSA_VREF pixel
Xpixel_6686 pixel_6686/gring pixel_6686/VDD pixel_6686/GND pixel_6686/VREF pixel_6686/ROW_SEL
+ pixel_6686/NB1 pixel_6686/VBIAS pixel_6686/NB2 pixel_6686/AMP_IN pixel_6686/SF_IB
+ pixel_6686/PIX_OUT pixel_6686/CSA_VREF pixel
Xpixel_6697 pixel_6697/gring pixel_6697/VDD pixel_6697/GND pixel_6697/VREF pixel_6697/ROW_SEL
+ pixel_6697/NB1 pixel_6697/VBIAS pixel_6697/NB2 pixel_6697/AMP_IN pixel_6697/SF_IB
+ pixel_6697/PIX_OUT pixel_6697/CSA_VREF pixel
Xpixel_5930 pixel_5930/gring pixel_5930/VDD pixel_5930/GND pixel_5930/VREF pixel_5930/ROW_SEL
+ pixel_5930/NB1 pixel_5930/VBIAS pixel_5930/NB2 pixel_5930/AMP_IN pixel_5930/SF_IB
+ pixel_5930/PIX_OUT pixel_5930/CSA_VREF pixel
Xpixel_5941 pixel_5941/gring pixel_5941/VDD pixel_5941/GND pixel_5941/VREF pixel_5941/ROW_SEL
+ pixel_5941/NB1 pixel_5941/VBIAS pixel_5941/NB2 pixel_5941/AMP_IN pixel_5941/SF_IB
+ pixel_5941/PIX_OUT pixel_5941/CSA_VREF pixel
Xpixel_5952 pixel_5952/gring pixel_5952/VDD pixel_5952/GND pixel_5952/VREF pixel_5952/ROW_SEL
+ pixel_5952/NB1 pixel_5952/VBIAS pixel_5952/NB2 pixel_5952/AMP_IN pixel_5952/SF_IB
+ pixel_5952/PIX_OUT pixel_5952/CSA_VREF pixel
Xpixel_5963 pixel_5963/gring pixel_5963/VDD pixel_5963/GND pixel_5963/VREF pixel_5963/ROW_SEL
+ pixel_5963/NB1 pixel_5963/VBIAS pixel_5963/NB2 pixel_5963/AMP_IN pixel_5963/SF_IB
+ pixel_5963/PIX_OUT pixel_5963/CSA_VREF pixel
Xpixel_5974 pixel_5974/gring pixel_5974/VDD pixel_5974/GND pixel_5974/VREF pixel_5974/ROW_SEL
+ pixel_5974/NB1 pixel_5974/VBIAS pixel_5974/NB2 pixel_5974/AMP_IN pixel_5974/SF_IB
+ pixel_5974/PIX_OUT pixel_5974/CSA_VREF pixel
Xpixel_5985 pixel_5985/gring pixel_5985/VDD pixel_5985/GND pixel_5985/VREF pixel_5985/ROW_SEL
+ pixel_5985/NB1 pixel_5985/VBIAS pixel_5985/NB2 pixel_5985/AMP_IN pixel_5985/SF_IB
+ pixel_5985/PIX_OUT pixel_5985/CSA_VREF pixel
Xpixel_5996 pixel_5996/gring pixel_5996/VDD pixel_5996/GND pixel_5996/VREF pixel_5996/ROW_SEL
+ pixel_5996/NB1 pixel_5996/VBIAS pixel_5996/NB2 pixel_5996/AMP_IN pixel_5996/SF_IB
+ pixel_5996/PIX_OUT pixel_5996/CSA_VREF pixel
Xpixel_9290 pixel_9290/gring pixel_9290/VDD pixel_9290/GND pixel_9290/VREF pixel_9290/ROW_SEL
+ pixel_9290/NB1 pixel_9290/VBIAS pixel_9290/NB2 pixel_9290/AMP_IN pixel_9290/SF_IB
+ pixel_9290/PIX_OUT pixel_9290/CSA_VREF pixel
Xpixel_5204 pixel_5204/gring pixel_5204/VDD pixel_5204/GND pixel_5204/VREF pixel_5204/ROW_SEL
+ pixel_5204/NB1 pixel_5204/VBIAS pixel_5204/NB2 pixel_5204/AMP_IN pixel_5204/SF_IB
+ pixel_5204/PIX_OUT pixel_5204/CSA_VREF pixel
Xpixel_5215 pixel_5215/gring pixel_5215/VDD pixel_5215/GND pixel_5215/VREF pixel_5215/ROW_SEL
+ pixel_5215/NB1 pixel_5215/VBIAS pixel_5215/NB2 pixel_5215/AMP_IN pixel_5215/SF_IB
+ pixel_5215/PIX_OUT pixel_5215/CSA_VREF pixel
Xpixel_5226 pixel_5226/gring pixel_5226/VDD pixel_5226/GND pixel_5226/VREF pixel_5226/ROW_SEL
+ pixel_5226/NB1 pixel_5226/VBIAS pixel_5226/NB2 pixel_5226/AMP_IN pixel_5226/SF_IB
+ pixel_5226/PIX_OUT pixel_5226/CSA_VREF pixel
Xpixel_5237 pixel_5237/gring pixel_5237/VDD pixel_5237/GND pixel_5237/VREF pixel_5237/ROW_SEL
+ pixel_5237/NB1 pixel_5237/VBIAS pixel_5237/NB2 pixel_5237/AMP_IN pixel_5237/SF_IB
+ pixel_5237/PIX_OUT pixel_5237/CSA_VREF pixel
Xpixel_5248 pixel_5248/gring pixel_5248/VDD pixel_5248/GND pixel_5248/VREF pixel_5248/ROW_SEL
+ pixel_5248/NB1 pixel_5248/VBIAS pixel_5248/NB2 pixel_5248/AMP_IN pixel_5248/SF_IB
+ pixel_5248/PIX_OUT pixel_5248/CSA_VREF pixel
Xpixel_4503 pixel_4503/gring pixel_4503/VDD pixel_4503/GND pixel_4503/VREF pixel_4503/ROW_SEL
+ pixel_4503/NB1 pixel_4503/VBIAS pixel_4503/NB2 pixel_4503/AMP_IN pixel_4503/SF_IB
+ pixel_4503/PIX_OUT pixel_4503/CSA_VREF pixel
Xpixel_531 pixel_531/gring pixel_531/VDD pixel_531/GND pixel_531/VREF pixel_531/ROW_SEL
+ pixel_531/NB1 pixel_531/VBIAS pixel_531/NB2 pixel_531/AMP_IN pixel_531/SF_IB pixel_531/PIX_OUT
+ pixel_531/CSA_VREF pixel
Xpixel_520 pixel_520/gring pixel_520/VDD pixel_520/GND pixel_520/VREF pixel_520/ROW_SEL
+ pixel_520/NB1 pixel_520/VBIAS pixel_520/NB2 pixel_520/AMP_IN pixel_520/SF_IB pixel_520/PIX_OUT
+ pixel_520/CSA_VREF pixel
Xpixel_5259 pixel_5259/gring pixel_5259/VDD pixel_5259/GND pixel_5259/VREF pixel_5259/ROW_SEL
+ pixel_5259/NB1 pixel_5259/VBIAS pixel_5259/NB2 pixel_5259/AMP_IN pixel_5259/SF_IB
+ pixel_5259/PIX_OUT pixel_5259/CSA_VREF pixel
Xpixel_4514 pixel_4514/gring pixel_4514/VDD pixel_4514/GND pixel_4514/VREF pixel_4514/ROW_SEL
+ pixel_4514/NB1 pixel_4514/VBIAS pixel_4514/NB2 pixel_4514/AMP_IN pixel_4514/SF_IB
+ pixel_4514/PIX_OUT pixel_4514/CSA_VREF pixel
Xpixel_4525 pixel_4525/gring pixel_4525/VDD pixel_4525/GND pixel_4525/VREF pixel_4525/ROW_SEL
+ pixel_4525/NB1 pixel_4525/VBIAS pixel_4525/NB2 pixel_4525/AMP_IN pixel_4525/SF_IB
+ pixel_4525/PIX_OUT pixel_4525/CSA_VREF pixel
Xpixel_4536 pixel_4536/gring pixel_4536/VDD pixel_4536/GND pixel_4536/VREF pixel_4536/ROW_SEL
+ pixel_4536/NB1 pixel_4536/VBIAS pixel_4536/NB2 pixel_4536/AMP_IN pixel_4536/SF_IB
+ pixel_4536/PIX_OUT pixel_4536/CSA_VREF pixel
Xpixel_575 pixel_575/gring pixel_575/VDD pixel_575/GND pixel_575/VREF pixel_575/ROW_SEL
+ pixel_575/NB1 pixel_575/VBIAS pixel_575/NB2 pixel_575/AMP_IN pixel_575/SF_IB pixel_575/PIX_OUT
+ pixel_575/CSA_VREF pixel
Xpixel_564 pixel_564/gring pixel_564/VDD pixel_564/GND pixel_564/VREF pixel_564/ROW_SEL
+ pixel_564/NB1 pixel_564/VBIAS pixel_564/NB2 pixel_564/AMP_IN pixel_564/SF_IB pixel_564/PIX_OUT
+ pixel_564/CSA_VREF pixel
Xpixel_553 pixel_553/gring pixel_553/VDD pixel_553/GND pixel_553/VREF pixel_553/ROW_SEL
+ pixel_553/NB1 pixel_553/VBIAS pixel_553/NB2 pixel_553/AMP_IN pixel_553/SF_IB pixel_553/PIX_OUT
+ pixel_553/CSA_VREF pixel
Xpixel_542 pixel_542/gring pixel_542/VDD pixel_542/GND pixel_542/VREF pixel_542/ROW_SEL
+ pixel_542/NB1 pixel_542/VBIAS pixel_542/NB2 pixel_542/AMP_IN pixel_542/SF_IB pixel_542/PIX_OUT
+ pixel_542/CSA_VREF pixel
Xpixel_4547 pixel_4547/gring pixel_4547/VDD pixel_4547/GND pixel_4547/VREF pixel_4547/ROW_SEL
+ pixel_4547/NB1 pixel_4547/VBIAS pixel_4547/NB2 pixel_4547/AMP_IN pixel_4547/SF_IB
+ pixel_4547/PIX_OUT pixel_4547/CSA_VREF pixel
Xpixel_4558 pixel_4558/gring pixel_4558/VDD pixel_4558/GND pixel_4558/VREF pixel_4558/ROW_SEL
+ pixel_4558/NB1 pixel_4558/VBIAS pixel_4558/NB2 pixel_4558/AMP_IN pixel_4558/SF_IB
+ pixel_4558/PIX_OUT pixel_4558/CSA_VREF pixel
Xpixel_4569 pixel_4569/gring pixel_4569/VDD pixel_4569/GND pixel_4569/VREF pixel_4569/ROW_SEL
+ pixel_4569/NB1 pixel_4569/VBIAS pixel_4569/NB2 pixel_4569/AMP_IN pixel_4569/SF_IB
+ pixel_4569/PIX_OUT pixel_4569/CSA_VREF pixel
Xpixel_3802 pixel_3802/gring pixel_3802/VDD pixel_3802/GND pixel_3802/VREF pixel_3802/ROW_SEL
+ pixel_3802/NB1 pixel_3802/VBIAS pixel_3802/NB2 pixel_3802/AMP_IN pixel_3802/SF_IB
+ pixel_3802/PIX_OUT pixel_3802/CSA_VREF pixel
Xpixel_3813 pixel_3813/gring pixel_3813/VDD pixel_3813/GND pixel_3813/VREF pixel_3813/ROW_SEL
+ pixel_3813/NB1 pixel_3813/VBIAS pixel_3813/NB2 pixel_3813/AMP_IN pixel_3813/SF_IB
+ pixel_3813/PIX_OUT pixel_3813/CSA_VREF pixel
Xpixel_3824 pixel_3824/gring pixel_3824/VDD pixel_3824/GND pixel_3824/VREF pixel_3824/ROW_SEL
+ pixel_3824/NB1 pixel_3824/VBIAS pixel_3824/NB2 pixel_3824/AMP_IN pixel_3824/SF_IB
+ pixel_3824/PIX_OUT pixel_3824/CSA_VREF pixel
Xpixel_597 pixel_597/gring pixel_597/VDD pixel_597/GND pixel_597/VREF pixel_597/ROW_SEL
+ pixel_597/NB1 pixel_597/VBIAS pixel_597/NB2 pixel_597/AMP_IN pixel_597/SF_IB pixel_597/PIX_OUT
+ pixel_597/CSA_VREF pixel
Xpixel_586 pixel_586/gring pixel_586/VDD pixel_586/GND pixel_586/VREF pixel_586/ROW_SEL
+ pixel_586/NB1 pixel_586/VBIAS pixel_586/NB2 pixel_586/AMP_IN pixel_586/SF_IB pixel_586/PIX_OUT
+ pixel_586/CSA_VREF pixel
Xpixel_3868 pixel_3868/gring pixel_3868/VDD pixel_3868/GND pixel_3868/VREF pixel_3868/ROW_SEL
+ pixel_3868/NB1 pixel_3868/VBIAS pixel_3868/NB2 pixel_3868/AMP_IN pixel_3868/SF_IB
+ pixel_3868/PIX_OUT pixel_3868/CSA_VREF pixel
Xpixel_3857 pixel_3857/gring pixel_3857/VDD pixel_3857/GND pixel_3857/VREF pixel_3857/ROW_SEL
+ pixel_3857/NB1 pixel_3857/VBIAS pixel_3857/NB2 pixel_3857/AMP_IN pixel_3857/SF_IB
+ pixel_3857/PIX_OUT pixel_3857/CSA_VREF pixel
Xpixel_3846 pixel_3846/gring pixel_3846/VDD pixel_3846/GND pixel_3846/VREF pixel_3846/ROW_SEL
+ pixel_3846/NB1 pixel_3846/VBIAS pixel_3846/NB2 pixel_3846/AMP_IN pixel_3846/SF_IB
+ pixel_3846/PIX_OUT pixel_3846/CSA_VREF pixel
Xpixel_3835 pixel_3835/gring pixel_3835/VDD pixel_3835/GND pixel_3835/VREF pixel_3835/ROW_SEL
+ pixel_3835/NB1 pixel_3835/VBIAS pixel_3835/NB2 pixel_3835/AMP_IN pixel_3835/SF_IB
+ pixel_3835/PIX_OUT pixel_3835/CSA_VREF pixel
Xpixel_3879 pixel_3879/gring pixel_3879/VDD pixel_3879/GND pixel_3879/VREF pixel_3879/ROW_SEL
+ pixel_3879/NB1 pixel_3879/VBIAS pixel_3879/NB2 pixel_3879/AMP_IN pixel_3879/SF_IB
+ pixel_3879/PIX_OUT pixel_3879/CSA_VREF pixel
Xpixel_7140 pixel_7140/gring pixel_7140/VDD pixel_7140/GND pixel_7140/VREF pixel_7140/ROW_SEL
+ pixel_7140/NB1 pixel_7140/VBIAS pixel_7140/NB2 pixel_7140/AMP_IN pixel_7140/SF_IB
+ pixel_7140/PIX_OUT pixel_7140/CSA_VREF pixel
Xpixel_7151 pixel_7151/gring pixel_7151/VDD pixel_7151/GND pixel_7151/VREF pixel_7151/ROW_SEL
+ pixel_7151/NB1 pixel_7151/VBIAS pixel_7151/NB2 pixel_7151/AMP_IN pixel_7151/SF_IB
+ pixel_7151/PIX_OUT pixel_7151/CSA_VREF pixel
Xpixel_7162 pixel_7162/gring pixel_7162/VDD pixel_7162/GND pixel_7162/VREF pixel_7162/ROW_SEL
+ pixel_7162/NB1 pixel_7162/VBIAS pixel_7162/NB2 pixel_7162/AMP_IN pixel_7162/SF_IB
+ pixel_7162/PIX_OUT pixel_7162/CSA_VREF pixel
Xpixel_7173 pixel_7173/gring pixel_7173/VDD pixel_7173/GND pixel_7173/VREF pixel_7173/ROW_SEL
+ pixel_7173/NB1 pixel_7173/VBIAS pixel_7173/NB2 pixel_7173/AMP_IN pixel_7173/SF_IB
+ pixel_7173/PIX_OUT pixel_7173/CSA_VREF pixel
Xpixel_7184 pixel_7184/gring pixel_7184/VDD pixel_7184/GND pixel_7184/VREF pixel_7184/ROW_SEL
+ pixel_7184/NB1 pixel_7184/VBIAS pixel_7184/NB2 pixel_7184/AMP_IN pixel_7184/SF_IB
+ pixel_7184/PIX_OUT pixel_7184/CSA_VREF pixel
Xpixel_7195 pixel_7195/gring pixel_7195/VDD pixel_7195/GND pixel_7195/VREF pixel_7195/ROW_SEL
+ pixel_7195/NB1 pixel_7195/VBIAS pixel_7195/NB2 pixel_7195/AMP_IN pixel_7195/SF_IB
+ pixel_7195/PIX_OUT pixel_7195/CSA_VREF pixel
Xpixel_6450 pixel_6450/gring pixel_6450/VDD pixel_6450/GND pixel_6450/VREF pixel_6450/ROW_SEL
+ pixel_6450/NB1 pixel_6450/VBIAS pixel_6450/NB2 pixel_6450/AMP_IN pixel_6450/SF_IB
+ pixel_6450/PIX_OUT pixel_6450/CSA_VREF pixel
Xpixel_6461 pixel_6461/gring pixel_6461/VDD pixel_6461/GND pixel_6461/VREF pixel_6461/ROW_SEL
+ pixel_6461/NB1 pixel_6461/VBIAS pixel_6461/NB2 pixel_6461/AMP_IN pixel_6461/SF_IB
+ pixel_6461/PIX_OUT pixel_6461/CSA_VREF pixel
Xpixel_6472 pixel_6472/gring pixel_6472/VDD pixel_6472/GND pixel_6472/VREF pixel_6472/ROW_SEL
+ pixel_6472/NB1 pixel_6472/VBIAS pixel_6472/NB2 pixel_6472/AMP_IN pixel_6472/SF_IB
+ pixel_6472/PIX_OUT pixel_6472/CSA_VREF pixel
Xpixel_6483 pixel_6483/gring pixel_6483/VDD pixel_6483/GND pixel_6483/VREF pixel_6483/ROW_SEL
+ pixel_6483/NB1 pixel_6483/VBIAS pixel_6483/NB2 pixel_6483/AMP_IN pixel_6483/SF_IB
+ pixel_6483/PIX_OUT pixel_6483/CSA_VREF pixel
Xpixel_6494 pixel_6494/gring pixel_6494/VDD pixel_6494/GND pixel_6494/VREF pixel_6494/ROW_SEL
+ pixel_6494/NB1 pixel_6494/VBIAS pixel_6494/NB2 pixel_6494/AMP_IN pixel_6494/SF_IB
+ pixel_6494/PIX_OUT pixel_6494/CSA_VREF pixel
Xpixel_5760 pixel_5760/gring pixel_5760/VDD pixel_5760/GND pixel_5760/VREF pixel_5760/ROW_SEL
+ pixel_5760/NB1 pixel_5760/VBIAS pixel_5760/NB2 pixel_5760/AMP_IN pixel_5760/SF_IB
+ pixel_5760/PIX_OUT pixel_5760/CSA_VREF pixel
Xpixel_5771 pixel_5771/gring pixel_5771/VDD pixel_5771/GND pixel_5771/VREF pixel_5771/ROW_SEL
+ pixel_5771/NB1 pixel_5771/VBIAS pixel_5771/NB2 pixel_5771/AMP_IN pixel_5771/SF_IB
+ pixel_5771/PIX_OUT pixel_5771/CSA_VREF pixel
Xpixel_5782 pixel_5782/gring pixel_5782/VDD pixel_5782/GND pixel_5782/VREF pixel_5782/ROW_SEL
+ pixel_5782/NB1 pixel_5782/VBIAS pixel_5782/NB2 pixel_5782/AMP_IN pixel_5782/SF_IB
+ pixel_5782/PIX_OUT pixel_5782/CSA_VREF pixel
Xpixel_5793 pixel_5793/gring pixel_5793/VDD pixel_5793/GND pixel_5793/VREF pixel_5793/ROW_SEL
+ pixel_5793/NB1 pixel_5793/VBIAS pixel_5793/NB2 pixel_5793/AMP_IN pixel_5793/SF_IB
+ pixel_5793/PIX_OUT pixel_5793/CSA_VREF pixel
Xpixel_3109 pixel_3109/gring pixel_3109/VDD pixel_3109/GND pixel_3109/VREF pixel_3109/ROW_SEL
+ pixel_3109/NB1 pixel_3109/VBIAS pixel_3109/NB2 pixel_3109/AMP_IN pixel_3109/SF_IB
+ pixel_3109/PIX_OUT pixel_3109/CSA_VREF pixel
Xpixel_2419 pixel_2419/gring pixel_2419/VDD pixel_2419/GND pixel_2419/VREF pixel_2419/ROW_SEL
+ pixel_2419/NB1 pixel_2419/VBIAS pixel_2419/NB2 pixel_2419/AMP_IN pixel_2419/SF_IB
+ pixel_2419/PIX_OUT pixel_2419/CSA_VREF pixel
Xpixel_2408 pixel_2408/gring pixel_2408/VDD pixel_2408/GND pixel_2408/VREF pixel_2408/ROW_SEL
+ pixel_2408/NB1 pixel_2408/VBIAS pixel_2408/NB2 pixel_2408/AMP_IN pixel_2408/SF_IB
+ pixel_2408/PIX_OUT pixel_2408/CSA_VREF pixel
Xpixel_1707 pixel_1707/gring pixel_1707/VDD pixel_1707/GND pixel_1707/VREF pixel_1707/ROW_SEL
+ pixel_1707/NB1 pixel_1707/VBIAS pixel_1707/NB2 pixel_1707/AMP_IN pixel_1707/SF_IB
+ pixel_1707/PIX_OUT pixel_1707/CSA_VREF pixel
Xpixel_1729 pixel_1729/gring pixel_1729/VDD pixel_1729/GND pixel_1729/VREF pixel_1729/ROW_SEL
+ pixel_1729/NB1 pixel_1729/VBIAS pixel_1729/NB2 pixel_1729/AMP_IN pixel_1729/SF_IB
+ pixel_1729/PIX_OUT pixel_1729/CSA_VREF pixel
Xpixel_1718 pixel_1718/gring pixel_1718/VDD pixel_1718/GND pixel_1718/VREF pixel_1718/ROW_SEL
+ pixel_1718/NB1 pixel_1718/VBIAS pixel_1718/NB2 pixel_1718/AMP_IN pixel_1718/SF_IB
+ pixel_1718/PIX_OUT pixel_1718/CSA_VREF pixel
Xpixel_5001 pixel_5001/gring pixel_5001/VDD pixel_5001/GND pixel_5001/VREF pixel_5001/ROW_SEL
+ pixel_5001/NB1 pixel_5001/VBIAS pixel_5001/NB2 pixel_5001/AMP_IN pixel_5001/SF_IB
+ pixel_5001/PIX_OUT pixel_5001/CSA_VREF pixel
Xpixel_5012 pixel_5012/gring pixel_5012/VDD pixel_5012/GND pixel_5012/VREF pixel_5012/ROW_SEL
+ pixel_5012/NB1 pixel_5012/VBIAS pixel_5012/NB2 pixel_5012/AMP_IN pixel_5012/SF_IB
+ pixel_5012/PIX_OUT pixel_5012/CSA_VREF pixel
Xpixel_5023 pixel_5023/gring pixel_5023/VDD pixel_5023/GND pixel_5023/VREF pixel_5023/ROW_SEL
+ pixel_5023/NB1 pixel_5023/VBIAS pixel_5023/NB2 pixel_5023/AMP_IN pixel_5023/SF_IB
+ pixel_5023/PIX_OUT pixel_5023/CSA_VREF pixel
Xpixel_5034 pixel_5034/gring pixel_5034/VDD pixel_5034/GND pixel_5034/VREF pixel_5034/ROW_SEL
+ pixel_5034/NB1 pixel_5034/VBIAS pixel_5034/NB2 pixel_5034/AMP_IN pixel_5034/SF_IB
+ pixel_5034/PIX_OUT pixel_5034/CSA_VREF pixel
Xpixel_5045 pixel_5045/gring pixel_5045/VDD pixel_5045/GND pixel_5045/VREF pixel_5045/ROW_SEL
+ pixel_5045/NB1 pixel_5045/VBIAS pixel_5045/NB2 pixel_5045/AMP_IN pixel_5045/SF_IB
+ pixel_5045/PIX_OUT pixel_5045/CSA_VREF pixel
Xpixel_5056 pixel_5056/gring pixel_5056/VDD pixel_5056/GND pixel_5056/VREF pixel_5056/ROW_SEL
+ pixel_5056/NB1 pixel_5056/VBIAS pixel_5056/NB2 pixel_5056/AMP_IN pixel_5056/SF_IB
+ pixel_5056/PIX_OUT pixel_5056/CSA_VREF pixel
Xpixel_4300 pixel_4300/gring pixel_4300/VDD pixel_4300/GND pixel_4300/VREF pixel_4300/ROW_SEL
+ pixel_4300/NB1 pixel_4300/VBIAS pixel_4300/NB2 pixel_4300/AMP_IN pixel_4300/SF_IB
+ pixel_4300/PIX_OUT pixel_4300/CSA_VREF pixel
Xpixel_4311 pixel_4311/gring pixel_4311/VDD pixel_4311/GND pixel_4311/VREF pixel_4311/ROW_SEL
+ pixel_4311/NB1 pixel_4311/VBIAS pixel_4311/NB2 pixel_4311/AMP_IN pixel_4311/SF_IB
+ pixel_4311/PIX_OUT pixel_4311/CSA_VREF pixel
Xpixel_5067 pixel_5067/gring pixel_5067/VDD pixel_5067/GND pixel_5067/VREF pixel_5067/ROW_SEL
+ pixel_5067/NB1 pixel_5067/VBIAS pixel_5067/NB2 pixel_5067/AMP_IN pixel_5067/SF_IB
+ pixel_5067/PIX_OUT pixel_5067/CSA_VREF pixel
Xpixel_5078 pixel_5078/gring pixel_5078/VDD pixel_5078/GND pixel_5078/VREF pixel_5078/ROW_SEL
+ pixel_5078/NB1 pixel_5078/VBIAS pixel_5078/NB2 pixel_5078/AMP_IN pixel_5078/SF_IB
+ pixel_5078/PIX_OUT pixel_5078/CSA_VREF pixel
Xpixel_5089 pixel_5089/gring pixel_5089/VDD pixel_5089/GND pixel_5089/VREF pixel_5089/ROW_SEL
+ pixel_5089/NB1 pixel_5089/VBIAS pixel_5089/NB2 pixel_5089/AMP_IN pixel_5089/SF_IB
+ pixel_5089/PIX_OUT pixel_5089/CSA_VREF pixel
Xpixel_4322 pixel_4322/gring pixel_4322/VDD pixel_4322/GND pixel_4322/VREF pixel_4322/ROW_SEL
+ pixel_4322/NB1 pixel_4322/VBIAS pixel_4322/NB2 pixel_4322/AMP_IN pixel_4322/SF_IB
+ pixel_4322/PIX_OUT pixel_4322/CSA_VREF pixel
Xpixel_4333 pixel_4333/gring pixel_4333/VDD pixel_4333/GND pixel_4333/VREF pixel_4333/ROW_SEL
+ pixel_4333/NB1 pixel_4333/VBIAS pixel_4333/NB2 pixel_4333/AMP_IN pixel_4333/SF_IB
+ pixel_4333/PIX_OUT pixel_4333/CSA_VREF pixel
Xpixel_4344 pixel_4344/gring pixel_4344/VDD pixel_4344/GND pixel_4344/VREF pixel_4344/ROW_SEL
+ pixel_4344/NB1 pixel_4344/VBIAS pixel_4344/NB2 pixel_4344/AMP_IN pixel_4344/SF_IB
+ pixel_4344/PIX_OUT pixel_4344/CSA_VREF pixel
Xpixel_383 pixel_383/gring pixel_383/VDD pixel_383/GND pixel_383/VREF pixel_383/ROW_SEL
+ pixel_383/NB1 pixel_383/VBIAS pixel_383/NB2 pixel_383/AMP_IN pixel_383/SF_IB pixel_383/PIX_OUT
+ pixel_383/CSA_VREF pixel
Xpixel_372 pixel_372/gring pixel_372/VDD pixel_372/GND pixel_372/VREF pixel_372/ROW_SEL
+ pixel_372/NB1 pixel_372/VBIAS pixel_372/NB2 pixel_372/AMP_IN pixel_372/SF_IB pixel_372/PIX_OUT
+ pixel_372/CSA_VREF pixel
Xpixel_361 pixel_361/gring pixel_361/VDD pixel_361/GND pixel_361/VREF pixel_361/ROW_SEL
+ pixel_361/NB1 pixel_361/VBIAS pixel_361/NB2 pixel_361/AMP_IN pixel_361/SF_IB pixel_361/PIX_OUT
+ pixel_361/CSA_VREF pixel
Xpixel_350 pixel_350/gring pixel_350/VDD pixel_350/GND pixel_350/VREF pixel_350/ROW_SEL
+ pixel_350/NB1 pixel_350/VBIAS pixel_350/NB2 pixel_350/AMP_IN pixel_350/SF_IB pixel_350/PIX_OUT
+ pixel_350/CSA_VREF pixel
Xpixel_3643 pixel_3643/gring pixel_3643/VDD pixel_3643/GND pixel_3643/VREF pixel_3643/ROW_SEL
+ pixel_3643/NB1 pixel_3643/VBIAS pixel_3643/NB2 pixel_3643/AMP_IN pixel_3643/SF_IB
+ pixel_3643/PIX_OUT pixel_3643/CSA_VREF pixel
Xpixel_3632 pixel_3632/gring pixel_3632/VDD pixel_3632/GND pixel_3632/VREF pixel_3632/ROW_SEL
+ pixel_3632/NB1 pixel_3632/VBIAS pixel_3632/NB2 pixel_3632/AMP_IN pixel_3632/SF_IB
+ pixel_3632/PIX_OUT pixel_3632/CSA_VREF pixel
Xpixel_3621 pixel_3621/gring pixel_3621/VDD pixel_3621/GND pixel_3621/VREF pixel_3621/ROW_SEL
+ pixel_3621/NB1 pixel_3621/VBIAS pixel_3621/NB2 pixel_3621/AMP_IN pixel_3621/SF_IB
+ pixel_3621/PIX_OUT pixel_3621/CSA_VREF pixel
Xpixel_3610 pixel_3610/gring pixel_3610/VDD pixel_3610/GND pixel_3610/VREF pixel_3610/ROW_SEL
+ pixel_3610/NB1 pixel_3610/VBIAS pixel_3610/NB2 pixel_3610/AMP_IN pixel_3610/SF_IB
+ pixel_3610/PIX_OUT pixel_3610/CSA_VREF pixel
Xpixel_4355 pixel_4355/gring pixel_4355/VDD pixel_4355/GND pixel_4355/VREF pixel_4355/ROW_SEL
+ pixel_4355/NB1 pixel_4355/VBIAS pixel_4355/NB2 pixel_4355/AMP_IN pixel_4355/SF_IB
+ pixel_4355/PIX_OUT pixel_4355/CSA_VREF pixel
Xpixel_4366 pixel_4366/gring pixel_4366/VDD pixel_4366/GND pixel_4366/VREF pixel_4366/ROW_SEL
+ pixel_4366/NB1 pixel_4366/VBIAS pixel_4366/NB2 pixel_4366/AMP_IN pixel_4366/SF_IB
+ pixel_4366/PIX_OUT pixel_4366/CSA_VREF pixel
Xpixel_4377 pixel_4377/gring pixel_4377/VDD pixel_4377/GND pixel_4377/VREF pixel_4377/ROW_SEL
+ pixel_4377/NB1 pixel_4377/VBIAS pixel_4377/NB2 pixel_4377/AMP_IN pixel_4377/SF_IB
+ pixel_4377/PIX_OUT pixel_4377/CSA_VREF pixel
Xpixel_4388 pixel_4388/gring pixel_4388/VDD pixel_4388/GND pixel_4388/VREF pixel_4388/ROW_SEL
+ pixel_4388/NB1 pixel_4388/VBIAS pixel_4388/NB2 pixel_4388/AMP_IN pixel_4388/SF_IB
+ pixel_4388/PIX_OUT pixel_4388/CSA_VREF pixel
Xpixel_394 pixel_394/gring pixel_394/VDD pixel_394/GND pixel_394/VREF pixel_394/ROW_SEL
+ pixel_394/NB1 pixel_394/VBIAS pixel_394/NB2 pixel_394/AMP_IN pixel_394/SF_IB pixel_394/PIX_OUT
+ pixel_394/CSA_VREF pixel
Xpixel_2931 pixel_2931/gring pixel_2931/VDD pixel_2931/GND pixel_2931/VREF pixel_2931/ROW_SEL
+ pixel_2931/NB1 pixel_2931/VBIAS pixel_2931/NB2 pixel_2931/AMP_IN pixel_2931/SF_IB
+ pixel_2931/PIX_OUT pixel_2931/CSA_VREF pixel
Xpixel_2920 pixel_2920/gring pixel_2920/VDD pixel_2920/GND pixel_2920/VREF pixel_2920/ROW_SEL
+ pixel_2920/NB1 pixel_2920/VBIAS pixel_2920/NB2 pixel_2920/AMP_IN pixel_2920/SF_IB
+ pixel_2920/PIX_OUT pixel_2920/CSA_VREF pixel
Xpixel_3676 pixel_3676/gring pixel_3676/VDD pixel_3676/GND pixel_3676/VREF pixel_3676/ROW_SEL
+ pixel_3676/NB1 pixel_3676/VBIAS pixel_3676/NB2 pixel_3676/AMP_IN pixel_3676/SF_IB
+ pixel_3676/PIX_OUT pixel_3676/CSA_VREF pixel
Xpixel_3665 pixel_3665/gring pixel_3665/VDD pixel_3665/GND pixel_3665/VREF pixel_3665/ROW_SEL
+ pixel_3665/NB1 pixel_3665/VBIAS pixel_3665/NB2 pixel_3665/AMP_IN pixel_3665/SF_IB
+ pixel_3665/PIX_OUT pixel_3665/CSA_VREF pixel
Xpixel_3654 pixel_3654/gring pixel_3654/VDD pixel_3654/GND pixel_3654/VREF pixel_3654/ROW_SEL
+ pixel_3654/NB1 pixel_3654/VBIAS pixel_3654/NB2 pixel_3654/AMP_IN pixel_3654/SF_IB
+ pixel_3654/PIX_OUT pixel_3654/CSA_VREF pixel
Xpixel_4399 pixel_4399/gring pixel_4399/VDD pixel_4399/GND pixel_4399/VREF pixel_4399/ROW_SEL
+ pixel_4399/NB1 pixel_4399/VBIAS pixel_4399/NB2 pixel_4399/AMP_IN pixel_4399/SF_IB
+ pixel_4399/PIX_OUT pixel_4399/CSA_VREF pixel
Xpixel_2964 pixel_2964/gring pixel_2964/VDD pixel_2964/GND pixel_2964/VREF pixel_2964/ROW_SEL
+ pixel_2964/NB1 pixel_2964/VBIAS pixel_2964/NB2 pixel_2964/AMP_IN pixel_2964/SF_IB
+ pixel_2964/PIX_OUT pixel_2964/CSA_VREF pixel
Xpixel_2953 pixel_2953/gring pixel_2953/VDD pixel_2953/GND pixel_2953/VREF pixel_2953/ROW_SEL
+ pixel_2953/NB1 pixel_2953/VBIAS pixel_2953/NB2 pixel_2953/AMP_IN pixel_2953/SF_IB
+ pixel_2953/PIX_OUT pixel_2953/CSA_VREF pixel
Xpixel_2942 pixel_2942/gring pixel_2942/VDD pixel_2942/GND pixel_2942/VREF pixel_2942/ROW_SEL
+ pixel_2942/NB1 pixel_2942/VBIAS pixel_2942/NB2 pixel_2942/AMP_IN pixel_2942/SF_IB
+ pixel_2942/PIX_OUT pixel_2942/CSA_VREF pixel
Xpixel_3698 pixel_3698/gring pixel_3698/VDD pixel_3698/GND pixel_3698/VREF pixel_3698/ROW_SEL
+ pixel_3698/NB1 pixel_3698/VBIAS pixel_3698/NB2 pixel_3698/AMP_IN pixel_3698/SF_IB
+ pixel_3698/PIX_OUT pixel_3698/CSA_VREF pixel
Xpixel_3687 pixel_3687/gring pixel_3687/VDD pixel_3687/GND pixel_3687/VREF pixel_3687/ROW_SEL
+ pixel_3687/NB1 pixel_3687/VBIAS pixel_3687/NB2 pixel_3687/AMP_IN pixel_3687/SF_IB
+ pixel_3687/PIX_OUT pixel_3687/CSA_VREF pixel
Xpixel_2997 pixel_2997/gring pixel_2997/VDD pixel_2997/GND pixel_2997/VREF pixel_2997/ROW_SEL
+ pixel_2997/NB1 pixel_2997/VBIAS pixel_2997/NB2 pixel_2997/AMP_IN pixel_2997/SF_IB
+ pixel_2997/PIX_OUT pixel_2997/CSA_VREF pixel
Xpixel_2986 pixel_2986/gring pixel_2986/VDD pixel_2986/GND pixel_2986/VREF pixel_2986/ROW_SEL
+ pixel_2986/NB1 pixel_2986/VBIAS pixel_2986/NB2 pixel_2986/AMP_IN pixel_2986/SF_IB
+ pixel_2986/PIX_OUT pixel_2986/CSA_VREF pixel
Xpixel_2975 pixel_2975/gring pixel_2975/VDD pixel_2975/GND pixel_2975/VREF pixel_2975/ROW_SEL
+ pixel_2975/NB1 pixel_2975/VBIAS pixel_2975/NB2 pixel_2975/AMP_IN pixel_2975/SF_IB
+ pixel_2975/PIX_OUT pixel_2975/CSA_VREF pixel
Xpixel_6280 pixel_6280/gring pixel_6280/VDD pixel_6280/GND pixel_6280/VREF pixel_6280/ROW_SEL
+ pixel_6280/NB1 pixel_6280/VBIAS pixel_6280/NB2 pixel_6280/AMP_IN pixel_6280/SF_IB
+ pixel_6280/PIX_OUT pixel_6280/CSA_VREF pixel
Xpixel_6291 pixel_6291/gring pixel_6291/VDD pixel_6291/GND pixel_6291/VREF pixel_6291/ROW_SEL
+ pixel_6291/NB1 pixel_6291/VBIAS pixel_6291/NB2 pixel_6291/AMP_IN pixel_6291/SF_IB
+ pixel_6291/PIX_OUT pixel_6291/CSA_VREF pixel
Xpixel_5590 pixel_5590/gring pixel_5590/VDD pixel_5590/GND pixel_5590/VREF pixel_5590/ROW_SEL
+ pixel_5590/NB1 pixel_5590/VBIAS pixel_5590/NB2 pixel_5590/AMP_IN pixel_5590/SF_IB
+ pixel_5590/PIX_OUT pixel_5590/CSA_VREF pixel
Xpixel_7909 pixel_7909/gring pixel_7909/VDD pixel_7909/GND pixel_7909/VREF pixel_7909/ROW_SEL
+ pixel_7909/NB1 pixel_7909/VBIAS pixel_7909/NB2 pixel_7909/AMP_IN pixel_7909/SF_IB
+ pixel_7909/PIX_OUT pixel_7909/CSA_VREF pixel
Xpixel_2227 pixel_2227/gring pixel_2227/VDD pixel_2227/GND pixel_2227/VREF pixel_2227/ROW_SEL
+ pixel_2227/NB1 pixel_2227/VBIAS pixel_2227/NB2 pixel_2227/AMP_IN pixel_2227/SF_IB
+ pixel_2227/PIX_OUT pixel_2227/CSA_VREF pixel
Xpixel_2216 pixel_2216/gring pixel_2216/VDD pixel_2216/GND pixel_2216/VREF pixel_2216/ROW_SEL
+ pixel_2216/NB1 pixel_2216/VBIAS pixel_2216/NB2 pixel_2216/AMP_IN pixel_2216/SF_IB
+ pixel_2216/PIX_OUT pixel_2216/CSA_VREF pixel
Xpixel_2205 pixel_2205/gring pixel_2205/VDD pixel_2205/GND pixel_2205/VREF pixel_2205/ROW_SEL
+ pixel_2205/NB1 pixel_2205/VBIAS pixel_2205/NB2 pixel_2205/AMP_IN pixel_2205/SF_IB
+ pixel_2205/PIX_OUT pixel_2205/CSA_VREF pixel
Xpixel_1515 pixel_1515/gring pixel_1515/VDD pixel_1515/GND pixel_1515/VREF pixel_1515/ROW_SEL
+ pixel_1515/NB1 pixel_1515/VBIAS pixel_1515/NB2 pixel_1515/AMP_IN pixel_1515/SF_IB
+ pixel_1515/PIX_OUT pixel_1515/CSA_VREF pixel
Xpixel_1504 pixel_1504/gring pixel_1504/VDD pixel_1504/GND pixel_1504/VREF pixel_1504/ROW_SEL
+ pixel_1504/NB1 pixel_1504/VBIAS pixel_1504/NB2 pixel_1504/AMP_IN pixel_1504/SF_IB
+ pixel_1504/PIX_OUT pixel_1504/CSA_VREF pixel
Xpixel_2249 pixel_2249/gring pixel_2249/VDD pixel_2249/GND pixel_2249/VREF pixel_2249/ROW_SEL
+ pixel_2249/NB1 pixel_2249/VBIAS pixel_2249/NB2 pixel_2249/AMP_IN pixel_2249/SF_IB
+ pixel_2249/PIX_OUT pixel_2249/CSA_VREF pixel
Xpixel_2238 pixel_2238/gring pixel_2238/VDD pixel_2238/GND pixel_2238/VREF pixel_2238/ROW_SEL
+ pixel_2238/NB1 pixel_2238/VBIAS pixel_2238/NB2 pixel_2238/AMP_IN pixel_2238/SF_IB
+ pixel_2238/PIX_OUT pixel_2238/CSA_VREF pixel
Xpixel_1559 pixel_1559/gring pixel_1559/VDD pixel_1559/GND pixel_1559/VREF pixel_1559/ROW_SEL
+ pixel_1559/NB1 pixel_1559/VBIAS pixel_1559/NB2 pixel_1559/AMP_IN pixel_1559/SF_IB
+ pixel_1559/PIX_OUT pixel_1559/CSA_VREF pixel
Xpixel_1548 pixel_1548/gring pixel_1548/VDD pixel_1548/GND pixel_1548/VREF pixel_1548/ROW_SEL
+ pixel_1548/NB1 pixel_1548/VBIAS pixel_1548/NB2 pixel_1548/AMP_IN pixel_1548/SF_IB
+ pixel_1548/PIX_OUT pixel_1548/CSA_VREF pixel
Xpixel_1537 pixel_1537/gring pixel_1537/VDD pixel_1537/GND pixel_1537/VREF pixel_1537/ROW_SEL
+ pixel_1537/NB1 pixel_1537/VBIAS pixel_1537/NB2 pixel_1537/AMP_IN pixel_1537/SF_IB
+ pixel_1537/PIX_OUT pixel_1537/CSA_VREF pixel
Xpixel_1526 pixel_1526/gring pixel_1526/VDD pixel_1526/GND pixel_1526/VREF pixel_1526/ROW_SEL
+ pixel_1526/NB1 pixel_1526/VBIAS pixel_1526/NB2 pixel_1526/AMP_IN pixel_1526/SF_IB
+ pixel_1526/PIX_OUT pixel_1526/CSA_VREF pixel
Xpixel_9823 pixel_9823/gring pixel_9823/VDD pixel_9823/GND pixel_9823/VREF pixel_9823/ROW_SEL
+ pixel_9823/NB1 pixel_9823/VBIAS pixel_9823/NB2 pixel_9823/AMP_IN pixel_9823/SF_IB
+ pixel_9823/PIX_OUT pixel_9823/CSA_VREF pixel
Xpixel_9812 pixel_9812/gring pixel_9812/VDD pixel_9812/GND pixel_9812/VREF pixel_9812/ROW_SEL
+ pixel_9812/NB1 pixel_9812/VBIAS pixel_9812/NB2 pixel_9812/AMP_IN pixel_9812/SF_IB
+ pixel_9812/PIX_OUT pixel_9812/CSA_VREF pixel
Xpixel_9801 pixel_9801/gring pixel_9801/VDD pixel_9801/GND pixel_9801/VREF pixel_9801/ROW_SEL
+ pixel_9801/NB1 pixel_9801/VBIAS pixel_9801/NB2 pixel_9801/AMP_IN pixel_9801/SF_IB
+ pixel_9801/PIX_OUT pixel_9801/CSA_VREF pixel
Xpixel_9845 pixel_9845/gring pixel_9845/VDD pixel_9845/GND pixel_9845/VREF pixel_9845/ROW_SEL
+ pixel_9845/NB1 pixel_9845/VBIAS pixel_9845/NB2 pixel_9845/AMP_IN pixel_9845/SF_IB
+ pixel_9845/PIX_OUT pixel_9845/CSA_VREF pixel
Xpixel_9834 pixel_9834/gring pixel_9834/VDD pixel_9834/GND pixel_9834/VREF pixel_9834/ROW_SEL
+ pixel_9834/NB1 pixel_9834/VBIAS pixel_9834/NB2 pixel_9834/AMP_IN pixel_9834/SF_IB
+ pixel_9834/PIX_OUT pixel_9834/CSA_VREF pixel
Xpixel_9856 pixel_9856/gring pixel_9856/VDD pixel_9856/GND pixel_9856/VREF pixel_9856/ROW_SEL
+ pixel_9856/NB1 pixel_9856/VBIAS pixel_9856/NB2 pixel_9856/AMP_IN pixel_9856/SF_IB
+ pixel_9856/PIX_OUT pixel_9856/CSA_VREF pixel
Xpixel_9867 pixel_9867/gring pixel_9867/VDD pixel_9867/GND pixel_9867/VREF pixel_9867/ROW_SEL
+ pixel_9867/NB1 pixel_9867/VBIAS pixel_9867/NB2 pixel_9867/AMP_IN pixel_9867/SF_IB
+ pixel_9867/PIX_OUT pixel_9867/CSA_VREF pixel
Xpixel_9878 pixel_9878/gring pixel_9878/VDD pixel_9878/GND pixel_9878/VREF pixel_9878/ROW_SEL
+ pixel_9878/NB1 pixel_9878/VBIAS pixel_9878/NB2 pixel_9878/AMP_IN pixel_9878/SF_IB
+ pixel_9878/PIX_OUT pixel_9878/CSA_VREF pixel
Xpixel_9889 pixel_9889/gring pixel_9889/VDD pixel_9889/GND pixel_9889/VREF pixel_9889/ROW_SEL
+ pixel_9889/NB1 pixel_9889/VBIAS pixel_9889/NB2 pixel_9889/AMP_IN pixel_9889/SF_IB
+ pixel_9889/PIX_OUT pixel_9889/CSA_VREF pixel
Xpixel_4130 pixel_4130/gring pixel_4130/VDD pixel_4130/GND pixel_4130/VREF pixel_4130/ROW_SEL
+ pixel_4130/NB1 pixel_4130/VBIAS pixel_4130/NB2 pixel_4130/AMP_IN pixel_4130/SF_IB
+ pixel_4130/PIX_OUT pixel_4130/CSA_VREF pixel
Xpixel_4141 pixel_4141/gring pixel_4141/VDD pixel_4141/GND pixel_4141/VREF pixel_4141/ROW_SEL
+ pixel_4141/NB1 pixel_4141/VBIAS pixel_4141/NB2 pixel_4141/AMP_IN pixel_4141/SF_IB
+ pixel_4141/PIX_OUT pixel_4141/CSA_VREF pixel
Xpixel_4152 pixel_4152/gring pixel_4152/VDD pixel_4152/GND pixel_4152/VREF pixel_4152/ROW_SEL
+ pixel_4152/NB1 pixel_4152/VBIAS pixel_4152/NB2 pixel_4152/AMP_IN pixel_4152/SF_IB
+ pixel_4152/PIX_OUT pixel_4152/CSA_VREF pixel
Xpixel_191 pixel_191/gring pixel_191/VDD pixel_191/GND pixel_191/VREF pixel_191/ROW_SEL
+ pixel_191/NB1 pixel_191/VBIAS pixel_191/NB2 pixel_191/AMP_IN pixel_191/SF_IB pixel_191/PIX_OUT
+ pixel_191/CSA_VREF pixel
Xpixel_180 pixel_180/gring pixel_180/VDD pixel_180/GND pixel_180/VREF pixel_180/ROW_SEL
+ pixel_180/NB1 pixel_180/VBIAS pixel_180/NB2 pixel_180/AMP_IN pixel_180/SF_IB pixel_180/PIX_OUT
+ pixel_180/CSA_VREF pixel
Xpixel_3451 pixel_3451/gring pixel_3451/VDD pixel_3451/GND pixel_3451/VREF pixel_3451/ROW_SEL
+ pixel_3451/NB1 pixel_3451/VBIAS pixel_3451/NB2 pixel_3451/AMP_IN pixel_3451/SF_IB
+ pixel_3451/PIX_OUT pixel_3451/CSA_VREF pixel
Xpixel_3440 pixel_3440/gring pixel_3440/VDD pixel_3440/GND pixel_3440/VREF pixel_3440/ROW_SEL
+ pixel_3440/NB1 pixel_3440/VBIAS pixel_3440/NB2 pixel_3440/AMP_IN pixel_3440/SF_IB
+ pixel_3440/PIX_OUT pixel_3440/CSA_VREF pixel
Xpixel_4163 pixel_4163/gring pixel_4163/VDD pixel_4163/GND pixel_4163/VREF pixel_4163/ROW_SEL
+ pixel_4163/NB1 pixel_4163/VBIAS pixel_4163/NB2 pixel_4163/AMP_IN pixel_4163/SF_IB
+ pixel_4163/PIX_OUT pixel_4163/CSA_VREF pixel
Xpixel_4174 pixel_4174/gring pixel_4174/VDD pixel_4174/GND pixel_4174/VREF pixel_4174/ROW_SEL
+ pixel_4174/NB1 pixel_4174/VBIAS pixel_4174/NB2 pixel_4174/AMP_IN pixel_4174/SF_IB
+ pixel_4174/PIX_OUT pixel_4174/CSA_VREF pixel
Xpixel_4185 pixel_4185/gring pixel_4185/VDD pixel_4185/GND pixel_4185/VREF pixel_4185/ROW_SEL
+ pixel_4185/NB1 pixel_4185/VBIAS pixel_4185/NB2 pixel_4185/AMP_IN pixel_4185/SF_IB
+ pixel_4185/PIX_OUT pixel_4185/CSA_VREF pixel
Xpixel_4196 pixel_4196/gring pixel_4196/VDD pixel_4196/GND pixel_4196/VREF pixel_4196/ROW_SEL
+ pixel_4196/NB1 pixel_4196/VBIAS pixel_4196/NB2 pixel_4196/AMP_IN pixel_4196/SF_IB
+ pixel_4196/PIX_OUT pixel_4196/CSA_VREF pixel
Xpixel_3484 pixel_3484/gring pixel_3484/VDD pixel_3484/GND pixel_3484/VREF pixel_3484/ROW_SEL
+ pixel_3484/NB1 pixel_3484/VBIAS pixel_3484/NB2 pixel_3484/AMP_IN pixel_3484/SF_IB
+ pixel_3484/PIX_OUT pixel_3484/CSA_VREF pixel
Xpixel_3473 pixel_3473/gring pixel_3473/VDD pixel_3473/GND pixel_3473/VREF pixel_3473/ROW_SEL
+ pixel_3473/NB1 pixel_3473/VBIAS pixel_3473/NB2 pixel_3473/AMP_IN pixel_3473/SF_IB
+ pixel_3473/PIX_OUT pixel_3473/CSA_VREF pixel
Xpixel_3462 pixel_3462/gring pixel_3462/VDD pixel_3462/GND pixel_3462/VREF pixel_3462/ROW_SEL
+ pixel_3462/NB1 pixel_3462/VBIAS pixel_3462/NB2 pixel_3462/AMP_IN pixel_3462/SF_IB
+ pixel_3462/PIX_OUT pixel_3462/CSA_VREF pixel
Xpixel_2783 pixel_2783/gring pixel_2783/VDD pixel_2783/GND pixel_2783/VREF pixel_2783/ROW_SEL
+ pixel_2783/NB1 pixel_2783/VBIAS pixel_2783/NB2 pixel_2783/AMP_IN pixel_2783/SF_IB
+ pixel_2783/PIX_OUT pixel_2783/CSA_VREF pixel
Xpixel_2772 pixel_2772/gring pixel_2772/VDD pixel_2772/GND pixel_2772/VREF pixel_2772/ROW_SEL
+ pixel_2772/NB1 pixel_2772/VBIAS pixel_2772/NB2 pixel_2772/AMP_IN pixel_2772/SF_IB
+ pixel_2772/PIX_OUT pixel_2772/CSA_VREF pixel
Xpixel_2761 pixel_2761/gring pixel_2761/VDD pixel_2761/GND pixel_2761/VREF pixel_2761/ROW_SEL
+ pixel_2761/NB1 pixel_2761/VBIAS pixel_2761/NB2 pixel_2761/AMP_IN pixel_2761/SF_IB
+ pixel_2761/PIX_OUT pixel_2761/CSA_VREF pixel
Xpixel_2750 pixel_2750/gring pixel_2750/VDD pixel_2750/GND pixel_2750/VREF pixel_2750/ROW_SEL
+ pixel_2750/NB1 pixel_2750/VBIAS pixel_2750/NB2 pixel_2750/AMP_IN pixel_2750/SF_IB
+ pixel_2750/PIX_OUT pixel_2750/CSA_VREF pixel
Xpixel_3495 pixel_3495/gring pixel_3495/VDD pixel_3495/GND pixel_3495/VREF pixel_3495/ROW_SEL
+ pixel_3495/NB1 pixel_3495/VBIAS pixel_3495/NB2 pixel_3495/AMP_IN pixel_3495/SF_IB
+ pixel_3495/PIX_OUT pixel_3495/CSA_VREF pixel
Xpixel_2794 pixel_2794/gring pixel_2794/VDD pixel_2794/GND pixel_2794/VREF pixel_2794/ROW_SEL
+ pixel_2794/NB1 pixel_2794/VBIAS pixel_2794/NB2 pixel_2794/AMP_IN pixel_2794/SF_IB
+ pixel_2794/PIX_OUT pixel_2794/CSA_VREF pixel
Xpixel_9119 pixel_9119/gring pixel_9119/VDD pixel_9119/GND pixel_9119/VREF pixel_9119/ROW_SEL
+ pixel_9119/NB1 pixel_9119/VBIAS pixel_9119/NB2 pixel_9119/AMP_IN pixel_9119/SF_IB
+ pixel_9119/PIX_OUT pixel_9119/CSA_VREF pixel
Xpixel_9108 pixel_9108/gring pixel_9108/VDD pixel_9108/GND pixel_9108/VREF pixel_9108/ROW_SEL
+ pixel_9108/NB1 pixel_9108/VBIAS pixel_9108/NB2 pixel_9108/AMP_IN pixel_9108/SF_IB
+ pixel_9108/PIX_OUT pixel_9108/CSA_VREF pixel
Xpixel_8407 pixel_8407/gring pixel_8407/VDD pixel_8407/GND pixel_8407/VREF pixel_8407/ROW_SEL
+ pixel_8407/NB1 pixel_8407/VBIAS pixel_8407/NB2 pixel_8407/AMP_IN pixel_8407/SF_IB
+ pixel_8407/PIX_OUT pixel_8407/CSA_VREF pixel
Xpixel_8429 pixel_8429/gring pixel_8429/VDD pixel_8429/GND pixel_8429/VREF pixel_8429/ROW_SEL
+ pixel_8429/NB1 pixel_8429/VBIAS pixel_8429/NB2 pixel_8429/AMP_IN pixel_8429/SF_IB
+ pixel_8429/PIX_OUT pixel_8429/CSA_VREF pixel
Xpixel_8418 pixel_8418/gring pixel_8418/VDD pixel_8418/GND pixel_8418/VREF pixel_8418/ROW_SEL
+ pixel_8418/NB1 pixel_8418/VBIAS pixel_8418/NB2 pixel_8418/AMP_IN pixel_8418/SF_IB
+ pixel_8418/PIX_OUT pixel_8418/CSA_VREF pixel
Xpixel_7706 pixel_7706/gring pixel_7706/VDD pixel_7706/GND pixel_7706/VREF pixel_7706/ROW_SEL
+ pixel_7706/NB1 pixel_7706/VBIAS pixel_7706/NB2 pixel_7706/AMP_IN pixel_7706/SF_IB
+ pixel_7706/PIX_OUT pixel_7706/CSA_VREF pixel
Xpixel_7717 pixel_7717/gring pixel_7717/VDD pixel_7717/GND pixel_7717/VREF pixel_7717/ROW_SEL
+ pixel_7717/NB1 pixel_7717/VBIAS pixel_7717/NB2 pixel_7717/AMP_IN pixel_7717/SF_IB
+ pixel_7717/PIX_OUT pixel_7717/CSA_VREF pixel
Xpixel_7728 pixel_7728/gring pixel_7728/VDD pixel_7728/GND pixel_7728/VREF pixel_7728/ROW_SEL
+ pixel_7728/NB1 pixel_7728/VBIAS pixel_7728/NB2 pixel_7728/AMP_IN pixel_7728/SF_IB
+ pixel_7728/PIX_OUT pixel_7728/CSA_VREF pixel
Xpixel_7739 pixel_7739/gring pixel_7739/VDD pixel_7739/GND pixel_7739/VREF pixel_7739/ROW_SEL
+ pixel_7739/NB1 pixel_7739/VBIAS pixel_7739/NB2 pixel_7739/AMP_IN pixel_7739/SF_IB
+ pixel_7739/PIX_OUT pixel_7739/CSA_VREF pixel
Xpixel_2002 pixel_2002/gring pixel_2002/VDD pixel_2002/GND pixel_2002/VREF pixel_2002/ROW_SEL
+ pixel_2002/NB1 pixel_2002/VBIAS pixel_2002/NB2 pixel_2002/AMP_IN pixel_2002/SF_IB
+ pixel_2002/PIX_OUT pixel_2002/CSA_VREF pixel
Xpixel_2035 pixel_2035/gring pixel_2035/VDD pixel_2035/GND pixel_2035/VREF pixel_2035/ROW_SEL
+ pixel_2035/NB1 pixel_2035/VBIAS pixel_2035/NB2 pixel_2035/AMP_IN pixel_2035/SF_IB
+ pixel_2035/PIX_OUT pixel_2035/CSA_VREF pixel
Xpixel_2024 pixel_2024/gring pixel_2024/VDD pixel_2024/GND pixel_2024/VREF pixel_2024/ROW_SEL
+ pixel_2024/NB1 pixel_2024/VBIAS pixel_2024/NB2 pixel_2024/AMP_IN pixel_2024/SF_IB
+ pixel_2024/PIX_OUT pixel_2024/CSA_VREF pixel
Xpixel_2013 pixel_2013/gring pixel_2013/VDD pixel_2013/GND pixel_2013/VREF pixel_2013/ROW_SEL
+ pixel_2013/NB1 pixel_2013/VBIAS pixel_2013/NB2 pixel_2013/AMP_IN pixel_2013/SF_IB
+ pixel_2013/PIX_OUT pixel_2013/CSA_VREF pixel
Xpixel_1323 pixel_1323/gring pixel_1323/VDD pixel_1323/GND pixel_1323/VREF pixel_1323/ROW_SEL
+ pixel_1323/NB1 pixel_1323/VBIAS pixel_1323/NB2 pixel_1323/AMP_IN pixel_1323/SF_IB
+ pixel_1323/PIX_OUT pixel_1323/CSA_VREF pixel
Xpixel_1312 pixel_1312/gring pixel_1312/VDD pixel_1312/GND pixel_1312/VREF pixel_1312/ROW_SEL
+ pixel_1312/NB1 pixel_1312/VBIAS pixel_1312/NB2 pixel_1312/AMP_IN pixel_1312/SF_IB
+ pixel_1312/PIX_OUT pixel_1312/CSA_VREF pixel
Xpixel_1301 pixel_1301/gring pixel_1301/VDD pixel_1301/GND pixel_1301/VREF pixel_1301/ROW_SEL
+ pixel_1301/NB1 pixel_1301/VBIAS pixel_1301/NB2 pixel_1301/AMP_IN pixel_1301/SF_IB
+ pixel_1301/PIX_OUT pixel_1301/CSA_VREF pixel
Xpixel_2068 pixel_2068/gring pixel_2068/VDD pixel_2068/GND pixel_2068/VREF pixel_2068/ROW_SEL
+ pixel_2068/NB1 pixel_2068/VBIAS pixel_2068/NB2 pixel_2068/AMP_IN pixel_2068/SF_IB
+ pixel_2068/PIX_OUT pixel_2068/CSA_VREF pixel
Xpixel_2057 pixel_2057/gring pixel_2057/VDD pixel_2057/GND pixel_2057/VREF pixel_2057/ROW_SEL
+ pixel_2057/NB1 pixel_2057/VBIAS pixel_2057/NB2 pixel_2057/AMP_IN pixel_2057/SF_IB
+ pixel_2057/PIX_OUT pixel_2057/CSA_VREF pixel
Xpixel_2046 pixel_2046/gring pixel_2046/VDD pixel_2046/GND pixel_2046/VREF pixel_2046/ROW_SEL
+ pixel_2046/NB1 pixel_2046/VBIAS pixel_2046/NB2 pixel_2046/AMP_IN pixel_2046/SF_IB
+ pixel_2046/PIX_OUT pixel_2046/CSA_VREF pixel
Xpixel_1367 pixel_1367/gring pixel_1367/VDD pixel_1367/GND pixel_1367/VREF pixel_1367/ROW_SEL
+ pixel_1367/NB1 pixel_1367/VBIAS pixel_1367/NB2 pixel_1367/AMP_IN pixel_1367/SF_IB
+ pixel_1367/PIX_OUT pixel_1367/CSA_VREF pixel
Xpixel_1356 pixel_1356/gring pixel_1356/VDD pixel_1356/GND pixel_1356/VREF pixel_1356/ROW_SEL
+ pixel_1356/NB1 pixel_1356/VBIAS pixel_1356/NB2 pixel_1356/AMP_IN pixel_1356/SF_IB
+ pixel_1356/PIX_OUT pixel_1356/CSA_VREF pixel
Xpixel_1345 pixel_1345/gring pixel_1345/VDD pixel_1345/GND pixel_1345/VREF pixel_1345/ROW_SEL
+ pixel_1345/NB1 pixel_1345/VBIAS pixel_1345/NB2 pixel_1345/AMP_IN pixel_1345/SF_IB
+ pixel_1345/PIX_OUT pixel_1345/CSA_VREF pixel
Xpixel_1334 pixel_1334/gring pixel_1334/VDD pixel_1334/GND pixel_1334/VREF pixel_1334/ROW_SEL
+ pixel_1334/NB1 pixel_1334/VBIAS pixel_1334/NB2 pixel_1334/AMP_IN pixel_1334/SF_IB
+ pixel_1334/PIX_OUT pixel_1334/CSA_VREF pixel
Xpixel_2079 pixel_2079/gring pixel_2079/VDD pixel_2079/GND pixel_2079/VREF pixel_2079/ROW_SEL
+ pixel_2079/NB1 pixel_2079/VBIAS pixel_2079/NB2 pixel_2079/AMP_IN pixel_2079/SF_IB
+ pixel_2079/PIX_OUT pixel_2079/CSA_VREF pixel
Xpixel_1389 pixel_1389/gring pixel_1389/VDD pixel_1389/GND pixel_1389/VREF pixel_1389/ROW_SEL
+ pixel_1389/NB1 pixel_1389/VBIAS pixel_1389/NB2 pixel_1389/AMP_IN pixel_1389/SF_IB
+ pixel_1389/PIX_OUT pixel_1389/CSA_VREF pixel
Xpixel_1378 pixel_1378/gring pixel_1378/VDD pixel_1378/GND pixel_1378/VREF pixel_1378/ROW_SEL
+ pixel_1378/NB1 pixel_1378/VBIAS pixel_1378/NB2 pixel_1378/AMP_IN pixel_1378/SF_IB
+ pixel_1378/PIX_OUT pixel_1378/CSA_VREF pixel
Xpixel_9620 pixel_9620/gring pixel_9620/VDD pixel_9620/GND pixel_9620/VREF pixel_9620/ROW_SEL
+ pixel_9620/NB1 pixel_9620/VBIAS pixel_9620/NB2 pixel_9620/AMP_IN pixel_9620/SF_IB
+ pixel_9620/PIX_OUT pixel_9620/CSA_VREF pixel
Xpixel_9631 pixel_9631/gring pixel_9631/VDD pixel_9631/GND pixel_9631/VREF pixel_9631/ROW_SEL
+ pixel_9631/NB1 pixel_9631/VBIAS pixel_9631/NB2 pixel_9631/AMP_IN pixel_9631/SF_IB
+ pixel_9631/PIX_OUT pixel_9631/CSA_VREF pixel
Xpixel_8930 pixel_8930/gring pixel_8930/VDD pixel_8930/GND pixel_8930/VREF pixel_8930/ROW_SEL
+ pixel_8930/NB1 pixel_8930/VBIAS pixel_8930/NB2 pixel_8930/AMP_IN pixel_8930/SF_IB
+ pixel_8930/PIX_OUT pixel_8930/CSA_VREF pixel
Xpixel_9642 pixel_9642/gring pixel_9642/VDD pixel_9642/GND pixel_9642/VREF pixel_9642/ROW_SEL
+ pixel_9642/NB1 pixel_9642/VBIAS pixel_9642/NB2 pixel_9642/AMP_IN pixel_9642/SF_IB
+ pixel_9642/PIX_OUT pixel_9642/CSA_VREF pixel
Xpixel_9653 pixel_9653/gring pixel_9653/VDD pixel_9653/GND pixel_9653/VREF pixel_9653/ROW_SEL
+ pixel_9653/NB1 pixel_9653/VBIAS pixel_9653/NB2 pixel_9653/AMP_IN pixel_9653/SF_IB
+ pixel_9653/PIX_OUT pixel_9653/CSA_VREF pixel
Xpixel_9664 pixel_9664/gring pixel_9664/VDD pixel_9664/GND pixel_9664/VREF pixel_9664/ROW_SEL
+ pixel_9664/NB1 pixel_9664/VBIAS pixel_9664/NB2 pixel_9664/AMP_IN pixel_9664/SF_IB
+ pixel_9664/PIX_OUT pixel_9664/CSA_VREF pixel
Xpixel_9675 pixel_9675/gring pixel_9675/VDD pixel_9675/GND pixel_9675/VREF pixel_9675/ROW_SEL
+ pixel_9675/NB1 pixel_9675/VBIAS pixel_9675/NB2 pixel_9675/AMP_IN pixel_9675/SF_IB
+ pixel_9675/PIX_OUT pixel_9675/CSA_VREF pixel
Xpixel_8963 pixel_8963/gring pixel_8963/VDD pixel_8963/GND pixel_8963/VREF pixel_8963/ROW_SEL
+ pixel_8963/NB1 pixel_8963/VBIAS pixel_8963/NB2 pixel_8963/AMP_IN pixel_8963/SF_IB
+ pixel_8963/PIX_OUT pixel_8963/CSA_VREF pixel
Xpixel_8952 pixel_8952/gring pixel_8952/VDD pixel_8952/GND pixel_8952/VREF pixel_8952/ROW_SEL
+ pixel_8952/NB1 pixel_8952/VBIAS pixel_8952/NB2 pixel_8952/AMP_IN pixel_8952/SF_IB
+ pixel_8952/PIX_OUT pixel_8952/CSA_VREF pixel
Xpixel_8941 pixel_8941/gring pixel_8941/VDD pixel_8941/GND pixel_8941/VREF pixel_8941/ROW_SEL
+ pixel_8941/NB1 pixel_8941/VBIAS pixel_8941/NB2 pixel_8941/AMP_IN pixel_8941/SF_IB
+ pixel_8941/PIX_OUT pixel_8941/CSA_VREF pixel
Xpixel_9697 pixel_9697/gring pixel_9697/VDD pixel_9697/GND pixel_9697/VREF pixel_9697/ROW_SEL
+ pixel_9697/NB1 pixel_9697/VBIAS pixel_9697/NB2 pixel_9697/AMP_IN pixel_9697/SF_IB
+ pixel_9697/PIX_OUT pixel_9697/CSA_VREF pixel
Xpixel_9686 pixel_9686/gring pixel_9686/VDD pixel_9686/GND pixel_9686/VREF pixel_9686/ROW_SEL
+ pixel_9686/NB1 pixel_9686/VBIAS pixel_9686/NB2 pixel_9686/AMP_IN pixel_9686/SF_IB
+ pixel_9686/PIX_OUT pixel_9686/CSA_VREF pixel
Xpixel_8996 pixel_8996/gring pixel_8996/VDD pixel_8996/GND pixel_8996/VREF pixel_8996/ROW_SEL
+ pixel_8996/NB1 pixel_8996/VBIAS pixel_8996/NB2 pixel_8996/AMP_IN pixel_8996/SF_IB
+ pixel_8996/PIX_OUT pixel_8996/CSA_VREF pixel
Xpixel_8985 pixel_8985/gring pixel_8985/VDD pixel_8985/GND pixel_8985/VREF pixel_8985/ROW_SEL
+ pixel_8985/NB1 pixel_8985/VBIAS pixel_8985/NB2 pixel_8985/AMP_IN pixel_8985/SF_IB
+ pixel_8985/PIX_OUT pixel_8985/CSA_VREF pixel
Xpixel_8974 pixel_8974/gring pixel_8974/VDD pixel_8974/GND pixel_8974/VREF pixel_8974/ROW_SEL
+ pixel_8974/NB1 pixel_8974/VBIAS pixel_8974/NB2 pixel_8974/AMP_IN pixel_8974/SF_IB
+ pixel_8974/PIX_OUT pixel_8974/CSA_VREF pixel
Xpixel_3292 pixel_3292/gring pixel_3292/VDD pixel_3292/GND pixel_3292/VREF pixel_3292/ROW_SEL
+ pixel_3292/NB1 pixel_3292/VBIAS pixel_3292/NB2 pixel_3292/AMP_IN pixel_3292/SF_IB
+ pixel_3292/PIX_OUT pixel_3292/CSA_VREF pixel
Xpixel_3281 pixel_3281/gring pixel_3281/VDD pixel_3281/GND pixel_3281/VREF pixel_3281/ROW_SEL
+ pixel_3281/NB1 pixel_3281/VBIAS pixel_3281/NB2 pixel_3281/AMP_IN pixel_3281/SF_IB
+ pixel_3281/PIX_OUT pixel_3281/CSA_VREF pixel
Xpixel_3270 pixel_3270/gring pixel_3270/VDD pixel_3270/GND pixel_3270/VREF pixel_3270/ROW_SEL
+ pixel_3270/NB1 pixel_3270/VBIAS pixel_3270/NB2 pixel_3270/AMP_IN pixel_3270/SF_IB
+ pixel_3270/PIX_OUT pixel_3270/CSA_VREF pixel
Xpixel_2591 pixel_2591/gring pixel_2591/VDD pixel_2591/GND pixel_2591/VREF pixel_2591/ROW_SEL
+ pixel_2591/NB1 pixel_2591/VBIAS pixel_2591/NB2 pixel_2591/AMP_IN pixel_2591/SF_IB
+ pixel_2591/PIX_OUT pixel_2591/CSA_VREF pixel
Xpixel_2580 pixel_2580/gring pixel_2580/VDD pixel_2580/GND pixel_2580/VREF pixel_2580/ROW_SEL
+ pixel_2580/NB1 pixel_2580/VBIAS pixel_2580/NB2 pixel_2580/AMP_IN pixel_2580/SF_IB
+ pixel_2580/PIX_OUT pixel_2580/CSA_VREF pixel
Xpixel_1890 pixel_1890/gring pixel_1890/VDD pixel_1890/GND pixel_1890/VREF pixel_1890/ROW_SEL
+ pixel_1890/NB1 pixel_1890/VBIAS pixel_1890/NB2 pixel_1890/AMP_IN pixel_1890/SF_IB
+ pixel_1890/PIX_OUT pixel_1890/CSA_VREF pixel
Xpixel_905 pixel_905/gring pixel_905/VDD pixel_905/GND pixel_905/VREF pixel_905/ROW_SEL
+ pixel_905/NB1 pixel_905/VBIAS pixel_905/NB2 pixel_905/AMP_IN pixel_905/SF_IB pixel_905/PIX_OUT
+ pixel_905/CSA_VREF pixel
Xpixel_949 pixel_949/gring pixel_949/VDD pixel_949/GND pixel_949/VREF pixel_949/ROW_SEL
+ pixel_949/NB1 pixel_949/VBIAS pixel_949/NB2 pixel_949/AMP_IN pixel_949/SF_IB pixel_949/PIX_OUT
+ pixel_949/CSA_VREF pixel
Xpixel_938 pixel_938/gring pixel_938/VDD pixel_938/GND pixel_938/VREF pixel_938/ROW_SEL
+ pixel_938/NB1 pixel_938/VBIAS pixel_938/NB2 pixel_938/AMP_IN pixel_938/SF_IB pixel_938/PIX_OUT
+ pixel_938/CSA_VREF pixel
Xpixel_927 pixel_927/gring pixel_927/VDD pixel_927/GND pixel_927/VREF pixel_927/ROW_SEL
+ pixel_927/NB1 pixel_927/VBIAS pixel_927/NB2 pixel_927/AMP_IN pixel_927/SF_IB pixel_927/PIX_OUT
+ pixel_927/CSA_VREF pixel
Xpixel_916 pixel_916/gring pixel_916/VDD pixel_916/GND pixel_916/VREF pixel_916/ROW_SEL
+ pixel_916/NB1 pixel_916/VBIAS pixel_916/NB2 pixel_916/AMP_IN pixel_916/SF_IB pixel_916/PIX_OUT
+ pixel_916/CSA_VREF pixel
Xpixel_8204 pixel_8204/gring pixel_8204/VDD pixel_8204/GND pixel_8204/VREF pixel_8204/ROW_SEL
+ pixel_8204/NB1 pixel_8204/VBIAS pixel_8204/NB2 pixel_8204/AMP_IN pixel_8204/SF_IB
+ pixel_8204/PIX_OUT pixel_8204/CSA_VREF pixel
Xpixel_8215 pixel_8215/gring pixel_8215/VDD pixel_8215/GND pixel_8215/VREF pixel_8215/ROW_SEL
+ pixel_8215/NB1 pixel_8215/VBIAS pixel_8215/NB2 pixel_8215/AMP_IN pixel_8215/SF_IB
+ pixel_8215/PIX_OUT pixel_8215/CSA_VREF pixel
Xpixel_8226 pixel_8226/gring pixel_8226/VDD pixel_8226/GND pixel_8226/VREF pixel_8226/ROW_SEL
+ pixel_8226/NB1 pixel_8226/VBIAS pixel_8226/NB2 pixel_8226/AMP_IN pixel_8226/SF_IB
+ pixel_8226/PIX_OUT pixel_8226/CSA_VREF pixel
Xpixel_8237 pixel_8237/gring pixel_8237/VDD pixel_8237/GND pixel_8237/VREF pixel_8237/ROW_SEL
+ pixel_8237/NB1 pixel_8237/VBIAS pixel_8237/NB2 pixel_8237/AMP_IN pixel_8237/SF_IB
+ pixel_8237/PIX_OUT pixel_8237/CSA_VREF pixel
Xpixel_8248 pixel_8248/gring pixel_8248/VDD pixel_8248/GND pixel_8248/VREF pixel_8248/ROW_SEL
+ pixel_8248/NB1 pixel_8248/VBIAS pixel_8248/NB2 pixel_8248/AMP_IN pixel_8248/SF_IB
+ pixel_8248/PIX_OUT pixel_8248/CSA_VREF pixel
Xpixel_8259 pixel_8259/gring pixel_8259/VDD pixel_8259/GND pixel_8259/VREF pixel_8259/ROW_SEL
+ pixel_8259/NB1 pixel_8259/VBIAS pixel_8259/NB2 pixel_8259/AMP_IN pixel_8259/SF_IB
+ pixel_8259/PIX_OUT pixel_8259/CSA_VREF pixel
Xpixel_7503 pixel_7503/gring pixel_7503/VDD pixel_7503/GND pixel_7503/VREF pixel_7503/ROW_SEL
+ pixel_7503/NB1 pixel_7503/VBIAS pixel_7503/NB2 pixel_7503/AMP_IN pixel_7503/SF_IB
+ pixel_7503/PIX_OUT pixel_7503/CSA_VREF pixel
Xpixel_7514 pixel_7514/gring pixel_7514/VDD pixel_7514/GND pixel_7514/VREF pixel_7514/ROW_SEL
+ pixel_7514/NB1 pixel_7514/VBIAS pixel_7514/NB2 pixel_7514/AMP_IN pixel_7514/SF_IB
+ pixel_7514/PIX_OUT pixel_7514/CSA_VREF pixel
Xpixel_7525 pixel_7525/gring pixel_7525/VDD pixel_7525/GND pixel_7525/VREF pixel_7525/ROW_SEL
+ pixel_7525/NB1 pixel_7525/VBIAS pixel_7525/NB2 pixel_7525/AMP_IN pixel_7525/SF_IB
+ pixel_7525/PIX_OUT pixel_7525/CSA_VREF pixel
Xpixel_7536 pixel_7536/gring pixel_7536/VDD pixel_7536/GND pixel_7536/VREF pixel_7536/ROW_SEL
+ pixel_7536/NB1 pixel_7536/VBIAS pixel_7536/NB2 pixel_7536/AMP_IN pixel_7536/SF_IB
+ pixel_7536/PIX_OUT pixel_7536/CSA_VREF pixel
Xpixel_7547 pixel_7547/gring pixel_7547/VDD pixel_7547/GND pixel_7547/VREF pixel_7547/ROW_SEL
+ pixel_7547/NB1 pixel_7547/VBIAS pixel_7547/NB2 pixel_7547/AMP_IN pixel_7547/SF_IB
+ pixel_7547/PIX_OUT pixel_7547/CSA_VREF pixel
Xpixel_6802 pixel_6802/gring pixel_6802/VDD pixel_6802/GND pixel_6802/VREF pixel_6802/ROW_SEL
+ pixel_6802/NB1 pixel_6802/VBIAS pixel_6802/NB2 pixel_6802/AMP_IN pixel_6802/SF_IB
+ pixel_6802/PIX_OUT pixel_6802/CSA_VREF pixel
Xpixel_7558 pixel_7558/gring pixel_7558/VDD pixel_7558/GND pixel_7558/VREF pixel_7558/ROW_SEL
+ pixel_7558/NB1 pixel_7558/VBIAS pixel_7558/NB2 pixel_7558/AMP_IN pixel_7558/SF_IB
+ pixel_7558/PIX_OUT pixel_7558/CSA_VREF pixel
Xpixel_7569 pixel_7569/gring pixel_7569/VDD pixel_7569/GND pixel_7569/VREF pixel_7569/ROW_SEL
+ pixel_7569/NB1 pixel_7569/VBIAS pixel_7569/NB2 pixel_7569/AMP_IN pixel_7569/SF_IB
+ pixel_7569/PIX_OUT pixel_7569/CSA_VREF pixel
Xpixel_6813 pixel_6813/gring pixel_6813/VDD pixel_6813/GND pixel_6813/VREF pixel_6813/ROW_SEL
+ pixel_6813/NB1 pixel_6813/VBIAS pixel_6813/NB2 pixel_6813/AMP_IN pixel_6813/SF_IB
+ pixel_6813/PIX_OUT pixel_6813/CSA_VREF pixel
Xpixel_6824 pixel_6824/gring pixel_6824/VDD pixel_6824/GND pixel_6824/VREF pixel_6824/ROW_SEL
+ pixel_6824/NB1 pixel_6824/VBIAS pixel_6824/NB2 pixel_6824/AMP_IN pixel_6824/SF_IB
+ pixel_6824/PIX_OUT pixel_6824/CSA_VREF pixel
Xpixel_6835 pixel_6835/gring pixel_6835/VDD pixel_6835/GND pixel_6835/VREF pixel_6835/ROW_SEL
+ pixel_6835/NB1 pixel_6835/VBIAS pixel_6835/NB2 pixel_6835/AMP_IN pixel_6835/SF_IB
+ pixel_6835/PIX_OUT pixel_6835/CSA_VREF pixel
Xpixel_6846 pixel_6846/gring pixel_6846/VDD pixel_6846/GND pixel_6846/VREF pixel_6846/ROW_SEL
+ pixel_6846/NB1 pixel_6846/VBIAS pixel_6846/NB2 pixel_6846/AMP_IN pixel_6846/SF_IB
+ pixel_6846/PIX_OUT pixel_6846/CSA_VREF pixel
Xpixel_6857 pixel_6857/gring pixel_6857/VDD pixel_6857/GND pixel_6857/VREF pixel_6857/ROW_SEL
+ pixel_6857/NB1 pixel_6857/VBIAS pixel_6857/NB2 pixel_6857/AMP_IN pixel_6857/SF_IB
+ pixel_6857/PIX_OUT pixel_6857/CSA_VREF pixel
Xpixel_6868 pixel_6868/gring pixel_6868/VDD pixel_6868/GND pixel_6868/VREF pixel_6868/ROW_SEL
+ pixel_6868/NB1 pixel_6868/VBIAS pixel_6868/NB2 pixel_6868/AMP_IN pixel_6868/SF_IB
+ pixel_6868/PIX_OUT pixel_6868/CSA_VREF pixel
Xpixel_6879 pixel_6879/gring pixel_6879/VDD pixel_6879/GND pixel_6879/VREF pixel_6879/ROW_SEL
+ pixel_6879/NB1 pixel_6879/VBIAS pixel_6879/NB2 pixel_6879/AMP_IN pixel_6879/SF_IB
+ pixel_6879/PIX_OUT pixel_6879/CSA_VREF pixel
Xpixel_1142 pixel_1142/gring pixel_1142/VDD pixel_1142/GND pixel_1142/VREF pixel_1142/ROW_SEL
+ pixel_1142/NB1 pixel_1142/VBIAS pixel_1142/NB2 pixel_1142/AMP_IN pixel_1142/SF_IB
+ pixel_1142/PIX_OUT pixel_1142/CSA_VREF pixel
Xpixel_1131 pixel_1131/gring pixel_1131/VDD pixel_1131/GND pixel_1131/VREF pixel_1131/ROW_SEL
+ pixel_1131/NB1 pixel_1131/VBIAS pixel_1131/NB2 pixel_1131/AMP_IN pixel_1131/SF_IB
+ pixel_1131/PIX_OUT pixel_1131/CSA_VREF pixel
Xpixel_1120 pixel_1120/gring pixel_1120/VDD pixel_1120/GND pixel_1120/VREF pixel_1120/ROW_SEL
+ pixel_1120/NB1 pixel_1120/VBIAS pixel_1120/NB2 pixel_1120/AMP_IN pixel_1120/SF_IB
+ pixel_1120/PIX_OUT pixel_1120/CSA_VREF pixel
Xpixel_1175 pixel_1175/gring pixel_1175/VDD pixel_1175/GND pixel_1175/VREF pixel_1175/ROW_SEL
+ pixel_1175/NB1 pixel_1175/VBIAS pixel_1175/NB2 pixel_1175/AMP_IN pixel_1175/SF_IB
+ pixel_1175/PIX_OUT pixel_1175/CSA_VREF pixel
Xpixel_1164 pixel_1164/gring pixel_1164/VDD pixel_1164/GND pixel_1164/VREF pixel_1164/ROW_SEL
+ pixel_1164/NB1 pixel_1164/VBIAS pixel_1164/NB2 pixel_1164/AMP_IN pixel_1164/SF_IB
+ pixel_1164/PIX_OUT pixel_1164/CSA_VREF pixel
Xpixel_1153 pixel_1153/gring pixel_1153/VDD pixel_1153/GND pixel_1153/VREF pixel_1153/ROW_SEL
+ pixel_1153/NB1 pixel_1153/VBIAS pixel_1153/NB2 pixel_1153/AMP_IN pixel_1153/SF_IB
+ pixel_1153/PIX_OUT pixel_1153/CSA_VREF pixel
Xpixel_1197 pixel_1197/gring pixel_1197/VDD pixel_1197/GND pixel_1197/VREF pixel_1197/ROW_SEL
+ pixel_1197/NB1 pixel_1197/VBIAS pixel_1197/NB2 pixel_1197/AMP_IN pixel_1197/SF_IB
+ pixel_1197/PIX_OUT pixel_1197/CSA_VREF pixel
Xpixel_1186 pixel_1186/gring pixel_1186/VDD pixel_1186/GND pixel_1186/VREF pixel_1186/ROW_SEL
+ pixel_1186/NB1 pixel_1186/VBIAS pixel_1186/NB2 pixel_1186/AMP_IN pixel_1186/SF_IB
+ pixel_1186/PIX_OUT pixel_1186/CSA_VREF pixel
Xpixel_9450 pixel_9450/gring pixel_9450/VDD pixel_9450/GND pixel_9450/VREF pixel_9450/ROW_SEL
+ pixel_9450/NB1 pixel_9450/VBIAS pixel_9450/NB2 pixel_9450/AMP_IN pixel_9450/SF_IB
+ pixel_9450/PIX_OUT pixel_9450/CSA_VREF pixel
Xpixel_9483 pixel_9483/gring pixel_9483/VDD pixel_9483/GND pixel_9483/VREF pixel_9483/ROW_SEL
+ pixel_9483/NB1 pixel_9483/VBIAS pixel_9483/NB2 pixel_9483/AMP_IN pixel_9483/SF_IB
+ pixel_9483/PIX_OUT pixel_9483/CSA_VREF pixel
Xpixel_9472 pixel_9472/gring pixel_9472/VDD pixel_9472/GND pixel_9472/VREF pixel_9472/ROW_SEL
+ pixel_9472/NB1 pixel_9472/VBIAS pixel_9472/NB2 pixel_9472/AMP_IN pixel_9472/SF_IB
+ pixel_9472/PIX_OUT pixel_9472/CSA_VREF pixel
Xpixel_9461 pixel_9461/gring pixel_9461/VDD pixel_9461/GND pixel_9461/VREF pixel_9461/ROW_SEL
+ pixel_9461/NB1 pixel_9461/VBIAS pixel_9461/NB2 pixel_9461/AMP_IN pixel_9461/SF_IB
+ pixel_9461/PIX_OUT pixel_9461/CSA_VREF pixel
Xpixel_8771 pixel_8771/gring pixel_8771/VDD pixel_8771/GND pixel_8771/VREF pixel_8771/ROW_SEL
+ pixel_8771/NB1 pixel_8771/VBIAS pixel_8771/NB2 pixel_8771/AMP_IN pixel_8771/SF_IB
+ pixel_8771/PIX_OUT pixel_8771/CSA_VREF pixel
Xpixel_8760 pixel_8760/gring pixel_8760/VDD pixel_8760/GND pixel_8760/VREF pixel_8760/ROW_SEL
+ pixel_8760/NB1 pixel_8760/VBIAS pixel_8760/NB2 pixel_8760/AMP_IN pixel_8760/SF_IB
+ pixel_8760/PIX_OUT pixel_8760/CSA_VREF pixel
Xpixel_9494 pixel_9494/gring pixel_9494/VDD pixel_9494/GND pixel_9494/VREF pixel_9494/ROW_SEL
+ pixel_9494/NB1 pixel_9494/VBIAS pixel_9494/NB2 pixel_9494/AMP_IN pixel_9494/SF_IB
+ pixel_9494/PIX_OUT pixel_9494/CSA_VREF pixel
Xpixel_8793 pixel_8793/gring pixel_8793/VDD pixel_8793/GND pixel_8793/VREF pixel_8793/ROW_SEL
+ pixel_8793/NB1 pixel_8793/VBIAS pixel_8793/NB2 pixel_8793/AMP_IN pixel_8793/SF_IB
+ pixel_8793/PIX_OUT pixel_8793/CSA_VREF pixel
Xpixel_8782 pixel_8782/gring pixel_8782/VDD pixel_8782/GND pixel_8782/VREF pixel_8782/ROW_SEL
+ pixel_8782/NB1 pixel_8782/VBIAS pixel_8782/NB2 pixel_8782/AMP_IN pixel_8782/SF_IB
+ pixel_8782/PIX_OUT pixel_8782/CSA_VREF pixel
Xpixel_6109 pixel_6109/gring pixel_6109/VDD pixel_6109/GND pixel_6109/VREF pixel_6109/ROW_SEL
+ pixel_6109/NB1 pixel_6109/VBIAS pixel_6109/NB2 pixel_6109/AMP_IN pixel_6109/SF_IB
+ pixel_6109/PIX_OUT pixel_6109/CSA_VREF pixel
Xpixel_5408 pixel_5408/gring pixel_5408/VDD pixel_5408/GND pixel_5408/VREF pixel_5408/ROW_SEL
+ pixel_5408/NB1 pixel_5408/VBIAS pixel_5408/NB2 pixel_5408/AMP_IN pixel_5408/SF_IB
+ pixel_5408/PIX_OUT pixel_5408/CSA_VREF pixel
Xpixel_5419 pixel_5419/gring pixel_5419/VDD pixel_5419/GND pixel_5419/VREF pixel_5419/ROW_SEL
+ pixel_5419/NB1 pixel_5419/VBIAS pixel_5419/NB2 pixel_5419/AMP_IN pixel_5419/SF_IB
+ pixel_5419/PIX_OUT pixel_5419/CSA_VREF pixel
Xpixel_724 pixel_724/gring pixel_724/VDD pixel_724/GND pixel_724/VREF pixel_724/ROW_SEL
+ pixel_724/NB1 pixel_724/VBIAS pixel_724/NB2 pixel_724/AMP_IN pixel_724/SF_IB pixel_724/PIX_OUT
+ pixel_724/CSA_VREF pixel
Xpixel_713 pixel_713/gring pixel_713/VDD pixel_713/GND pixel_713/VREF pixel_713/ROW_SEL
+ pixel_713/NB1 pixel_713/VBIAS pixel_713/NB2 pixel_713/AMP_IN pixel_713/SF_IB pixel_713/PIX_OUT
+ pixel_713/CSA_VREF pixel
Xpixel_702 pixel_702/gring pixel_702/VDD pixel_702/GND pixel_702/VREF pixel_702/ROW_SEL
+ pixel_702/NB1 pixel_702/VBIAS pixel_702/NB2 pixel_702/AMP_IN pixel_702/SF_IB pixel_702/PIX_OUT
+ pixel_702/CSA_VREF pixel
Xpixel_4707 pixel_4707/gring pixel_4707/VDD pixel_4707/GND pixel_4707/VREF pixel_4707/ROW_SEL
+ pixel_4707/NB1 pixel_4707/VBIAS pixel_4707/NB2 pixel_4707/AMP_IN pixel_4707/SF_IB
+ pixel_4707/PIX_OUT pixel_4707/CSA_VREF pixel
Xpixel_4718 pixel_4718/gring pixel_4718/VDD pixel_4718/GND pixel_4718/VREF pixel_4718/ROW_SEL
+ pixel_4718/NB1 pixel_4718/VBIAS pixel_4718/NB2 pixel_4718/AMP_IN pixel_4718/SF_IB
+ pixel_4718/PIX_OUT pixel_4718/CSA_VREF pixel
Xpixel_757 pixel_757/gring pixel_757/VDD pixel_757/GND pixel_757/VREF pixel_757/ROW_SEL
+ pixel_757/NB1 pixel_757/VBIAS pixel_757/NB2 pixel_757/AMP_IN pixel_757/SF_IB pixel_757/PIX_OUT
+ pixel_757/CSA_VREF pixel
Xpixel_746 pixel_746/gring pixel_746/VDD pixel_746/GND pixel_746/VREF pixel_746/ROW_SEL
+ pixel_746/NB1 pixel_746/VBIAS pixel_746/NB2 pixel_746/AMP_IN pixel_746/SF_IB pixel_746/PIX_OUT
+ pixel_746/CSA_VREF pixel
Xpixel_735 pixel_735/gring pixel_735/VDD pixel_735/GND pixel_735/VREF pixel_735/ROW_SEL
+ pixel_735/NB1 pixel_735/VBIAS pixel_735/NB2 pixel_735/AMP_IN pixel_735/SF_IB pixel_735/PIX_OUT
+ pixel_735/CSA_VREF pixel
Xpixel_4729 pixel_4729/gring pixel_4729/VDD pixel_4729/GND pixel_4729/VREF pixel_4729/ROW_SEL
+ pixel_4729/NB1 pixel_4729/VBIAS pixel_4729/NB2 pixel_4729/AMP_IN pixel_4729/SF_IB
+ pixel_4729/PIX_OUT pixel_4729/CSA_VREF pixel
Xpixel_779 pixel_779/gring pixel_779/VDD pixel_779/GND pixel_779/VREF pixel_779/ROW_SEL
+ pixel_779/NB1 pixel_779/VBIAS pixel_779/NB2 pixel_779/AMP_IN pixel_779/SF_IB pixel_779/PIX_OUT
+ pixel_779/CSA_VREF pixel
Xpixel_768 pixel_768/gring pixel_768/VDD pixel_768/GND pixel_768/VREF pixel_768/ROW_SEL
+ pixel_768/NB1 pixel_768/VBIAS pixel_768/NB2 pixel_768/AMP_IN pixel_768/SF_IB pixel_768/PIX_OUT
+ pixel_768/CSA_VREF pixel
Xpixel_8001 pixel_8001/gring pixel_8001/VDD pixel_8001/GND pixel_8001/VREF pixel_8001/ROW_SEL
+ pixel_8001/NB1 pixel_8001/VBIAS pixel_8001/NB2 pixel_8001/AMP_IN pixel_8001/SF_IB
+ pixel_8001/PIX_OUT pixel_8001/CSA_VREF pixel
Xpixel_8012 pixel_8012/gring pixel_8012/VDD pixel_8012/GND pixel_8012/VREF pixel_8012/ROW_SEL
+ pixel_8012/NB1 pixel_8012/VBIAS pixel_8012/NB2 pixel_8012/AMP_IN pixel_8012/SF_IB
+ pixel_8012/PIX_OUT pixel_8012/CSA_VREF pixel
Xpixel_8023 pixel_8023/gring pixel_8023/VDD pixel_8023/GND pixel_8023/VREF pixel_8023/ROW_SEL
+ pixel_8023/NB1 pixel_8023/VBIAS pixel_8023/NB2 pixel_8023/AMP_IN pixel_8023/SF_IB
+ pixel_8023/PIX_OUT pixel_8023/CSA_VREF pixel
Xpixel_8034 pixel_8034/gring pixel_8034/VDD pixel_8034/GND pixel_8034/VREF pixel_8034/ROW_SEL
+ pixel_8034/NB1 pixel_8034/VBIAS pixel_8034/NB2 pixel_8034/AMP_IN pixel_8034/SF_IB
+ pixel_8034/PIX_OUT pixel_8034/CSA_VREF pixel
Xpixel_8045 pixel_8045/gring pixel_8045/VDD pixel_8045/GND pixel_8045/VREF pixel_8045/ROW_SEL
+ pixel_8045/NB1 pixel_8045/VBIAS pixel_8045/NB2 pixel_8045/AMP_IN pixel_8045/SF_IB
+ pixel_8045/PIX_OUT pixel_8045/CSA_VREF pixel
Xpixel_8056 pixel_8056/gring pixel_8056/VDD pixel_8056/GND pixel_8056/VREF pixel_8056/ROW_SEL
+ pixel_8056/NB1 pixel_8056/VBIAS pixel_8056/NB2 pixel_8056/AMP_IN pixel_8056/SF_IB
+ pixel_8056/PIX_OUT pixel_8056/CSA_VREF pixel
Xpixel_8067 pixel_8067/gring pixel_8067/VDD pixel_8067/GND pixel_8067/VREF pixel_8067/ROW_SEL
+ pixel_8067/NB1 pixel_8067/VBIAS pixel_8067/NB2 pixel_8067/AMP_IN pixel_8067/SF_IB
+ pixel_8067/PIX_OUT pixel_8067/CSA_VREF pixel
Xpixel_7300 pixel_7300/gring pixel_7300/VDD pixel_7300/GND pixel_7300/VREF pixel_7300/ROW_SEL
+ pixel_7300/NB1 pixel_7300/VBIAS pixel_7300/NB2 pixel_7300/AMP_IN pixel_7300/SF_IB
+ pixel_7300/PIX_OUT pixel_7300/CSA_VREF pixel
Xpixel_7311 pixel_7311/gring pixel_7311/VDD pixel_7311/GND pixel_7311/VREF pixel_7311/ROW_SEL
+ pixel_7311/NB1 pixel_7311/VBIAS pixel_7311/NB2 pixel_7311/AMP_IN pixel_7311/SF_IB
+ pixel_7311/PIX_OUT pixel_7311/CSA_VREF pixel
Xpixel_7322 pixel_7322/gring pixel_7322/VDD pixel_7322/GND pixel_7322/VREF pixel_7322/ROW_SEL
+ pixel_7322/NB1 pixel_7322/VBIAS pixel_7322/NB2 pixel_7322/AMP_IN pixel_7322/SF_IB
+ pixel_7322/PIX_OUT pixel_7322/CSA_VREF pixel
Xpixel_8078 pixel_8078/gring pixel_8078/VDD pixel_8078/GND pixel_8078/VREF pixel_8078/ROW_SEL
+ pixel_8078/NB1 pixel_8078/VBIAS pixel_8078/NB2 pixel_8078/AMP_IN pixel_8078/SF_IB
+ pixel_8078/PIX_OUT pixel_8078/CSA_VREF pixel
Xpixel_8089 pixel_8089/gring pixel_8089/VDD pixel_8089/GND pixel_8089/VREF pixel_8089/ROW_SEL
+ pixel_8089/NB1 pixel_8089/VBIAS pixel_8089/NB2 pixel_8089/AMP_IN pixel_8089/SF_IB
+ pixel_8089/PIX_OUT pixel_8089/CSA_VREF pixel
Xpixel_7333 pixel_7333/gring pixel_7333/VDD pixel_7333/GND pixel_7333/VREF pixel_7333/ROW_SEL
+ pixel_7333/NB1 pixel_7333/VBIAS pixel_7333/NB2 pixel_7333/AMP_IN pixel_7333/SF_IB
+ pixel_7333/PIX_OUT pixel_7333/CSA_VREF pixel
Xpixel_7344 pixel_7344/gring pixel_7344/VDD pixel_7344/GND pixel_7344/VREF pixel_7344/ROW_SEL
+ pixel_7344/NB1 pixel_7344/VBIAS pixel_7344/NB2 pixel_7344/AMP_IN pixel_7344/SF_IB
+ pixel_7344/PIX_OUT pixel_7344/CSA_VREF pixel
Xpixel_7355 pixel_7355/gring pixel_7355/VDD pixel_7355/GND pixel_7355/VREF pixel_7355/ROW_SEL
+ pixel_7355/NB1 pixel_7355/VBIAS pixel_7355/NB2 pixel_7355/AMP_IN pixel_7355/SF_IB
+ pixel_7355/PIX_OUT pixel_7355/CSA_VREF pixel
Xpixel_7366 pixel_7366/gring pixel_7366/VDD pixel_7366/GND pixel_7366/VREF pixel_7366/ROW_SEL
+ pixel_7366/NB1 pixel_7366/VBIAS pixel_7366/NB2 pixel_7366/AMP_IN pixel_7366/SF_IB
+ pixel_7366/PIX_OUT pixel_7366/CSA_VREF pixel
Xpixel_6610 pixel_6610/gring pixel_6610/VDD pixel_6610/GND pixel_6610/VREF pixel_6610/ROW_SEL
+ pixel_6610/NB1 pixel_6610/VBIAS pixel_6610/NB2 pixel_6610/AMP_IN pixel_6610/SF_IB
+ pixel_6610/PIX_OUT pixel_6610/CSA_VREF pixel
Xpixel_6621 pixel_6621/gring pixel_6621/VDD pixel_6621/GND pixel_6621/VREF pixel_6621/ROW_SEL
+ pixel_6621/NB1 pixel_6621/VBIAS pixel_6621/NB2 pixel_6621/AMP_IN pixel_6621/SF_IB
+ pixel_6621/PIX_OUT pixel_6621/CSA_VREF pixel
Xpixel_7377 pixel_7377/gring pixel_7377/VDD pixel_7377/GND pixel_7377/VREF pixel_7377/ROW_SEL
+ pixel_7377/NB1 pixel_7377/VBIAS pixel_7377/NB2 pixel_7377/AMP_IN pixel_7377/SF_IB
+ pixel_7377/PIX_OUT pixel_7377/CSA_VREF pixel
Xpixel_7388 pixel_7388/gring pixel_7388/VDD pixel_7388/GND pixel_7388/VREF pixel_7388/ROW_SEL
+ pixel_7388/NB1 pixel_7388/VBIAS pixel_7388/NB2 pixel_7388/AMP_IN pixel_7388/SF_IB
+ pixel_7388/PIX_OUT pixel_7388/CSA_VREF pixel
Xpixel_7399 pixel_7399/gring pixel_7399/VDD pixel_7399/GND pixel_7399/VREF pixel_7399/ROW_SEL
+ pixel_7399/NB1 pixel_7399/VBIAS pixel_7399/NB2 pixel_7399/AMP_IN pixel_7399/SF_IB
+ pixel_7399/PIX_OUT pixel_7399/CSA_VREF pixel
Xpixel_6632 pixel_6632/gring pixel_6632/VDD pixel_6632/GND pixel_6632/VREF pixel_6632/ROW_SEL
+ pixel_6632/NB1 pixel_6632/VBIAS pixel_6632/NB2 pixel_6632/AMP_IN pixel_6632/SF_IB
+ pixel_6632/PIX_OUT pixel_6632/CSA_VREF pixel
Xpixel_6643 pixel_6643/gring pixel_6643/VDD pixel_6643/GND pixel_6643/VREF pixel_6643/ROW_SEL
+ pixel_6643/NB1 pixel_6643/VBIAS pixel_6643/NB2 pixel_6643/AMP_IN pixel_6643/SF_IB
+ pixel_6643/PIX_OUT pixel_6643/CSA_VREF pixel
Xpixel_6654 pixel_6654/gring pixel_6654/VDD pixel_6654/GND pixel_6654/VREF pixel_6654/ROW_SEL
+ pixel_6654/NB1 pixel_6654/VBIAS pixel_6654/NB2 pixel_6654/AMP_IN pixel_6654/SF_IB
+ pixel_6654/PIX_OUT pixel_6654/CSA_VREF pixel
Xpixel_6665 pixel_6665/gring pixel_6665/VDD pixel_6665/GND pixel_6665/VREF pixel_6665/ROW_SEL
+ pixel_6665/NB1 pixel_6665/VBIAS pixel_6665/NB2 pixel_6665/AMP_IN pixel_6665/SF_IB
+ pixel_6665/PIX_OUT pixel_6665/CSA_VREF pixel
Xpixel_6676 pixel_6676/gring pixel_6676/VDD pixel_6676/GND pixel_6676/VREF pixel_6676/ROW_SEL
+ pixel_6676/NB1 pixel_6676/VBIAS pixel_6676/NB2 pixel_6676/AMP_IN pixel_6676/SF_IB
+ pixel_6676/PIX_OUT pixel_6676/CSA_VREF pixel
Xpixel_6687 pixel_6687/gring pixel_6687/VDD pixel_6687/GND pixel_6687/VREF pixel_6687/ROW_SEL
+ pixel_6687/NB1 pixel_6687/VBIAS pixel_6687/NB2 pixel_6687/AMP_IN pixel_6687/SF_IB
+ pixel_6687/PIX_OUT pixel_6687/CSA_VREF pixel
Xpixel_5920 pixel_5920/gring pixel_5920/VDD pixel_5920/GND pixel_5920/VREF pixel_5920/ROW_SEL
+ pixel_5920/NB1 pixel_5920/VBIAS pixel_5920/NB2 pixel_5920/AMP_IN pixel_5920/SF_IB
+ pixel_5920/PIX_OUT pixel_5920/CSA_VREF pixel
Xpixel_5931 pixel_5931/gring pixel_5931/VDD pixel_5931/GND pixel_5931/VREF pixel_5931/ROW_SEL
+ pixel_5931/NB1 pixel_5931/VBIAS pixel_5931/NB2 pixel_5931/AMP_IN pixel_5931/SF_IB
+ pixel_5931/PIX_OUT pixel_5931/CSA_VREF pixel
Xpixel_5942 pixel_5942/gring pixel_5942/VDD pixel_5942/GND pixel_5942/VREF pixel_5942/ROW_SEL
+ pixel_5942/NB1 pixel_5942/VBIAS pixel_5942/NB2 pixel_5942/AMP_IN pixel_5942/SF_IB
+ pixel_5942/PIX_OUT pixel_5942/CSA_VREF pixel
Xpixel_6698 pixel_6698/gring pixel_6698/VDD pixel_6698/GND pixel_6698/VREF pixel_6698/ROW_SEL
+ pixel_6698/NB1 pixel_6698/VBIAS pixel_6698/NB2 pixel_6698/AMP_IN pixel_6698/SF_IB
+ pixel_6698/PIX_OUT pixel_6698/CSA_VREF pixel
Xpixel_5953 pixel_5953/gring pixel_5953/VDD pixel_5953/GND pixel_5953/VREF pixel_5953/ROW_SEL
+ pixel_5953/NB1 pixel_5953/VBIAS pixel_5953/NB2 pixel_5953/AMP_IN pixel_5953/SF_IB
+ pixel_5953/PIX_OUT pixel_5953/CSA_VREF pixel
Xpixel_5964 pixel_5964/gring pixel_5964/VDD pixel_5964/GND pixel_5964/VREF pixel_5964/ROW_SEL
+ pixel_5964/NB1 pixel_5964/VBIAS pixel_5964/NB2 pixel_5964/AMP_IN pixel_5964/SF_IB
+ pixel_5964/PIX_OUT pixel_5964/CSA_VREF pixel
Xpixel_5975 pixel_5975/gring pixel_5975/VDD pixel_5975/GND pixel_5975/VREF pixel_5975/ROW_SEL
+ pixel_5975/NB1 pixel_5975/VBIAS pixel_5975/NB2 pixel_5975/AMP_IN pixel_5975/SF_IB
+ pixel_5975/PIX_OUT pixel_5975/CSA_VREF pixel
Xpixel_5986 pixel_5986/gring pixel_5986/VDD pixel_5986/GND pixel_5986/VREF pixel_5986/ROW_SEL
+ pixel_5986/NB1 pixel_5986/VBIAS pixel_5986/NB2 pixel_5986/AMP_IN pixel_5986/SF_IB
+ pixel_5986/PIX_OUT pixel_5986/CSA_VREF pixel
Xpixel_5997 pixel_5997/gring pixel_5997/VDD pixel_5997/GND pixel_5997/VREF pixel_5997/ROW_SEL
+ pixel_5997/NB1 pixel_5997/VBIAS pixel_5997/NB2 pixel_5997/AMP_IN pixel_5997/SF_IB
+ pixel_5997/PIX_OUT pixel_5997/CSA_VREF pixel
Xpixel_9291 pixel_9291/gring pixel_9291/VDD pixel_9291/GND pixel_9291/VREF pixel_9291/ROW_SEL
+ pixel_9291/NB1 pixel_9291/VBIAS pixel_9291/NB2 pixel_9291/AMP_IN pixel_9291/SF_IB
+ pixel_9291/PIX_OUT pixel_9291/CSA_VREF pixel
Xpixel_9280 pixel_9280/gring pixel_9280/VDD pixel_9280/GND pixel_9280/VREF pixel_9280/ROW_SEL
+ pixel_9280/NB1 pixel_9280/VBIAS pixel_9280/NB2 pixel_9280/AMP_IN pixel_9280/SF_IB
+ pixel_9280/PIX_OUT pixel_9280/CSA_VREF pixel
Xpixel_8590 pixel_8590/gring pixel_8590/VDD pixel_8590/GND pixel_8590/VREF pixel_8590/ROW_SEL
+ pixel_8590/NB1 pixel_8590/VBIAS pixel_8590/NB2 pixel_8590/AMP_IN pixel_8590/SF_IB
+ pixel_8590/PIX_OUT pixel_8590/CSA_VREF pixel
Xpixel_5205 pixel_5205/gring pixel_5205/VDD pixel_5205/GND pixel_5205/VREF pixel_5205/ROW_SEL
+ pixel_5205/NB1 pixel_5205/VBIAS pixel_5205/NB2 pixel_5205/AMP_IN pixel_5205/SF_IB
+ pixel_5205/PIX_OUT pixel_5205/CSA_VREF pixel
Xpixel_5216 pixel_5216/gring pixel_5216/VDD pixel_5216/GND pixel_5216/VREF pixel_5216/ROW_SEL
+ pixel_5216/NB1 pixel_5216/VBIAS pixel_5216/NB2 pixel_5216/AMP_IN pixel_5216/SF_IB
+ pixel_5216/PIX_OUT pixel_5216/CSA_VREF pixel
Xpixel_5227 pixel_5227/gring pixel_5227/VDD pixel_5227/GND pixel_5227/VREF pixel_5227/ROW_SEL
+ pixel_5227/NB1 pixel_5227/VBIAS pixel_5227/NB2 pixel_5227/AMP_IN pixel_5227/SF_IB
+ pixel_5227/PIX_OUT pixel_5227/CSA_VREF pixel
Xpixel_5238 pixel_5238/gring pixel_5238/VDD pixel_5238/GND pixel_5238/VREF pixel_5238/ROW_SEL
+ pixel_5238/NB1 pixel_5238/VBIAS pixel_5238/NB2 pixel_5238/AMP_IN pixel_5238/SF_IB
+ pixel_5238/PIX_OUT pixel_5238/CSA_VREF pixel
Xpixel_532 pixel_532/gring pixel_532/VDD pixel_532/GND pixel_532/VREF pixel_532/ROW_SEL
+ pixel_532/NB1 pixel_532/VBIAS pixel_532/NB2 pixel_532/AMP_IN pixel_532/SF_IB pixel_532/PIX_OUT
+ pixel_532/CSA_VREF pixel
Xpixel_521 pixel_521/gring pixel_521/VDD pixel_521/GND pixel_521/VREF pixel_521/ROW_SEL
+ pixel_521/NB1 pixel_521/VBIAS pixel_521/NB2 pixel_521/AMP_IN pixel_521/SF_IB pixel_521/PIX_OUT
+ pixel_521/CSA_VREF pixel
Xpixel_510 pixel_510/gring pixel_510/VDD pixel_510/GND pixel_510/VREF pixel_510/ROW_SEL
+ pixel_510/NB1 pixel_510/VBIAS pixel_510/NB2 pixel_510/AMP_IN pixel_510/SF_IB pixel_510/PIX_OUT
+ pixel_510/CSA_VREF pixel
Xpixel_5249 pixel_5249/gring pixel_5249/VDD pixel_5249/GND pixel_5249/VREF pixel_5249/ROW_SEL
+ pixel_5249/NB1 pixel_5249/VBIAS pixel_5249/NB2 pixel_5249/AMP_IN pixel_5249/SF_IB
+ pixel_5249/PIX_OUT pixel_5249/CSA_VREF pixel
Xpixel_4504 pixel_4504/gring pixel_4504/VDD pixel_4504/GND pixel_4504/VREF pixel_4504/ROW_SEL
+ pixel_4504/NB1 pixel_4504/VBIAS pixel_4504/NB2 pixel_4504/AMP_IN pixel_4504/SF_IB
+ pixel_4504/PIX_OUT pixel_4504/CSA_VREF pixel
Xpixel_4515 pixel_4515/gring pixel_4515/VDD pixel_4515/GND pixel_4515/VREF pixel_4515/ROW_SEL
+ pixel_4515/NB1 pixel_4515/VBIAS pixel_4515/NB2 pixel_4515/AMP_IN pixel_4515/SF_IB
+ pixel_4515/PIX_OUT pixel_4515/CSA_VREF pixel
Xpixel_4526 pixel_4526/gring pixel_4526/VDD pixel_4526/GND pixel_4526/VREF pixel_4526/ROW_SEL
+ pixel_4526/NB1 pixel_4526/VBIAS pixel_4526/NB2 pixel_4526/AMP_IN pixel_4526/SF_IB
+ pixel_4526/PIX_OUT pixel_4526/CSA_VREF pixel
Xpixel_4537 pixel_4537/gring pixel_4537/VDD pixel_4537/GND pixel_4537/VREF pixel_4537/ROW_SEL
+ pixel_4537/NB1 pixel_4537/VBIAS pixel_4537/NB2 pixel_4537/AMP_IN pixel_4537/SF_IB
+ pixel_4537/PIX_OUT pixel_4537/CSA_VREF pixel
Xpixel_565 pixel_565/gring pixel_565/VDD pixel_565/GND pixel_565/VREF pixel_565/ROW_SEL
+ pixel_565/NB1 pixel_565/VBIAS pixel_565/NB2 pixel_565/AMP_IN pixel_565/SF_IB pixel_565/PIX_OUT
+ pixel_565/CSA_VREF pixel
Xpixel_554 pixel_554/gring pixel_554/VDD pixel_554/GND pixel_554/VREF pixel_554/ROW_SEL
+ pixel_554/NB1 pixel_554/VBIAS pixel_554/NB2 pixel_554/AMP_IN pixel_554/SF_IB pixel_554/PIX_OUT
+ pixel_554/CSA_VREF pixel
Xpixel_543 pixel_543/gring pixel_543/VDD pixel_543/GND pixel_543/VREF pixel_543/ROW_SEL
+ pixel_543/NB1 pixel_543/VBIAS pixel_543/NB2 pixel_543/AMP_IN pixel_543/SF_IB pixel_543/PIX_OUT
+ pixel_543/CSA_VREF pixel
Xpixel_4548 pixel_4548/gring pixel_4548/VDD pixel_4548/GND pixel_4548/VREF pixel_4548/ROW_SEL
+ pixel_4548/NB1 pixel_4548/VBIAS pixel_4548/NB2 pixel_4548/AMP_IN pixel_4548/SF_IB
+ pixel_4548/PIX_OUT pixel_4548/CSA_VREF pixel
Xpixel_4559 pixel_4559/gring pixel_4559/VDD pixel_4559/GND pixel_4559/VREF pixel_4559/ROW_SEL
+ pixel_4559/NB1 pixel_4559/VBIAS pixel_4559/NB2 pixel_4559/AMP_IN pixel_4559/SF_IB
+ pixel_4559/PIX_OUT pixel_4559/CSA_VREF pixel
Xpixel_3803 pixel_3803/gring pixel_3803/VDD pixel_3803/GND pixel_3803/VREF pixel_3803/ROW_SEL
+ pixel_3803/NB1 pixel_3803/VBIAS pixel_3803/NB2 pixel_3803/AMP_IN pixel_3803/SF_IB
+ pixel_3803/PIX_OUT pixel_3803/CSA_VREF pixel
Xpixel_3814 pixel_3814/gring pixel_3814/VDD pixel_3814/GND pixel_3814/VREF pixel_3814/ROW_SEL
+ pixel_3814/NB1 pixel_3814/VBIAS pixel_3814/NB2 pixel_3814/AMP_IN pixel_3814/SF_IB
+ pixel_3814/PIX_OUT pixel_3814/CSA_VREF pixel
Xpixel_3825 pixel_3825/gring pixel_3825/VDD pixel_3825/GND pixel_3825/VREF pixel_3825/ROW_SEL
+ pixel_3825/NB1 pixel_3825/VBIAS pixel_3825/NB2 pixel_3825/AMP_IN pixel_3825/SF_IB
+ pixel_3825/PIX_OUT pixel_3825/CSA_VREF pixel
Xpixel_598 pixel_598/gring pixel_598/VDD pixel_598/GND pixel_598/VREF pixel_598/ROW_SEL
+ pixel_598/NB1 pixel_598/VBIAS pixel_598/NB2 pixel_598/AMP_IN pixel_598/SF_IB pixel_598/PIX_OUT
+ pixel_598/CSA_VREF pixel
Xpixel_587 pixel_587/gring pixel_587/VDD pixel_587/GND pixel_587/VREF pixel_587/ROW_SEL
+ pixel_587/NB1 pixel_587/VBIAS pixel_587/NB2 pixel_587/AMP_IN pixel_587/SF_IB pixel_587/PIX_OUT
+ pixel_587/CSA_VREF pixel
Xpixel_576 pixel_576/gring pixel_576/VDD pixel_576/GND pixel_576/VREF pixel_576/ROW_SEL
+ pixel_576/NB1 pixel_576/VBIAS pixel_576/NB2 pixel_576/AMP_IN pixel_576/SF_IB pixel_576/PIX_OUT
+ pixel_576/CSA_VREF pixel
Xpixel_3858 pixel_3858/gring pixel_3858/VDD pixel_3858/GND pixel_3858/VREF pixel_3858/ROW_SEL
+ pixel_3858/NB1 pixel_3858/VBIAS pixel_3858/NB2 pixel_3858/AMP_IN pixel_3858/SF_IB
+ pixel_3858/PIX_OUT pixel_3858/CSA_VREF pixel
Xpixel_3847 pixel_3847/gring pixel_3847/VDD pixel_3847/GND pixel_3847/VREF pixel_3847/ROW_SEL
+ pixel_3847/NB1 pixel_3847/VBIAS pixel_3847/NB2 pixel_3847/AMP_IN pixel_3847/SF_IB
+ pixel_3847/PIX_OUT pixel_3847/CSA_VREF pixel
Xpixel_3836 pixel_3836/gring pixel_3836/VDD pixel_3836/GND pixel_3836/VREF pixel_3836/ROW_SEL
+ pixel_3836/NB1 pixel_3836/VBIAS pixel_3836/NB2 pixel_3836/AMP_IN pixel_3836/SF_IB
+ pixel_3836/PIX_OUT pixel_3836/CSA_VREF pixel
Xpixel_3869 pixel_3869/gring pixel_3869/VDD pixel_3869/GND pixel_3869/VREF pixel_3869/ROW_SEL
+ pixel_3869/NB1 pixel_3869/VBIAS pixel_3869/NB2 pixel_3869/AMP_IN pixel_3869/SF_IB
+ pixel_3869/PIX_OUT pixel_3869/CSA_VREF pixel
Xpixel_7130 pixel_7130/gring pixel_7130/VDD pixel_7130/GND pixel_7130/VREF pixel_7130/ROW_SEL
+ pixel_7130/NB1 pixel_7130/VBIAS pixel_7130/NB2 pixel_7130/AMP_IN pixel_7130/SF_IB
+ pixel_7130/PIX_OUT pixel_7130/CSA_VREF pixel
Xpixel_7141 pixel_7141/gring pixel_7141/VDD pixel_7141/GND pixel_7141/VREF pixel_7141/ROW_SEL
+ pixel_7141/NB1 pixel_7141/VBIAS pixel_7141/NB2 pixel_7141/AMP_IN pixel_7141/SF_IB
+ pixel_7141/PIX_OUT pixel_7141/CSA_VREF pixel
Xpixel_7152 pixel_7152/gring pixel_7152/VDD pixel_7152/GND pixel_7152/VREF pixel_7152/ROW_SEL
+ pixel_7152/NB1 pixel_7152/VBIAS pixel_7152/NB2 pixel_7152/AMP_IN pixel_7152/SF_IB
+ pixel_7152/PIX_OUT pixel_7152/CSA_VREF pixel
Xpixel_7163 pixel_7163/gring pixel_7163/VDD pixel_7163/GND pixel_7163/VREF pixel_7163/ROW_SEL
+ pixel_7163/NB1 pixel_7163/VBIAS pixel_7163/NB2 pixel_7163/AMP_IN pixel_7163/SF_IB
+ pixel_7163/PIX_OUT pixel_7163/CSA_VREF pixel
Xpixel_7174 pixel_7174/gring pixel_7174/VDD pixel_7174/GND pixel_7174/VREF pixel_7174/ROW_SEL
+ pixel_7174/NB1 pixel_7174/VBIAS pixel_7174/NB2 pixel_7174/AMP_IN pixel_7174/SF_IB
+ pixel_7174/PIX_OUT pixel_7174/CSA_VREF pixel
Xpixel_7185 pixel_7185/gring pixel_7185/VDD pixel_7185/GND pixel_7185/VREF pixel_7185/ROW_SEL
+ pixel_7185/NB1 pixel_7185/VBIAS pixel_7185/NB2 pixel_7185/AMP_IN pixel_7185/SF_IB
+ pixel_7185/PIX_OUT pixel_7185/CSA_VREF pixel
Xpixel_7196 pixel_7196/gring pixel_7196/VDD pixel_7196/GND pixel_7196/VREF pixel_7196/ROW_SEL
+ pixel_7196/NB1 pixel_7196/VBIAS pixel_7196/NB2 pixel_7196/AMP_IN pixel_7196/SF_IB
+ pixel_7196/PIX_OUT pixel_7196/CSA_VREF pixel
Xpixel_6440 pixel_6440/gring pixel_6440/VDD pixel_6440/GND pixel_6440/VREF pixel_6440/ROW_SEL
+ pixel_6440/NB1 pixel_6440/VBIAS pixel_6440/NB2 pixel_6440/AMP_IN pixel_6440/SF_IB
+ pixel_6440/PIX_OUT pixel_6440/CSA_VREF pixel
Xpixel_6451 pixel_6451/gring pixel_6451/VDD pixel_6451/GND pixel_6451/VREF pixel_6451/ROW_SEL
+ pixel_6451/NB1 pixel_6451/VBIAS pixel_6451/NB2 pixel_6451/AMP_IN pixel_6451/SF_IB
+ pixel_6451/PIX_OUT pixel_6451/CSA_VREF pixel
Xpixel_6462 pixel_6462/gring pixel_6462/VDD pixel_6462/GND pixel_6462/VREF pixel_6462/ROW_SEL
+ pixel_6462/NB1 pixel_6462/VBIAS pixel_6462/NB2 pixel_6462/AMP_IN pixel_6462/SF_IB
+ pixel_6462/PIX_OUT pixel_6462/CSA_VREF pixel
Xpixel_6473 pixel_6473/gring pixel_6473/VDD pixel_6473/GND pixel_6473/VREF pixel_6473/ROW_SEL
+ pixel_6473/NB1 pixel_6473/VBIAS pixel_6473/NB2 pixel_6473/AMP_IN pixel_6473/SF_IB
+ pixel_6473/PIX_OUT pixel_6473/CSA_VREF pixel
Xpixel_6484 pixel_6484/gring pixel_6484/VDD pixel_6484/GND pixel_6484/VREF pixel_6484/ROW_SEL
+ pixel_6484/NB1 pixel_6484/VBIAS pixel_6484/NB2 pixel_6484/AMP_IN pixel_6484/SF_IB
+ pixel_6484/PIX_OUT pixel_6484/CSA_VREF pixel
Xpixel_6495 pixel_6495/gring pixel_6495/VDD pixel_6495/GND pixel_6495/VREF pixel_6495/ROW_SEL
+ pixel_6495/NB1 pixel_6495/VBIAS pixel_6495/NB2 pixel_6495/AMP_IN pixel_6495/SF_IB
+ pixel_6495/PIX_OUT pixel_6495/CSA_VREF pixel
Xpixel_5750 pixel_5750/gring pixel_5750/VDD pixel_5750/GND pixel_5750/VREF pixel_5750/ROW_SEL
+ pixel_5750/NB1 pixel_5750/VBIAS pixel_5750/NB2 pixel_5750/AMP_IN pixel_5750/SF_IB
+ pixel_5750/PIX_OUT pixel_5750/CSA_VREF pixel
Xpixel_5761 pixel_5761/gring pixel_5761/VDD pixel_5761/GND pixel_5761/VREF pixel_5761/ROW_SEL
+ pixel_5761/NB1 pixel_5761/VBIAS pixel_5761/NB2 pixel_5761/AMP_IN pixel_5761/SF_IB
+ pixel_5761/PIX_OUT pixel_5761/CSA_VREF pixel
Xpixel_5772 pixel_5772/gring pixel_5772/VDD pixel_5772/GND pixel_5772/VREF pixel_5772/ROW_SEL
+ pixel_5772/NB1 pixel_5772/VBIAS pixel_5772/NB2 pixel_5772/AMP_IN pixel_5772/SF_IB
+ pixel_5772/PIX_OUT pixel_5772/CSA_VREF pixel
Xpixel_5783 pixel_5783/gring pixel_5783/VDD pixel_5783/GND pixel_5783/VREF pixel_5783/ROW_SEL
+ pixel_5783/NB1 pixel_5783/VBIAS pixel_5783/NB2 pixel_5783/AMP_IN pixel_5783/SF_IB
+ pixel_5783/PIX_OUT pixel_5783/CSA_VREF pixel
Xpixel_5794 pixel_5794/gring pixel_5794/VDD pixel_5794/GND pixel_5794/VREF pixel_5794/ROW_SEL
+ pixel_5794/NB1 pixel_5794/VBIAS pixel_5794/NB2 pixel_5794/AMP_IN pixel_5794/SF_IB
+ pixel_5794/PIX_OUT pixel_5794/CSA_VREF pixel
Xpixel_2409 pixel_2409/gring pixel_2409/VDD pixel_2409/GND pixel_2409/VREF pixel_2409/ROW_SEL
+ pixel_2409/NB1 pixel_2409/VBIAS pixel_2409/NB2 pixel_2409/AMP_IN pixel_2409/SF_IB
+ pixel_2409/PIX_OUT pixel_2409/CSA_VREF pixel
Xpixel_1708 pixel_1708/gring pixel_1708/VDD pixel_1708/GND pixel_1708/VREF pixel_1708/ROW_SEL
+ pixel_1708/NB1 pixel_1708/VBIAS pixel_1708/NB2 pixel_1708/AMP_IN pixel_1708/SF_IB
+ pixel_1708/PIX_OUT pixel_1708/CSA_VREF pixel
Xpixel_1719 pixel_1719/gring pixel_1719/VDD pixel_1719/GND pixel_1719/VREF pixel_1719/ROW_SEL
+ pixel_1719/NB1 pixel_1719/VBIAS pixel_1719/NB2 pixel_1719/AMP_IN pixel_1719/SF_IB
+ pixel_1719/PIX_OUT pixel_1719/CSA_VREF pixel
Xpixel_5002 pixel_5002/gring pixel_5002/VDD pixel_5002/GND pixel_5002/VREF pixel_5002/ROW_SEL
+ pixel_5002/NB1 pixel_5002/VBIAS pixel_5002/NB2 pixel_5002/AMP_IN pixel_5002/SF_IB
+ pixel_5002/PIX_OUT pixel_5002/CSA_VREF pixel
Xpixel_5013 pixel_5013/gring pixel_5013/VDD pixel_5013/GND pixel_5013/VREF pixel_5013/ROW_SEL
+ pixel_5013/NB1 pixel_5013/VBIAS pixel_5013/NB2 pixel_5013/AMP_IN pixel_5013/SF_IB
+ pixel_5013/PIX_OUT pixel_5013/CSA_VREF pixel
Xpixel_5024 pixel_5024/gring pixel_5024/VDD pixel_5024/GND pixel_5024/VREF pixel_5024/ROW_SEL
+ pixel_5024/NB1 pixel_5024/VBIAS pixel_5024/NB2 pixel_5024/AMP_IN pixel_5024/SF_IB
+ pixel_5024/PIX_OUT pixel_5024/CSA_VREF pixel
Xpixel_5035 pixel_5035/gring pixel_5035/VDD pixel_5035/GND pixel_5035/VREF pixel_5035/ROW_SEL
+ pixel_5035/NB1 pixel_5035/VBIAS pixel_5035/NB2 pixel_5035/AMP_IN pixel_5035/SF_IB
+ pixel_5035/PIX_OUT pixel_5035/CSA_VREF pixel
Xpixel_5046 pixel_5046/gring pixel_5046/VDD pixel_5046/GND pixel_5046/VREF pixel_5046/ROW_SEL
+ pixel_5046/NB1 pixel_5046/VBIAS pixel_5046/NB2 pixel_5046/AMP_IN pixel_5046/SF_IB
+ pixel_5046/PIX_OUT pixel_5046/CSA_VREF pixel
Xpixel_4301 pixel_4301/gring pixel_4301/VDD pixel_4301/GND pixel_4301/VREF pixel_4301/ROW_SEL
+ pixel_4301/NB1 pixel_4301/VBIAS pixel_4301/NB2 pixel_4301/AMP_IN pixel_4301/SF_IB
+ pixel_4301/PIX_OUT pixel_4301/CSA_VREF pixel
Xpixel_340 pixel_340/gring pixel_340/VDD pixel_340/GND pixel_340/VREF pixel_340/ROW_SEL
+ pixel_340/NB1 pixel_340/VBIAS pixel_340/NB2 pixel_340/AMP_IN pixel_340/SF_IB pixel_340/PIX_OUT
+ pixel_340/CSA_VREF pixel
Xpixel_3600 pixel_3600/gring pixel_3600/VDD pixel_3600/GND pixel_3600/VREF pixel_3600/ROW_SEL
+ pixel_3600/NB1 pixel_3600/VBIAS pixel_3600/NB2 pixel_3600/AMP_IN pixel_3600/SF_IB
+ pixel_3600/PIX_OUT pixel_3600/CSA_VREF pixel
Xpixel_5057 pixel_5057/gring pixel_5057/VDD pixel_5057/GND pixel_5057/VREF pixel_5057/ROW_SEL
+ pixel_5057/NB1 pixel_5057/VBIAS pixel_5057/NB2 pixel_5057/AMP_IN pixel_5057/SF_IB
+ pixel_5057/PIX_OUT pixel_5057/CSA_VREF pixel
Xpixel_5068 pixel_5068/gring pixel_5068/VDD pixel_5068/GND pixel_5068/VREF pixel_5068/ROW_SEL
+ pixel_5068/NB1 pixel_5068/VBIAS pixel_5068/NB2 pixel_5068/AMP_IN pixel_5068/SF_IB
+ pixel_5068/PIX_OUT pixel_5068/CSA_VREF pixel
Xpixel_5079 pixel_5079/gring pixel_5079/VDD pixel_5079/GND pixel_5079/VREF pixel_5079/ROW_SEL
+ pixel_5079/NB1 pixel_5079/VBIAS pixel_5079/NB2 pixel_5079/AMP_IN pixel_5079/SF_IB
+ pixel_5079/PIX_OUT pixel_5079/CSA_VREF pixel
Xpixel_4312 pixel_4312/gring pixel_4312/VDD pixel_4312/GND pixel_4312/VREF pixel_4312/ROW_SEL
+ pixel_4312/NB1 pixel_4312/VBIAS pixel_4312/NB2 pixel_4312/AMP_IN pixel_4312/SF_IB
+ pixel_4312/PIX_OUT pixel_4312/CSA_VREF pixel
Xpixel_4323 pixel_4323/gring pixel_4323/VDD pixel_4323/GND pixel_4323/VREF pixel_4323/ROW_SEL
+ pixel_4323/NB1 pixel_4323/VBIAS pixel_4323/NB2 pixel_4323/AMP_IN pixel_4323/SF_IB
+ pixel_4323/PIX_OUT pixel_4323/CSA_VREF pixel
Xpixel_4334 pixel_4334/gring pixel_4334/VDD pixel_4334/GND pixel_4334/VREF pixel_4334/ROW_SEL
+ pixel_4334/NB1 pixel_4334/VBIAS pixel_4334/NB2 pixel_4334/AMP_IN pixel_4334/SF_IB
+ pixel_4334/PIX_OUT pixel_4334/CSA_VREF pixel
Xpixel_4345 pixel_4345/gring pixel_4345/VDD pixel_4345/GND pixel_4345/VREF pixel_4345/ROW_SEL
+ pixel_4345/NB1 pixel_4345/VBIAS pixel_4345/NB2 pixel_4345/AMP_IN pixel_4345/SF_IB
+ pixel_4345/PIX_OUT pixel_4345/CSA_VREF pixel
Xpixel_373 pixel_373/gring pixel_373/VDD pixel_373/GND pixel_373/VREF pixel_373/ROW_SEL
+ pixel_373/NB1 pixel_373/VBIAS pixel_373/NB2 pixel_373/AMP_IN pixel_373/SF_IB pixel_373/PIX_OUT
+ pixel_373/CSA_VREF pixel
Xpixel_362 pixel_362/gring pixel_362/VDD pixel_362/GND pixel_362/VREF pixel_362/ROW_SEL
+ pixel_362/NB1 pixel_362/VBIAS pixel_362/NB2 pixel_362/AMP_IN pixel_362/SF_IB pixel_362/PIX_OUT
+ pixel_362/CSA_VREF pixel
Xpixel_351 pixel_351/gring pixel_351/VDD pixel_351/GND pixel_351/VREF pixel_351/ROW_SEL
+ pixel_351/NB1 pixel_351/VBIAS pixel_351/NB2 pixel_351/AMP_IN pixel_351/SF_IB pixel_351/PIX_OUT
+ pixel_351/CSA_VREF pixel
Xpixel_3633 pixel_3633/gring pixel_3633/VDD pixel_3633/GND pixel_3633/VREF pixel_3633/ROW_SEL
+ pixel_3633/NB1 pixel_3633/VBIAS pixel_3633/NB2 pixel_3633/AMP_IN pixel_3633/SF_IB
+ pixel_3633/PIX_OUT pixel_3633/CSA_VREF pixel
Xpixel_3622 pixel_3622/gring pixel_3622/VDD pixel_3622/GND pixel_3622/VREF pixel_3622/ROW_SEL
+ pixel_3622/NB1 pixel_3622/VBIAS pixel_3622/NB2 pixel_3622/AMP_IN pixel_3622/SF_IB
+ pixel_3622/PIX_OUT pixel_3622/CSA_VREF pixel
Xpixel_3611 pixel_3611/gring pixel_3611/VDD pixel_3611/GND pixel_3611/VREF pixel_3611/ROW_SEL
+ pixel_3611/NB1 pixel_3611/VBIAS pixel_3611/NB2 pixel_3611/AMP_IN pixel_3611/SF_IB
+ pixel_3611/PIX_OUT pixel_3611/CSA_VREF pixel
Xpixel_4356 pixel_4356/gring pixel_4356/VDD pixel_4356/GND pixel_4356/VREF pixel_4356/ROW_SEL
+ pixel_4356/NB1 pixel_4356/VBIAS pixel_4356/NB2 pixel_4356/AMP_IN pixel_4356/SF_IB
+ pixel_4356/PIX_OUT pixel_4356/CSA_VREF pixel
Xpixel_4367 pixel_4367/gring pixel_4367/VDD pixel_4367/GND pixel_4367/VREF pixel_4367/ROW_SEL
+ pixel_4367/NB1 pixel_4367/VBIAS pixel_4367/NB2 pixel_4367/AMP_IN pixel_4367/SF_IB
+ pixel_4367/PIX_OUT pixel_4367/CSA_VREF pixel
Xpixel_4378 pixel_4378/gring pixel_4378/VDD pixel_4378/GND pixel_4378/VREF pixel_4378/ROW_SEL
+ pixel_4378/NB1 pixel_4378/VBIAS pixel_4378/NB2 pixel_4378/AMP_IN pixel_4378/SF_IB
+ pixel_4378/PIX_OUT pixel_4378/CSA_VREF pixel
Xpixel_395 pixel_395/gring pixel_395/VDD pixel_395/GND pixel_395/VREF pixel_395/ROW_SEL
+ pixel_395/NB1 pixel_395/VBIAS pixel_395/NB2 pixel_395/AMP_IN pixel_395/SF_IB pixel_395/PIX_OUT
+ pixel_395/CSA_VREF pixel
Xpixel_384 pixel_384/gring pixel_384/VDD pixel_384/GND pixel_384/VREF pixel_384/ROW_SEL
+ pixel_384/NB1 pixel_384/VBIAS pixel_384/NB2 pixel_384/AMP_IN pixel_384/SF_IB pixel_384/PIX_OUT
+ pixel_384/CSA_VREF pixel
Xpixel_2932 pixel_2932/gring pixel_2932/VDD pixel_2932/GND pixel_2932/VREF pixel_2932/ROW_SEL
+ pixel_2932/NB1 pixel_2932/VBIAS pixel_2932/NB2 pixel_2932/AMP_IN pixel_2932/SF_IB
+ pixel_2932/PIX_OUT pixel_2932/CSA_VREF pixel
Xpixel_2921 pixel_2921/gring pixel_2921/VDD pixel_2921/GND pixel_2921/VREF pixel_2921/ROW_SEL
+ pixel_2921/NB1 pixel_2921/VBIAS pixel_2921/NB2 pixel_2921/AMP_IN pixel_2921/SF_IB
+ pixel_2921/PIX_OUT pixel_2921/CSA_VREF pixel
Xpixel_2910 pixel_2910/gring pixel_2910/VDD pixel_2910/GND pixel_2910/VREF pixel_2910/ROW_SEL
+ pixel_2910/NB1 pixel_2910/VBIAS pixel_2910/NB2 pixel_2910/AMP_IN pixel_2910/SF_IB
+ pixel_2910/PIX_OUT pixel_2910/CSA_VREF pixel
Xpixel_3666 pixel_3666/gring pixel_3666/VDD pixel_3666/GND pixel_3666/VREF pixel_3666/ROW_SEL
+ pixel_3666/NB1 pixel_3666/VBIAS pixel_3666/NB2 pixel_3666/AMP_IN pixel_3666/SF_IB
+ pixel_3666/PIX_OUT pixel_3666/CSA_VREF pixel
Xpixel_3655 pixel_3655/gring pixel_3655/VDD pixel_3655/GND pixel_3655/VREF pixel_3655/ROW_SEL
+ pixel_3655/NB1 pixel_3655/VBIAS pixel_3655/NB2 pixel_3655/AMP_IN pixel_3655/SF_IB
+ pixel_3655/PIX_OUT pixel_3655/CSA_VREF pixel
Xpixel_3644 pixel_3644/gring pixel_3644/VDD pixel_3644/GND pixel_3644/VREF pixel_3644/ROW_SEL
+ pixel_3644/NB1 pixel_3644/VBIAS pixel_3644/NB2 pixel_3644/AMP_IN pixel_3644/SF_IB
+ pixel_3644/PIX_OUT pixel_3644/CSA_VREF pixel
Xpixel_4389 pixel_4389/gring pixel_4389/VDD pixel_4389/GND pixel_4389/VREF pixel_4389/ROW_SEL
+ pixel_4389/NB1 pixel_4389/VBIAS pixel_4389/NB2 pixel_4389/AMP_IN pixel_4389/SF_IB
+ pixel_4389/PIX_OUT pixel_4389/CSA_VREF pixel
Xpixel_2965 pixel_2965/gring pixel_2965/VDD pixel_2965/GND pixel_2965/VREF pixel_2965/ROW_SEL
+ pixel_2965/NB1 pixel_2965/VBIAS pixel_2965/NB2 pixel_2965/AMP_IN pixel_2965/SF_IB
+ pixel_2965/PIX_OUT pixel_2965/CSA_VREF pixel
Xpixel_2954 pixel_2954/gring pixel_2954/VDD pixel_2954/GND pixel_2954/VREF pixel_2954/ROW_SEL
+ pixel_2954/NB1 pixel_2954/VBIAS pixel_2954/NB2 pixel_2954/AMP_IN pixel_2954/SF_IB
+ pixel_2954/PIX_OUT pixel_2954/CSA_VREF pixel
Xpixel_2943 pixel_2943/gring pixel_2943/VDD pixel_2943/GND pixel_2943/VREF pixel_2943/ROW_SEL
+ pixel_2943/NB1 pixel_2943/VBIAS pixel_2943/NB2 pixel_2943/AMP_IN pixel_2943/SF_IB
+ pixel_2943/PIX_OUT pixel_2943/CSA_VREF pixel
Xpixel_3699 pixel_3699/gring pixel_3699/VDD pixel_3699/GND pixel_3699/VREF pixel_3699/ROW_SEL
+ pixel_3699/NB1 pixel_3699/VBIAS pixel_3699/NB2 pixel_3699/AMP_IN pixel_3699/SF_IB
+ pixel_3699/PIX_OUT pixel_3699/CSA_VREF pixel
Xpixel_3688 pixel_3688/gring pixel_3688/VDD pixel_3688/GND pixel_3688/VREF pixel_3688/ROW_SEL
+ pixel_3688/NB1 pixel_3688/VBIAS pixel_3688/NB2 pixel_3688/AMP_IN pixel_3688/SF_IB
+ pixel_3688/PIX_OUT pixel_3688/CSA_VREF pixel
Xpixel_3677 pixel_3677/gring pixel_3677/VDD pixel_3677/GND pixel_3677/VREF pixel_3677/ROW_SEL
+ pixel_3677/NB1 pixel_3677/VBIAS pixel_3677/NB2 pixel_3677/AMP_IN pixel_3677/SF_IB
+ pixel_3677/PIX_OUT pixel_3677/CSA_VREF pixel
Xpixel_2998 pixel_2998/gring pixel_2998/VDD pixel_2998/GND pixel_2998/VREF pixel_2998/ROW_SEL
+ pixel_2998/NB1 pixel_2998/VBIAS pixel_2998/NB2 pixel_2998/AMP_IN pixel_2998/SF_IB
+ pixel_2998/PIX_OUT pixel_2998/CSA_VREF pixel
Xpixel_2987 pixel_2987/gring pixel_2987/VDD pixel_2987/GND pixel_2987/VREF pixel_2987/ROW_SEL
+ pixel_2987/NB1 pixel_2987/VBIAS pixel_2987/NB2 pixel_2987/AMP_IN pixel_2987/SF_IB
+ pixel_2987/PIX_OUT pixel_2987/CSA_VREF pixel
Xpixel_2976 pixel_2976/gring pixel_2976/VDD pixel_2976/GND pixel_2976/VREF pixel_2976/ROW_SEL
+ pixel_2976/NB1 pixel_2976/VBIAS pixel_2976/NB2 pixel_2976/AMP_IN pixel_2976/SF_IB
+ pixel_2976/PIX_OUT pixel_2976/CSA_VREF pixel
Xpixel_6270 pixel_6270/gring pixel_6270/VDD pixel_6270/GND pixel_6270/VREF pixel_6270/ROW_SEL
+ pixel_6270/NB1 pixel_6270/VBIAS pixel_6270/NB2 pixel_6270/AMP_IN pixel_6270/SF_IB
+ pixel_6270/PIX_OUT pixel_6270/CSA_VREF pixel
Xpixel_6281 pixel_6281/gring pixel_6281/VDD pixel_6281/GND pixel_6281/VREF pixel_6281/ROW_SEL
+ pixel_6281/NB1 pixel_6281/VBIAS pixel_6281/NB2 pixel_6281/AMP_IN pixel_6281/SF_IB
+ pixel_6281/PIX_OUT pixel_6281/CSA_VREF pixel
Xpixel_6292 pixel_6292/gring pixel_6292/VDD pixel_6292/GND pixel_6292/VREF pixel_6292/ROW_SEL
+ pixel_6292/NB1 pixel_6292/VBIAS pixel_6292/NB2 pixel_6292/AMP_IN pixel_6292/SF_IB
+ pixel_6292/PIX_OUT pixel_6292/CSA_VREF pixel
Xpixel_5580 pixel_5580/gring pixel_5580/VDD pixel_5580/GND pixel_5580/VREF pixel_5580/ROW_SEL
+ pixel_5580/NB1 pixel_5580/VBIAS pixel_5580/NB2 pixel_5580/AMP_IN pixel_5580/SF_IB
+ pixel_5580/PIX_OUT pixel_5580/CSA_VREF pixel
Xpixel_5591 pixel_5591/gring pixel_5591/VDD pixel_5591/GND pixel_5591/VREF pixel_5591/ROW_SEL
+ pixel_5591/NB1 pixel_5591/VBIAS pixel_5591/NB2 pixel_5591/AMP_IN pixel_5591/SF_IB
+ pixel_5591/PIX_OUT pixel_5591/CSA_VREF pixel
Xpixel_4890 pixel_4890/gring pixel_4890/VDD pixel_4890/GND pixel_4890/VREF pixel_4890/ROW_SEL
+ pixel_4890/NB1 pixel_4890/VBIAS pixel_4890/NB2 pixel_4890/AMP_IN pixel_4890/SF_IB
+ pixel_4890/PIX_OUT pixel_4890/CSA_VREF pixel
Xpixel_2217 pixel_2217/gring pixel_2217/VDD pixel_2217/GND pixel_2217/VREF pixel_2217/ROW_SEL
+ pixel_2217/NB1 pixel_2217/VBIAS pixel_2217/NB2 pixel_2217/AMP_IN pixel_2217/SF_IB
+ pixel_2217/PIX_OUT pixel_2217/CSA_VREF pixel
Xpixel_2206 pixel_2206/gring pixel_2206/VDD pixel_2206/GND pixel_2206/VREF pixel_2206/ROW_SEL
+ pixel_2206/NB1 pixel_2206/VBIAS pixel_2206/NB2 pixel_2206/AMP_IN pixel_2206/SF_IB
+ pixel_2206/PIX_OUT pixel_2206/CSA_VREF pixel
Xpixel_1516 pixel_1516/gring pixel_1516/VDD pixel_1516/GND pixel_1516/VREF pixel_1516/ROW_SEL
+ pixel_1516/NB1 pixel_1516/VBIAS pixel_1516/NB2 pixel_1516/AMP_IN pixel_1516/SF_IB
+ pixel_1516/PIX_OUT pixel_1516/CSA_VREF pixel
Xpixel_1505 pixel_1505/gring pixel_1505/VDD pixel_1505/GND pixel_1505/VREF pixel_1505/ROW_SEL
+ pixel_1505/NB1 pixel_1505/VBIAS pixel_1505/NB2 pixel_1505/AMP_IN pixel_1505/SF_IB
+ pixel_1505/PIX_OUT pixel_1505/CSA_VREF pixel
Xpixel_2239 pixel_2239/gring pixel_2239/VDD pixel_2239/GND pixel_2239/VREF pixel_2239/ROW_SEL
+ pixel_2239/NB1 pixel_2239/VBIAS pixel_2239/NB2 pixel_2239/AMP_IN pixel_2239/SF_IB
+ pixel_2239/PIX_OUT pixel_2239/CSA_VREF pixel
Xpixel_2228 pixel_2228/gring pixel_2228/VDD pixel_2228/GND pixel_2228/VREF pixel_2228/ROW_SEL
+ pixel_2228/NB1 pixel_2228/VBIAS pixel_2228/NB2 pixel_2228/AMP_IN pixel_2228/SF_IB
+ pixel_2228/PIX_OUT pixel_2228/CSA_VREF pixel
Xpixel_1549 pixel_1549/gring pixel_1549/VDD pixel_1549/GND pixel_1549/VREF pixel_1549/ROW_SEL
+ pixel_1549/NB1 pixel_1549/VBIAS pixel_1549/NB2 pixel_1549/AMP_IN pixel_1549/SF_IB
+ pixel_1549/PIX_OUT pixel_1549/CSA_VREF pixel
Xpixel_1538 pixel_1538/gring pixel_1538/VDD pixel_1538/GND pixel_1538/VREF pixel_1538/ROW_SEL
+ pixel_1538/NB1 pixel_1538/VBIAS pixel_1538/NB2 pixel_1538/AMP_IN pixel_1538/SF_IB
+ pixel_1538/PIX_OUT pixel_1538/CSA_VREF pixel
Xpixel_1527 pixel_1527/gring pixel_1527/VDD pixel_1527/GND pixel_1527/VREF pixel_1527/ROW_SEL
+ pixel_1527/NB1 pixel_1527/VBIAS pixel_1527/NB2 pixel_1527/AMP_IN pixel_1527/SF_IB
+ pixel_1527/PIX_OUT pixel_1527/CSA_VREF pixel
Xpixel_9824 pixel_9824/gring pixel_9824/VDD pixel_9824/GND pixel_9824/VREF pixel_9824/ROW_SEL
+ pixel_9824/NB1 pixel_9824/VBIAS pixel_9824/NB2 pixel_9824/AMP_IN pixel_9824/SF_IB
+ pixel_9824/PIX_OUT pixel_9824/CSA_VREF pixel
Xpixel_9813 pixel_9813/gring pixel_9813/VDD pixel_9813/GND pixel_9813/VREF pixel_9813/ROW_SEL
+ pixel_9813/NB1 pixel_9813/VBIAS pixel_9813/NB2 pixel_9813/AMP_IN pixel_9813/SF_IB
+ pixel_9813/PIX_OUT pixel_9813/CSA_VREF pixel
Xpixel_9802 pixel_9802/gring pixel_9802/VDD pixel_9802/GND pixel_9802/VREF pixel_9802/ROW_SEL
+ pixel_9802/NB1 pixel_9802/VBIAS pixel_9802/NB2 pixel_9802/AMP_IN pixel_9802/SF_IB
+ pixel_9802/PIX_OUT pixel_9802/CSA_VREF pixel
Xpixel_9846 pixel_9846/gring pixel_9846/VDD pixel_9846/GND pixel_9846/VREF pixel_9846/ROW_SEL
+ pixel_9846/NB1 pixel_9846/VBIAS pixel_9846/NB2 pixel_9846/AMP_IN pixel_9846/SF_IB
+ pixel_9846/PIX_OUT pixel_9846/CSA_VREF pixel
Xpixel_9835 pixel_9835/gring pixel_9835/VDD pixel_9835/GND pixel_9835/VREF pixel_9835/ROW_SEL
+ pixel_9835/NB1 pixel_9835/VBIAS pixel_9835/NB2 pixel_9835/AMP_IN pixel_9835/SF_IB
+ pixel_9835/PIX_OUT pixel_9835/CSA_VREF pixel
Xpixel_9857 pixel_9857/gring pixel_9857/VDD pixel_9857/GND pixel_9857/VREF pixel_9857/ROW_SEL
+ pixel_9857/NB1 pixel_9857/VBIAS pixel_9857/NB2 pixel_9857/AMP_IN pixel_9857/SF_IB
+ pixel_9857/PIX_OUT pixel_9857/CSA_VREF pixel
Xpixel_9868 pixel_9868/gring pixel_9868/VDD pixel_9868/GND pixel_9868/VREF pixel_9868/ROW_SEL
+ pixel_9868/NB1 pixel_9868/VBIAS pixel_9868/NB2 pixel_9868/AMP_IN pixel_9868/SF_IB
+ pixel_9868/PIX_OUT pixel_9868/CSA_VREF pixel
Xpixel_9879 pixel_9879/gring pixel_9879/VDD pixel_9879/GND pixel_9879/VREF pixel_9879/ROW_SEL
+ pixel_9879/NB1 pixel_9879/VBIAS pixel_9879/NB2 pixel_9879/AMP_IN pixel_9879/SF_IB
+ pixel_9879/PIX_OUT pixel_9879/CSA_VREF pixel
Xpixel_4120 pixel_4120/gring pixel_4120/VDD pixel_4120/GND pixel_4120/VREF pixel_4120/ROW_SEL
+ pixel_4120/NB1 pixel_4120/VBIAS pixel_4120/NB2 pixel_4120/AMP_IN pixel_4120/SF_IB
+ pixel_4120/PIX_OUT pixel_4120/CSA_VREF pixel
Xpixel_4131 pixel_4131/gring pixel_4131/VDD pixel_4131/GND pixel_4131/VREF pixel_4131/ROW_SEL
+ pixel_4131/NB1 pixel_4131/VBIAS pixel_4131/NB2 pixel_4131/AMP_IN pixel_4131/SF_IB
+ pixel_4131/PIX_OUT pixel_4131/CSA_VREF pixel
Xpixel_4142 pixel_4142/gring pixel_4142/VDD pixel_4142/GND pixel_4142/VREF pixel_4142/ROW_SEL
+ pixel_4142/NB1 pixel_4142/VBIAS pixel_4142/NB2 pixel_4142/AMP_IN pixel_4142/SF_IB
+ pixel_4142/PIX_OUT pixel_4142/CSA_VREF pixel
Xpixel_4153 pixel_4153/gring pixel_4153/VDD pixel_4153/GND pixel_4153/VREF pixel_4153/ROW_SEL
+ pixel_4153/NB1 pixel_4153/VBIAS pixel_4153/NB2 pixel_4153/AMP_IN pixel_4153/SF_IB
+ pixel_4153/PIX_OUT pixel_4153/CSA_VREF pixel
Xpixel_181 pixel_181/gring pixel_181/VDD pixel_181/GND pixel_181/VREF pixel_181/ROW_SEL
+ pixel_181/NB1 pixel_181/VBIAS pixel_181/NB2 pixel_181/AMP_IN pixel_181/SF_IB pixel_181/PIX_OUT
+ pixel_181/CSA_VREF pixel
Xpixel_170 pixel_170/gring pixel_170/VDD pixel_170/GND pixel_170/VREF pixel_170/ROW_SEL
+ pixel_170/NB1 pixel_170/VBIAS pixel_170/NB2 pixel_170/AMP_IN pixel_170/SF_IB pixel_170/PIX_OUT
+ pixel_170/CSA_VREF pixel
Xpixel_3441 pixel_3441/gring pixel_3441/VDD pixel_3441/GND pixel_3441/VREF pixel_3441/ROW_SEL
+ pixel_3441/NB1 pixel_3441/VBIAS pixel_3441/NB2 pixel_3441/AMP_IN pixel_3441/SF_IB
+ pixel_3441/PIX_OUT pixel_3441/CSA_VREF pixel
Xpixel_3430 pixel_3430/gring pixel_3430/VDD pixel_3430/GND pixel_3430/VREF pixel_3430/ROW_SEL
+ pixel_3430/NB1 pixel_3430/VBIAS pixel_3430/NB2 pixel_3430/AMP_IN pixel_3430/SF_IB
+ pixel_3430/PIX_OUT pixel_3430/CSA_VREF pixel
Xpixel_4164 pixel_4164/gring pixel_4164/VDD pixel_4164/GND pixel_4164/VREF pixel_4164/ROW_SEL
+ pixel_4164/NB1 pixel_4164/VBIAS pixel_4164/NB2 pixel_4164/AMP_IN pixel_4164/SF_IB
+ pixel_4164/PIX_OUT pixel_4164/CSA_VREF pixel
Xpixel_4175 pixel_4175/gring pixel_4175/VDD pixel_4175/GND pixel_4175/VREF pixel_4175/ROW_SEL
+ pixel_4175/NB1 pixel_4175/VBIAS pixel_4175/NB2 pixel_4175/AMP_IN pixel_4175/SF_IB
+ pixel_4175/PIX_OUT pixel_4175/CSA_VREF pixel
Xpixel_4186 pixel_4186/gring pixel_4186/VDD pixel_4186/GND pixel_4186/VREF pixel_4186/ROW_SEL
+ pixel_4186/NB1 pixel_4186/VBIAS pixel_4186/NB2 pixel_4186/AMP_IN pixel_4186/SF_IB
+ pixel_4186/PIX_OUT pixel_4186/CSA_VREF pixel
Xpixel_192 pixel_192/gring pixel_192/VDD pixel_192/GND pixel_192/VREF pixel_192/ROW_SEL
+ pixel_192/NB1 pixel_192/VBIAS pixel_192/NB2 pixel_192/AMP_IN pixel_192/SF_IB pixel_192/PIX_OUT
+ pixel_192/CSA_VREF pixel
Xpixel_2740 pixel_2740/gring pixel_2740/VDD pixel_2740/GND pixel_2740/VREF pixel_2740/ROW_SEL
+ pixel_2740/NB1 pixel_2740/VBIAS pixel_2740/NB2 pixel_2740/AMP_IN pixel_2740/SF_IB
+ pixel_2740/PIX_OUT pixel_2740/CSA_VREF pixel
Xpixel_3485 pixel_3485/gring pixel_3485/VDD pixel_3485/GND pixel_3485/VREF pixel_3485/ROW_SEL
+ pixel_3485/NB1 pixel_3485/VBIAS pixel_3485/NB2 pixel_3485/AMP_IN pixel_3485/SF_IB
+ pixel_3485/PIX_OUT pixel_3485/CSA_VREF pixel
Xpixel_3474 pixel_3474/gring pixel_3474/VDD pixel_3474/GND pixel_3474/VREF pixel_3474/ROW_SEL
+ pixel_3474/NB1 pixel_3474/VBIAS pixel_3474/NB2 pixel_3474/AMP_IN pixel_3474/SF_IB
+ pixel_3474/PIX_OUT pixel_3474/CSA_VREF pixel
Xpixel_3463 pixel_3463/gring pixel_3463/VDD pixel_3463/GND pixel_3463/VREF pixel_3463/ROW_SEL
+ pixel_3463/NB1 pixel_3463/VBIAS pixel_3463/NB2 pixel_3463/AMP_IN pixel_3463/SF_IB
+ pixel_3463/PIX_OUT pixel_3463/CSA_VREF pixel
Xpixel_3452 pixel_3452/gring pixel_3452/VDD pixel_3452/GND pixel_3452/VREF pixel_3452/ROW_SEL
+ pixel_3452/NB1 pixel_3452/VBIAS pixel_3452/NB2 pixel_3452/AMP_IN pixel_3452/SF_IB
+ pixel_3452/PIX_OUT pixel_3452/CSA_VREF pixel
Xpixel_4197 pixel_4197/gring pixel_4197/VDD pixel_4197/GND pixel_4197/VREF pixel_4197/ROW_SEL
+ pixel_4197/NB1 pixel_4197/VBIAS pixel_4197/NB2 pixel_4197/AMP_IN pixel_4197/SF_IB
+ pixel_4197/PIX_OUT pixel_4197/CSA_VREF pixel
Xpixel_2773 pixel_2773/gring pixel_2773/VDD pixel_2773/GND pixel_2773/VREF pixel_2773/ROW_SEL
+ pixel_2773/NB1 pixel_2773/VBIAS pixel_2773/NB2 pixel_2773/AMP_IN pixel_2773/SF_IB
+ pixel_2773/PIX_OUT pixel_2773/CSA_VREF pixel
Xpixel_2762 pixel_2762/gring pixel_2762/VDD pixel_2762/GND pixel_2762/VREF pixel_2762/ROW_SEL
+ pixel_2762/NB1 pixel_2762/VBIAS pixel_2762/NB2 pixel_2762/AMP_IN pixel_2762/SF_IB
+ pixel_2762/PIX_OUT pixel_2762/CSA_VREF pixel
Xpixel_2751 pixel_2751/gring pixel_2751/VDD pixel_2751/GND pixel_2751/VREF pixel_2751/ROW_SEL
+ pixel_2751/NB1 pixel_2751/VBIAS pixel_2751/NB2 pixel_2751/AMP_IN pixel_2751/SF_IB
+ pixel_2751/PIX_OUT pixel_2751/CSA_VREF pixel
Xpixel_3496 pixel_3496/gring pixel_3496/VDD pixel_3496/GND pixel_3496/VREF pixel_3496/ROW_SEL
+ pixel_3496/NB1 pixel_3496/VBIAS pixel_3496/NB2 pixel_3496/AMP_IN pixel_3496/SF_IB
+ pixel_3496/PIX_OUT pixel_3496/CSA_VREF pixel
Xpixel_2795 pixel_2795/gring pixel_2795/VDD pixel_2795/GND pixel_2795/VREF pixel_2795/ROW_SEL
+ pixel_2795/NB1 pixel_2795/VBIAS pixel_2795/NB2 pixel_2795/AMP_IN pixel_2795/SF_IB
+ pixel_2795/PIX_OUT pixel_2795/CSA_VREF pixel
Xpixel_2784 pixel_2784/gring pixel_2784/VDD pixel_2784/GND pixel_2784/VREF pixel_2784/ROW_SEL
+ pixel_2784/NB1 pixel_2784/VBIAS pixel_2784/NB2 pixel_2784/AMP_IN pixel_2784/SF_IB
+ pixel_2784/PIX_OUT pixel_2784/CSA_VREF pixel
Xpixel_9109 pixel_9109/gring pixel_9109/VDD pixel_9109/GND pixel_9109/VREF pixel_9109/ROW_SEL
+ pixel_9109/NB1 pixel_9109/VBIAS pixel_9109/NB2 pixel_9109/AMP_IN pixel_9109/SF_IB
+ pixel_9109/PIX_OUT pixel_9109/CSA_VREF pixel
Xpixel_8408 pixel_8408/gring pixel_8408/VDD pixel_8408/GND pixel_8408/VREF pixel_8408/ROW_SEL
+ pixel_8408/NB1 pixel_8408/VBIAS pixel_8408/NB2 pixel_8408/AMP_IN pixel_8408/SF_IB
+ pixel_8408/PIX_OUT pixel_8408/CSA_VREF pixel
Xpixel_8419 pixel_8419/gring pixel_8419/VDD pixel_8419/GND pixel_8419/VREF pixel_8419/ROW_SEL
+ pixel_8419/NB1 pixel_8419/VBIAS pixel_8419/NB2 pixel_8419/AMP_IN pixel_8419/SF_IB
+ pixel_8419/PIX_OUT pixel_8419/CSA_VREF pixel
Xpixel_7707 pixel_7707/gring pixel_7707/VDD pixel_7707/GND pixel_7707/VREF pixel_7707/ROW_SEL
+ pixel_7707/NB1 pixel_7707/VBIAS pixel_7707/NB2 pixel_7707/AMP_IN pixel_7707/SF_IB
+ pixel_7707/PIX_OUT pixel_7707/CSA_VREF pixel
Xpixel_7718 pixel_7718/gring pixel_7718/VDD pixel_7718/GND pixel_7718/VREF pixel_7718/ROW_SEL
+ pixel_7718/NB1 pixel_7718/VBIAS pixel_7718/NB2 pixel_7718/AMP_IN pixel_7718/SF_IB
+ pixel_7718/PIX_OUT pixel_7718/CSA_VREF pixel
Xpixel_7729 pixel_7729/gring pixel_7729/VDD pixel_7729/GND pixel_7729/VREF pixel_7729/ROW_SEL
+ pixel_7729/NB1 pixel_7729/VBIAS pixel_7729/NB2 pixel_7729/AMP_IN pixel_7729/SF_IB
+ pixel_7729/PIX_OUT pixel_7729/CSA_VREF pixel
Xpixel_2036 pixel_2036/gring pixel_2036/VDD pixel_2036/GND pixel_2036/VREF pixel_2036/ROW_SEL
+ pixel_2036/NB1 pixel_2036/VBIAS pixel_2036/NB2 pixel_2036/AMP_IN pixel_2036/SF_IB
+ pixel_2036/PIX_OUT pixel_2036/CSA_VREF pixel
Xpixel_2025 pixel_2025/gring pixel_2025/VDD pixel_2025/GND pixel_2025/VREF pixel_2025/ROW_SEL
+ pixel_2025/NB1 pixel_2025/VBIAS pixel_2025/NB2 pixel_2025/AMP_IN pixel_2025/SF_IB
+ pixel_2025/PIX_OUT pixel_2025/CSA_VREF pixel
Xpixel_2014 pixel_2014/gring pixel_2014/VDD pixel_2014/GND pixel_2014/VREF pixel_2014/ROW_SEL
+ pixel_2014/NB1 pixel_2014/VBIAS pixel_2014/NB2 pixel_2014/AMP_IN pixel_2014/SF_IB
+ pixel_2014/PIX_OUT pixel_2014/CSA_VREF pixel
Xpixel_2003 pixel_2003/gring pixel_2003/VDD pixel_2003/GND pixel_2003/VREF pixel_2003/ROW_SEL
+ pixel_2003/NB1 pixel_2003/VBIAS pixel_2003/NB2 pixel_2003/AMP_IN pixel_2003/SF_IB
+ pixel_2003/PIX_OUT pixel_2003/CSA_VREF pixel
Xpixel_1324 pixel_1324/gring pixel_1324/VDD pixel_1324/GND pixel_1324/VREF pixel_1324/ROW_SEL
+ pixel_1324/NB1 pixel_1324/VBIAS pixel_1324/NB2 pixel_1324/AMP_IN pixel_1324/SF_IB
+ pixel_1324/PIX_OUT pixel_1324/CSA_VREF pixel
Xpixel_1313 pixel_1313/gring pixel_1313/VDD pixel_1313/GND pixel_1313/VREF pixel_1313/ROW_SEL
+ pixel_1313/NB1 pixel_1313/VBIAS pixel_1313/NB2 pixel_1313/AMP_IN pixel_1313/SF_IB
+ pixel_1313/PIX_OUT pixel_1313/CSA_VREF pixel
Xpixel_1302 pixel_1302/gring pixel_1302/VDD pixel_1302/GND pixel_1302/VREF pixel_1302/ROW_SEL
+ pixel_1302/NB1 pixel_1302/VBIAS pixel_1302/NB2 pixel_1302/AMP_IN pixel_1302/SF_IB
+ pixel_1302/PIX_OUT pixel_1302/CSA_VREF pixel
Xpixel_2069 pixel_2069/gring pixel_2069/VDD pixel_2069/GND pixel_2069/VREF pixel_2069/ROW_SEL
+ pixel_2069/NB1 pixel_2069/VBIAS pixel_2069/NB2 pixel_2069/AMP_IN pixel_2069/SF_IB
+ pixel_2069/PIX_OUT pixel_2069/CSA_VREF pixel
Xpixel_2058 pixel_2058/gring pixel_2058/VDD pixel_2058/GND pixel_2058/VREF pixel_2058/ROW_SEL
+ pixel_2058/NB1 pixel_2058/VBIAS pixel_2058/NB2 pixel_2058/AMP_IN pixel_2058/SF_IB
+ pixel_2058/PIX_OUT pixel_2058/CSA_VREF pixel
Xpixel_2047 pixel_2047/gring pixel_2047/VDD pixel_2047/GND pixel_2047/VREF pixel_2047/ROW_SEL
+ pixel_2047/NB1 pixel_2047/VBIAS pixel_2047/NB2 pixel_2047/AMP_IN pixel_2047/SF_IB
+ pixel_2047/PIX_OUT pixel_2047/CSA_VREF pixel
Xpixel_1357 pixel_1357/gring pixel_1357/VDD pixel_1357/GND pixel_1357/VREF pixel_1357/ROW_SEL
+ pixel_1357/NB1 pixel_1357/VBIAS pixel_1357/NB2 pixel_1357/AMP_IN pixel_1357/SF_IB
+ pixel_1357/PIX_OUT pixel_1357/CSA_VREF pixel
Xpixel_1346 pixel_1346/gring pixel_1346/VDD pixel_1346/GND pixel_1346/VREF pixel_1346/ROW_SEL
+ pixel_1346/NB1 pixel_1346/VBIAS pixel_1346/NB2 pixel_1346/AMP_IN pixel_1346/SF_IB
+ pixel_1346/PIX_OUT pixel_1346/CSA_VREF pixel
Xpixel_1335 pixel_1335/gring pixel_1335/VDD pixel_1335/GND pixel_1335/VREF pixel_1335/ROW_SEL
+ pixel_1335/NB1 pixel_1335/VBIAS pixel_1335/NB2 pixel_1335/AMP_IN pixel_1335/SF_IB
+ pixel_1335/PIX_OUT pixel_1335/CSA_VREF pixel
Xpixel_1379 pixel_1379/gring pixel_1379/VDD pixel_1379/GND pixel_1379/VREF pixel_1379/ROW_SEL
+ pixel_1379/NB1 pixel_1379/VBIAS pixel_1379/NB2 pixel_1379/AMP_IN pixel_1379/SF_IB
+ pixel_1379/PIX_OUT pixel_1379/CSA_VREF pixel
Xpixel_1368 pixel_1368/gring pixel_1368/VDD pixel_1368/GND pixel_1368/VREF pixel_1368/ROW_SEL
+ pixel_1368/NB1 pixel_1368/VBIAS pixel_1368/NB2 pixel_1368/AMP_IN pixel_1368/SF_IB
+ pixel_1368/PIX_OUT pixel_1368/CSA_VREF pixel
Xpixel_9610 pixel_9610/gring pixel_9610/VDD pixel_9610/GND pixel_9610/VREF pixel_9610/ROW_SEL
+ pixel_9610/NB1 pixel_9610/VBIAS pixel_9610/NB2 pixel_9610/AMP_IN pixel_9610/SF_IB
+ pixel_9610/PIX_OUT pixel_9610/CSA_VREF pixel
Xpixel_9621 pixel_9621/gring pixel_9621/VDD pixel_9621/GND pixel_9621/VREF pixel_9621/ROW_SEL
+ pixel_9621/NB1 pixel_9621/VBIAS pixel_9621/NB2 pixel_9621/AMP_IN pixel_9621/SF_IB
+ pixel_9621/PIX_OUT pixel_9621/CSA_VREF pixel
Xpixel_9632 pixel_9632/gring pixel_9632/VDD pixel_9632/GND pixel_9632/VREF pixel_9632/ROW_SEL
+ pixel_9632/NB1 pixel_9632/VBIAS pixel_9632/NB2 pixel_9632/AMP_IN pixel_9632/SF_IB
+ pixel_9632/PIX_OUT pixel_9632/CSA_VREF pixel
Xpixel_8920 pixel_8920/gring pixel_8920/VDD pixel_8920/GND pixel_8920/VREF pixel_8920/ROW_SEL
+ pixel_8920/NB1 pixel_8920/VBIAS pixel_8920/NB2 pixel_8920/AMP_IN pixel_8920/SF_IB
+ pixel_8920/PIX_OUT pixel_8920/CSA_VREF pixel
Xpixel_9643 pixel_9643/gring pixel_9643/VDD pixel_9643/GND pixel_9643/VREF pixel_9643/ROW_SEL
+ pixel_9643/NB1 pixel_9643/VBIAS pixel_9643/NB2 pixel_9643/AMP_IN pixel_9643/SF_IB
+ pixel_9643/PIX_OUT pixel_9643/CSA_VREF pixel
Xpixel_9654 pixel_9654/gring pixel_9654/VDD pixel_9654/GND pixel_9654/VREF pixel_9654/ROW_SEL
+ pixel_9654/NB1 pixel_9654/VBIAS pixel_9654/NB2 pixel_9654/AMP_IN pixel_9654/SF_IB
+ pixel_9654/PIX_OUT pixel_9654/CSA_VREF pixel
Xpixel_9665 pixel_9665/gring pixel_9665/VDD pixel_9665/GND pixel_9665/VREF pixel_9665/ROW_SEL
+ pixel_9665/NB1 pixel_9665/VBIAS pixel_9665/NB2 pixel_9665/AMP_IN pixel_9665/SF_IB
+ pixel_9665/PIX_OUT pixel_9665/CSA_VREF pixel
Xpixel_8964 pixel_8964/gring pixel_8964/VDD pixel_8964/GND pixel_8964/VREF pixel_8964/ROW_SEL
+ pixel_8964/NB1 pixel_8964/VBIAS pixel_8964/NB2 pixel_8964/AMP_IN pixel_8964/SF_IB
+ pixel_8964/PIX_OUT pixel_8964/CSA_VREF pixel
Xpixel_8953 pixel_8953/gring pixel_8953/VDD pixel_8953/GND pixel_8953/VREF pixel_8953/ROW_SEL
+ pixel_8953/NB1 pixel_8953/VBIAS pixel_8953/NB2 pixel_8953/AMP_IN pixel_8953/SF_IB
+ pixel_8953/PIX_OUT pixel_8953/CSA_VREF pixel
Xpixel_8942 pixel_8942/gring pixel_8942/VDD pixel_8942/GND pixel_8942/VREF pixel_8942/ROW_SEL
+ pixel_8942/NB1 pixel_8942/VBIAS pixel_8942/NB2 pixel_8942/AMP_IN pixel_8942/SF_IB
+ pixel_8942/PIX_OUT pixel_8942/CSA_VREF pixel
Xpixel_8931 pixel_8931/gring pixel_8931/VDD pixel_8931/GND pixel_8931/VREF pixel_8931/ROW_SEL
+ pixel_8931/NB1 pixel_8931/VBIAS pixel_8931/NB2 pixel_8931/AMP_IN pixel_8931/SF_IB
+ pixel_8931/PIX_OUT pixel_8931/CSA_VREF pixel
Xpixel_9698 pixel_9698/gring pixel_9698/VDD pixel_9698/GND pixel_9698/VREF pixel_9698/ROW_SEL
+ pixel_9698/NB1 pixel_9698/VBIAS pixel_9698/NB2 pixel_9698/AMP_IN pixel_9698/SF_IB
+ pixel_9698/PIX_OUT pixel_9698/CSA_VREF pixel
Xpixel_9687 pixel_9687/gring pixel_9687/VDD pixel_9687/GND pixel_9687/VREF pixel_9687/ROW_SEL
+ pixel_9687/NB1 pixel_9687/VBIAS pixel_9687/NB2 pixel_9687/AMP_IN pixel_9687/SF_IB
+ pixel_9687/PIX_OUT pixel_9687/CSA_VREF pixel
Xpixel_9676 pixel_9676/gring pixel_9676/VDD pixel_9676/GND pixel_9676/VREF pixel_9676/ROW_SEL
+ pixel_9676/NB1 pixel_9676/VBIAS pixel_9676/NB2 pixel_9676/AMP_IN pixel_9676/SF_IB
+ pixel_9676/PIX_OUT pixel_9676/CSA_VREF pixel
Xpixel_8997 pixel_8997/gring pixel_8997/VDD pixel_8997/GND pixel_8997/VREF pixel_8997/ROW_SEL
+ pixel_8997/NB1 pixel_8997/VBIAS pixel_8997/NB2 pixel_8997/AMP_IN pixel_8997/SF_IB
+ pixel_8997/PIX_OUT pixel_8997/CSA_VREF pixel
Xpixel_8986 pixel_8986/gring pixel_8986/VDD pixel_8986/GND pixel_8986/VREF pixel_8986/ROW_SEL
+ pixel_8986/NB1 pixel_8986/VBIAS pixel_8986/NB2 pixel_8986/AMP_IN pixel_8986/SF_IB
+ pixel_8986/PIX_OUT pixel_8986/CSA_VREF pixel
Xpixel_8975 pixel_8975/gring pixel_8975/VDD pixel_8975/GND pixel_8975/VREF pixel_8975/ROW_SEL
+ pixel_8975/NB1 pixel_8975/VBIAS pixel_8975/NB2 pixel_8975/AMP_IN pixel_8975/SF_IB
+ pixel_8975/PIX_OUT pixel_8975/CSA_VREF pixel
Xpixel_3260 pixel_3260/gring pixel_3260/VDD pixel_3260/GND pixel_3260/VREF pixel_3260/ROW_SEL
+ pixel_3260/NB1 pixel_3260/VBIAS pixel_3260/NB2 pixel_3260/AMP_IN pixel_3260/SF_IB
+ pixel_3260/PIX_OUT pixel_3260/CSA_VREF pixel
Xpixel_3293 pixel_3293/gring pixel_3293/VDD pixel_3293/GND pixel_3293/VREF pixel_3293/ROW_SEL
+ pixel_3293/NB1 pixel_3293/VBIAS pixel_3293/NB2 pixel_3293/AMP_IN pixel_3293/SF_IB
+ pixel_3293/PIX_OUT pixel_3293/CSA_VREF pixel
Xpixel_3282 pixel_3282/gring pixel_3282/VDD pixel_3282/GND pixel_3282/VREF pixel_3282/ROW_SEL
+ pixel_3282/NB1 pixel_3282/VBIAS pixel_3282/NB2 pixel_3282/AMP_IN pixel_3282/SF_IB
+ pixel_3282/PIX_OUT pixel_3282/CSA_VREF pixel
Xpixel_3271 pixel_3271/gring pixel_3271/VDD pixel_3271/GND pixel_3271/VREF pixel_3271/ROW_SEL
+ pixel_3271/NB1 pixel_3271/VBIAS pixel_3271/NB2 pixel_3271/AMP_IN pixel_3271/SF_IB
+ pixel_3271/PIX_OUT pixel_3271/CSA_VREF pixel
Xpixel_2581 pixel_2581/gring pixel_2581/VDD pixel_2581/GND pixel_2581/VREF pixel_2581/ROW_SEL
+ pixel_2581/NB1 pixel_2581/VBIAS pixel_2581/NB2 pixel_2581/AMP_IN pixel_2581/SF_IB
+ pixel_2581/PIX_OUT pixel_2581/CSA_VREF pixel
Xpixel_2570 pixel_2570/gring pixel_2570/VDD pixel_2570/GND pixel_2570/VREF pixel_2570/ROW_SEL
+ pixel_2570/NB1 pixel_2570/VBIAS pixel_2570/NB2 pixel_2570/AMP_IN pixel_2570/SF_IB
+ pixel_2570/PIX_OUT pixel_2570/CSA_VREF pixel
Xpixel_1880 pixel_1880/gring pixel_1880/VDD pixel_1880/GND pixel_1880/VREF pixel_1880/ROW_SEL
+ pixel_1880/NB1 pixel_1880/VBIAS pixel_1880/NB2 pixel_1880/AMP_IN pixel_1880/SF_IB
+ pixel_1880/PIX_OUT pixel_1880/CSA_VREF pixel
Xpixel_2592 pixel_2592/gring pixel_2592/VDD pixel_2592/GND pixel_2592/VREF pixel_2592/ROW_SEL
+ pixel_2592/NB1 pixel_2592/VBIAS pixel_2592/NB2 pixel_2592/AMP_IN pixel_2592/SF_IB
+ pixel_2592/PIX_OUT pixel_2592/CSA_VREF pixel
Xpixel_1891 pixel_1891/gring pixel_1891/VDD pixel_1891/GND pixel_1891/VREF pixel_1891/ROW_SEL
+ pixel_1891/NB1 pixel_1891/VBIAS pixel_1891/NB2 pixel_1891/AMP_IN pixel_1891/SF_IB
+ pixel_1891/PIX_OUT pixel_1891/CSA_VREF pixel
Xpixel_906 pixel_906/gring pixel_906/VDD pixel_906/GND pixel_906/VREF pixel_906/ROW_SEL
+ pixel_906/NB1 pixel_906/VBIAS pixel_906/NB2 pixel_906/AMP_IN pixel_906/SF_IB pixel_906/PIX_OUT
+ pixel_906/CSA_VREF pixel
Xpixel_939 pixel_939/gring pixel_939/VDD pixel_939/GND pixel_939/VREF pixel_939/ROW_SEL
+ pixel_939/NB1 pixel_939/VBIAS pixel_939/NB2 pixel_939/AMP_IN pixel_939/SF_IB pixel_939/PIX_OUT
+ pixel_939/CSA_VREF pixel
Xpixel_928 pixel_928/gring pixel_928/VDD pixel_928/GND pixel_928/VREF pixel_928/ROW_SEL
+ pixel_928/NB1 pixel_928/VBIAS pixel_928/NB2 pixel_928/AMP_IN pixel_928/SF_IB pixel_928/PIX_OUT
+ pixel_928/CSA_VREF pixel
Xpixel_917 pixel_917/gring pixel_917/VDD pixel_917/GND pixel_917/VREF pixel_917/ROW_SEL
+ pixel_917/NB1 pixel_917/VBIAS pixel_917/NB2 pixel_917/AMP_IN pixel_917/SF_IB pixel_917/PIX_OUT
+ pixel_917/CSA_VREF pixel
Xpixel_8205 pixel_8205/gring pixel_8205/VDD pixel_8205/GND pixel_8205/VREF pixel_8205/ROW_SEL
+ pixel_8205/NB1 pixel_8205/VBIAS pixel_8205/NB2 pixel_8205/AMP_IN pixel_8205/SF_IB
+ pixel_8205/PIX_OUT pixel_8205/CSA_VREF pixel
Xpixel_8216 pixel_8216/gring pixel_8216/VDD pixel_8216/GND pixel_8216/VREF pixel_8216/ROW_SEL
+ pixel_8216/NB1 pixel_8216/VBIAS pixel_8216/NB2 pixel_8216/AMP_IN pixel_8216/SF_IB
+ pixel_8216/PIX_OUT pixel_8216/CSA_VREF pixel
Xpixel_8227 pixel_8227/gring pixel_8227/VDD pixel_8227/GND pixel_8227/VREF pixel_8227/ROW_SEL
+ pixel_8227/NB1 pixel_8227/VBIAS pixel_8227/NB2 pixel_8227/AMP_IN pixel_8227/SF_IB
+ pixel_8227/PIX_OUT pixel_8227/CSA_VREF pixel
Xpixel_8238 pixel_8238/gring pixel_8238/VDD pixel_8238/GND pixel_8238/VREF pixel_8238/ROW_SEL
+ pixel_8238/NB1 pixel_8238/VBIAS pixel_8238/NB2 pixel_8238/AMP_IN pixel_8238/SF_IB
+ pixel_8238/PIX_OUT pixel_8238/CSA_VREF pixel
Xpixel_8249 pixel_8249/gring pixel_8249/VDD pixel_8249/GND pixel_8249/VREF pixel_8249/ROW_SEL
+ pixel_8249/NB1 pixel_8249/VBIAS pixel_8249/NB2 pixel_8249/AMP_IN pixel_8249/SF_IB
+ pixel_8249/PIX_OUT pixel_8249/CSA_VREF pixel
Xpixel_7504 pixel_7504/gring pixel_7504/VDD pixel_7504/GND pixel_7504/VREF pixel_7504/ROW_SEL
+ pixel_7504/NB1 pixel_7504/VBIAS pixel_7504/NB2 pixel_7504/AMP_IN pixel_7504/SF_IB
+ pixel_7504/PIX_OUT pixel_7504/CSA_VREF pixel
Xpixel_7515 pixel_7515/gring pixel_7515/VDD pixel_7515/GND pixel_7515/VREF pixel_7515/ROW_SEL
+ pixel_7515/NB1 pixel_7515/VBIAS pixel_7515/NB2 pixel_7515/AMP_IN pixel_7515/SF_IB
+ pixel_7515/PIX_OUT pixel_7515/CSA_VREF pixel
Xpixel_7526 pixel_7526/gring pixel_7526/VDD pixel_7526/GND pixel_7526/VREF pixel_7526/ROW_SEL
+ pixel_7526/NB1 pixel_7526/VBIAS pixel_7526/NB2 pixel_7526/AMP_IN pixel_7526/SF_IB
+ pixel_7526/PIX_OUT pixel_7526/CSA_VREF pixel
Xpixel_7537 pixel_7537/gring pixel_7537/VDD pixel_7537/GND pixel_7537/VREF pixel_7537/ROW_SEL
+ pixel_7537/NB1 pixel_7537/VBIAS pixel_7537/NB2 pixel_7537/AMP_IN pixel_7537/SF_IB
+ pixel_7537/PIX_OUT pixel_7537/CSA_VREF pixel
Xpixel_7548 pixel_7548/gring pixel_7548/VDD pixel_7548/GND pixel_7548/VREF pixel_7548/ROW_SEL
+ pixel_7548/NB1 pixel_7548/VBIAS pixel_7548/NB2 pixel_7548/AMP_IN pixel_7548/SF_IB
+ pixel_7548/PIX_OUT pixel_7548/CSA_VREF pixel
Xpixel_6803 pixel_6803/gring pixel_6803/VDD pixel_6803/GND pixel_6803/VREF pixel_6803/ROW_SEL
+ pixel_6803/NB1 pixel_6803/VBIAS pixel_6803/NB2 pixel_6803/AMP_IN pixel_6803/SF_IB
+ pixel_6803/PIX_OUT pixel_6803/CSA_VREF pixel
Xpixel_7559 pixel_7559/gring pixel_7559/VDD pixel_7559/GND pixel_7559/VREF pixel_7559/ROW_SEL
+ pixel_7559/NB1 pixel_7559/VBIAS pixel_7559/NB2 pixel_7559/AMP_IN pixel_7559/SF_IB
+ pixel_7559/PIX_OUT pixel_7559/CSA_VREF pixel
Xpixel_6814 pixel_6814/gring pixel_6814/VDD pixel_6814/GND pixel_6814/VREF pixel_6814/ROW_SEL
+ pixel_6814/NB1 pixel_6814/VBIAS pixel_6814/NB2 pixel_6814/AMP_IN pixel_6814/SF_IB
+ pixel_6814/PIX_OUT pixel_6814/CSA_VREF pixel
Xpixel_6825 pixel_6825/gring pixel_6825/VDD pixel_6825/GND pixel_6825/VREF pixel_6825/ROW_SEL
+ pixel_6825/NB1 pixel_6825/VBIAS pixel_6825/NB2 pixel_6825/AMP_IN pixel_6825/SF_IB
+ pixel_6825/PIX_OUT pixel_6825/CSA_VREF pixel
Xpixel_6836 pixel_6836/gring pixel_6836/VDD pixel_6836/GND pixel_6836/VREF pixel_6836/ROW_SEL
+ pixel_6836/NB1 pixel_6836/VBIAS pixel_6836/NB2 pixel_6836/AMP_IN pixel_6836/SF_IB
+ pixel_6836/PIX_OUT pixel_6836/CSA_VREF pixel
Xpixel_6847 pixel_6847/gring pixel_6847/VDD pixel_6847/GND pixel_6847/VREF pixel_6847/ROW_SEL
+ pixel_6847/NB1 pixel_6847/VBIAS pixel_6847/NB2 pixel_6847/AMP_IN pixel_6847/SF_IB
+ pixel_6847/PIX_OUT pixel_6847/CSA_VREF pixel
Xpixel_6858 pixel_6858/gring pixel_6858/VDD pixel_6858/GND pixel_6858/VREF pixel_6858/ROW_SEL
+ pixel_6858/NB1 pixel_6858/VBIAS pixel_6858/NB2 pixel_6858/AMP_IN pixel_6858/SF_IB
+ pixel_6858/PIX_OUT pixel_6858/CSA_VREF pixel
Xpixel_6869 pixel_6869/gring pixel_6869/VDD pixel_6869/GND pixel_6869/VREF pixel_6869/ROW_SEL
+ pixel_6869/NB1 pixel_6869/VBIAS pixel_6869/NB2 pixel_6869/AMP_IN pixel_6869/SF_IB
+ pixel_6869/PIX_OUT pixel_6869/CSA_VREF pixel
Xpixel_1132 pixel_1132/gring pixel_1132/VDD pixel_1132/GND pixel_1132/VREF pixel_1132/ROW_SEL
+ pixel_1132/NB1 pixel_1132/VBIAS pixel_1132/NB2 pixel_1132/AMP_IN pixel_1132/SF_IB
+ pixel_1132/PIX_OUT pixel_1132/CSA_VREF pixel
Xpixel_1121 pixel_1121/gring pixel_1121/VDD pixel_1121/GND pixel_1121/VREF pixel_1121/ROW_SEL
+ pixel_1121/NB1 pixel_1121/VBIAS pixel_1121/NB2 pixel_1121/AMP_IN pixel_1121/SF_IB
+ pixel_1121/PIX_OUT pixel_1121/CSA_VREF pixel
Xpixel_1110 pixel_1110/gring pixel_1110/VDD pixel_1110/GND pixel_1110/VREF pixel_1110/ROW_SEL
+ pixel_1110/NB1 pixel_1110/VBIAS pixel_1110/NB2 pixel_1110/AMP_IN pixel_1110/SF_IB
+ pixel_1110/PIX_OUT pixel_1110/CSA_VREF pixel
Xpixel_1165 pixel_1165/gring pixel_1165/VDD pixel_1165/GND pixel_1165/VREF pixel_1165/ROW_SEL
+ pixel_1165/NB1 pixel_1165/VBIAS pixel_1165/NB2 pixel_1165/AMP_IN pixel_1165/SF_IB
+ pixel_1165/PIX_OUT pixel_1165/CSA_VREF pixel
Xpixel_1154 pixel_1154/gring pixel_1154/VDD pixel_1154/GND pixel_1154/VREF pixel_1154/ROW_SEL
+ pixel_1154/NB1 pixel_1154/VBIAS pixel_1154/NB2 pixel_1154/AMP_IN pixel_1154/SF_IB
+ pixel_1154/PIX_OUT pixel_1154/CSA_VREF pixel
Xpixel_1143 pixel_1143/gring pixel_1143/VDD pixel_1143/GND pixel_1143/VREF pixel_1143/ROW_SEL
+ pixel_1143/NB1 pixel_1143/VBIAS pixel_1143/NB2 pixel_1143/AMP_IN pixel_1143/SF_IB
+ pixel_1143/PIX_OUT pixel_1143/CSA_VREF pixel
Xpixel_1198 pixel_1198/gring pixel_1198/VDD pixel_1198/GND pixel_1198/VREF pixel_1198/ROW_SEL
+ pixel_1198/NB1 pixel_1198/VBIAS pixel_1198/NB2 pixel_1198/AMP_IN pixel_1198/SF_IB
+ pixel_1198/PIX_OUT pixel_1198/CSA_VREF pixel
Xpixel_1187 pixel_1187/gring pixel_1187/VDD pixel_1187/GND pixel_1187/VREF pixel_1187/ROW_SEL
+ pixel_1187/NB1 pixel_1187/VBIAS pixel_1187/NB2 pixel_1187/AMP_IN pixel_1187/SF_IB
+ pixel_1187/PIX_OUT pixel_1187/CSA_VREF pixel
Xpixel_1176 pixel_1176/gring pixel_1176/VDD pixel_1176/GND pixel_1176/VREF pixel_1176/ROW_SEL
+ pixel_1176/NB1 pixel_1176/VBIAS pixel_1176/NB2 pixel_1176/AMP_IN pixel_1176/SF_IB
+ pixel_1176/PIX_OUT pixel_1176/CSA_VREF pixel
Xpixel_9440 pixel_9440/gring pixel_9440/VDD pixel_9440/GND pixel_9440/VREF pixel_9440/ROW_SEL
+ pixel_9440/NB1 pixel_9440/VBIAS pixel_9440/NB2 pixel_9440/AMP_IN pixel_9440/SF_IB
+ pixel_9440/PIX_OUT pixel_9440/CSA_VREF pixel
Xpixel_9473 pixel_9473/gring pixel_9473/VDD pixel_9473/GND pixel_9473/VREF pixel_9473/ROW_SEL
+ pixel_9473/NB1 pixel_9473/VBIAS pixel_9473/NB2 pixel_9473/AMP_IN pixel_9473/SF_IB
+ pixel_9473/PIX_OUT pixel_9473/CSA_VREF pixel
Xpixel_9462 pixel_9462/gring pixel_9462/VDD pixel_9462/GND pixel_9462/VREF pixel_9462/ROW_SEL
+ pixel_9462/NB1 pixel_9462/VBIAS pixel_9462/NB2 pixel_9462/AMP_IN pixel_9462/SF_IB
+ pixel_9462/PIX_OUT pixel_9462/CSA_VREF pixel
Xpixel_9451 pixel_9451/gring pixel_9451/VDD pixel_9451/GND pixel_9451/VREF pixel_9451/ROW_SEL
+ pixel_9451/NB1 pixel_9451/VBIAS pixel_9451/NB2 pixel_9451/AMP_IN pixel_9451/SF_IB
+ pixel_9451/PIX_OUT pixel_9451/CSA_VREF pixel
Xpixel_8772 pixel_8772/gring pixel_8772/VDD pixel_8772/GND pixel_8772/VREF pixel_8772/ROW_SEL
+ pixel_8772/NB1 pixel_8772/VBIAS pixel_8772/NB2 pixel_8772/AMP_IN pixel_8772/SF_IB
+ pixel_8772/PIX_OUT pixel_8772/CSA_VREF pixel
Xpixel_8761 pixel_8761/gring pixel_8761/VDD pixel_8761/GND pixel_8761/VREF pixel_8761/ROW_SEL
+ pixel_8761/NB1 pixel_8761/VBIAS pixel_8761/NB2 pixel_8761/AMP_IN pixel_8761/SF_IB
+ pixel_8761/PIX_OUT pixel_8761/CSA_VREF pixel
Xpixel_8750 pixel_8750/gring pixel_8750/VDD pixel_8750/GND pixel_8750/VREF pixel_8750/ROW_SEL
+ pixel_8750/NB1 pixel_8750/VBIAS pixel_8750/NB2 pixel_8750/AMP_IN pixel_8750/SF_IB
+ pixel_8750/PIX_OUT pixel_8750/CSA_VREF pixel
Xpixel_9495 pixel_9495/gring pixel_9495/VDD pixel_9495/GND pixel_9495/VREF pixel_9495/ROW_SEL
+ pixel_9495/NB1 pixel_9495/VBIAS pixel_9495/NB2 pixel_9495/AMP_IN pixel_9495/SF_IB
+ pixel_9495/PIX_OUT pixel_9495/CSA_VREF pixel
Xpixel_9484 pixel_9484/gring pixel_9484/VDD pixel_9484/GND pixel_9484/VREF pixel_9484/ROW_SEL
+ pixel_9484/NB1 pixel_9484/VBIAS pixel_9484/NB2 pixel_9484/AMP_IN pixel_9484/SF_IB
+ pixel_9484/PIX_OUT pixel_9484/CSA_VREF pixel
Xpixel_8794 pixel_8794/gring pixel_8794/VDD pixel_8794/GND pixel_8794/VREF pixel_8794/ROW_SEL
+ pixel_8794/NB1 pixel_8794/VBIAS pixel_8794/NB2 pixel_8794/AMP_IN pixel_8794/SF_IB
+ pixel_8794/PIX_OUT pixel_8794/CSA_VREF pixel
Xpixel_8783 pixel_8783/gring pixel_8783/VDD pixel_8783/GND pixel_8783/VREF pixel_8783/ROW_SEL
+ pixel_8783/NB1 pixel_8783/VBIAS pixel_8783/NB2 pixel_8783/AMP_IN pixel_8783/SF_IB
+ pixel_8783/PIX_OUT pixel_8783/CSA_VREF pixel
Xpixel_3090 pixel_3090/gring pixel_3090/VDD pixel_3090/GND pixel_3090/VREF pixel_3090/ROW_SEL
+ pixel_3090/NB1 pixel_3090/VBIAS pixel_3090/NB2 pixel_3090/AMP_IN pixel_3090/SF_IB
+ pixel_3090/PIX_OUT pixel_3090/CSA_VREF pixel
Xpixel_5409 pixel_5409/gring pixel_5409/VDD pixel_5409/GND pixel_5409/VREF pixel_5409/ROW_SEL
+ pixel_5409/NB1 pixel_5409/VBIAS pixel_5409/NB2 pixel_5409/AMP_IN pixel_5409/SF_IB
+ pixel_5409/PIX_OUT pixel_5409/CSA_VREF pixel
Xpixel_714 pixel_714/gring pixel_714/VDD pixel_714/GND pixel_714/VREF pixel_714/ROW_SEL
+ pixel_714/NB1 pixel_714/VBIAS pixel_714/NB2 pixel_714/AMP_IN pixel_714/SF_IB pixel_714/PIX_OUT
+ pixel_714/CSA_VREF pixel
Xpixel_703 pixel_703/gring pixel_703/VDD pixel_703/GND pixel_703/VREF pixel_703/ROW_SEL
+ pixel_703/NB1 pixel_703/VBIAS pixel_703/NB2 pixel_703/AMP_IN pixel_703/SF_IB pixel_703/PIX_OUT
+ pixel_703/CSA_VREF pixel
Xpixel_4708 pixel_4708/gring pixel_4708/VDD pixel_4708/GND pixel_4708/VREF pixel_4708/ROW_SEL
+ pixel_4708/NB1 pixel_4708/VBIAS pixel_4708/NB2 pixel_4708/AMP_IN pixel_4708/SF_IB
+ pixel_4708/PIX_OUT pixel_4708/CSA_VREF pixel
Xpixel_4719 pixel_4719/gring pixel_4719/VDD pixel_4719/GND pixel_4719/VREF pixel_4719/ROW_SEL
+ pixel_4719/NB1 pixel_4719/VBIAS pixel_4719/NB2 pixel_4719/AMP_IN pixel_4719/SF_IB
+ pixel_4719/PIX_OUT pixel_4719/CSA_VREF pixel
Xpixel_747 pixel_747/gring pixel_747/VDD pixel_747/GND pixel_747/VREF pixel_747/ROW_SEL
+ pixel_747/NB1 pixel_747/VBIAS pixel_747/NB2 pixel_747/AMP_IN pixel_747/SF_IB pixel_747/PIX_OUT
+ pixel_747/CSA_VREF pixel
Xpixel_736 pixel_736/gring pixel_736/VDD pixel_736/GND pixel_736/VREF pixel_736/ROW_SEL
+ pixel_736/NB1 pixel_736/VBIAS pixel_736/NB2 pixel_736/AMP_IN pixel_736/SF_IB pixel_736/PIX_OUT
+ pixel_736/CSA_VREF pixel
Xpixel_725 pixel_725/gring pixel_725/VDD pixel_725/GND pixel_725/VREF pixel_725/ROW_SEL
+ pixel_725/NB1 pixel_725/VBIAS pixel_725/NB2 pixel_725/AMP_IN pixel_725/SF_IB pixel_725/PIX_OUT
+ pixel_725/CSA_VREF pixel
Xpixel_769 pixel_769/gring pixel_769/VDD pixel_769/GND pixel_769/VREF pixel_769/ROW_SEL
+ pixel_769/NB1 pixel_769/VBIAS pixel_769/NB2 pixel_769/AMP_IN pixel_769/SF_IB pixel_769/PIX_OUT
+ pixel_769/CSA_VREF pixel
Xpixel_758 pixel_758/gring pixel_758/VDD pixel_758/GND pixel_758/VREF pixel_758/ROW_SEL
+ pixel_758/NB1 pixel_758/VBIAS pixel_758/NB2 pixel_758/AMP_IN pixel_758/SF_IB pixel_758/PIX_OUT
+ pixel_758/CSA_VREF pixel
Xpixel_8002 pixel_8002/gring pixel_8002/VDD pixel_8002/GND pixel_8002/VREF pixel_8002/ROW_SEL
+ pixel_8002/NB1 pixel_8002/VBIAS pixel_8002/NB2 pixel_8002/AMP_IN pixel_8002/SF_IB
+ pixel_8002/PIX_OUT pixel_8002/CSA_VREF pixel
Xpixel_8013 pixel_8013/gring pixel_8013/VDD pixel_8013/GND pixel_8013/VREF pixel_8013/ROW_SEL
+ pixel_8013/NB1 pixel_8013/VBIAS pixel_8013/NB2 pixel_8013/AMP_IN pixel_8013/SF_IB
+ pixel_8013/PIX_OUT pixel_8013/CSA_VREF pixel
Xpixel_8024 pixel_8024/gring pixel_8024/VDD pixel_8024/GND pixel_8024/VREF pixel_8024/ROW_SEL
+ pixel_8024/NB1 pixel_8024/VBIAS pixel_8024/NB2 pixel_8024/AMP_IN pixel_8024/SF_IB
+ pixel_8024/PIX_OUT pixel_8024/CSA_VREF pixel
Xpixel_8035 pixel_8035/gring pixel_8035/VDD pixel_8035/GND pixel_8035/VREF pixel_8035/ROW_SEL
+ pixel_8035/NB1 pixel_8035/VBIAS pixel_8035/NB2 pixel_8035/AMP_IN pixel_8035/SF_IB
+ pixel_8035/PIX_OUT pixel_8035/CSA_VREF pixel
Xpixel_8046 pixel_8046/gring pixel_8046/VDD pixel_8046/GND pixel_8046/VREF pixel_8046/ROW_SEL
+ pixel_8046/NB1 pixel_8046/VBIAS pixel_8046/NB2 pixel_8046/AMP_IN pixel_8046/SF_IB
+ pixel_8046/PIX_OUT pixel_8046/CSA_VREF pixel
Xpixel_8057 pixel_8057/gring pixel_8057/VDD pixel_8057/GND pixel_8057/VREF pixel_8057/ROW_SEL
+ pixel_8057/NB1 pixel_8057/VBIAS pixel_8057/NB2 pixel_8057/AMP_IN pixel_8057/SF_IB
+ pixel_8057/PIX_OUT pixel_8057/CSA_VREF pixel
Xpixel_8068 pixel_8068/gring pixel_8068/VDD pixel_8068/GND pixel_8068/VREF pixel_8068/ROW_SEL
+ pixel_8068/NB1 pixel_8068/VBIAS pixel_8068/NB2 pixel_8068/AMP_IN pixel_8068/SF_IB
+ pixel_8068/PIX_OUT pixel_8068/CSA_VREF pixel
Xpixel_7301 pixel_7301/gring pixel_7301/VDD pixel_7301/GND pixel_7301/VREF pixel_7301/ROW_SEL
+ pixel_7301/NB1 pixel_7301/VBIAS pixel_7301/NB2 pixel_7301/AMP_IN pixel_7301/SF_IB
+ pixel_7301/PIX_OUT pixel_7301/CSA_VREF pixel
Xpixel_7312 pixel_7312/gring pixel_7312/VDD pixel_7312/GND pixel_7312/VREF pixel_7312/ROW_SEL
+ pixel_7312/NB1 pixel_7312/VBIAS pixel_7312/NB2 pixel_7312/AMP_IN pixel_7312/SF_IB
+ pixel_7312/PIX_OUT pixel_7312/CSA_VREF pixel
Xpixel_7323 pixel_7323/gring pixel_7323/VDD pixel_7323/GND pixel_7323/VREF pixel_7323/ROW_SEL
+ pixel_7323/NB1 pixel_7323/VBIAS pixel_7323/NB2 pixel_7323/AMP_IN pixel_7323/SF_IB
+ pixel_7323/PIX_OUT pixel_7323/CSA_VREF pixel
Xpixel_8079 pixel_8079/gring pixel_8079/VDD pixel_8079/GND pixel_8079/VREF pixel_8079/ROW_SEL
+ pixel_8079/NB1 pixel_8079/VBIAS pixel_8079/NB2 pixel_8079/AMP_IN pixel_8079/SF_IB
+ pixel_8079/PIX_OUT pixel_8079/CSA_VREF pixel
Xpixel_7334 pixel_7334/gring pixel_7334/VDD pixel_7334/GND pixel_7334/VREF pixel_7334/ROW_SEL
+ pixel_7334/NB1 pixel_7334/VBIAS pixel_7334/NB2 pixel_7334/AMP_IN pixel_7334/SF_IB
+ pixel_7334/PIX_OUT pixel_7334/CSA_VREF pixel
Xpixel_7345 pixel_7345/gring pixel_7345/VDD pixel_7345/GND pixel_7345/VREF pixel_7345/ROW_SEL
+ pixel_7345/NB1 pixel_7345/VBIAS pixel_7345/NB2 pixel_7345/AMP_IN pixel_7345/SF_IB
+ pixel_7345/PIX_OUT pixel_7345/CSA_VREF pixel
Xpixel_7356 pixel_7356/gring pixel_7356/VDD pixel_7356/GND pixel_7356/VREF pixel_7356/ROW_SEL
+ pixel_7356/NB1 pixel_7356/VBIAS pixel_7356/NB2 pixel_7356/AMP_IN pixel_7356/SF_IB
+ pixel_7356/PIX_OUT pixel_7356/CSA_VREF pixel
Xpixel_6600 pixel_6600/gring pixel_6600/VDD pixel_6600/GND pixel_6600/VREF pixel_6600/ROW_SEL
+ pixel_6600/NB1 pixel_6600/VBIAS pixel_6600/NB2 pixel_6600/AMP_IN pixel_6600/SF_IB
+ pixel_6600/PIX_OUT pixel_6600/CSA_VREF pixel
Xpixel_6611 pixel_6611/gring pixel_6611/VDD pixel_6611/GND pixel_6611/VREF pixel_6611/ROW_SEL
+ pixel_6611/NB1 pixel_6611/VBIAS pixel_6611/NB2 pixel_6611/AMP_IN pixel_6611/SF_IB
+ pixel_6611/PIX_OUT pixel_6611/CSA_VREF pixel
Xpixel_7367 pixel_7367/gring pixel_7367/VDD pixel_7367/GND pixel_7367/VREF pixel_7367/ROW_SEL
+ pixel_7367/NB1 pixel_7367/VBIAS pixel_7367/NB2 pixel_7367/AMP_IN pixel_7367/SF_IB
+ pixel_7367/PIX_OUT pixel_7367/CSA_VREF pixel
Xpixel_7378 pixel_7378/gring pixel_7378/VDD pixel_7378/GND pixel_7378/VREF pixel_7378/ROW_SEL
+ pixel_7378/NB1 pixel_7378/VBIAS pixel_7378/NB2 pixel_7378/AMP_IN pixel_7378/SF_IB
+ pixel_7378/PIX_OUT pixel_7378/CSA_VREF pixel
Xpixel_7389 pixel_7389/gring pixel_7389/VDD pixel_7389/GND pixel_7389/VREF pixel_7389/ROW_SEL
+ pixel_7389/NB1 pixel_7389/VBIAS pixel_7389/NB2 pixel_7389/AMP_IN pixel_7389/SF_IB
+ pixel_7389/PIX_OUT pixel_7389/CSA_VREF pixel
Xpixel_6622 pixel_6622/gring pixel_6622/VDD pixel_6622/GND pixel_6622/VREF pixel_6622/ROW_SEL
+ pixel_6622/NB1 pixel_6622/VBIAS pixel_6622/NB2 pixel_6622/AMP_IN pixel_6622/SF_IB
+ pixel_6622/PIX_OUT pixel_6622/CSA_VREF pixel
Xpixel_6633 pixel_6633/gring pixel_6633/VDD pixel_6633/GND pixel_6633/VREF pixel_6633/ROW_SEL
+ pixel_6633/NB1 pixel_6633/VBIAS pixel_6633/NB2 pixel_6633/AMP_IN pixel_6633/SF_IB
+ pixel_6633/PIX_OUT pixel_6633/CSA_VREF pixel
Xpixel_6644 pixel_6644/gring pixel_6644/VDD pixel_6644/GND pixel_6644/VREF pixel_6644/ROW_SEL
+ pixel_6644/NB1 pixel_6644/VBIAS pixel_6644/NB2 pixel_6644/AMP_IN pixel_6644/SF_IB
+ pixel_6644/PIX_OUT pixel_6644/CSA_VREF pixel
Xpixel_5910 pixel_5910/gring pixel_5910/VDD pixel_5910/GND pixel_5910/VREF pixel_5910/ROW_SEL
+ pixel_5910/NB1 pixel_5910/VBIAS pixel_5910/NB2 pixel_5910/AMP_IN pixel_5910/SF_IB
+ pixel_5910/PIX_OUT pixel_5910/CSA_VREF pixel
Xpixel_6655 pixel_6655/gring pixel_6655/VDD pixel_6655/GND pixel_6655/VREF pixel_6655/ROW_SEL
+ pixel_6655/NB1 pixel_6655/VBIAS pixel_6655/NB2 pixel_6655/AMP_IN pixel_6655/SF_IB
+ pixel_6655/PIX_OUT pixel_6655/CSA_VREF pixel
Xpixel_6666 pixel_6666/gring pixel_6666/VDD pixel_6666/GND pixel_6666/VREF pixel_6666/ROW_SEL
+ pixel_6666/NB1 pixel_6666/VBIAS pixel_6666/NB2 pixel_6666/AMP_IN pixel_6666/SF_IB
+ pixel_6666/PIX_OUT pixel_6666/CSA_VREF pixel
Xpixel_6677 pixel_6677/gring pixel_6677/VDD pixel_6677/GND pixel_6677/VREF pixel_6677/ROW_SEL
+ pixel_6677/NB1 pixel_6677/VBIAS pixel_6677/NB2 pixel_6677/AMP_IN pixel_6677/SF_IB
+ pixel_6677/PIX_OUT pixel_6677/CSA_VREF pixel
Xpixel_6688 pixel_6688/gring pixel_6688/VDD pixel_6688/GND pixel_6688/VREF pixel_6688/ROW_SEL
+ pixel_6688/NB1 pixel_6688/VBIAS pixel_6688/NB2 pixel_6688/AMP_IN pixel_6688/SF_IB
+ pixel_6688/PIX_OUT pixel_6688/CSA_VREF pixel
Xpixel_5921 pixel_5921/gring pixel_5921/VDD pixel_5921/GND pixel_5921/VREF pixel_5921/ROW_SEL
+ pixel_5921/NB1 pixel_5921/VBIAS pixel_5921/NB2 pixel_5921/AMP_IN pixel_5921/SF_IB
+ pixel_5921/PIX_OUT pixel_5921/CSA_VREF pixel
Xpixel_5932 pixel_5932/gring pixel_5932/VDD pixel_5932/GND pixel_5932/VREF pixel_5932/ROW_SEL
+ pixel_5932/NB1 pixel_5932/VBIAS pixel_5932/NB2 pixel_5932/AMP_IN pixel_5932/SF_IB
+ pixel_5932/PIX_OUT pixel_5932/CSA_VREF pixel
Xpixel_5943 pixel_5943/gring pixel_5943/VDD pixel_5943/GND pixel_5943/VREF pixel_5943/ROW_SEL
+ pixel_5943/NB1 pixel_5943/VBIAS pixel_5943/NB2 pixel_5943/AMP_IN pixel_5943/SF_IB
+ pixel_5943/PIX_OUT pixel_5943/CSA_VREF pixel
Xpixel_6699 pixel_6699/gring pixel_6699/VDD pixel_6699/GND pixel_6699/VREF pixel_6699/ROW_SEL
+ pixel_6699/NB1 pixel_6699/VBIAS pixel_6699/NB2 pixel_6699/AMP_IN pixel_6699/SF_IB
+ pixel_6699/PIX_OUT pixel_6699/CSA_VREF pixel
Xpixel_5954 pixel_5954/gring pixel_5954/VDD pixel_5954/GND pixel_5954/VREF pixel_5954/ROW_SEL
+ pixel_5954/NB1 pixel_5954/VBIAS pixel_5954/NB2 pixel_5954/AMP_IN pixel_5954/SF_IB
+ pixel_5954/PIX_OUT pixel_5954/CSA_VREF pixel
Xpixel_5965 pixel_5965/gring pixel_5965/VDD pixel_5965/GND pixel_5965/VREF pixel_5965/ROW_SEL
+ pixel_5965/NB1 pixel_5965/VBIAS pixel_5965/NB2 pixel_5965/AMP_IN pixel_5965/SF_IB
+ pixel_5965/PIX_OUT pixel_5965/CSA_VREF pixel
Xpixel_5976 pixel_5976/gring pixel_5976/VDD pixel_5976/GND pixel_5976/VREF pixel_5976/ROW_SEL
+ pixel_5976/NB1 pixel_5976/VBIAS pixel_5976/NB2 pixel_5976/AMP_IN pixel_5976/SF_IB
+ pixel_5976/PIX_OUT pixel_5976/CSA_VREF pixel
Xpixel_5987 pixel_5987/gring pixel_5987/VDD pixel_5987/GND pixel_5987/VREF pixel_5987/ROW_SEL
+ pixel_5987/NB1 pixel_5987/VBIAS pixel_5987/NB2 pixel_5987/AMP_IN pixel_5987/SF_IB
+ pixel_5987/PIX_OUT pixel_5987/CSA_VREF pixel
Xpixel_5998 pixel_5998/gring pixel_5998/VDD pixel_5998/GND pixel_5998/VREF pixel_5998/ROW_SEL
+ pixel_5998/NB1 pixel_5998/VBIAS pixel_5998/NB2 pixel_5998/AMP_IN pixel_5998/SF_IB
+ pixel_5998/PIX_OUT pixel_5998/CSA_VREF pixel
Xpixel_9292 pixel_9292/gring pixel_9292/VDD pixel_9292/GND pixel_9292/VREF pixel_9292/ROW_SEL
+ pixel_9292/NB1 pixel_9292/VBIAS pixel_9292/NB2 pixel_9292/AMP_IN pixel_9292/SF_IB
+ pixel_9292/PIX_OUT pixel_9292/CSA_VREF pixel
Xpixel_9281 pixel_9281/gring pixel_9281/VDD pixel_9281/GND pixel_9281/VREF pixel_9281/ROW_SEL
+ pixel_9281/NB1 pixel_9281/VBIAS pixel_9281/NB2 pixel_9281/AMP_IN pixel_9281/SF_IB
+ pixel_9281/PIX_OUT pixel_9281/CSA_VREF pixel
Xpixel_9270 pixel_9270/gring pixel_9270/VDD pixel_9270/GND pixel_9270/VREF pixel_9270/ROW_SEL
+ pixel_9270/NB1 pixel_9270/VBIAS pixel_9270/NB2 pixel_9270/AMP_IN pixel_9270/SF_IB
+ pixel_9270/PIX_OUT pixel_9270/CSA_VREF pixel
Xpixel_8580 pixel_8580/gring pixel_8580/VDD pixel_8580/GND pixel_8580/VREF pixel_8580/ROW_SEL
+ pixel_8580/NB1 pixel_8580/VBIAS pixel_8580/NB2 pixel_8580/AMP_IN pixel_8580/SF_IB
+ pixel_8580/PIX_OUT pixel_8580/CSA_VREF pixel
Xpixel_8591 pixel_8591/gring pixel_8591/VDD pixel_8591/GND pixel_8591/VREF pixel_8591/ROW_SEL
+ pixel_8591/NB1 pixel_8591/VBIAS pixel_8591/NB2 pixel_8591/AMP_IN pixel_8591/SF_IB
+ pixel_8591/PIX_OUT pixel_8591/CSA_VREF pixel
Xpixel_7890 pixel_7890/gring pixel_7890/VDD pixel_7890/GND pixel_7890/VREF pixel_7890/ROW_SEL
+ pixel_7890/NB1 pixel_7890/VBIAS pixel_7890/NB2 pixel_7890/AMP_IN pixel_7890/SF_IB
+ pixel_7890/PIX_OUT pixel_7890/CSA_VREF pixel
Xpixel_5206 pixel_5206/gring pixel_5206/VDD pixel_5206/GND pixel_5206/VREF pixel_5206/ROW_SEL
+ pixel_5206/NB1 pixel_5206/VBIAS pixel_5206/NB2 pixel_5206/AMP_IN pixel_5206/SF_IB
+ pixel_5206/PIX_OUT pixel_5206/CSA_VREF pixel
Xpixel_5217 pixel_5217/gring pixel_5217/VDD pixel_5217/GND pixel_5217/VREF pixel_5217/ROW_SEL
+ pixel_5217/NB1 pixel_5217/VBIAS pixel_5217/NB2 pixel_5217/AMP_IN pixel_5217/SF_IB
+ pixel_5217/PIX_OUT pixel_5217/CSA_VREF pixel
Xpixel_5228 pixel_5228/gring pixel_5228/VDD pixel_5228/GND pixel_5228/VREF pixel_5228/ROW_SEL
+ pixel_5228/NB1 pixel_5228/VBIAS pixel_5228/NB2 pixel_5228/AMP_IN pixel_5228/SF_IB
+ pixel_5228/PIX_OUT pixel_5228/CSA_VREF pixel
Xpixel_5239 pixel_5239/gring pixel_5239/VDD pixel_5239/GND pixel_5239/VREF pixel_5239/ROW_SEL
+ pixel_5239/NB1 pixel_5239/VBIAS pixel_5239/NB2 pixel_5239/AMP_IN pixel_5239/SF_IB
+ pixel_5239/PIX_OUT pixel_5239/CSA_VREF pixel
Xpixel_522 pixel_522/gring pixel_522/VDD pixel_522/GND pixel_522/VREF pixel_522/ROW_SEL
+ pixel_522/NB1 pixel_522/VBIAS pixel_522/NB2 pixel_522/AMP_IN pixel_522/SF_IB pixel_522/PIX_OUT
+ pixel_522/CSA_VREF pixel
Xpixel_511 pixel_511/gring pixel_511/VDD pixel_511/GND pixel_511/VREF pixel_511/ROW_SEL
+ pixel_511/NB1 pixel_511/VBIAS pixel_511/NB2 pixel_511/AMP_IN pixel_511/SF_IB pixel_511/PIX_OUT
+ pixel_511/CSA_VREF pixel
Xpixel_500 pixel_500/gring pixel_500/VDD pixel_500/GND pixel_500/VREF pixel_500/ROW_SEL
+ pixel_500/NB1 pixel_500/VBIAS pixel_500/NB2 pixel_500/AMP_IN pixel_500/SF_IB pixel_500/PIX_OUT
+ pixel_500/CSA_VREF pixel
Xpixel_4505 pixel_4505/gring pixel_4505/VDD pixel_4505/GND pixel_4505/VREF pixel_4505/ROW_SEL
+ pixel_4505/NB1 pixel_4505/VBIAS pixel_4505/NB2 pixel_4505/AMP_IN pixel_4505/SF_IB
+ pixel_4505/PIX_OUT pixel_4505/CSA_VREF pixel
Xpixel_4516 pixel_4516/gring pixel_4516/VDD pixel_4516/GND pixel_4516/VREF pixel_4516/ROW_SEL
+ pixel_4516/NB1 pixel_4516/VBIAS pixel_4516/NB2 pixel_4516/AMP_IN pixel_4516/SF_IB
+ pixel_4516/PIX_OUT pixel_4516/CSA_VREF pixel
Xpixel_4527 pixel_4527/gring pixel_4527/VDD pixel_4527/GND pixel_4527/VREF pixel_4527/ROW_SEL
+ pixel_4527/NB1 pixel_4527/VBIAS pixel_4527/NB2 pixel_4527/AMP_IN pixel_4527/SF_IB
+ pixel_4527/PIX_OUT pixel_4527/CSA_VREF pixel
Xpixel_566 pixel_566/gring pixel_566/VDD pixel_566/GND pixel_566/VREF pixel_566/ROW_SEL
+ pixel_566/NB1 pixel_566/VBIAS pixel_566/NB2 pixel_566/AMP_IN pixel_566/SF_IB pixel_566/PIX_OUT
+ pixel_566/CSA_VREF pixel
Xpixel_555 pixel_555/gring pixel_555/VDD pixel_555/GND pixel_555/VREF pixel_555/ROW_SEL
+ pixel_555/NB1 pixel_555/VBIAS pixel_555/NB2 pixel_555/AMP_IN pixel_555/SF_IB pixel_555/PIX_OUT
+ pixel_555/CSA_VREF pixel
Xpixel_544 pixel_544/gring pixel_544/VDD pixel_544/GND pixel_544/VREF pixel_544/ROW_SEL
+ pixel_544/NB1 pixel_544/VBIAS pixel_544/NB2 pixel_544/AMP_IN pixel_544/SF_IB pixel_544/PIX_OUT
+ pixel_544/CSA_VREF pixel
Xpixel_533 pixel_533/gring pixel_533/VDD pixel_533/GND pixel_533/VREF pixel_533/ROW_SEL
+ pixel_533/NB1 pixel_533/VBIAS pixel_533/NB2 pixel_533/AMP_IN pixel_533/SF_IB pixel_533/PIX_OUT
+ pixel_533/CSA_VREF pixel
Xpixel_4538 pixel_4538/gring pixel_4538/VDD pixel_4538/GND pixel_4538/VREF pixel_4538/ROW_SEL
+ pixel_4538/NB1 pixel_4538/VBIAS pixel_4538/NB2 pixel_4538/AMP_IN pixel_4538/SF_IB
+ pixel_4538/PIX_OUT pixel_4538/CSA_VREF pixel
Xpixel_4549 pixel_4549/gring pixel_4549/VDD pixel_4549/GND pixel_4549/VREF pixel_4549/ROW_SEL
+ pixel_4549/NB1 pixel_4549/VBIAS pixel_4549/NB2 pixel_4549/AMP_IN pixel_4549/SF_IB
+ pixel_4549/PIX_OUT pixel_4549/CSA_VREF pixel
Xpixel_3804 pixel_3804/gring pixel_3804/VDD pixel_3804/GND pixel_3804/VREF pixel_3804/ROW_SEL
+ pixel_3804/NB1 pixel_3804/VBIAS pixel_3804/NB2 pixel_3804/AMP_IN pixel_3804/SF_IB
+ pixel_3804/PIX_OUT pixel_3804/CSA_VREF pixel
Xpixel_3815 pixel_3815/gring pixel_3815/VDD pixel_3815/GND pixel_3815/VREF pixel_3815/ROW_SEL
+ pixel_3815/NB1 pixel_3815/VBIAS pixel_3815/NB2 pixel_3815/AMP_IN pixel_3815/SF_IB
+ pixel_3815/PIX_OUT pixel_3815/CSA_VREF pixel
Xpixel_599 pixel_599/gring pixel_599/VDD pixel_599/GND pixel_599/VREF pixel_599/ROW_SEL
+ pixel_599/NB1 pixel_599/VBIAS pixel_599/NB2 pixel_599/AMP_IN pixel_599/SF_IB pixel_599/PIX_OUT
+ pixel_599/CSA_VREF pixel
Xpixel_588 pixel_588/gring pixel_588/VDD pixel_588/GND pixel_588/VREF pixel_588/ROW_SEL
+ pixel_588/NB1 pixel_588/VBIAS pixel_588/NB2 pixel_588/AMP_IN pixel_588/SF_IB pixel_588/PIX_OUT
+ pixel_588/CSA_VREF pixel
Xpixel_577 pixel_577/gring pixel_577/VDD pixel_577/GND pixel_577/VREF pixel_577/ROW_SEL
+ pixel_577/NB1 pixel_577/VBIAS pixel_577/NB2 pixel_577/AMP_IN pixel_577/SF_IB pixel_577/PIX_OUT
+ pixel_577/CSA_VREF pixel
Xpixel_3859 pixel_3859/gring pixel_3859/VDD pixel_3859/GND pixel_3859/VREF pixel_3859/ROW_SEL
+ pixel_3859/NB1 pixel_3859/VBIAS pixel_3859/NB2 pixel_3859/AMP_IN pixel_3859/SF_IB
+ pixel_3859/PIX_OUT pixel_3859/CSA_VREF pixel
Xpixel_3848 pixel_3848/gring pixel_3848/VDD pixel_3848/GND pixel_3848/VREF pixel_3848/ROW_SEL
+ pixel_3848/NB1 pixel_3848/VBIAS pixel_3848/NB2 pixel_3848/AMP_IN pixel_3848/SF_IB
+ pixel_3848/PIX_OUT pixel_3848/CSA_VREF pixel
Xpixel_3826 pixel_3826/gring pixel_3826/VDD pixel_3826/GND pixel_3826/VREF pixel_3826/ROW_SEL
+ pixel_3826/NB1 pixel_3826/VBIAS pixel_3826/NB2 pixel_3826/AMP_IN pixel_3826/SF_IB
+ pixel_3826/PIX_OUT pixel_3826/CSA_VREF pixel
Xpixel_3837 pixel_3837/gring pixel_3837/VDD pixel_3837/GND pixel_3837/VREF pixel_3837/ROW_SEL
+ pixel_3837/NB1 pixel_3837/VBIAS pixel_3837/NB2 pixel_3837/AMP_IN pixel_3837/SF_IB
+ pixel_3837/PIX_OUT pixel_3837/CSA_VREF pixel
Xpixel_7120 pixel_7120/gring pixel_7120/VDD pixel_7120/GND pixel_7120/VREF pixel_7120/ROW_SEL
+ pixel_7120/NB1 pixel_7120/VBIAS pixel_7120/NB2 pixel_7120/AMP_IN pixel_7120/SF_IB
+ pixel_7120/PIX_OUT pixel_7120/CSA_VREF pixel
Xpixel_7131 pixel_7131/gring pixel_7131/VDD pixel_7131/GND pixel_7131/VREF pixel_7131/ROW_SEL
+ pixel_7131/NB1 pixel_7131/VBIAS pixel_7131/NB2 pixel_7131/AMP_IN pixel_7131/SF_IB
+ pixel_7131/PIX_OUT pixel_7131/CSA_VREF pixel
Xpixel_7142 pixel_7142/gring pixel_7142/VDD pixel_7142/GND pixel_7142/VREF pixel_7142/ROW_SEL
+ pixel_7142/NB1 pixel_7142/VBIAS pixel_7142/NB2 pixel_7142/AMP_IN pixel_7142/SF_IB
+ pixel_7142/PIX_OUT pixel_7142/CSA_VREF pixel
Xpixel_7153 pixel_7153/gring pixel_7153/VDD pixel_7153/GND pixel_7153/VREF pixel_7153/ROW_SEL
+ pixel_7153/NB1 pixel_7153/VBIAS pixel_7153/NB2 pixel_7153/AMP_IN pixel_7153/SF_IB
+ pixel_7153/PIX_OUT pixel_7153/CSA_VREF pixel
Xpixel_7164 pixel_7164/gring pixel_7164/VDD pixel_7164/GND pixel_7164/VREF pixel_7164/ROW_SEL
+ pixel_7164/NB1 pixel_7164/VBIAS pixel_7164/NB2 pixel_7164/AMP_IN pixel_7164/SF_IB
+ pixel_7164/PIX_OUT pixel_7164/CSA_VREF pixel
Xpixel_7175 pixel_7175/gring pixel_7175/VDD pixel_7175/GND pixel_7175/VREF pixel_7175/ROW_SEL
+ pixel_7175/NB1 pixel_7175/VBIAS pixel_7175/NB2 pixel_7175/AMP_IN pixel_7175/SF_IB
+ pixel_7175/PIX_OUT pixel_7175/CSA_VREF pixel
Xpixel_7186 pixel_7186/gring pixel_7186/VDD pixel_7186/GND pixel_7186/VREF pixel_7186/ROW_SEL
+ pixel_7186/NB1 pixel_7186/VBIAS pixel_7186/NB2 pixel_7186/AMP_IN pixel_7186/SF_IB
+ pixel_7186/PIX_OUT pixel_7186/CSA_VREF pixel
Xpixel_7197 pixel_7197/gring pixel_7197/VDD pixel_7197/GND pixel_7197/VREF pixel_7197/ROW_SEL
+ pixel_7197/NB1 pixel_7197/VBIAS pixel_7197/NB2 pixel_7197/AMP_IN pixel_7197/SF_IB
+ pixel_7197/PIX_OUT pixel_7197/CSA_VREF pixel
Xpixel_6430 pixel_6430/gring pixel_6430/VDD pixel_6430/GND pixel_6430/VREF pixel_6430/ROW_SEL
+ pixel_6430/NB1 pixel_6430/VBIAS pixel_6430/NB2 pixel_6430/AMP_IN pixel_6430/SF_IB
+ pixel_6430/PIX_OUT pixel_6430/CSA_VREF pixel
Xpixel_6441 pixel_6441/gring pixel_6441/VDD pixel_6441/GND pixel_6441/VREF pixel_6441/ROW_SEL
+ pixel_6441/NB1 pixel_6441/VBIAS pixel_6441/NB2 pixel_6441/AMP_IN pixel_6441/SF_IB
+ pixel_6441/PIX_OUT pixel_6441/CSA_VREF pixel
Xpixel_6452 pixel_6452/gring pixel_6452/VDD pixel_6452/GND pixel_6452/VREF pixel_6452/ROW_SEL
+ pixel_6452/NB1 pixel_6452/VBIAS pixel_6452/NB2 pixel_6452/AMP_IN pixel_6452/SF_IB
+ pixel_6452/PIX_OUT pixel_6452/CSA_VREF pixel
Xpixel_6463 pixel_6463/gring pixel_6463/VDD pixel_6463/GND pixel_6463/VREF pixel_6463/ROW_SEL
+ pixel_6463/NB1 pixel_6463/VBIAS pixel_6463/NB2 pixel_6463/AMP_IN pixel_6463/SF_IB
+ pixel_6463/PIX_OUT pixel_6463/CSA_VREF pixel
Xpixel_6474 pixel_6474/gring pixel_6474/VDD pixel_6474/GND pixel_6474/VREF pixel_6474/ROW_SEL
+ pixel_6474/NB1 pixel_6474/VBIAS pixel_6474/NB2 pixel_6474/AMP_IN pixel_6474/SF_IB
+ pixel_6474/PIX_OUT pixel_6474/CSA_VREF pixel
Xpixel_6485 pixel_6485/gring pixel_6485/VDD pixel_6485/GND pixel_6485/VREF pixel_6485/ROW_SEL
+ pixel_6485/NB1 pixel_6485/VBIAS pixel_6485/NB2 pixel_6485/AMP_IN pixel_6485/SF_IB
+ pixel_6485/PIX_OUT pixel_6485/CSA_VREF pixel
Xpixel_6496 pixel_6496/gring pixel_6496/VDD pixel_6496/GND pixel_6496/VREF pixel_6496/ROW_SEL
+ pixel_6496/NB1 pixel_6496/VBIAS pixel_6496/NB2 pixel_6496/AMP_IN pixel_6496/SF_IB
+ pixel_6496/PIX_OUT pixel_6496/CSA_VREF pixel
Xpixel_5740 pixel_5740/gring pixel_5740/VDD pixel_5740/GND pixel_5740/VREF pixel_5740/ROW_SEL
+ pixel_5740/NB1 pixel_5740/VBIAS pixel_5740/NB2 pixel_5740/AMP_IN pixel_5740/SF_IB
+ pixel_5740/PIX_OUT pixel_5740/CSA_VREF pixel
Xpixel_5751 pixel_5751/gring pixel_5751/VDD pixel_5751/GND pixel_5751/VREF pixel_5751/ROW_SEL
+ pixel_5751/NB1 pixel_5751/VBIAS pixel_5751/NB2 pixel_5751/AMP_IN pixel_5751/SF_IB
+ pixel_5751/PIX_OUT pixel_5751/CSA_VREF pixel
Xpixel_5762 pixel_5762/gring pixel_5762/VDD pixel_5762/GND pixel_5762/VREF pixel_5762/ROW_SEL
+ pixel_5762/NB1 pixel_5762/VBIAS pixel_5762/NB2 pixel_5762/AMP_IN pixel_5762/SF_IB
+ pixel_5762/PIX_OUT pixel_5762/CSA_VREF pixel
Xpixel_5773 pixel_5773/gring pixel_5773/VDD pixel_5773/GND pixel_5773/VREF pixel_5773/ROW_SEL
+ pixel_5773/NB1 pixel_5773/VBIAS pixel_5773/NB2 pixel_5773/AMP_IN pixel_5773/SF_IB
+ pixel_5773/PIX_OUT pixel_5773/CSA_VREF pixel
Xpixel_5784 pixel_5784/gring pixel_5784/VDD pixel_5784/GND pixel_5784/VREF pixel_5784/ROW_SEL
+ pixel_5784/NB1 pixel_5784/VBIAS pixel_5784/NB2 pixel_5784/AMP_IN pixel_5784/SF_IB
+ pixel_5784/PIX_OUT pixel_5784/CSA_VREF pixel
Xpixel_5795 pixel_5795/gring pixel_5795/VDD pixel_5795/GND pixel_5795/VREF pixel_5795/ROW_SEL
+ pixel_5795/NB1 pixel_5795/VBIAS pixel_5795/NB2 pixel_5795/AMP_IN pixel_5795/SF_IB
+ pixel_5795/PIX_OUT pixel_5795/CSA_VREF pixel
Xpixel_1709 pixel_1709/gring pixel_1709/VDD pixel_1709/GND pixel_1709/VREF pixel_1709/ROW_SEL
+ pixel_1709/NB1 pixel_1709/VBIAS pixel_1709/NB2 pixel_1709/AMP_IN pixel_1709/SF_IB
+ pixel_1709/PIX_OUT pixel_1709/CSA_VREF pixel
Xpixel_5003 pixel_5003/gring pixel_5003/VDD pixel_5003/GND pixel_5003/VREF pixel_5003/ROW_SEL
+ pixel_5003/NB1 pixel_5003/VBIAS pixel_5003/NB2 pixel_5003/AMP_IN pixel_5003/SF_IB
+ pixel_5003/PIX_OUT pixel_5003/CSA_VREF pixel
Xpixel_5014 pixel_5014/gring pixel_5014/VDD pixel_5014/GND pixel_5014/VREF pixel_5014/ROW_SEL
+ pixel_5014/NB1 pixel_5014/VBIAS pixel_5014/NB2 pixel_5014/AMP_IN pixel_5014/SF_IB
+ pixel_5014/PIX_OUT pixel_5014/CSA_VREF pixel
Xpixel_5025 pixel_5025/gring pixel_5025/VDD pixel_5025/GND pixel_5025/VREF pixel_5025/ROW_SEL
+ pixel_5025/NB1 pixel_5025/VBIAS pixel_5025/NB2 pixel_5025/AMP_IN pixel_5025/SF_IB
+ pixel_5025/PIX_OUT pixel_5025/CSA_VREF pixel
Xpixel_5036 pixel_5036/gring pixel_5036/VDD pixel_5036/GND pixel_5036/VREF pixel_5036/ROW_SEL
+ pixel_5036/NB1 pixel_5036/VBIAS pixel_5036/NB2 pixel_5036/AMP_IN pixel_5036/SF_IB
+ pixel_5036/PIX_OUT pixel_5036/CSA_VREF pixel
Xpixel_5047 pixel_5047/gring pixel_5047/VDD pixel_5047/GND pixel_5047/VREF pixel_5047/ROW_SEL
+ pixel_5047/NB1 pixel_5047/VBIAS pixel_5047/NB2 pixel_5047/AMP_IN pixel_5047/SF_IB
+ pixel_5047/PIX_OUT pixel_5047/CSA_VREF pixel
Xpixel_4302 pixel_4302/gring pixel_4302/VDD pixel_4302/GND pixel_4302/VREF pixel_4302/ROW_SEL
+ pixel_4302/NB1 pixel_4302/VBIAS pixel_4302/NB2 pixel_4302/AMP_IN pixel_4302/SF_IB
+ pixel_4302/PIX_OUT pixel_4302/CSA_VREF pixel
Xpixel_330 pixel_330/gring pixel_330/VDD pixel_330/GND pixel_330/VREF pixel_330/ROW_SEL
+ pixel_330/NB1 pixel_330/VBIAS pixel_330/NB2 pixel_330/AMP_IN pixel_330/SF_IB pixel_330/PIX_OUT
+ pixel_330/CSA_VREF pixel
Xpixel_5058 pixel_5058/gring pixel_5058/VDD pixel_5058/GND pixel_5058/VREF pixel_5058/ROW_SEL
+ pixel_5058/NB1 pixel_5058/VBIAS pixel_5058/NB2 pixel_5058/AMP_IN pixel_5058/SF_IB
+ pixel_5058/PIX_OUT pixel_5058/CSA_VREF pixel
Xpixel_5069 pixel_5069/gring pixel_5069/VDD pixel_5069/GND pixel_5069/VREF pixel_5069/ROW_SEL
+ pixel_5069/NB1 pixel_5069/VBIAS pixel_5069/NB2 pixel_5069/AMP_IN pixel_5069/SF_IB
+ pixel_5069/PIX_OUT pixel_5069/CSA_VREF pixel
Xpixel_4313 pixel_4313/gring pixel_4313/VDD pixel_4313/GND pixel_4313/VREF pixel_4313/ROW_SEL
+ pixel_4313/NB1 pixel_4313/VBIAS pixel_4313/NB2 pixel_4313/AMP_IN pixel_4313/SF_IB
+ pixel_4313/PIX_OUT pixel_4313/CSA_VREF pixel
Xpixel_4324 pixel_4324/gring pixel_4324/VDD pixel_4324/GND pixel_4324/VREF pixel_4324/ROW_SEL
+ pixel_4324/NB1 pixel_4324/VBIAS pixel_4324/NB2 pixel_4324/AMP_IN pixel_4324/SF_IB
+ pixel_4324/PIX_OUT pixel_4324/CSA_VREF pixel
Xpixel_4335 pixel_4335/gring pixel_4335/VDD pixel_4335/GND pixel_4335/VREF pixel_4335/ROW_SEL
+ pixel_4335/NB1 pixel_4335/VBIAS pixel_4335/NB2 pixel_4335/AMP_IN pixel_4335/SF_IB
+ pixel_4335/PIX_OUT pixel_4335/CSA_VREF pixel
Xpixel_374 pixel_374/gring pixel_374/VDD pixel_374/GND pixel_374/VREF pixel_374/ROW_SEL
+ pixel_374/NB1 pixel_374/VBIAS pixel_374/NB2 pixel_374/AMP_IN pixel_374/SF_IB pixel_374/PIX_OUT
+ pixel_374/CSA_VREF pixel
Xpixel_363 pixel_363/gring pixel_363/VDD pixel_363/GND pixel_363/VREF pixel_363/ROW_SEL
+ pixel_363/NB1 pixel_363/VBIAS pixel_363/NB2 pixel_363/AMP_IN pixel_363/SF_IB pixel_363/PIX_OUT
+ pixel_363/CSA_VREF pixel
Xpixel_352 pixel_352/gring pixel_352/VDD pixel_352/GND pixel_352/VREF pixel_352/ROW_SEL
+ pixel_352/NB1 pixel_352/VBIAS pixel_352/NB2 pixel_352/AMP_IN pixel_352/SF_IB pixel_352/PIX_OUT
+ pixel_352/CSA_VREF pixel
Xpixel_341 pixel_341/gring pixel_341/VDD pixel_341/GND pixel_341/VREF pixel_341/ROW_SEL
+ pixel_341/NB1 pixel_341/VBIAS pixel_341/NB2 pixel_341/AMP_IN pixel_341/SF_IB pixel_341/PIX_OUT
+ pixel_341/CSA_VREF pixel
Xpixel_3634 pixel_3634/gring pixel_3634/VDD pixel_3634/GND pixel_3634/VREF pixel_3634/ROW_SEL
+ pixel_3634/NB1 pixel_3634/VBIAS pixel_3634/NB2 pixel_3634/AMP_IN pixel_3634/SF_IB
+ pixel_3634/PIX_OUT pixel_3634/CSA_VREF pixel
Xpixel_3623 pixel_3623/gring pixel_3623/VDD pixel_3623/GND pixel_3623/VREF pixel_3623/ROW_SEL
+ pixel_3623/NB1 pixel_3623/VBIAS pixel_3623/NB2 pixel_3623/AMP_IN pixel_3623/SF_IB
+ pixel_3623/PIX_OUT pixel_3623/CSA_VREF pixel
Xpixel_3612 pixel_3612/gring pixel_3612/VDD pixel_3612/GND pixel_3612/VREF pixel_3612/ROW_SEL
+ pixel_3612/NB1 pixel_3612/VBIAS pixel_3612/NB2 pixel_3612/AMP_IN pixel_3612/SF_IB
+ pixel_3612/PIX_OUT pixel_3612/CSA_VREF pixel
Xpixel_3601 pixel_3601/gring pixel_3601/VDD pixel_3601/GND pixel_3601/VREF pixel_3601/ROW_SEL
+ pixel_3601/NB1 pixel_3601/VBIAS pixel_3601/NB2 pixel_3601/AMP_IN pixel_3601/SF_IB
+ pixel_3601/PIX_OUT pixel_3601/CSA_VREF pixel
Xpixel_4346 pixel_4346/gring pixel_4346/VDD pixel_4346/GND pixel_4346/VREF pixel_4346/ROW_SEL
+ pixel_4346/NB1 pixel_4346/VBIAS pixel_4346/NB2 pixel_4346/AMP_IN pixel_4346/SF_IB
+ pixel_4346/PIX_OUT pixel_4346/CSA_VREF pixel
Xpixel_4357 pixel_4357/gring pixel_4357/VDD pixel_4357/GND pixel_4357/VREF pixel_4357/ROW_SEL
+ pixel_4357/NB1 pixel_4357/VBIAS pixel_4357/NB2 pixel_4357/AMP_IN pixel_4357/SF_IB
+ pixel_4357/PIX_OUT pixel_4357/CSA_VREF pixel
Xpixel_4368 pixel_4368/gring pixel_4368/VDD pixel_4368/GND pixel_4368/VREF pixel_4368/ROW_SEL
+ pixel_4368/NB1 pixel_4368/VBIAS pixel_4368/NB2 pixel_4368/AMP_IN pixel_4368/SF_IB
+ pixel_4368/PIX_OUT pixel_4368/CSA_VREF pixel
Xpixel_4379 pixel_4379/gring pixel_4379/VDD pixel_4379/GND pixel_4379/VREF pixel_4379/ROW_SEL
+ pixel_4379/NB1 pixel_4379/VBIAS pixel_4379/NB2 pixel_4379/AMP_IN pixel_4379/SF_IB
+ pixel_4379/PIX_OUT pixel_4379/CSA_VREF pixel
Xpixel_396 pixel_396/gring pixel_396/VDD pixel_396/GND pixel_396/VREF pixel_396/ROW_SEL
+ pixel_396/NB1 pixel_396/VBIAS pixel_396/NB2 pixel_396/AMP_IN pixel_396/SF_IB pixel_396/PIX_OUT
+ pixel_396/CSA_VREF pixel
Xpixel_385 pixel_385/gring pixel_385/VDD pixel_385/GND pixel_385/VREF pixel_385/ROW_SEL
+ pixel_385/NB1 pixel_385/VBIAS pixel_385/NB2 pixel_385/AMP_IN pixel_385/SF_IB pixel_385/PIX_OUT
+ pixel_385/CSA_VREF pixel
Xpixel_2922 pixel_2922/gring pixel_2922/VDD pixel_2922/GND pixel_2922/VREF pixel_2922/ROW_SEL
+ pixel_2922/NB1 pixel_2922/VBIAS pixel_2922/NB2 pixel_2922/AMP_IN pixel_2922/SF_IB
+ pixel_2922/PIX_OUT pixel_2922/CSA_VREF pixel
Xpixel_2911 pixel_2911/gring pixel_2911/VDD pixel_2911/GND pixel_2911/VREF pixel_2911/ROW_SEL
+ pixel_2911/NB1 pixel_2911/VBIAS pixel_2911/NB2 pixel_2911/AMP_IN pixel_2911/SF_IB
+ pixel_2911/PIX_OUT pixel_2911/CSA_VREF pixel
Xpixel_2900 pixel_2900/gring pixel_2900/VDD pixel_2900/GND pixel_2900/VREF pixel_2900/ROW_SEL
+ pixel_2900/NB1 pixel_2900/VBIAS pixel_2900/NB2 pixel_2900/AMP_IN pixel_2900/SF_IB
+ pixel_2900/PIX_OUT pixel_2900/CSA_VREF pixel
Xpixel_3667 pixel_3667/gring pixel_3667/VDD pixel_3667/GND pixel_3667/VREF pixel_3667/ROW_SEL
+ pixel_3667/NB1 pixel_3667/VBIAS pixel_3667/NB2 pixel_3667/AMP_IN pixel_3667/SF_IB
+ pixel_3667/PIX_OUT pixel_3667/CSA_VREF pixel
Xpixel_3656 pixel_3656/gring pixel_3656/VDD pixel_3656/GND pixel_3656/VREF pixel_3656/ROW_SEL
+ pixel_3656/NB1 pixel_3656/VBIAS pixel_3656/NB2 pixel_3656/AMP_IN pixel_3656/SF_IB
+ pixel_3656/PIX_OUT pixel_3656/CSA_VREF pixel
Xpixel_3645 pixel_3645/gring pixel_3645/VDD pixel_3645/GND pixel_3645/VREF pixel_3645/ROW_SEL
+ pixel_3645/NB1 pixel_3645/VBIAS pixel_3645/NB2 pixel_3645/AMP_IN pixel_3645/SF_IB
+ pixel_3645/PIX_OUT pixel_3645/CSA_VREF pixel
Xpixel_2955 pixel_2955/gring pixel_2955/VDD pixel_2955/GND pixel_2955/VREF pixel_2955/ROW_SEL
+ pixel_2955/NB1 pixel_2955/VBIAS pixel_2955/NB2 pixel_2955/AMP_IN pixel_2955/SF_IB
+ pixel_2955/PIX_OUT pixel_2955/CSA_VREF pixel
Xpixel_2944 pixel_2944/gring pixel_2944/VDD pixel_2944/GND pixel_2944/VREF pixel_2944/ROW_SEL
+ pixel_2944/NB1 pixel_2944/VBIAS pixel_2944/NB2 pixel_2944/AMP_IN pixel_2944/SF_IB
+ pixel_2944/PIX_OUT pixel_2944/CSA_VREF pixel
Xpixel_2933 pixel_2933/gring pixel_2933/VDD pixel_2933/GND pixel_2933/VREF pixel_2933/ROW_SEL
+ pixel_2933/NB1 pixel_2933/VBIAS pixel_2933/NB2 pixel_2933/AMP_IN pixel_2933/SF_IB
+ pixel_2933/PIX_OUT pixel_2933/CSA_VREF pixel
Xpixel_3689 pixel_3689/gring pixel_3689/VDD pixel_3689/GND pixel_3689/VREF pixel_3689/ROW_SEL
+ pixel_3689/NB1 pixel_3689/VBIAS pixel_3689/NB2 pixel_3689/AMP_IN pixel_3689/SF_IB
+ pixel_3689/PIX_OUT pixel_3689/CSA_VREF pixel
Xpixel_3678 pixel_3678/gring pixel_3678/VDD pixel_3678/GND pixel_3678/VREF pixel_3678/ROW_SEL
+ pixel_3678/NB1 pixel_3678/VBIAS pixel_3678/NB2 pixel_3678/AMP_IN pixel_3678/SF_IB
+ pixel_3678/PIX_OUT pixel_3678/CSA_VREF pixel
Xpixel_2999 pixel_2999/gring pixel_2999/VDD pixel_2999/GND pixel_2999/VREF pixel_2999/ROW_SEL
+ pixel_2999/NB1 pixel_2999/VBIAS pixel_2999/NB2 pixel_2999/AMP_IN pixel_2999/SF_IB
+ pixel_2999/PIX_OUT pixel_2999/CSA_VREF pixel
Xpixel_2988 pixel_2988/gring pixel_2988/VDD pixel_2988/GND pixel_2988/VREF pixel_2988/ROW_SEL
+ pixel_2988/NB1 pixel_2988/VBIAS pixel_2988/NB2 pixel_2988/AMP_IN pixel_2988/SF_IB
+ pixel_2988/PIX_OUT pixel_2988/CSA_VREF pixel
Xpixel_2977 pixel_2977/gring pixel_2977/VDD pixel_2977/GND pixel_2977/VREF pixel_2977/ROW_SEL
+ pixel_2977/NB1 pixel_2977/VBIAS pixel_2977/NB2 pixel_2977/AMP_IN pixel_2977/SF_IB
+ pixel_2977/PIX_OUT pixel_2977/CSA_VREF pixel
Xpixel_2966 pixel_2966/gring pixel_2966/VDD pixel_2966/GND pixel_2966/VREF pixel_2966/ROW_SEL
+ pixel_2966/NB1 pixel_2966/VBIAS pixel_2966/NB2 pixel_2966/AMP_IN pixel_2966/SF_IB
+ pixel_2966/PIX_OUT pixel_2966/CSA_VREF pixel
Xpixel_6260 pixel_6260/gring pixel_6260/VDD pixel_6260/GND pixel_6260/VREF pixel_6260/ROW_SEL
+ pixel_6260/NB1 pixel_6260/VBIAS pixel_6260/NB2 pixel_6260/AMP_IN pixel_6260/SF_IB
+ pixel_6260/PIX_OUT pixel_6260/CSA_VREF pixel
Xpixel_6271 pixel_6271/gring pixel_6271/VDD pixel_6271/GND pixel_6271/VREF pixel_6271/ROW_SEL
+ pixel_6271/NB1 pixel_6271/VBIAS pixel_6271/NB2 pixel_6271/AMP_IN pixel_6271/SF_IB
+ pixel_6271/PIX_OUT pixel_6271/CSA_VREF pixel
Xpixel_6282 pixel_6282/gring pixel_6282/VDD pixel_6282/GND pixel_6282/VREF pixel_6282/ROW_SEL
+ pixel_6282/NB1 pixel_6282/VBIAS pixel_6282/NB2 pixel_6282/AMP_IN pixel_6282/SF_IB
+ pixel_6282/PIX_OUT pixel_6282/CSA_VREF pixel
Xpixel_6293 pixel_6293/gring pixel_6293/VDD pixel_6293/GND pixel_6293/VREF pixel_6293/ROW_SEL
+ pixel_6293/NB1 pixel_6293/VBIAS pixel_6293/NB2 pixel_6293/AMP_IN pixel_6293/SF_IB
+ pixel_6293/PIX_OUT pixel_6293/CSA_VREF pixel
Xpixel_5570 pixel_5570/gring pixel_5570/VDD pixel_5570/GND pixel_5570/VREF pixel_5570/ROW_SEL
+ pixel_5570/NB1 pixel_5570/VBIAS pixel_5570/NB2 pixel_5570/AMP_IN pixel_5570/SF_IB
+ pixel_5570/PIX_OUT pixel_5570/CSA_VREF pixel
Xpixel_5581 pixel_5581/gring pixel_5581/VDD pixel_5581/GND pixel_5581/VREF pixel_5581/ROW_SEL
+ pixel_5581/NB1 pixel_5581/VBIAS pixel_5581/NB2 pixel_5581/AMP_IN pixel_5581/SF_IB
+ pixel_5581/PIX_OUT pixel_5581/CSA_VREF pixel
Xpixel_5592 pixel_5592/gring pixel_5592/VDD pixel_5592/GND pixel_5592/VREF pixel_5592/ROW_SEL
+ pixel_5592/NB1 pixel_5592/VBIAS pixel_5592/NB2 pixel_5592/AMP_IN pixel_5592/SF_IB
+ pixel_5592/PIX_OUT pixel_5592/CSA_VREF pixel
Xpixel_4880 pixel_4880/gring pixel_4880/VDD pixel_4880/GND pixel_4880/VREF pixel_4880/ROW_SEL
+ pixel_4880/NB1 pixel_4880/VBIAS pixel_4880/NB2 pixel_4880/AMP_IN pixel_4880/SF_IB
+ pixel_4880/PIX_OUT pixel_4880/CSA_VREF pixel
Xpixel_4891 pixel_4891/gring pixel_4891/VDD pixel_4891/GND pixel_4891/VREF pixel_4891/ROW_SEL
+ pixel_4891/NB1 pixel_4891/VBIAS pixel_4891/NB2 pixel_4891/AMP_IN pixel_4891/SF_IB
+ pixel_4891/PIX_OUT pixel_4891/CSA_VREF pixel
Xpixel_2218 pixel_2218/gring pixel_2218/VDD pixel_2218/GND pixel_2218/VREF pixel_2218/ROW_SEL
+ pixel_2218/NB1 pixel_2218/VBIAS pixel_2218/NB2 pixel_2218/AMP_IN pixel_2218/SF_IB
+ pixel_2218/PIX_OUT pixel_2218/CSA_VREF pixel
Xpixel_2207 pixel_2207/gring pixel_2207/VDD pixel_2207/GND pixel_2207/VREF pixel_2207/ROW_SEL
+ pixel_2207/NB1 pixel_2207/VBIAS pixel_2207/NB2 pixel_2207/AMP_IN pixel_2207/SF_IB
+ pixel_2207/PIX_OUT pixel_2207/CSA_VREF pixel
Xpixel_1506 pixel_1506/gring pixel_1506/VDD pixel_1506/GND pixel_1506/VREF pixel_1506/ROW_SEL
+ pixel_1506/NB1 pixel_1506/VBIAS pixel_1506/NB2 pixel_1506/AMP_IN pixel_1506/SF_IB
+ pixel_1506/PIX_OUT pixel_1506/CSA_VREF pixel
Xpixel_2229 pixel_2229/gring pixel_2229/VDD pixel_2229/GND pixel_2229/VREF pixel_2229/ROW_SEL
+ pixel_2229/NB1 pixel_2229/VBIAS pixel_2229/NB2 pixel_2229/AMP_IN pixel_2229/SF_IB
+ pixel_2229/PIX_OUT pixel_2229/CSA_VREF pixel
Xpixel_1539 pixel_1539/gring pixel_1539/VDD pixel_1539/GND pixel_1539/VREF pixel_1539/ROW_SEL
+ pixel_1539/NB1 pixel_1539/VBIAS pixel_1539/NB2 pixel_1539/AMP_IN pixel_1539/SF_IB
+ pixel_1539/PIX_OUT pixel_1539/CSA_VREF pixel
Xpixel_1528 pixel_1528/gring pixel_1528/VDD pixel_1528/GND pixel_1528/VREF pixel_1528/ROW_SEL
+ pixel_1528/NB1 pixel_1528/VBIAS pixel_1528/NB2 pixel_1528/AMP_IN pixel_1528/SF_IB
+ pixel_1528/PIX_OUT pixel_1528/CSA_VREF pixel
Xpixel_1517 pixel_1517/gring pixel_1517/VDD pixel_1517/GND pixel_1517/VREF pixel_1517/ROW_SEL
+ pixel_1517/NB1 pixel_1517/VBIAS pixel_1517/NB2 pixel_1517/AMP_IN pixel_1517/SF_IB
+ pixel_1517/PIX_OUT pixel_1517/CSA_VREF pixel
Xpixel_9814 pixel_9814/gring pixel_9814/VDD pixel_9814/GND pixel_9814/VREF pixel_9814/ROW_SEL
+ pixel_9814/NB1 pixel_9814/VBIAS pixel_9814/NB2 pixel_9814/AMP_IN pixel_9814/SF_IB
+ pixel_9814/PIX_OUT pixel_9814/CSA_VREF pixel
Xpixel_9803 pixel_9803/gring pixel_9803/VDD pixel_9803/GND pixel_9803/VREF pixel_9803/ROW_SEL
+ pixel_9803/NB1 pixel_9803/VBIAS pixel_9803/NB2 pixel_9803/AMP_IN pixel_9803/SF_IB
+ pixel_9803/PIX_OUT pixel_9803/CSA_VREF pixel
Xpixel_9847 pixel_9847/gring pixel_9847/VDD pixel_9847/GND pixel_9847/VREF pixel_9847/ROW_SEL
+ pixel_9847/NB1 pixel_9847/VBIAS pixel_9847/NB2 pixel_9847/AMP_IN pixel_9847/SF_IB
+ pixel_9847/PIX_OUT pixel_9847/CSA_VREF pixel
Xpixel_9836 pixel_9836/gring pixel_9836/VDD pixel_9836/GND pixel_9836/VREF pixel_9836/ROW_SEL
+ pixel_9836/NB1 pixel_9836/VBIAS pixel_9836/NB2 pixel_9836/AMP_IN pixel_9836/SF_IB
+ pixel_9836/PIX_OUT pixel_9836/CSA_VREF pixel
Xpixel_9825 pixel_9825/gring pixel_9825/VDD pixel_9825/GND pixel_9825/VREF pixel_9825/ROW_SEL
+ pixel_9825/NB1 pixel_9825/VBIAS pixel_9825/NB2 pixel_9825/AMP_IN pixel_9825/SF_IB
+ pixel_9825/PIX_OUT pixel_9825/CSA_VREF pixel
Xpixel_9858 pixel_9858/gring pixel_9858/VDD pixel_9858/GND pixel_9858/VREF pixel_9858/ROW_SEL
+ pixel_9858/NB1 pixel_9858/VBIAS pixel_9858/NB2 pixel_9858/AMP_IN pixel_9858/SF_IB
+ pixel_9858/PIX_OUT pixel_9858/CSA_VREF pixel
Xpixel_9869 pixel_9869/gring pixel_9869/VDD pixel_9869/GND pixel_9869/VREF pixel_9869/ROW_SEL
+ pixel_9869/NB1 pixel_9869/VBIAS pixel_9869/NB2 pixel_9869/AMP_IN pixel_9869/SF_IB
+ pixel_9869/PIX_OUT pixel_9869/CSA_VREF pixel
Xpixel_4110 pixel_4110/gring pixel_4110/VDD pixel_4110/GND pixel_4110/VREF pixel_4110/ROW_SEL
+ pixel_4110/NB1 pixel_4110/VBIAS pixel_4110/NB2 pixel_4110/AMP_IN pixel_4110/SF_IB
+ pixel_4110/PIX_OUT pixel_4110/CSA_VREF pixel
Xpixel_4121 pixel_4121/gring pixel_4121/VDD pixel_4121/GND pixel_4121/VREF pixel_4121/ROW_SEL
+ pixel_4121/NB1 pixel_4121/VBIAS pixel_4121/NB2 pixel_4121/AMP_IN pixel_4121/SF_IB
+ pixel_4121/PIX_OUT pixel_4121/CSA_VREF pixel
Xpixel_4132 pixel_4132/gring pixel_4132/VDD pixel_4132/GND pixel_4132/VREF pixel_4132/ROW_SEL
+ pixel_4132/NB1 pixel_4132/VBIAS pixel_4132/NB2 pixel_4132/AMP_IN pixel_4132/SF_IB
+ pixel_4132/PIX_OUT pixel_4132/CSA_VREF pixel
Xpixel_4143 pixel_4143/gring pixel_4143/VDD pixel_4143/GND pixel_4143/VREF pixel_4143/ROW_SEL
+ pixel_4143/NB1 pixel_4143/VBIAS pixel_4143/NB2 pixel_4143/AMP_IN pixel_4143/SF_IB
+ pixel_4143/PIX_OUT pixel_4143/CSA_VREF pixel
Xpixel_182 pixel_182/gring pixel_182/VDD pixel_182/GND pixel_182/VREF pixel_182/ROW_SEL
+ pixel_182/NB1 pixel_182/VBIAS pixel_182/NB2 pixel_182/AMP_IN pixel_182/SF_IB pixel_182/PIX_OUT
+ pixel_182/CSA_VREF pixel
Xpixel_171 pixel_171/gring pixel_171/VDD pixel_171/GND pixel_171/VREF pixel_171/ROW_SEL
+ pixel_171/NB1 pixel_171/VBIAS pixel_171/NB2 pixel_171/AMP_IN pixel_171/SF_IB pixel_171/PIX_OUT
+ pixel_171/CSA_VREF pixel
Xpixel_160 pixel_160/gring pixel_160/VDD pixel_160/GND pixel_160/VREF pixel_160/ROW_SEL
+ pixel_160/NB1 pixel_160/VBIAS pixel_160/NB2 pixel_160/AMP_IN pixel_160/SF_IB pixel_160/PIX_OUT
+ pixel_160/CSA_VREF pixel
Xpixel_3442 pixel_3442/gring pixel_3442/VDD pixel_3442/GND pixel_3442/VREF pixel_3442/ROW_SEL
+ pixel_3442/NB1 pixel_3442/VBIAS pixel_3442/NB2 pixel_3442/AMP_IN pixel_3442/SF_IB
+ pixel_3442/PIX_OUT pixel_3442/CSA_VREF pixel
Xpixel_3431 pixel_3431/gring pixel_3431/VDD pixel_3431/GND pixel_3431/VREF pixel_3431/ROW_SEL
+ pixel_3431/NB1 pixel_3431/VBIAS pixel_3431/NB2 pixel_3431/AMP_IN pixel_3431/SF_IB
+ pixel_3431/PIX_OUT pixel_3431/CSA_VREF pixel
Xpixel_3420 pixel_3420/gring pixel_3420/VDD pixel_3420/GND pixel_3420/VREF pixel_3420/ROW_SEL
+ pixel_3420/NB1 pixel_3420/VBIAS pixel_3420/NB2 pixel_3420/AMP_IN pixel_3420/SF_IB
+ pixel_3420/PIX_OUT pixel_3420/CSA_VREF pixel
Xpixel_4154 pixel_4154/gring pixel_4154/VDD pixel_4154/GND pixel_4154/VREF pixel_4154/ROW_SEL
+ pixel_4154/NB1 pixel_4154/VBIAS pixel_4154/NB2 pixel_4154/AMP_IN pixel_4154/SF_IB
+ pixel_4154/PIX_OUT pixel_4154/CSA_VREF pixel
Xpixel_4165 pixel_4165/gring pixel_4165/VDD pixel_4165/GND pixel_4165/VREF pixel_4165/ROW_SEL
+ pixel_4165/NB1 pixel_4165/VBIAS pixel_4165/NB2 pixel_4165/AMP_IN pixel_4165/SF_IB
+ pixel_4165/PIX_OUT pixel_4165/CSA_VREF pixel
Xpixel_4176 pixel_4176/gring pixel_4176/VDD pixel_4176/GND pixel_4176/VREF pixel_4176/ROW_SEL
+ pixel_4176/NB1 pixel_4176/VBIAS pixel_4176/NB2 pixel_4176/AMP_IN pixel_4176/SF_IB
+ pixel_4176/PIX_OUT pixel_4176/CSA_VREF pixel
Xpixel_4187 pixel_4187/gring pixel_4187/VDD pixel_4187/GND pixel_4187/VREF pixel_4187/ROW_SEL
+ pixel_4187/NB1 pixel_4187/VBIAS pixel_4187/NB2 pixel_4187/AMP_IN pixel_4187/SF_IB
+ pixel_4187/PIX_OUT pixel_4187/CSA_VREF pixel
Xpixel_193 pixel_193/gring pixel_193/VDD pixel_193/GND pixel_193/VREF pixel_193/ROW_SEL
+ pixel_193/NB1 pixel_193/VBIAS pixel_193/NB2 pixel_193/AMP_IN pixel_193/SF_IB pixel_193/PIX_OUT
+ pixel_193/CSA_VREF pixel
Xpixel_2730 pixel_2730/gring pixel_2730/VDD pixel_2730/GND pixel_2730/VREF pixel_2730/ROW_SEL
+ pixel_2730/NB1 pixel_2730/VBIAS pixel_2730/NB2 pixel_2730/AMP_IN pixel_2730/SF_IB
+ pixel_2730/PIX_OUT pixel_2730/CSA_VREF pixel
Xpixel_3475 pixel_3475/gring pixel_3475/VDD pixel_3475/GND pixel_3475/VREF pixel_3475/ROW_SEL
+ pixel_3475/NB1 pixel_3475/VBIAS pixel_3475/NB2 pixel_3475/AMP_IN pixel_3475/SF_IB
+ pixel_3475/PIX_OUT pixel_3475/CSA_VREF pixel
Xpixel_3464 pixel_3464/gring pixel_3464/VDD pixel_3464/GND pixel_3464/VREF pixel_3464/ROW_SEL
+ pixel_3464/NB1 pixel_3464/VBIAS pixel_3464/NB2 pixel_3464/AMP_IN pixel_3464/SF_IB
+ pixel_3464/PIX_OUT pixel_3464/CSA_VREF pixel
Xpixel_3453 pixel_3453/gring pixel_3453/VDD pixel_3453/GND pixel_3453/VREF pixel_3453/ROW_SEL
+ pixel_3453/NB1 pixel_3453/VBIAS pixel_3453/NB2 pixel_3453/AMP_IN pixel_3453/SF_IB
+ pixel_3453/PIX_OUT pixel_3453/CSA_VREF pixel
Xpixel_4198 pixel_4198/gring pixel_4198/VDD pixel_4198/GND pixel_4198/VREF pixel_4198/ROW_SEL
+ pixel_4198/NB1 pixel_4198/VBIAS pixel_4198/NB2 pixel_4198/AMP_IN pixel_4198/SF_IB
+ pixel_4198/PIX_OUT pixel_4198/CSA_VREF pixel
Xpixel_2774 pixel_2774/gring pixel_2774/VDD pixel_2774/GND pixel_2774/VREF pixel_2774/ROW_SEL
+ pixel_2774/NB1 pixel_2774/VBIAS pixel_2774/NB2 pixel_2774/AMP_IN pixel_2774/SF_IB
+ pixel_2774/PIX_OUT pixel_2774/CSA_VREF pixel
Xpixel_2763 pixel_2763/gring pixel_2763/VDD pixel_2763/GND pixel_2763/VREF pixel_2763/ROW_SEL
+ pixel_2763/NB1 pixel_2763/VBIAS pixel_2763/NB2 pixel_2763/AMP_IN pixel_2763/SF_IB
+ pixel_2763/PIX_OUT pixel_2763/CSA_VREF pixel
Xpixel_2752 pixel_2752/gring pixel_2752/VDD pixel_2752/GND pixel_2752/VREF pixel_2752/ROW_SEL
+ pixel_2752/NB1 pixel_2752/VBIAS pixel_2752/NB2 pixel_2752/AMP_IN pixel_2752/SF_IB
+ pixel_2752/PIX_OUT pixel_2752/CSA_VREF pixel
Xpixel_2741 pixel_2741/gring pixel_2741/VDD pixel_2741/GND pixel_2741/VREF pixel_2741/ROW_SEL
+ pixel_2741/NB1 pixel_2741/VBIAS pixel_2741/NB2 pixel_2741/AMP_IN pixel_2741/SF_IB
+ pixel_2741/PIX_OUT pixel_2741/CSA_VREF pixel
Xpixel_3497 pixel_3497/gring pixel_3497/VDD pixel_3497/GND pixel_3497/VREF pixel_3497/ROW_SEL
+ pixel_3497/NB1 pixel_3497/VBIAS pixel_3497/NB2 pixel_3497/AMP_IN pixel_3497/SF_IB
+ pixel_3497/PIX_OUT pixel_3497/CSA_VREF pixel
Xpixel_3486 pixel_3486/gring pixel_3486/VDD pixel_3486/GND pixel_3486/VREF pixel_3486/ROW_SEL
+ pixel_3486/NB1 pixel_3486/VBIAS pixel_3486/NB2 pixel_3486/AMP_IN pixel_3486/SF_IB
+ pixel_3486/PIX_OUT pixel_3486/CSA_VREF pixel
Xpixel_2796 pixel_2796/gring pixel_2796/VDD pixel_2796/GND pixel_2796/VREF pixel_2796/ROW_SEL
+ pixel_2796/NB1 pixel_2796/VBIAS pixel_2796/NB2 pixel_2796/AMP_IN pixel_2796/SF_IB
+ pixel_2796/PIX_OUT pixel_2796/CSA_VREF pixel
Xpixel_2785 pixel_2785/gring pixel_2785/VDD pixel_2785/GND pixel_2785/VREF pixel_2785/ROW_SEL
+ pixel_2785/NB1 pixel_2785/VBIAS pixel_2785/NB2 pixel_2785/AMP_IN pixel_2785/SF_IB
+ pixel_2785/PIX_OUT pixel_2785/CSA_VREF pixel
Xpixel_6090 pixel_6090/gring pixel_6090/VDD pixel_6090/GND pixel_6090/VREF pixel_6090/ROW_SEL
+ pixel_6090/NB1 pixel_6090/VBIAS pixel_6090/NB2 pixel_6090/AMP_IN pixel_6090/SF_IB
+ pixel_6090/PIX_OUT pixel_6090/CSA_VREF pixel
Xpixel_8409 pixel_8409/gring pixel_8409/VDD pixel_8409/GND pixel_8409/VREF pixel_8409/ROW_SEL
+ pixel_8409/NB1 pixel_8409/VBIAS pixel_8409/NB2 pixel_8409/AMP_IN pixel_8409/SF_IB
+ pixel_8409/PIX_OUT pixel_8409/CSA_VREF pixel
Xpixel_7708 pixel_7708/gring pixel_7708/VDD pixel_7708/GND pixel_7708/VREF pixel_7708/ROW_SEL
+ pixel_7708/NB1 pixel_7708/VBIAS pixel_7708/NB2 pixel_7708/AMP_IN pixel_7708/SF_IB
+ pixel_7708/PIX_OUT pixel_7708/CSA_VREF pixel
Xpixel_7719 pixel_7719/gring pixel_7719/VDD pixel_7719/GND pixel_7719/VREF pixel_7719/ROW_SEL
+ pixel_7719/NB1 pixel_7719/VBIAS pixel_7719/NB2 pixel_7719/AMP_IN pixel_7719/SF_IB
+ pixel_7719/PIX_OUT pixel_7719/CSA_VREF pixel
Xpixel_2026 pixel_2026/gring pixel_2026/VDD pixel_2026/GND pixel_2026/VREF pixel_2026/ROW_SEL
+ pixel_2026/NB1 pixel_2026/VBIAS pixel_2026/NB2 pixel_2026/AMP_IN pixel_2026/SF_IB
+ pixel_2026/PIX_OUT pixel_2026/CSA_VREF pixel
Xpixel_2015 pixel_2015/gring pixel_2015/VDD pixel_2015/GND pixel_2015/VREF pixel_2015/ROW_SEL
+ pixel_2015/NB1 pixel_2015/VBIAS pixel_2015/NB2 pixel_2015/AMP_IN pixel_2015/SF_IB
+ pixel_2015/PIX_OUT pixel_2015/CSA_VREF pixel
Xpixel_2004 pixel_2004/gring pixel_2004/VDD pixel_2004/GND pixel_2004/VREF pixel_2004/ROW_SEL
+ pixel_2004/NB1 pixel_2004/VBIAS pixel_2004/NB2 pixel_2004/AMP_IN pixel_2004/SF_IB
+ pixel_2004/PIX_OUT pixel_2004/CSA_VREF pixel
Xpixel_1314 pixel_1314/gring pixel_1314/VDD pixel_1314/GND pixel_1314/VREF pixel_1314/ROW_SEL
+ pixel_1314/NB1 pixel_1314/VBIAS pixel_1314/NB2 pixel_1314/AMP_IN pixel_1314/SF_IB
+ pixel_1314/PIX_OUT pixel_1314/CSA_VREF pixel
Xpixel_1303 pixel_1303/gring pixel_1303/VDD pixel_1303/GND pixel_1303/VREF pixel_1303/ROW_SEL
+ pixel_1303/NB1 pixel_1303/VBIAS pixel_1303/NB2 pixel_1303/AMP_IN pixel_1303/SF_IB
+ pixel_1303/PIX_OUT pixel_1303/CSA_VREF pixel
Xpixel_2059 pixel_2059/gring pixel_2059/VDD pixel_2059/GND pixel_2059/VREF pixel_2059/ROW_SEL
+ pixel_2059/NB1 pixel_2059/VBIAS pixel_2059/NB2 pixel_2059/AMP_IN pixel_2059/SF_IB
+ pixel_2059/PIX_OUT pixel_2059/CSA_VREF pixel
Xpixel_2048 pixel_2048/gring pixel_2048/VDD pixel_2048/GND pixel_2048/VREF pixel_2048/ROW_SEL
+ pixel_2048/NB1 pixel_2048/VBIAS pixel_2048/NB2 pixel_2048/AMP_IN pixel_2048/SF_IB
+ pixel_2048/PIX_OUT pixel_2048/CSA_VREF pixel
Xpixel_2037 pixel_2037/gring pixel_2037/VDD pixel_2037/GND pixel_2037/VREF pixel_2037/ROW_SEL
+ pixel_2037/NB1 pixel_2037/VBIAS pixel_2037/NB2 pixel_2037/AMP_IN pixel_2037/SF_IB
+ pixel_2037/PIX_OUT pixel_2037/CSA_VREF pixel
Xpixel_1358 pixel_1358/gring pixel_1358/VDD pixel_1358/GND pixel_1358/VREF pixel_1358/ROW_SEL
+ pixel_1358/NB1 pixel_1358/VBIAS pixel_1358/NB2 pixel_1358/AMP_IN pixel_1358/SF_IB
+ pixel_1358/PIX_OUT pixel_1358/CSA_VREF pixel
Xpixel_1347 pixel_1347/gring pixel_1347/VDD pixel_1347/GND pixel_1347/VREF pixel_1347/ROW_SEL
+ pixel_1347/NB1 pixel_1347/VBIAS pixel_1347/NB2 pixel_1347/AMP_IN pixel_1347/SF_IB
+ pixel_1347/PIX_OUT pixel_1347/CSA_VREF pixel
Xpixel_1336 pixel_1336/gring pixel_1336/VDD pixel_1336/GND pixel_1336/VREF pixel_1336/ROW_SEL
+ pixel_1336/NB1 pixel_1336/VBIAS pixel_1336/NB2 pixel_1336/AMP_IN pixel_1336/SF_IB
+ pixel_1336/PIX_OUT pixel_1336/CSA_VREF pixel
Xpixel_1325 pixel_1325/gring pixel_1325/VDD pixel_1325/GND pixel_1325/VREF pixel_1325/ROW_SEL
+ pixel_1325/NB1 pixel_1325/VBIAS pixel_1325/NB2 pixel_1325/AMP_IN pixel_1325/SF_IB
+ pixel_1325/PIX_OUT pixel_1325/CSA_VREF pixel
Xpixel_1369 pixel_1369/gring pixel_1369/VDD pixel_1369/GND pixel_1369/VREF pixel_1369/ROW_SEL
+ pixel_1369/NB1 pixel_1369/VBIAS pixel_1369/NB2 pixel_1369/AMP_IN pixel_1369/SF_IB
+ pixel_1369/PIX_OUT pixel_1369/CSA_VREF pixel
Xpixel_9600 pixel_9600/gring pixel_9600/VDD pixel_9600/GND pixel_9600/VREF pixel_9600/ROW_SEL
+ pixel_9600/NB1 pixel_9600/VBIAS pixel_9600/NB2 pixel_9600/AMP_IN pixel_9600/SF_IB
+ pixel_9600/PIX_OUT pixel_9600/CSA_VREF pixel
Xpixel_9611 pixel_9611/gring pixel_9611/VDD pixel_9611/GND pixel_9611/VREF pixel_9611/ROW_SEL
+ pixel_9611/NB1 pixel_9611/VBIAS pixel_9611/NB2 pixel_9611/AMP_IN pixel_9611/SF_IB
+ pixel_9611/PIX_OUT pixel_9611/CSA_VREF pixel
Xpixel_9622 pixel_9622/gring pixel_9622/VDD pixel_9622/GND pixel_9622/VREF pixel_9622/ROW_SEL
+ pixel_9622/NB1 pixel_9622/VBIAS pixel_9622/NB2 pixel_9622/AMP_IN pixel_9622/SF_IB
+ pixel_9622/PIX_OUT pixel_9622/CSA_VREF pixel
Xpixel_8921 pixel_8921/gring pixel_8921/VDD pixel_8921/GND pixel_8921/VREF pixel_8921/ROW_SEL
+ pixel_8921/NB1 pixel_8921/VBIAS pixel_8921/NB2 pixel_8921/AMP_IN pixel_8921/SF_IB
+ pixel_8921/PIX_OUT pixel_8921/CSA_VREF pixel
Xpixel_8910 pixel_8910/gring pixel_8910/VDD pixel_8910/GND pixel_8910/VREF pixel_8910/ROW_SEL
+ pixel_8910/NB1 pixel_8910/VBIAS pixel_8910/NB2 pixel_8910/AMP_IN pixel_8910/SF_IB
+ pixel_8910/PIX_OUT pixel_8910/CSA_VREF pixel
Xpixel_9633 pixel_9633/gring pixel_9633/VDD pixel_9633/GND pixel_9633/VREF pixel_9633/ROW_SEL
+ pixel_9633/NB1 pixel_9633/VBIAS pixel_9633/NB2 pixel_9633/AMP_IN pixel_9633/SF_IB
+ pixel_9633/PIX_OUT pixel_9633/CSA_VREF pixel
Xpixel_9644 pixel_9644/gring pixel_9644/VDD pixel_9644/GND pixel_9644/VREF pixel_9644/ROW_SEL
+ pixel_9644/NB1 pixel_9644/VBIAS pixel_9644/NB2 pixel_9644/AMP_IN pixel_9644/SF_IB
+ pixel_9644/PIX_OUT pixel_9644/CSA_VREF pixel
Xpixel_9655 pixel_9655/gring pixel_9655/VDD pixel_9655/GND pixel_9655/VREF pixel_9655/ROW_SEL
+ pixel_9655/NB1 pixel_9655/VBIAS pixel_9655/NB2 pixel_9655/AMP_IN pixel_9655/SF_IB
+ pixel_9655/PIX_OUT pixel_9655/CSA_VREF pixel
Xpixel_9666 pixel_9666/gring pixel_9666/VDD pixel_9666/GND pixel_9666/VREF pixel_9666/ROW_SEL
+ pixel_9666/NB1 pixel_9666/VBIAS pixel_9666/NB2 pixel_9666/AMP_IN pixel_9666/SF_IB
+ pixel_9666/PIX_OUT pixel_9666/CSA_VREF pixel
Xpixel_8954 pixel_8954/gring pixel_8954/VDD pixel_8954/GND pixel_8954/VREF pixel_8954/ROW_SEL
+ pixel_8954/NB1 pixel_8954/VBIAS pixel_8954/NB2 pixel_8954/AMP_IN pixel_8954/SF_IB
+ pixel_8954/PIX_OUT pixel_8954/CSA_VREF pixel
Xpixel_8943 pixel_8943/gring pixel_8943/VDD pixel_8943/GND pixel_8943/VREF pixel_8943/ROW_SEL
+ pixel_8943/NB1 pixel_8943/VBIAS pixel_8943/NB2 pixel_8943/AMP_IN pixel_8943/SF_IB
+ pixel_8943/PIX_OUT pixel_8943/CSA_VREF pixel
Xpixel_8932 pixel_8932/gring pixel_8932/VDD pixel_8932/GND pixel_8932/VREF pixel_8932/ROW_SEL
+ pixel_8932/NB1 pixel_8932/VBIAS pixel_8932/NB2 pixel_8932/AMP_IN pixel_8932/SF_IB
+ pixel_8932/PIX_OUT pixel_8932/CSA_VREF pixel
Xpixel_9699 pixel_9699/gring pixel_9699/VDD pixel_9699/GND pixel_9699/VREF pixel_9699/ROW_SEL
+ pixel_9699/NB1 pixel_9699/VBIAS pixel_9699/NB2 pixel_9699/AMP_IN pixel_9699/SF_IB
+ pixel_9699/PIX_OUT pixel_9699/CSA_VREF pixel
Xpixel_9688 pixel_9688/gring pixel_9688/VDD pixel_9688/GND pixel_9688/VREF pixel_9688/ROW_SEL
+ pixel_9688/NB1 pixel_9688/VBIAS pixel_9688/NB2 pixel_9688/AMP_IN pixel_9688/SF_IB
+ pixel_9688/PIX_OUT pixel_9688/CSA_VREF pixel
Xpixel_9677 pixel_9677/gring pixel_9677/VDD pixel_9677/GND pixel_9677/VREF pixel_9677/ROW_SEL
+ pixel_9677/NB1 pixel_9677/VBIAS pixel_9677/NB2 pixel_9677/AMP_IN pixel_9677/SF_IB
+ pixel_9677/PIX_OUT pixel_9677/CSA_VREF pixel
Xpixel_8987 pixel_8987/gring pixel_8987/VDD pixel_8987/GND pixel_8987/VREF pixel_8987/ROW_SEL
+ pixel_8987/NB1 pixel_8987/VBIAS pixel_8987/NB2 pixel_8987/AMP_IN pixel_8987/SF_IB
+ pixel_8987/PIX_OUT pixel_8987/CSA_VREF pixel
Xpixel_8976 pixel_8976/gring pixel_8976/VDD pixel_8976/GND pixel_8976/VREF pixel_8976/ROW_SEL
+ pixel_8976/NB1 pixel_8976/VBIAS pixel_8976/NB2 pixel_8976/AMP_IN pixel_8976/SF_IB
+ pixel_8976/PIX_OUT pixel_8976/CSA_VREF pixel
Xpixel_8965 pixel_8965/gring pixel_8965/VDD pixel_8965/GND pixel_8965/VREF pixel_8965/ROW_SEL
+ pixel_8965/NB1 pixel_8965/VBIAS pixel_8965/NB2 pixel_8965/AMP_IN pixel_8965/SF_IB
+ pixel_8965/PIX_OUT pixel_8965/CSA_VREF pixel
Xpixel_8998 pixel_8998/gring pixel_8998/VDD pixel_8998/GND pixel_8998/VREF pixel_8998/ROW_SEL
+ pixel_8998/NB1 pixel_8998/VBIAS pixel_8998/NB2 pixel_8998/AMP_IN pixel_8998/SF_IB
+ pixel_8998/PIX_OUT pixel_8998/CSA_VREF pixel
Xpixel_3250 pixel_3250/gring pixel_3250/VDD pixel_3250/GND pixel_3250/VREF pixel_3250/ROW_SEL
+ pixel_3250/NB1 pixel_3250/VBIAS pixel_3250/NB2 pixel_3250/AMP_IN pixel_3250/SF_IB
+ pixel_3250/PIX_OUT pixel_3250/CSA_VREF pixel
Xpixel_3283 pixel_3283/gring pixel_3283/VDD pixel_3283/GND pixel_3283/VREF pixel_3283/ROW_SEL
+ pixel_3283/NB1 pixel_3283/VBIAS pixel_3283/NB2 pixel_3283/AMP_IN pixel_3283/SF_IB
+ pixel_3283/PIX_OUT pixel_3283/CSA_VREF pixel
Xpixel_3272 pixel_3272/gring pixel_3272/VDD pixel_3272/GND pixel_3272/VREF pixel_3272/ROW_SEL
+ pixel_3272/NB1 pixel_3272/VBIAS pixel_3272/NB2 pixel_3272/AMP_IN pixel_3272/SF_IB
+ pixel_3272/PIX_OUT pixel_3272/CSA_VREF pixel
Xpixel_3261 pixel_3261/gring pixel_3261/VDD pixel_3261/GND pixel_3261/VREF pixel_3261/ROW_SEL
+ pixel_3261/NB1 pixel_3261/VBIAS pixel_3261/NB2 pixel_3261/AMP_IN pixel_3261/SF_IB
+ pixel_3261/PIX_OUT pixel_3261/CSA_VREF pixel
Xpixel_2582 pixel_2582/gring pixel_2582/VDD pixel_2582/GND pixel_2582/VREF pixel_2582/ROW_SEL
+ pixel_2582/NB1 pixel_2582/VBIAS pixel_2582/NB2 pixel_2582/AMP_IN pixel_2582/SF_IB
+ pixel_2582/PIX_OUT pixel_2582/CSA_VREF pixel
Xpixel_2571 pixel_2571/gring pixel_2571/VDD pixel_2571/GND pixel_2571/VREF pixel_2571/ROW_SEL
+ pixel_2571/NB1 pixel_2571/VBIAS pixel_2571/NB2 pixel_2571/AMP_IN pixel_2571/SF_IB
+ pixel_2571/PIX_OUT pixel_2571/CSA_VREF pixel
Xpixel_2560 pixel_2560/gring pixel_2560/VDD pixel_2560/GND pixel_2560/VREF pixel_2560/ROW_SEL
+ pixel_2560/NB1 pixel_2560/VBIAS pixel_2560/NB2 pixel_2560/AMP_IN pixel_2560/SF_IB
+ pixel_2560/PIX_OUT pixel_2560/CSA_VREF pixel
Xpixel_3294 pixel_3294/gring pixel_3294/VDD pixel_3294/GND pixel_3294/VREF pixel_3294/ROW_SEL
+ pixel_3294/NB1 pixel_3294/VBIAS pixel_3294/NB2 pixel_3294/AMP_IN pixel_3294/SF_IB
+ pixel_3294/PIX_OUT pixel_3294/CSA_VREF pixel
Xpixel_1870 pixel_1870/gring pixel_1870/VDD pixel_1870/GND pixel_1870/VREF pixel_1870/ROW_SEL
+ pixel_1870/NB1 pixel_1870/VBIAS pixel_1870/NB2 pixel_1870/AMP_IN pixel_1870/SF_IB
+ pixel_1870/PIX_OUT pixel_1870/CSA_VREF pixel
Xpixel_2593 pixel_2593/gring pixel_2593/VDD pixel_2593/GND pixel_2593/VREF pixel_2593/ROW_SEL
+ pixel_2593/NB1 pixel_2593/VBIAS pixel_2593/NB2 pixel_2593/AMP_IN pixel_2593/SF_IB
+ pixel_2593/PIX_OUT pixel_2593/CSA_VREF pixel
Xpixel_1892 pixel_1892/gring pixel_1892/VDD pixel_1892/GND pixel_1892/VREF pixel_1892/ROW_SEL
+ pixel_1892/NB1 pixel_1892/VBIAS pixel_1892/NB2 pixel_1892/AMP_IN pixel_1892/SF_IB
+ pixel_1892/PIX_OUT pixel_1892/CSA_VREF pixel
Xpixel_1881 pixel_1881/gring pixel_1881/VDD pixel_1881/GND pixel_1881/VREF pixel_1881/ROW_SEL
+ pixel_1881/NB1 pixel_1881/VBIAS pixel_1881/NB2 pixel_1881/AMP_IN pixel_1881/SF_IB
+ pixel_1881/PIX_OUT pixel_1881/CSA_VREF pixel
Xpixel_929 pixel_929/gring pixel_929/VDD pixel_929/GND pixel_929/VREF pixel_929/ROW_SEL
+ pixel_929/NB1 pixel_929/VBIAS pixel_929/NB2 pixel_929/AMP_IN pixel_929/SF_IB pixel_929/PIX_OUT
+ pixel_929/CSA_VREF pixel
Xpixel_918 pixel_918/gring pixel_918/VDD pixel_918/GND pixel_918/VREF pixel_918/ROW_SEL
+ pixel_918/NB1 pixel_918/VBIAS pixel_918/NB2 pixel_918/AMP_IN pixel_918/SF_IB pixel_918/PIX_OUT
+ pixel_918/CSA_VREF pixel
Xpixel_907 pixel_907/gring pixel_907/VDD pixel_907/GND pixel_907/VREF pixel_907/ROW_SEL
+ pixel_907/NB1 pixel_907/VBIAS pixel_907/NB2 pixel_907/AMP_IN pixel_907/SF_IB pixel_907/PIX_OUT
+ pixel_907/CSA_VREF pixel
Xpixel_8206 pixel_8206/gring pixel_8206/VDD pixel_8206/GND pixel_8206/VREF pixel_8206/ROW_SEL
+ pixel_8206/NB1 pixel_8206/VBIAS pixel_8206/NB2 pixel_8206/AMP_IN pixel_8206/SF_IB
+ pixel_8206/PIX_OUT pixel_8206/CSA_VREF pixel
Xpixel_8217 pixel_8217/gring pixel_8217/VDD pixel_8217/GND pixel_8217/VREF pixel_8217/ROW_SEL
+ pixel_8217/NB1 pixel_8217/VBIAS pixel_8217/NB2 pixel_8217/AMP_IN pixel_8217/SF_IB
+ pixel_8217/PIX_OUT pixel_8217/CSA_VREF pixel
Xpixel_8228 pixel_8228/gring pixel_8228/VDD pixel_8228/GND pixel_8228/VREF pixel_8228/ROW_SEL
+ pixel_8228/NB1 pixel_8228/VBIAS pixel_8228/NB2 pixel_8228/AMP_IN pixel_8228/SF_IB
+ pixel_8228/PIX_OUT pixel_8228/CSA_VREF pixel
Xpixel_8239 pixel_8239/gring pixel_8239/VDD pixel_8239/GND pixel_8239/VREF pixel_8239/ROW_SEL
+ pixel_8239/NB1 pixel_8239/VBIAS pixel_8239/NB2 pixel_8239/AMP_IN pixel_8239/SF_IB
+ pixel_8239/PIX_OUT pixel_8239/CSA_VREF pixel
Xpixel_7505 pixel_7505/gring pixel_7505/VDD pixel_7505/GND pixel_7505/VREF pixel_7505/ROW_SEL
+ pixel_7505/NB1 pixel_7505/VBIAS pixel_7505/NB2 pixel_7505/AMP_IN pixel_7505/SF_IB
+ pixel_7505/PIX_OUT pixel_7505/CSA_VREF pixel
Xpixel_7516 pixel_7516/gring pixel_7516/VDD pixel_7516/GND pixel_7516/VREF pixel_7516/ROW_SEL
+ pixel_7516/NB1 pixel_7516/VBIAS pixel_7516/NB2 pixel_7516/AMP_IN pixel_7516/SF_IB
+ pixel_7516/PIX_OUT pixel_7516/CSA_VREF pixel
Xpixel_7527 pixel_7527/gring pixel_7527/VDD pixel_7527/GND pixel_7527/VREF pixel_7527/ROW_SEL
+ pixel_7527/NB1 pixel_7527/VBIAS pixel_7527/NB2 pixel_7527/AMP_IN pixel_7527/SF_IB
+ pixel_7527/PIX_OUT pixel_7527/CSA_VREF pixel
Xpixel_7538 pixel_7538/gring pixel_7538/VDD pixel_7538/GND pixel_7538/VREF pixel_7538/ROW_SEL
+ pixel_7538/NB1 pixel_7538/VBIAS pixel_7538/NB2 pixel_7538/AMP_IN pixel_7538/SF_IB
+ pixel_7538/PIX_OUT pixel_7538/CSA_VREF pixel
Xpixel_7549 pixel_7549/gring pixel_7549/VDD pixel_7549/GND pixel_7549/VREF pixel_7549/ROW_SEL
+ pixel_7549/NB1 pixel_7549/VBIAS pixel_7549/NB2 pixel_7549/AMP_IN pixel_7549/SF_IB
+ pixel_7549/PIX_OUT pixel_7549/CSA_VREF pixel
Xpixel_6804 pixel_6804/gring pixel_6804/VDD pixel_6804/GND pixel_6804/VREF pixel_6804/ROW_SEL
+ pixel_6804/NB1 pixel_6804/VBIAS pixel_6804/NB2 pixel_6804/AMP_IN pixel_6804/SF_IB
+ pixel_6804/PIX_OUT pixel_6804/CSA_VREF pixel
Xpixel_6815 pixel_6815/gring pixel_6815/VDD pixel_6815/GND pixel_6815/VREF pixel_6815/ROW_SEL
+ pixel_6815/NB1 pixel_6815/VBIAS pixel_6815/NB2 pixel_6815/AMP_IN pixel_6815/SF_IB
+ pixel_6815/PIX_OUT pixel_6815/CSA_VREF pixel
Xpixel_6826 pixel_6826/gring pixel_6826/VDD pixel_6826/GND pixel_6826/VREF pixel_6826/ROW_SEL
+ pixel_6826/NB1 pixel_6826/VBIAS pixel_6826/NB2 pixel_6826/AMP_IN pixel_6826/SF_IB
+ pixel_6826/PIX_OUT pixel_6826/CSA_VREF pixel
Xpixel_6837 pixel_6837/gring pixel_6837/VDD pixel_6837/GND pixel_6837/VREF pixel_6837/ROW_SEL
+ pixel_6837/NB1 pixel_6837/VBIAS pixel_6837/NB2 pixel_6837/AMP_IN pixel_6837/SF_IB
+ pixel_6837/PIX_OUT pixel_6837/CSA_VREF pixel
Xpixel_6848 pixel_6848/gring pixel_6848/VDD pixel_6848/GND pixel_6848/VREF pixel_6848/ROW_SEL
+ pixel_6848/NB1 pixel_6848/VBIAS pixel_6848/NB2 pixel_6848/AMP_IN pixel_6848/SF_IB
+ pixel_6848/PIX_OUT pixel_6848/CSA_VREF pixel
Xpixel_6859 pixel_6859/gring pixel_6859/VDD pixel_6859/GND pixel_6859/VREF pixel_6859/ROW_SEL
+ pixel_6859/NB1 pixel_6859/VBIAS pixel_6859/NB2 pixel_6859/AMP_IN pixel_6859/SF_IB
+ pixel_6859/PIX_OUT pixel_6859/CSA_VREF pixel
Xpixel_1133 pixel_1133/gring pixel_1133/VDD pixel_1133/GND pixel_1133/VREF pixel_1133/ROW_SEL
+ pixel_1133/NB1 pixel_1133/VBIAS pixel_1133/NB2 pixel_1133/AMP_IN pixel_1133/SF_IB
+ pixel_1133/PIX_OUT pixel_1133/CSA_VREF pixel
Xpixel_1122 pixel_1122/gring pixel_1122/VDD pixel_1122/GND pixel_1122/VREF pixel_1122/ROW_SEL
+ pixel_1122/NB1 pixel_1122/VBIAS pixel_1122/NB2 pixel_1122/AMP_IN pixel_1122/SF_IB
+ pixel_1122/PIX_OUT pixel_1122/CSA_VREF pixel
Xpixel_1111 pixel_1111/gring pixel_1111/VDD pixel_1111/GND pixel_1111/VREF pixel_1111/ROW_SEL
+ pixel_1111/NB1 pixel_1111/VBIAS pixel_1111/NB2 pixel_1111/AMP_IN pixel_1111/SF_IB
+ pixel_1111/PIX_OUT pixel_1111/CSA_VREF pixel
Xpixel_1100 pixel_1100/gring pixel_1100/VDD pixel_1100/GND pixel_1100/VREF pixel_1100/ROW_SEL
+ pixel_1100/NB1 pixel_1100/VBIAS pixel_1100/NB2 pixel_1100/AMP_IN pixel_1100/SF_IB
+ pixel_1100/PIX_OUT pixel_1100/CSA_VREF pixel
Xpixel_1166 pixel_1166/gring pixel_1166/VDD pixel_1166/GND pixel_1166/VREF pixel_1166/ROW_SEL
+ pixel_1166/NB1 pixel_1166/VBIAS pixel_1166/NB2 pixel_1166/AMP_IN pixel_1166/SF_IB
+ pixel_1166/PIX_OUT pixel_1166/CSA_VREF pixel
Xpixel_1155 pixel_1155/gring pixel_1155/VDD pixel_1155/GND pixel_1155/VREF pixel_1155/ROW_SEL
+ pixel_1155/NB1 pixel_1155/VBIAS pixel_1155/NB2 pixel_1155/AMP_IN pixel_1155/SF_IB
+ pixel_1155/PIX_OUT pixel_1155/CSA_VREF pixel
Xpixel_1144 pixel_1144/gring pixel_1144/VDD pixel_1144/GND pixel_1144/VREF pixel_1144/ROW_SEL
+ pixel_1144/NB1 pixel_1144/VBIAS pixel_1144/NB2 pixel_1144/AMP_IN pixel_1144/SF_IB
+ pixel_1144/PIX_OUT pixel_1144/CSA_VREF pixel
Xpixel_1199 pixel_1199/gring pixel_1199/VDD pixel_1199/GND pixel_1199/VREF pixel_1199/ROW_SEL
+ pixel_1199/NB1 pixel_1199/VBIAS pixel_1199/NB2 pixel_1199/AMP_IN pixel_1199/SF_IB
+ pixel_1199/PIX_OUT pixel_1199/CSA_VREF pixel
Xpixel_1188 pixel_1188/gring pixel_1188/VDD pixel_1188/GND pixel_1188/VREF pixel_1188/ROW_SEL
+ pixel_1188/NB1 pixel_1188/VBIAS pixel_1188/NB2 pixel_1188/AMP_IN pixel_1188/SF_IB
+ pixel_1188/PIX_OUT pixel_1188/CSA_VREF pixel
Xpixel_1177 pixel_1177/gring pixel_1177/VDD pixel_1177/GND pixel_1177/VREF pixel_1177/ROW_SEL
+ pixel_1177/NB1 pixel_1177/VBIAS pixel_1177/NB2 pixel_1177/AMP_IN pixel_1177/SF_IB
+ pixel_1177/PIX_OUT pixel_1177/CSA_VREF pixel
Xpixel_9441 pixel_9441/gring pixel_9441/VDD pixel_9441/GND pixel_9441/VREF pixel_9441/ROW_SEL
+ pixel_9441/NB1 pixel_9441/VBIAS pixel_9441/NB2 pixel_9441/AMP_IN pixel_9441/SF_IB
+ pixel_9441/PIX_OUT pixel_9441/CSA_VREF pixel
Xpixel_9430 pixel_9430/gring pixel_9430/VDD pixel_9430/GND pixel_9430/VREF pixel_9430/ROW_SEL
+ pixel_9430/NB1 pixel_9430/VBIAS pixel_9430/NB2 pixel_9430/AMP_IN pixel_9430/SF_IB
+ pixel_9430/PIX_OUT pixel_9430/CSA_VREF pixel
Xpixel_9474 pixel_9474/gring pixel_9474/VDD pixel_9474/GND pixel_9474/VREF pixel_9474/ROW_SEL
+ pixel_9474/NB1 pixel_9474/VBIAS pixel_9474/NB2 pixel_9474/AMP_IN pixel_9474/SF_IB
+ pixel_9474/PIX_OUT pixel_9474/CSA_VREF pixel
Xpixel_9463 pixel_9463/gring pixel_9463/VDD pixel_9463/GND pixel_9463/VREF pixel_9463/ROW_SEL
+ pixel_9463/NB1 pixel_9463/VBIAS pixel_9463/NB2 pixel_9463/AMP_IN pixel_9463/SF_IB
+ pixel_9463/PIX_OUT pixel_9463/CSA_VREF pixel
Xpixel_9452 pixel_9452/gring pixel_9452/VDD pixel_9452/GND pixel_9452/VREF pixel_9452/ROW_SEL
+ pixel_9452/NB1 pixel_9452/VBIAS pixel_9452/NB2 pixel_9452/AMP_IN pixel_9452/SF_IB
+ pixel_9452/PIX_OUT pixel_9452/CSA_VREF pixel
Xpixel_8762 pixel_8762/gring pixel_8762/VDD pixel_8762/GND pixel_8762/VREF pixel_8762/ROW_SEL
+ pixel_8762/NB1 pixel_8762/VBIAS pixel_8762/NB2 pixel_8762/AMP_IN pixel_8762/SF_IB
+ pixel_8762/PIX_OUT pixel_8762/CSA_VREF pixel
Xpixel_8751 pixel_8751/gring pixel_8751/VDD pixel_8751/GND pixel_8751/VREF pixel_8751/ROW_SEL
+ pixel_8751/NB1 pixel_8751/VBIAS pixel_8751/NB2 pixel_8751/AMP_IN pixel_8751/SF_IB
+ pixel_8751/PIX_OUT pixel_8751/CSA_VREF pixel
Xpixel_8740 pixel_8740/gring pixel_8740/VDD pixel_8740/GND pixel_8740/VREF pixel_8740/ROW_SEL
+ pixel_8740/NB1 pixel_8740/VBIAS pixel_8740/NB2 pixel_8740/AMP_IN pixel_8740/SF_IB
+ pixel_8740/PIX_OUT pixel_8740/CSA_VREF pixel
Xpixel_9496 pixel_9496/gring pixel_9496/VDD pixel_9496/GND pixel_9496/VREF pixel_9496/ROW_SEL
+ pixel_9496/NB1 pixel_9496/VBIAS pixel_9496/NB2 pixel_9496/AMP_IN pixel_9496/SF_IB
+ pixel_9496/PIX_OUT pixel_9496/CSA_VREF pixel
Xpixel_9485 pixel_9485/gring pixel_9485/VDD pixel_9485/GND pixel_9485/VREF pixel_9485/ROW_SEL
+ pixel_9485/NB1 pixel_9485/VBIAS pixel_9485/NB2 pixel_9485/AMP_IN pixel_9485/SF_IB
+ pixel_9485/PIX_OUT pixel_9485/CSA_VREF pixel
Xpixel_8795 pixel_8795/gring pixel_8795/VDD pixel_8795/GND pixel_8795/VREF pixel_8795/ROW_SEL
+ pixel_8795/NB1 pixel_8795/VBIAS pixel_8795/NB2 pixel_8795/AMP_IN pixel_8795/SF_IB
+ pixel_8795/PIX_OUT pixel_8795/CSA_VREF pixel
Xpixel_8784 pixel_8784/gring pixel_8784/VDD pixel_8784/GND pixel_8784/VREF pixel_8784/ROW_SEL
+ pixel_8784/NB1 pixel_8784/VBIAS pixel_8784/NB2 pixel_8784/AMP_IN pixel_8784/SF_IB
+ pixel_8784/PIX_OUT pixel_8784/CSA_VREF pixel
Xpixel_8773 pixel_8773/gring pixel_8773/VDD pixel_8773/GND pixel_8773/VREF pixel_8773/ROW_SEL
+ pixel_8773/NB1 pixel_8773/VBIAS pixel_8773/NB2 pixel_8773/AMP_IN pixel_8773/SF_IB
+ pixel_8773/PIX_OUT pixel_8773/CSA_VREF pixel
Xpixel_3091 pixel_3091/gring pixel_3091/VDD pixel_3091/GND pixel_3091/VREF pixel_3091/ROW_SEL
+ pixel_3091/NB1 pixel_3091/VBIAS pixel_3091/NB2 pixel_3091/AMP_IN pixel_3091/SF_IB
+ pixel_3091/PIX_OUT pixel_3091/CSA_VREF pixel
Xpixel_3080 pixel_3080/gring pixel_3080/VDD pixel_3080/GND pixel_3080/VREF pixel_3080/ROW_SEL
+ pixel_3080/NB1 pixel_3080/VBIAS pixel_3080/NB2 pixel_3080/AMP_IN pixel_3080/SF_IB
+ pixel_3080/PIX_OUT pixel_3080/CSA_VREF pixel
Xpixel_2390 pixel_2390/gring pixel_2390/VDD pixel_2390/GND pixel_2390/VREF pixel_2390/ROW_SEL
+ pixel_2390/NB1 pixel_2390/VBIAS pixel_2390/NB2 pixel_2390/AMP_IN pixel_2390/SF_IB
+ pixel_2390/PIX_OUT pixel_2390/CSA_VREF pixel
Xpixel_715 pixel_715/gring pixel_715/VDD pixel_715/GND pixel_715/VREF pixel_715/ROW_SEL
+ pixel_715/NB1 pixel_715/VBIAS pixel_715/NB2 pixel_715/AMP_IN pixel_715/SF_IB pixel_715/PIX_OUT
+ pixel_715/CSA_VREF pixel
Xpixel_704 pixel_704/gring pixel_704/VDD pixel_704/GND pixel_704/VREF pixel_704/ROW_SEL
+ pixel_704/NB1 pixel_704/VBIAS pixel_704/NB2 pixel_704/AMP_IN pixel_704/SF_IB pixel_704/PIX_OUT
+ pixel_704/CSA_VREF pixel
Xpixel_4709 pixel_4709/gring pixel_4709/VDD pixel_4709/GND pixel_4709/VREF pixel_4709/ROW_SEL
+ pixel_4709/NB1 pixel_4709/VBIAS pixel_4709/NB2 pixel_4709/AMP_IN pixel_4709/SF_IB
+ pixel_4709/PIX_OUT pixel_4709/CSA_VREF pixel
Xpixel_748 pixel_748/gring pixel_748/VDD pixel_748/GND pixel_748/VREF pixel_748/ROW_SEL
+ pixel_748/NB1 pixel_748/VBIAS pixel_748/NB2 pixel_748/AMP_IN pixel_748/SF_IB pixel_748/PIX_OUT
+ pixel_748/CSA_VREF pixel
Xpixel_737 pixel_737/gring pixel_737/VDD pixel_737/GND pixel_737/VREF pixel_737/ROW_SEL
+ pixel_737/NB1 pixel_737/VBIAS pixel_737/NB2 pixel_737/AMP_IN pixel_737/SF_IB pixel_737/PIX_OUT
+ pixel_737/CSA_VREF pixel
Xpixel_726 pixel_726/gring pixel_726/VDD pixel_726/GND pixel_726/VREF pixel_726/ROW_SEL
+ pixel_726/NB1 pixel_726/VBIAS pixel_726/NB2 pixel_726/AMP_IN pixel_726/SF_IB pixel_726/PIX_OUT
+ pixel_726/CSA_VREF pixel
Xpixel_759 pixel_759/gring pixel_759/VDD pixel_759/GND pixel_759/VREF pixel_759/ROW_SEL
+ pixel_759/NB1 pixel_759/VBIAS pixel_759/NB2 pixel_759/AMP_IN pixel_759/SF_IB pixel_759/PIX_OUT
+ pixel_759/CSA_VREF pixel
Xpixel_8003 pixel_8003/gring pixel_8003/VDD pixel_8003/GND pixel_8003/VREF pixel_8003/ROW_SEL
+ pixel_8003/NB1 pixel_8003/VBIAS pixel_8003/NB2 pixel_8003/AMP_IN pixel_8003/SF_IB
+ pixel_8003/PIX_OUT pixel_8003/CSA_VREF pixel
Xpixel_8014 pixel_8014/gring pixel_8014/VDD pixel_8014/GND pixel_8014/VREF pixel_8014/ROW_SEL
+ pixel_8014/NB1 pixel_8014/VBIAS pixel_8014/NB2 pixel_8014/AMP_IN pixel_8014/SF_IB
+ pixel_8014/PIX_OUT pixel_8014/CSA_VREF pixel
Xpixel_8025 pixel_8025/gring pixel_8025/VDD pixel_8025/GND pixel_8025/VREF pixel_8025/ROW_SEL
+ pixel_8025/NB1 pixel_8025/VBIAS pixel_8025/NB2 pixel_8025/AMP_IN pixel_8025/SF_IB
+ pixel_8025/PIX_OUT pixel_8025/CSA_VREF pixel
Xpixel_8036 pixel_8036/gring pixel_8036/VDD pixel_8036/GND pixel_8036/VREF pixel_8036/ROW_SEL
+ pixel_8036/NB1 pixel_8036/VBIAS pixel_8036/NB2 pixel_8036/AMP_IN pixel_8036/SF_IB
+ pixel_8036/PIX_OUT pixel_8036/CSA_VREF pixel
Xpixel_8047 pixel_8047/gring pixel_8047/VDD pixel_8047/GND pixel_8047/VREF pixel_8047/ROW_SEL
+ pixel_8047/NB1 pixel_8047/VBIAS pixel_8047/NB2 pixel_8047/AMP_IN pixel_8047/SF_IB
+ pixel_8047/PIX_OUT pixel_8047/CSA_VREF pixel
Xpixel_8058 pixel_8058/gring pixel_8058/VDD pixel_8058/GND pixel_8058/VREF pixel_8058/ROW_SEL
+ pixel_8058/NB1 pixel_8058/VBIAS pixel_8058/NB2 pixel_8058/AMP_IN pixel_8058/SF_IB
+ pixel_8058/PIX_OUT pixel_8058/CSA_VREF pixel
Xpixel_7302 pixel_7302/gring pixel_7302/VDD pixel_7302/GND pixel_7302/VREF pixel_7302/ROW_SEL
+ pixel_7302/NB1 pixel_7302/VBIAS pixel_7302/NB2 pixel_7302/AMP_IN pixel_7302/SF_IB
+ pixel_7302/PIX_OUT pixel_7302/CSA_VREF pixel
Xpixel_7313 pixel_7313/gring pixel_7313/VDD pixel_7313/GND pixel_7313/VREF pixel_7313/ROW_SEL
+ pixel_7313/NB1 pixel_7313/VBIAS pixel_7313/NB2 pixel_7313/AMP_IN pixel_7313/SF_IB
+ pixel_7313/PIX_OUT pixel_7313/CSA_VREF pixel
Xpixel_8069 pixel_8069/gring pixel_8069/VDD pixel_8069/GND pixel_8069/VREF pixel_8069/ROW_SEL
+ pixel_8069/NB1 pixel_8069/VBIAS pixel_8069/NB2 pixel_8069/AMP_IN pixel_8069/SF_IB
+ pixel_8069/PIX_OUT pixel_8069/CSA_VREF pixel
Xpixel_7324 pixel_7324/gring pixel_7324/VDD pixel_7324/GND pixel_7324/VREF pixel_7324/ROW_SEL
+ pixel_7324/NB1 pixel_7324/VBIAS pixel_7324/NB2 pixel_7324/AMP_IN pixel_7324/SF_IB
+ pixel_7324/PIX_OUT pixel_7324/CSA_VREF pixel
Xpixel_7335 pixel_7335/gring pixel_7335/VDD pixel_7335/GND pixel_7335/VREF pixel_7335/ROW_SEL
+ pixel_7335/NB1 pixel_7335/VBIAS pixel_7335/NB2 pixel_7335/AMP_IN pixel_7335/SF_IB
+ pixel_7335/PIX_OUT pixel_7335/CSA_VREF pixel
Xpixel_7346 pixel_7346/gring pixel_7346/VDD pixel_7346/GND pixel_7346/VREF pixel_7346/ROW_SEL
+ pixel_7346/NB1 pixel_7346/VBIAS pixel_7346/NB2 pixel_7346/AMP_IN pixel_7346/SF_IB
+ pixel_7346/PIX_OUT pixel_7346/CSA_VREF pixel
Xpixel_7357 pixel_7357/gring pixel_7357/VDD pixel_7357/GND pixel_7357/VREF pixel_7357/ROW_SEL
+ pixel_7357/NB1 pixel_7357/VBIAS pixel_7357/NB2 pixel_7357/AMP_IN pixel_7357/SF_IB
+ pixel_7357/PIX_OUT pixel_7357/CSA_VREF pixel
Xpixel_6601 pixel_6601/gring pixel_6601/VDD pixel_6601/GND pixel_6601/VREF pixel_6601/ROW_SEL
+ pixel_6601/NB1 pixel_6601/VBIAS pixel_6601/NB2 pixel_6601/AMP_IN pixel_6601/SF_IB
+ pixel_6601/PIX_OUT pixel_6601/CSA_VREF pixel
Xpixel_6612 pixel_6612/gring pixel_6612/VDD pixel_6612/GND pixel_6612/VREF pixel_6612/ROW_SEL
+ pixel_6612/NB1 pixel_6612/VBIAS pixel_6612/NB2 pixel_6612/AMP_IN pixel_6612/SF_IB
+ pixel_6612/PIX_OUT pixel_6612/CSA_VREF pixel
Xpixel_7368 pixel_7368/gring pixel_7368/VDD pixel_7368/GND pixel_7368/VREF pixel_7368/ROW_SEL
+ pixel_7368/NB1 pixel_7368/VBIAS pixel_7368/NB2 pixel_7368/AMP_IN pixel_7368/SF_IB
+ pixel_7368/PIX_OUT pixel_7368/CSA_VREF pixel
Xpixel_7379 pixel_7379/gring pixel_7379/VDD pixel_7379/GND pixel_7379/VREF pixel_7379/ROW_SEL
+ pixel_7379/NB1 pixel_7379/VBIAS pixel_7379/NB2 pixel_7379/AMP_IN pixel_7379/SF_IB
+ pixel_7379/PIX_OUT pixel_7379/CSA_VREF pixel
Xpixel_6623 pixel_6623/gring pixel_6623/VDD pixel_6623/GND pixel_6623/VREF pixel_6623/ROW_SEL
+ pixel_6623/NB1 pixel_6623/VBIAS pixel_6623/NB2 pixel_6623/AMP_IN pixel_6623/SF_IB
+ pixel_6623/PIX_OUT pixel_6623/CSA_VREF pixel
Xpixel_6634 pixel_6634/gring pixel_6634/VDD pixel_6634/GND pixel_6634/VREF pixel_6634/ROW_SEL
+ pixel_6634/NB1 pixel_6634/VBIAS pixel_6634/NB2 pixel_6634/AMP_IN pixel_6634/SF_IB
+ pixel_6634/PIX_OUT pixel_6634/CSA_VREF pixel
Xpixel_6645 pixel_6645/gring pixel_6645/VDD pixel_6645/GND pixel_6645/VREF pixel_6645/ROW_SEL
+ pixel_6645/NB1 pixel_6645/VBIAS pixel_6645/NB2 pixel_6645/AMP_IN pixel_6645/SF_IB
+ pixel_6645/PIX_OUT pixel_6645/CSA_VREF pixel
Xpixel_5900 pixel_5900/gring pixel_5900/VDD pixel_5900/GND pixel_5900/VREF pixel_5900/ROW_SEL
+ pixel_5900/NB1 pixel_5900/VBIAS pixel_5900/NB2 pixel_5900/AMP_IN pixel_5900/SF_IB
+ pixel_5900/PIX_OUT pixel_5900/CSA_VREF pixel
Xpixel_6656 pixel_6656/gring pixel_6656/VDD pixel_6656/GND pixel_6656/VREF pixel_6656/ROW_SEL
+ pixel_6656/NB1 pixel_6656/VBIAS pixel_6656/NB2 pixel_6656/AMP_IN pixel_6656/SF_IB
+ pixel_6656/PIX_OUT pixel_6656/CSA_VREF pixel
Xpixel_6667 pixel_6667/gring pixel_6667/VDD pixel_6667/GND pixel_6667/VREF pixel_6667/ROW_SEL
+ pixel_6667/NB1 pixel_6667/VBIAS pixel_6667/NB2 pixel_6667/AMP_IN pixel_6667/SF_IB
+ pixel_6667/PIX_OUT pixel_6667/CSA_VREF pixel
Xpixel_6678 pixel_6678/gring pixel_6678/VDD pixel_6678/GND pixel_6678/VREF pixel_6678/ROW_SEL
+ pixel_6678/NB1 pixel_6678/VBIAS pixel_6678/NB2 pixel_6678/AMP_IN pixel_6678/SF_IB
+ pixel_6678/PIX_OUT pixel_6678/CSA_VREF pixel
Xpixel_5911 pixel_5911/gring pixel_5911/VDD pixel_5911/GND pixel_5911/VREF pixel_5911/ROW_SEL
+ pixel_5911/NB1 pixel_5911/VBIAS pixel_5911/NB2 pixel_5911/AMP_IN pixel_5911/SF_IB
+ pixel_5911/PIX_OUT pixel_5911/CSA_VREF pixel
Xpixel_5922 pixel_5922/gring pixel_5922/VDD pixel_5922/GND pixel_5922/VREF pixel_5922/ROW_SEL
+ pixel_5922/NB1 pixel_5922/VBIAS pixel_5922/NB2 pixel_5922/AMP_IN pixel_5922/SF_IB
+ pixel_5922/PIX_OUT pixel_5922/CSA_VREF pixel
Xpixel_5933 pixel_5933/gring pixel_5933/VDD pixel_5933/GND pixel_5933/VREF pixel_5933/ROW_SEL
+ pixel_5933/NB1 pixel_5933/VBIAS pixel_5933/NB2 pixel_5933/AMP_IN pixel_5933/SF_IB
+ pixel_5933/PIX_OUT pixel_5933/CSA_VREF pixel
Xpixel_6689 pixel_6689/gring pixel_6689/VDD pixel_6689/GND pixel_6689/VREF pixel_6689/ROW_SEL
+ pixel_6689/NB1 pixel_6689/VBIAS pixel_6689/NB2 pixel_6689/AMP_IN pixel_6689/SF_IB
+ pixel_6689/PIX_OUT pixel_6689/CSA_VREF pixel
Xpixel_5944 pixel_5944/gring pixel_5944/VDD pixel_5944/GND pixel_5944/VREF pixel_5944/ROW_SEL
+ pixel_5944/NB1 pixel_5944/VBIAS pixel_5944/NB2 pixel_5944/AMP_IN pixel_5944/SF_IB
+ pixel_5944/PIX_OUT pixel_5944/CSA_VREF pixel
Xpixel_5955 pixel_5955/gring pixel_5955/VDD pixel_5955/GND pixel_5955/VREF pixel_5955/ROW_SEL
+ pixel_5955/NB1 pixel_5955/VBIAS pixel_5955/NB2 pixel_5955/AMP_IN pixel_5955/SF_IB
+ pixel_5955/PIX_OUT pixel_5955/CSA_VREF pixel
Xpixel_5966 pixel_5966/gring pixel_5966/VDD pixel_5966/GND pixel_5966/VREF pixel_5966/ROW_SEL
+ pixel_5966/NB1 pixel_5966/VBIAS pixel_5966/NB2 pixel_5966/AMP_IN pixel_5966/SF_IB
+ pixel_5966/PIX_OUT pixel_5966/CSA_VREF pixel
Xpixel_5977 pixel_5977/gring pixel_5977/VDD pixel_5977/GND pixel_5977/VREF pixel_5977/ROW_SEL
+ pixel_5977/NB1 pixel_5977/VBIAS pixel_5977/NB2 pixel_5977/AMP_IN pixel_5977/SF_IB
+ pixel_5977/PIX_OUT pixel_5977/CSA_VREF pixel
Xpixel_5988 pixel_5988/gring pixel_5988/VDD pixel_5988/GND pixel_5988/VREF pixel_5988/ROW_SEL
+ pixel_5988/NB1 pixel_5988/VBIAS pixel_5988/NB2 pixel_5988/AMP_IN pixel_5988/SF_IB
+ pixel_5988/PIX_OUT pixel_5988/CSA_VREF pixel
Xpixel_5999 pixel_5999/gring pixel_5999/VDD pixel_5999/GND pixel_5999/VREF pixel_5999/ROW_SEL
+ pixel_5999/NB1 pixel_5999/VBIAS pixel_5999/NB2 pixel_5999/AMP_IN pixel_5999/SF_IB
+ pixel_5999/PIX_OUT pixel_5999/CSA_VREF pixel
Xpixel_9282 pixel_9282/gring pixel_9282/VDD pixel_9282/GND pixel_9282/VREF pixel_9282/ROW_SEL
+ pixel_9282/NB1 pixel_9282/VBIAS pixel_9282/NB2 pixel_9282/AMP_IN pixel_9282/SF_IB
+ pixel_9282/PIX_OUT pixel_9282/CSA_VREF pixel
Xpixel_9271 pixel_9271/gring pixel_9271/VDD pixel_9271/GND pixel_9271/VREF pixel_9271/ROW_SEL
+ pixel_9271/NB1 pixel_9271/VBIAS pixel_9271/NB2 pixel_9271/AMP_IN pixel_9271/SF_IB
+ pixel_9271/PIX_OUT pixel_9271/CSA_VREF pixel
Xpixel_9260 pixel_9260/gring pixel_9260/VDD pixel_9260/GND pixel_9260/VREF pixel_9260/ROW_SEL
+ pixel_9260/NB1 pixel_9260/VBIAS pixel_9260/NB2 pixel_9260/AMP_IN pixel_9260/SF_IB
+ pixel_9260/PIX_OUT pixel_9260/CSA_VREF pixel
Xpixel_8581 pixel_8581/gring pixel_8581/VDD pixel_8581/GND pixel_8581/VREF pixel_8581/ROW_SEL
+ pixel_8581/NB1 pixel_8581/VBIAS pixel_8581/NB2 pixel_8581/AMP_IN pixel_8581/SF_IB
+ pixel_8581/PIX_OUT pixel_8581/CSA_VREF pixel
Xpixel_8570 pixel_8570/gring pixel_8570/VDD pixel_8570/GND pixel_8570/VREF pixel_8570/ROW_SEL
+ pixel_8570/NB1 pixel_8570/VBIAS pixel_8570/NB2 pixel_8570/AMP_IN pixel_8570/SF_IB
+ pixel_8570/PIX_OUT pixel_8570/CSA_VREF pixel
Xpixel_9293 pixel_9293/gring pixel_9293/VDD pixel_9293/GND pixel_9293/VREF pixel_9293/ROW_SEL
+ pixel_9293/NB1 pixel_9293/VBIAS pixel_9293/NB2 pixel_9293/AMP_IN pixel_9293/SF_IB
+ pixel_9293/PIX_OUT pixel_9293/CSA_VREF pixel
Xpixel_8592 pixel_8592/gring pixel_8592/VDD pixel_8592/GND pixel_8592/VREF pixel_8592/ROW_SEL
+ pixel_8592/NB1 pixel_8592/VBIAS pixel_8592/NB2 pixel_8592/AMP_IN pixel_8592/SF_IB
+ pixel_8592/PIX_OUT pixel_8592/CSA_VREF pixel
Xpixel_7880 pixel_7880/gring pixel_7880/VDD pixel_7880/GND pixel_7880/VREF pixel_7880/ROW_SEL
+ pixel_7880/NB1 pixel_7880/VBIAS pixel_7880/NB2 pixel_7880/AMP_IN pixel_7880/SF_IB
+ pixel_7880/PIX_OUT pixel_7880/CSA_VREF pixel
Xpixel_7891 pixel_7891/gring pixel_7891/VDD pixel_7891/GND pixel_7891/VREF pixel_7891/ROW_SEL
+ pixel_7891/NB1 pixel_7891/VBIAS pixel_7891/NB2 pixel_7891/AMP_IN pixel_7891/SF_IB
+ pixel_7891/PIX_OUT pixel_7891/CSA_VREF pixel
Xpixel_5207 pixel_5207/gring pixel_5207/VDD pixel_5207/GND pixel_5207/VREF pixel_5207/ROW_SEL
+ pixel_5207/NB1 pixel_5207/VBIAS pixel_5207/NB2 pixel_5207/AMP_IN pixel_5207/SF_IB
+ pixel_5207/PIX_OUT pixel_5207/CSA_VREF pixel
Xpixel_5218 pixel_5218/gring pixel_5218/VDD pixel_5218/GND pixel_5218/VREF pixel_5218/ROW_SEL
+ pixel_5218/NB1 pixel_5218/VBIAS pixel_5218/NB2 pixel_5218/AMP_IN pixel_5218/SF_IB
+ pixel_5218/PIX_OUT pixel_5218/CSA_VREF pixel
Xpixel_5229 pixel_5229/gring pixel_5229/VDD pixel_5229/GND pixel_5229/VREF pixel_5229/ROW_SEL
+ pixel_5229/NB1 pixel_5229/VBIAS pixel_5229/NB2 pixel_5229/AMP_IN pixel_5229/SF_IB
+ pixel_5229/PIX_OUT pixel_5229/CSA_VREF pixel
Xpixel_523 pixel_523/gring pixel_523/VDD pixel_523/GND pixel_523/VREF pixel_523/ROW_SEL
+ pixel_523/NB1 pixel_523/VBIAS pixel_523/NB2 pixel_523/AMP_IN pixel_523/SF_IB pixel_523/PIX_OUT
+ pixel_523/CSA_VREF pixel
Xpixel_512 pixel_512/gring pixel_512/VDD pixel_512/GND pixel_512/VREF pixel_512/ROW_SEL
+ pixel_512/NB1 pixel_512/VBIAS pixel_512/NB2 pixel_512/AMP_IN pixel_512/SF_IB pixel_512/PIX_OUT
+ pixel_512/CSA_VREF pixel
Xpixel_501 pixel_501/gring pixel_501/VDD pixel_501/GND pixel_501/VREF pixel_501/ROW_SEL
+ pixel_501/NB1 pixel_501/VBIAS pixel_501/NB2 pixel_501/AMP_IN pixel_501/SF_IB pixel_501/PIX_OUT
+ pixel_501/CSA_VREF pixel
Xpixel_4506 pixel_4506/gring pixel_4506/VDD pixel_4506/GND pixel_4506/VREF pixel_4506/ROW_SEL
+ pixel_4506/NB1 pixel_4506/VBIAS pixel_4506/NB2 pixel_4506/AMP_IN pixel_4506/SF_IB
+ pixel_4506/PIX_OUT pixel_4506/CSA_VREF pixel
Xpixel_4517 pixel_4517/gring pixel_4517/VDD pixel_4517/GND pixel_4517/VREF pixel_4517/ROW_SEL
+ pixel_4517/NB1 pixel_4517/VBIAS pixel_4517/NB2 pixel_4517/AMP_IN pixel_4517/SF_IB
+ pixel_4517/PIX_OUT pixel_4517/CSA_VREF pixel
Xpixel_4528 pixel_4528/gring pixel_4528/VDD pixel_4528/GND pixel_4528/VREF pixel_4528/ROW_SEL
+ pixel_4528/NB1 pixel_4528/VBIAS pixel_4528/NB2 pixel_4528/AMP_IN pixel_4528/SF_IB
+ pixel_4528/PIX_OUT pixel_4528/CSA_VREF pixel
Xpixel_556 pixel_556/gring pixel_556/VDD pixel_556/GND pixel_556/VREF pixel_556/ROW_SEL
+ pixel_556/NB1 pixel_556/VBIAS pixel_556/NB2 pixel_556/AMP_IN pixel_556/SF_IB pixel_556/PIX_OUT
+ pixel_556/CSA_VREF pixel
Xpixel_545 pixel_545/gring pixel_545/VDD pixel_545/GND pixel_545/VREF pixel_545/ROW_SEL
+ pixel_545/NB1 pixel_545/VBIAS pixel_545/NB2 pixel_545/AMP_IN pixel_545/SF_IB pixel_545/PIX_OUT
+ pixel_545/CSA_VREF pixel
Xpixel_534 pixel_534/gring pixel_534/VDD pixel_534/GND pixel_534/VREF pixel_534/ROW_SEL
+ pixel_534/NB1 pixel_534/VBIAS pixel_534/NB2 pixel_534/AMP_IN pixel_534/SF_IB pixel_534/PIX_OUT
+ pixel_534/CSA_VREF pixel
Xpixel_4539 pixel_4539/gring pixel_4539/VDD pixel_4539/GND pixel_4539/VREF pixel_4539/ROW_SEL
+ pixel_4539/NB1 pixel_4539/VBIAS pixel_4539/NB2 pixel_4539/AMP_IN pixel_4539/SF_IB
+ pixel_4539/PIX_OUT pixel_4539/CSA_VREF pixel
Xpixel_3805 pixel_3805/gring pixel_3805/VDD pixel_3805/GND pixel_3805/VREF pixel_3805/ROW_SEL
+ pixel_3805/NB1 pixel_3805/VBIAS pixel_3805/NB2 pixel_3805/AMP_IN pixel_3805/SF_IB
+ pixel_3805/PIX_OUT pixel_3805/CSA_VREF pixel
Xpixel_3816 pixel_3816/gring pixel_3816/VDD pixel_3816/GND pixel_3816/VREF pixel_3816/ROW_SEL
+ pixel_3816/NB1 pixel_3816/VBIAS pixel_3816/NB2 pixel_3816/AMP_IN pixel_3816/SF_IB
+ pixel_3816/PIX_OUT pixel_3816/CSA_VREF pixel
Xpixel_589 pixel_589/gring pixel_589/VDD pixel_589/GND pixel_589/VREF pixel_589/ROW_SEL
+ pixel_589/NB1 pixel_589/VBIAS pixel_589/NB2 pixel_589/AMP_IN pixel_589/SF_IB pixel_589/PIX_OUT
+ pixel_589/CSA_VREF pixel
Xpixel_578 pixel_578/gring pixel_578/VDD pixel_578/GND pixel_578/VREF pixel_578/ROW_SEL
+ pixel_578/NB1 pixel_578/VBIAS pixel_578/NB2 pixel_578/AMP_IN pixel_578/SF_IB pixel_578/PIX_OUT
+ pixel_578/CSA_VREF pixel
Xpixel_567 pixel_567/gring pixel_567/VDD pixel_567/GND pixel_567/VREF pixel_567/ROW_SEL
+ pixel_567/NB1 pixel_567/VBIAS pixel_567/NB2 pixel_567/AMP_IN pixel_567/SF_IB pixel_567/PIX_OUT
+ pixel_567/CSA_VREF pixel
Xpixel_3849 pixel_3849/gring pixel_3849/VDD pixel_3849/GND pixel_3849/VREF pixel_3849/ROW_SEL
+ pixel_3849/NB1 pixel_3849/VBIAS pixel_3849/NB2 pixel_3849/AMP_IN pixel_3849/SF_IB
+ pixel_3849/PIX_OUT pixel_3849/CSA_VREF pixel
Xpixel_3827 pixel_3827/gring pixel_3827/VDD pixel_3827/GND pixel_3827/VREF pixel_3827/ROW_SEL
+ pixel_3827/NB1 pixel_3827/VBIAS pixel_3827/NB2 pixel_3827/AMP_IN pixel_3827/SF_IB
+ pixel_3827/PIX_OUT pixel_3827/CSA_VREF pixel
Xpixel_3838 pixel_3838/gring pixel_3838/VDD pixel_3838/GND pixel_3838/VREF pixel_3838/ROW_SEL
+ pixel_3838/NB1 pixel_3838/VBIAS pixel_3838/NB2 pixel_3838/AMP_IN pixel_3838/SF_IB
+ pixel_3838/PIX_OUT pixel_3838/CSA_VREF pixel
Xpixel_7110 pixel_7110/gring pixel_7110/VDD pixel_7110/GND pixel_7110/VREF pixel_7110/ROW_SEL
+ pixel_7110/NB1 pixel_7110/VBIAS pixel_7110/NB2 pixel_7110/AMP_IN pixel_7110/SF_IB
+ pixel_7110/PIX_OUT pixel_7110/CSA_VREF pixel
Xpixel_7121 pixel_7121/gring pixel_7121/VDD pixel_7121/GND pixel_7121/VREF pixel_7121/ROW_SEL
+ pixel_7121/NB1 pixel_7121/VBIAS pixel_7121/NB2 pixel_7121/AMP_IN pixel_7121/SF_IB
+ pixel_7121/PIX_OUT pixel_7121/CSA_VREF pixel
Xpixel_7132 pixel_7132/gring pixel_7132/VDD pixel_7132/GND pixel_7132/VREF pixel_7132/ROW_SEL
+ pixel_7132/NB1 pixel_7132/VBIAS pixel_7132/NB2 pixel_7132/AMP_IN pixel_7132/SF_IB
+ pixel_7132/PIX_OUT pixel_7132/CSA_VREF pixel
Xpixel_7143 pixel_7143/gring pixel_7143/VDD pixel_7143/GND pixel_7143/VREF pixel_7143/ROW_SEL
+ pixel_7143/NB1 pixel_7143/VBIAS pixel_7143/NB2 pixel_7143/AMP_IN pixel_7143/SF_IB
+ pixel_7143/PIX_OUT pixel_7143/CSA_VREF pixel
Xpixel_7154 pixel_7154/gring pixel_7154/VDD pixel_7154/GND pixel_7154/VREF pixel_7154/ROW_SEL
+ pixel_7154/NB1 pixel_7154/VBIAS pixel_7154/NB2 pixel_7154/AMP_IN pixel_7154/SF_IB
+ pixel_7154/PIX_OUT pixel_7154/CSA_VREF pixel
Xpixel_7165 pixel_7165/gring pixel_7165/VDD pixel_7165/GND pixel_7165/VREF pixel_7165/ROW_SEL
+ pixel_7165/NB1 pixel_7165/VBIAS pixel_7165/NB2 pixel_7165/AMP_IN pixel_7165/SF_IB
+ pixel_7165/PIX_OUT pixel_7165/CSA_VREF pixel
Xpixel_6420 pixel_6420/gring pixel_6420/VDD pixel_6420/GND pixel_6420/VREF pixel_6420/ROW_SEL
+ pixel_6420/NB1 pixel_6420/VBIAS pixel_6420/NB2 pixel_6420/AMP_IN pixel_6420/SF_IB
+ pixel_6420/PIX_OUT pixel_6420/CSA_VREF pixel
Xpixel_7176 pixel_7176/gring pixel_7176/VDD pixel_7176/GND pixel_7176/VREF pixel_7176/ROW_SEL
+ pixel_7176/NB1 pixel_7176/VBIAS pixel_7176/NB2 pixel_7176/AMP_IN pixel_7176/SF_IB
+ pixel_7176/PIX_OUT pixel_7176/CSA_VREF pixel
Xpixel_7187 pixel_7187/gring pixel_7187/VDD pixel_7187/GND pixel_7187/VREF pixel_7187/ROW_SEL
+ pixel_7187/NB1 pixel_7187/VBIAS pixel_7187/NB2 pixel_7187/AMP_IN pixel_7187/SF_IB
+ pixel_7187/PIX_OUT pixel_7187/CSA_VREF pixel
Xpixel_7198 pixel_7198/gring pixel_7198/VDD pixel_7198/GND pixel_7198/VREF pixel_7198/ROW_SEL
+ pixel_7198/NB1 pixel_7198/VBIAS pixel_7198/NB2 pixel_7198/AMP_IN pixel_7198/SF_IB
+ pixel_7198/PIX_OUT pixel_7198/CSA_VREF pixel
Xpixel_6431 pixel_6431/gring pixel_6431/VDD pixel_6431/GND pixel_6431/VREF pixel_6431/ROW_SEL
+ pixel_6431/NB1 pixel_6431/VBIAS pixel_6431/NB2 pixel_6431/AMP_IN pixel_6431/SF_IB
+ pixel_6431/PIX_OUT pixel_6431/CSA_VREF pixel
Xpixel_6442 pixel_6442/gring pixel_6442/VDD pixel_6442/GND pixel_6442/VREF pixel_6442/ROW_SEL
+ pixel_6442/NB1 pixel_6442/VBIAS pixel_6442/NB2 pixel_6442/AMP_IN pixel_6442/SF_IB
+ pixel_6442/PIX_OUT pixel_6442/CSA_VREF pixel
Xpixel_6453 pixel_6453/gring pixel_6453/VDD pixel_6453/GND pixel_6453/VREF pixel_6453/ROW_SEL
+ pixel_6453/NB1 pixel_6453/VBIAS pixel_6453/NB2 pixel_6453/AMP_IN pixel_6453/SF_IB
+ pixel_6453/PIX_OUT pixel_6453/CSA_VREF pixel
Xpixel_6464 pixel_6464/gring pixel_6464/VDD pixel_6464/GND pixel_6464/VREF pixel_6464/ROW_SEL
+ pixel_6464/NB1 pixel_6464/VBIAS pixel_6464/NB2 pixel_6464/AMP_IN pixel_6464/SF_IB
+ pixel_6464/PIX_OUT pixel_6464/CSA_VREF pixel
Xpixel_6475 pixel_6475/gring pixel_6475/VDD pixel_6475/GND pixel_6475/VREF pixel_6475/ROW_SEL
+ pixel_6475/NB1 pixel_6475/VBIAS pixel_6475/NB2 pixel_6475/AMP_IN pixel_6475/SF_IB
+ pixel_6475/PIX_OUT pixel_6475/CSA_VREF pixel
Xpixel_6486 pixel_6486/gring pixel_6486/VDD pixel_6486/GND pixel_6486/VREF pixel_6486/ROW_SEL
+ pixel_6486/NB1 pixel_6486/VBIAS pixel_6486/NB2 pixel_6486/AMP_IN pixel_6486/SF_IB
+ pixel_6486/PIX_OUT pixel_6486/CSA_VREF pixel
Xpixel_5730 pixel_5730/gring pixel_5730/VDD pixel_5730/GND pixel_5730/VREF pixel_5730/ROW_SEL
+ pixel_5730/NB1 pixel_5730/VBIAS pixel_5730/NB2 pixel_5730/AMP_IN pixel_5730/SF_IB
+ pixel_5730/PIX_OUT pixel_5730/CSA_VREF pixel
Xpixel_5741 pixel_5741/gring pixel_5741/VDD pixel_5741/GND pixel_5741/VREF pixel_5741/ROW_SEL
+ pixel_5741/NB1 pixel_5741/VBIAS pixel_5741/NB2 pixel_5741/AMP_IN pixel_5741/SF_IB
+ pixel_5741/PIX_OUT pixel_5741/CSA_VREF pixel
Xpixel_5752 pixel_5752/gring pixel_5752/VDD pixel_5752/GND pixel_5752/VREF pixel_5752/ROW_SEL
+ pixel_5752/NB1 pixel_5752/VBIAS pixel_5752/NB2 pixel_5752/AMP_IN pixel_5752/SF_IB
+ pixel_5752/PIX_OUT pixel_5752/CSA_VREF pixel
Xpixel_6497 pixel_6497/gring pixel_6497/VDD pixel_6497/GND pixel_6497/VREF pixel_6497/ROW_SEL
+ pixel_6497/NB1 pixel_6497/VBIAS pixel_6497/NB2 pixel_6497/AMP_IN pixel_6497/SF_IB
+ pixel_6497/PIX_OUT pixel_6497/CSA_VREF pixel
Xpixel_5763 pixel_5763/gring pixel_5763/VDD pixel_5763/GND pixel_5763/VREF pixel_5763/ROW_SEL
+ pixel_5763/NB1 pixel_5763/VBIAS pixel_5763/NB2 pixel_5763/AMP_IN pixel_5763/SF_IB
+ pixel_5763/PIX_OUT pixel_5763/CSA_VREF pixel
Xpixel_5774 pixel_5774/gring pixel_5774/VDD pixel_5774/GND pixel_5774/VREF pixel_5774/ROW_SEL
+ pixel_5774/NB1 pixel_5774/VBIAS pixel_5774/NB2 pixel_5774/AMP_IN pixel_5774/SF_IB
+ pixel_5774/PIX_OUT pixel_5774/CSA_VREF pixel
Xpixel_5785 pixel_5785/gring pixel_5785/VDD pixel_5785/GND pixel_5785/VREF pixel_5785/ROW_SEL
+ pixel_5785/NB1 pixel_5785/VBIAS pixel_5785/NB2 pixel_5785/AMP_IN pixel_5785/SF_IB
+ pixel_5785/PIX_OUT pixel_5785/CSA_VREF pixel
Xpixel_5796 pixel_5796/gring pixel_5796/VDD pixel_5796/GND pixel_5796/VREF pixel_5796/ROW_SEL
+ pixel_5796/NB1 pixel_5796/VBIAS pixel_5796/NB2 pixel_5796/AMP_IN pixel_5796/SF_IB
+ pixel_5796/PIX_OUT pixel_5796/CSA_VREF pixel
Xpixel_9090 pixel_9090/gring pixel_9090/VDD pixel_9090/GND pixel_9090/VREF pixel_9090/ROW_SEL
+ pixel_9090/NB1 pixel_9090/VBIAS pixel_9090/NB2 pixel_9090/AMP_IN pixel_9090/SF_IB
+ pixel_9090/PIX_OUT pixel_9090/CSA_VREF pixel
Xpixel_90 pixel_90/gring pixel_90/VDD pixel_90/GND pixel_90/VREF pixel_90/ROW_SEL
+ pixel_90/NB1 pixel_90/VBIAS pixel_90/NB2 pixel_90/AMP_IN pixel_90/SF_IB pixel_90/PIX_OUT
+ pixel_90/CSA_VREF pixel
Xpixel_5004 pixel_5004/gring pixel_5004/VDD pixel_5004/GND pixel_5004/VREF pixel_5004/ROW_SEL
+ pixel_5004/NB1 pixel_5004/VBIAS pixel_5004/NB2 pixel_5004/AMP_IN pixel_5004/SF_IB
+ pixel_5004/PIX_OUT pixel_5004/CSA_VREF pixel
Xpixel_5015 pixel_5015/gring pixel_5015/VDD pixel_5015/GND pixel_5015/VREF pixel_5015/ROW_SEL
+ pixel_5015/NB1 pixel_5015/VBIAS pixel_5015/NB2 pixel_5015/AMP_IN pixel_5015/SF_IB
+ pixel_5015/PIX_OUT pixel_5015/CSA_VREF pixel
Xpixel_5026 pixel_5026/gring pixel_5026/VDD pixel_5026/GND pixel_5026/VREF pixel_5026/ROW_SEL
+ pixel_5026/NB1 pixel_5026/VBIAS pixel_5026/NB2 pixel_5026/AMP_IN pixel_5026/SF_IB
+ pixel_5026/PIX_OUT pixel_5026/CSA_VREF pixel
Xpixel_5037 pixel_5037/gring pixel_5037/VDD pixel_5037/GND pixel_5037/VREF pixel_5037/ROW_SEL
+ pixel_5037/NB1 pixel_5037/VBIAS pixel_5037/NB2 pixel_5037/AMP_IN pixel_5037/SF_IB
+ pixel_5037/PIX_OUT pixel_5037/CSA_VREF pixel
Xpixel_331 pixel_331/gring pixel_331/VDD pixel_331/GND pixel_331/VREF pixel_331/ROW_SEL
+ pixel_331/NB1 pixel_331/VBIAS pixel_331/NB2 pixel_331/AMP_IN pixel_331/SF_IB pixel_331/PIX_OUT
+ pixel_331/CSA_VREF pixel
Xpixel_320 pixel_320/gring pixel_320/VDD pixel_320/GND pixel_320/VREF pixel_320/ROW_SEL
+ pixel_320/NB1 pixel_320/VBIAS pixel_320/NB2 pixel_320/AMP_IN pixel_320/SF_IB pixel_320/PIX_OUT
+ pixel_320/CSA_VREF pixel
Xpixel_5048 pixel_5048/gring pixel_5048/VDD pixel_5048/GND pixel_5048/VREF pixel_5048/ROW_SEL
+ pixel_5048/NB1 pixel_5048/VBIAS pixel_5048/NB2 pixel_5048/AMP_IN pixel_5048/SF_IB
+ pixel_5048/PIX_OUT pixel_5048/CSA_VREF pixel
Xpixel_5059 pixel_5059/gring pixel_5059/VDD pixel_5059/GND pixel_5059/VREF pixel_5059/ROW_SEL
+ pixel_5059/NB1 pixel_5059/VBIAS pixel_5059/NB2 pixel_5059/AMP_IN pixel_5059/SF_IB
+ pixel_5059/PIX_OUT pixel_5059/CSA_VREF pixel
Xpixel_4303 pixel_4303/gring pixel_4303/VDD pixel_4303/GND pixel_4303/VREF pixel_4303/ROW_SEL
+ pixel_4303/NB1 pixel_4303/VBIAS pixel_4303/NB2 pixel_4303/AMP_IN pixel_4303/SF_IB
+ pixel_4303/PIX_OUT pixel_4303/CSA_VREF pixel
Xpixel_4314 pixel_4314/gring pixel_4314/VDD pixel_4314/GND pixel_4314/VREF pixel_4314/ROW_SEL
+ pixel_4314/NB1 pixel_4314/VBIAS pixel_4314/NB2 pixel_4314/AMP_IN pixel_4314/SF_IB
+ pixel_4314/PIX_OUT pixel_4314/CSA_VREF pixel
Xpixel_4325 pixel_4325/gring pixel_4325/VDD pixel_4325/GND pixel_4325/VREF pixel_4325/ROW_SEL
+ pixel_4325/NB1 pixel_4325/VBIAS pixel_4325/NB2 pixel_4325/AMP_IN pixel_4325/SF_IB
+ pixel_4325/PIX_OUT pixel_4325/CSA_VREF pixel
Xpixel_4336 pixel_4336/gring pixel_4336/VDD pixel_4336/GND pixel_4336/VREF pixel_4336/ROW_SEL
+ pixel_4336/NB1 pixel_4336/VBIAS pixel_4336/NB2 pixel_4336/AMP_IN pixel_4336/SF_IB
+ pixel_4336/PIX_OUT pixel_4336/CSA_VREF pixel
Xpixel_364 pixel_364/gring pixel_364/VDD pixel_364/GND pixel_364/VREF pixel_364/ROW_SEL
+ pixel_364/NB1 pixel_364/VBIAS pixel_364/NB2 pixel_364/AMP_IN pixel_364/SF_IB pixel_364/PIX_OUT
+ pixel_364/CSA_VREF pixel
Xpixel_353 pixel_353/gring pixel_353/VDD pixel_353/GND pixel_353/VREF pixel_353/ROW_SEL
+ pixel_353/NB1 pixel_353/VBIAS pixel_353/NB2 pixel_353/AMP_IN pixel_353/SF_IB pixel_353/PIX_OUT
+ pixel_353/CSA_VREF pixel
Xpixel_342 pixel_342/gring pixel_342/VDD pixel_342/GND pixel_342/VREF pixel_342/ROW_SEL
+ pixel_342/NB1 pixel_342/VBIAS pixel_342/NB2 pixel_342/AMP_IN pixel_342/SF_IB pixel_342/PIX_OUT
+ pixel_342/CSA_VREF pixel
Xpixel_3624 pixel_3624/gring pixel_3624/VDD pixel_3624/GND pixel_3624/VREF pixel_3624/ROW_SEL
+ pixel_3624/NB1 pixel_3624/VBIAS pixel_3624/NB2 pixel_3624/AMP_IN pixel_3624/SF_IB
+ pixel_3624/PIX_OUT pixel_3624/CSA_VREF pixel
Xpixel_3613 pixel_3613/gring pixel_3613/VDD pixel_3613/GND pixel_3613/VREF pixel_3613/ROW_SEL
+ pixel_3613/NB1 pixel_3613/VBIAS pixel_3613/NB2 pixel_3613/AMP_IN pixel_3613/SF_IB
+ pixel_3613/PIX_OUT pixel_3613/CSA_VREF pixel
Xpixel_3602 pixel_3602/gring pixel_3602/VDD pixel_3602/GND pixel_3602/VREF pixel_3602/ROW_SEL
+ pixel_3602/NB1 pixel_3602/VBIAS pixel_3602/NB2 pixel_3602/AMP_IN pixel_3602/SF_IB
+ pixel_3602/PIX_OUT pixel_3602/CSA_VREF pixel
Xpixel_4347 pixel_4347/gring pixel_4347/VDD pixel_4347/GND pixel_4347/VREF pixel_4347/ROW_SEL
+ pixel_4347/NB1 pixel_4347/VBIAS pixel_4347/NB2 pixel_4347/AMP_IN pixel_4347/SF_IB
+ pixel_4347/PIX_OUT pixel_4347/CSA_VREF pixel
Xpixel_4358 pixel_4358/gring pixel_4358/VDD pixel_4358/GND pixel_4358/VREF pixel_4358/ROW_SEL
+ pixel_4358/NB1 pixel_4358/VBIAS pixel_4358/NB2 pixel_4358/AMP_IN pixel_4358/SF_IB
+ pixel_4358/PIX_OUT pixel_4358/CSA_VREF pixel
Xpixel_4369 pixel_4369/gring pixel_4369/VDD pixel_4369/GND pixel_4369/VREF pixel_4369/ROW_SEL
+ pixel_4369/NB1 pixel_4369/VBIAS pixel_4369/NB2 pixel_4369/AMP_IN pixel_4369/SF_IB
+ pixel_4369/PIX_OUT pixel_4369/CSA_VREF pixel
Xpixel_397 pixel_397/gring pixel_397/VDD pixel_397/GND pixel_397/VREF pixel_397/ROW_SEL
+ pixel_397/NB1 pixel_397/VBIAS pixel_397/NB2 pixel_397/AMP_IN pixel_397/SF_IB pixel_397/PIX_OUT
+ pixel_397/CSA_VREF pixel
Xpixel_386 pixel_386/gring pixel_386/VDD pixel_386/GND pixel_386/VREF pixel_386/ROW_SEL
+ pixel_386/NB1 pixel_386/VBIAS pixel_386/NB2 pixel_386/AMP_IN pixel_386/SF_IB pixel_386/PIX_OUT
+ pixel_386/CSA_VREF pixel
Xpixel_375 pixel_375/gring pixel_375/VDD pixel_375/GND pixel_375/VREF pixel_375/ROW_SEL
+ pixel_375/NB1 pixel_375/VBIAS pixel_375/NB2 pixel_375/AMP_IN pixel_375/SF_IB pixel_375/PIX_OUT
+ pixel_375/CSA_VREF pixel
Xpixel_2923 pixel_2923/gring pixel_2923/VDD pixel_2923/GND pixel_2923/VREF pixel_2923/ROW_SEL
+ pixel_2923/NB1 pixel_2923/VBIAS pixel_2923/NB2 pixel_2923/AMP_IN pixel_2923/SF_IB
+ pixel_2923/PIX_OUT pixel_2923/CSA_VREF pixel
Xpixel_2912 pixel_2912/gring pixel_2912/VDD pixel_2912/GND pixel_2912/VREF pixel_2912/ROW_SEL
+ pixel_2912/NB1 pixel_2912/VBIAS pixel_2912/NB2 pixel_2912/AMP_IN pixel_2912/SF_IB
+ pixel_2912/PIX_OUT pixel_2912/CSA_VREF pixel
Xpixel_2901 pixel_2901/gring pixel_2901/VDD pixel_2901/GND pixel_2901/VREF pixel_2901/ROW_SEL
+ pixel_2901/NB1 pixel_2901/VBIAS pixel_2901/NB2 pixel_2901/AMP_IN pixel_2901/SF_IB
+ pixel_2901/PIX_OUT pixel_2901/CSA_VREF pixel
Xpixel_3657 pixel_3657/gring pixel_3657/VDD pixel_3657/GND pixel_3657/VREF pixel_3657/ROW_SEL
+ pixel_3657/NB1 pixel_3657/VBIAS pixel_3657/NB2 pixel_3657/AMP_IN pixel_3657/SF_IB
+ pixel_3657/PIX_OUT pixel_3657/CSA_VREF pixel
Xpixel_3646 pixel_3646/gring pixel_3646/VDD pixel_3646/GND pixel_3646/VREF pixel_3646/ROW_SEL
+ pixel_3646/NB1 pixel_3646/VBIAS pixel_3646/NB2 pixel_3646/AMP_IN pixel_3646/SF_IB
+ pixel_3646/PIX_OUT pixel_3646/CSA_VREF pixel
Xpixel_3635 pixel_3635/gring pixel_3635/VDD pixel_3635/GND pixel_3635/VREF pixel_3635/ROW_SEL
+ pixel_3635/NB1 pixel_3635/VBIAS pixel_3635/NB2 pixel_3635/AMP_IN pixel_3635/SF_IB
+ pixel_3635/PIX_OUT pixel_3635/CSA_VREF pixel
Xpixel_2956 pixel_2956/gring pixel_2956/VDD pixel_2956/GND pixel_2956/VREF pixel_2956/ROW_SEL
+ pixel_2956/NB1 pixel_2956/VBIAS pixel_2956/NB2 pixel_2956/AMP_IN pixel_2956/SF_IB
+ pixel_2956/PIX_OUT pixel_2956/CSA_VREF pixel
Xpixel_2945 pixel_2945/gring pixel_2945/VDD pixel_2945/GND pixel_2945/VREF pixel_2945/ROW_SEL
+ pixel_2945/NB1 pixel_2945/VBIAS pixel_2945/NB2 pixel_2945/AMP_IN pixel_2945/SF_IB
+ pixel_2945/PIX_OUT pixel_2945/CSA_VREF pixel
Xpixel_2934 pixel_2934/gring pixel_2934/VDD pixel_2934/GND pixel_2934/VREF pixel_2934/ROW_SEL
+ pixel_2934/NB1 pixel_2934/VBIAS pixel_2934/NB2 pixel_2934/AMP_IN pixel_2934/SF_IB
+ pixel_2934/PIX_OUT pixel_2934/CSA_VREF pixel
Xpixel_3679 pixel_3679/gring pixel_3679/VDD pixel_3679/GND pixel_3679/VREF pixel_3679/ROW_SEL
+ pixel_3679/NB1 pixel_3679/VBIAS pixel_3679/NB2 pixel_3679/AMP_IN pixel_3679/SF_IB
+ pixel_3679/PIX_OUT pixel_3679/CSA_VREF pixel
Xpixel_3668 pixel_3668/gring pixel_3668/VDD pixel_3668/GND pixel_3668/VREF pixel_3668/ROW_SEL
+ pixel_3668/NB1 pixel_3668/VBIAS pixel_3668/NB2 pixel_3668/AMP_IN pixel_3668/SF_IB
+ pixel_3668/PIX_OUT pixel_3668/CSA_VREF pixel
Xpixel_2989 pixel_2989/gring pixel_2989/VDD pixel_2989/GND pixel_2989/VREF pixel_2989/ROW_SEL
+ pixel_2989/NB1 pixel_2989/VBIAS pixel_2989/NB2 pixel_2989/AMP_IN pixel_2989/SF_IB
+ pixel_2989/PIX_OUT pixel_2989/CSA_VREF pixel
Xpixel_2978 pixel_2978/gring pixel_2978/VDD pixel_2978/GND pixel_2978/VREF pixel_2978/ROW_SEL
+ pixel_2978/NB1 pixel_2978/VBIAS pixel_2978/NB2 pixel_2978/AMP_IN pixel_2978/SF_IB
+ pixel_2978/PIX_OUT pixel_2978/CSA_VREF pixel
Xpixel_2967 pixel_2967/gring pixel_2967/VDD pixel_2967/GND pixel_2967/VREF pixel_2967/ROW_SEL
+ pixel_2967/NB1 pixel_2967/VBIAS pixel_2967/NB2 pixel_2967/AMP_IN pixel_2967/SF_IB
+ pixel_2967/PIX_OUT pixel_2967/CSA_VREF pixel
Xpixel_6250 pixel_6250/gring pixel_6250/VDD pixel_6250/GND pixel_6250/VREF pixel_6250/ROW_SEL
+ pixel_6250/NB1 pixel_6250/VBIAS pixel_6250/NB2 pixel_6250/AMP_IN pixel_6250/SF_IB
+ pixel_6250/PIX_OUT pixel_6250/CSA_VREF pixel
Xpixel_6261 pixel_6261/gring pixel_6261/VDD pixel_6261/GND pixel_6261/VREF pixel_6261/ROW_SEL
+ pixel_6261/NB1 pixel_6261/VBIAS pixel_6261/NB2 pixel_6261/AMP_IN pixel_6261/SF_IB
+ pixel_6261/PIX_OUT pixel_6261/CSA_VREF pixel
Xpixel_6272 pixel_6272/gring pixel_6272/VDD pixel_6272/GND pixel_6272/VREF pixel_6272/ROW_SEL
+ pixel_6272/NB1 pixel_6272/VBIAS pixel_6272/NB2 pixel_6272/AMP_IN pixel_6272/SF_IB
+ pixel_6272/PIX_OUT pixel_6272/CSA_VREF pixel
Xpixel_6283 pixel_6283/gring pixel_6283/VDD pixel_6283/GND pixel_6283/VREF pixel_6283/ROW_SEL
+ pixel_6283/NB1 pixel_6283/VBIAS pixel_6283/NB2 pixel_6283/AMP_IN pixel_6283/SF_IB
+ pixel_6283/PIX_OUT pixel_6283/CSA_VREF pixel
Xpixel_6294 pixel_6294/gring pixel_6294/VDD pixel_6294/GND pixel_6294/VREF pixel_6294/ROW_SEL
+ pixel_6294/NB1 pixel_6294/VBIAS pixel_6294/NB2 pixel_6294/AMP_IN pixel_6294/SF_IB
+ pixel_6294/PIX_OUT pixel_6294/CSA_VREF pixel
Xpixel_5560 pixel_5560/gring pixel_5560/VDD pixel_5560/GND pixel_5560/VREF pixel_5560/ROW_SEL
+ pixel_5560/NB1 pixel_5560/VBIAS pixel_5560/NB2 pixel_5560/AMP_IN pixel_5560/SF_IB
+ pixel_5560/PIX_OUT pixel_5560/CSA_VREF pixel
Xpixel_5571 pixel_5571/gring pixel_5571/VDD pixel_5571/GND pixel_5571/VREF pixel_5571/ROW_SEL
+ pixel_5571/NB1 pixel_5571/VBIAS pixel_5571/NB2 pixel_5571/AMP_IN pixel_5571/SF_IB
+ pixel_5571/PIX_OUT pixel_5571/CSA_VREF pixel
Xpixel_5582 pixel_5582/gring pixel_5582/VDD pixel_5582/GND pixel_5582/VREF pixel_5582/ROW_SEL
+ pixel_5582/NB1 pixel_5582/VBIAS pixel_5582/NB2 pixel_5582/AMP_IN pixel_5582/SF_IB
+ pixel_5582/PIX_OUT pixel_5582/CSA_VREF pixel
Xpixel_5593 pixel_5593/gring pixel_5593/VDD pixel_5593/GND pixel_5593/VREF pixel_5593/ROW_SEL
+ pixel_5593/NB1 pixel_5593/VBIAS pixel_5593/NB2 pixel_5593/AMP_IN pixel_5593/SF_IB
+ pixel_5593/PIX_OUT pixel_5593/CSA_VREF pixel
Xpixel_4870 pixel_4870/gring pixel_4870/VDD pixel_4870/GND pixel_4870/VREF pixel_4870/ROW_SEL
+ pixel_4870/NB1 pixel_4870/VBIAS pixel_4870/NB2 pixel_4870/AMP_IN pixel_4870/SF_IB
+ pixel_4870/PIX_OUT pixel_4870/CSA_VREF pixel
Xpixel_4881 pixel_4881/gring pixel_4881/VDD pixel_4881/GND pixel_4881/VREF pixel_4881/ROW_SEL
+ pixel_4881/NB1 pixel_4881/VBIAS pixel_4881/NB2 pixel_4881/AMP_IN pixel_4881/SF_IB
+ pixel_4881/PIX_OUT pixel_4881/CSA_VREF pixel
Xpixel_4892 pixel_4892/gring pixel_4892/VDD pixel_4892/GND pixel_4892/VREF pixel_4892/ROW_SEL
+ pixel_4892/NB1 pixel_4892/VBIAS pixel_4892/NB2 pixel_4892/AMP_IN pixel_4892/SF_IB
+ pixel_4892/PIX_OUT pixel_4892/CSA_VREF pixel
Xpixel_2208 pixel_2208/gring pixel_2208/VDD pixel_2208/GND pixel_2208/VREF pixel_2208/ROW_SEL
+ pixel_2208/NB1 pixel_2208/VBIAS pixel_2208/NB2 pixel_2208/AMP_IN pixel_2208/SF_IB
+ pixel_2208/PIX_OUT pixel_2208/CSA_VREF pixel
Xpixel_1507 pixel_1507/gring pixel_1507/VDD pixel_1507/GND pixel_1507/VREF pixel_1507/ROW_SEL
+ pixel_1507/NB1 pixel_1507/VBIAS pixel_1507/NB2 pixel_1507/AMP_IN pixel_1507/SF_IB
+ pixel_1507/PIX_OUT pixel_1507/CSA_VREF pixel
Xpixel_2219 pixel_2219/gring pixel_2219/VDD pixel_2219/GND pixel_2219/VREF pixel_2219/ROW_SEL
+ pixel_2219/NB1 pixel_2219/VBIAS pixel_2219/NB2 pixel_2219/AMP_IN pixel_2219/SF_IB
+ pixel_2219/PIX_OUT pixel_2219/CSA_VREF pixel
Xpixel_1529 pixel_1529/gring pixel_1529/VDD pixel_1529/GND pixel_1529/VREF pixel_1529/ROW_SEL
+ pixel_1529/NB1 pixel_1529/VBIAS pixel_1529/NB2 pixel_1529/AMP_IN pixel_1529/SF_IB
+ pixel_1529/PIX_OUT pixel_1529/CSA_VREF pixel
Xpixel_1518 pixel_1518/gring pixel_1518/VDD pixel_1518/GND pixel_1518/VREF pixel_1518/ROW_SEL
+ pixel_1518/NB1 pixel_1518/VBIAS pixel_1518/NB2 pixel_1518/AMP_IN pixel_1518/SF_IB
+ pixel_1518/PIX_OUT pixel_1518/CSA_VREF pixel
Xpixel_9815 pixel_9815/gring pixel_9815/VDD pixel_9815/GND pixel_9815/VREF pixel_9815/ROW_SEL
+ pixel_9815/NB1 pixel_9815/VBIAS pixel_9815/NB2 pixel_9815/AMP_IN pixel_9815/SF_IB
+ pixel_9815/PIX_OUT pixel_9815/CSA_VREF pixel
Xpixel_9804 pixel_9804/gring pixel_9804/VDD pixel_9804/GND pixel_9804/VREF pixel_9804/ROW_SEL
+ pixel_9804/NB1 pixel_9804/VBIAS pixel_9804/NB2 pixel_9804/AMP_IN pixel_9804/SF_IB
+ pixel_9804/PIX_OUT pixel_9804/CSA_VREF pixel
Xpixel_9837 pixel_9837/gring pixel_9837/VDD pixel_9837/GND pixel_9837/VREF pixel_9837/ROW_SEL
+ pixel_9837/NB1 pixel_9837/VBIAS pixel_9837/NB2 pixel_9837/AMP_IN pixel_9837/SF_IB
+ pixel_9837/PIX_OUT pixel_9837/CSA_VREF pixel
Xpixel_9826 pixel_9826/gring pixel_9826/VDD pixel_9826/GND pixel_9826/VREF pixel_9826/ROW_SEL
+ pixel_9826/NB1 pixel_9826/VBIAS pixel_9826/NB2 pixel_9826/AMP_IN pixel_9826/SF_IB
+ pixel_9826/PIX_OUT pixel_9826/CSA_VREF pixel
Xpixel_9848 pixel_9848/gring pixel_9848/VDD pixel_9848/GND pixel_9848/VREF pixel_9848/ROW_SEL
+ pixel_9848/NB1 pixel_9848/VBIAS pixel_9848/NB2 pixel_9848/AMP_IN pixel_9848/SF_IB
+ pixel_9848/PIX_OUT pixel_9848/CSA_VREF pixel
Xpixel_9859 pixel_9859/gring pixel_9859/VDD pixel_9859/GND pixel_9859/VREF pixel_9859/ROW_SEL
+ pixel_9859/NB1 pixel_9859/VBIAS pixel_9859/NB2 pixel_9859/AMP_IN pixel_9859/SF_IB
+ pixel_9859/PIX_OUT pixel_9859/CSA_VREF pixel
Xpixel_4100 pixel_4100/gring pixel_4100/VDD pixel_4100/GND pixel_4100/VREF pixel_4100/ROW_SEL
+ pixel_4100/NB1 pixel_4100/VBIAS pixel_4100/NB2 pixel_4100/AMP_IN pixel_4100/SF_IB
+ pixel_4100/PIX_OUT pixel_4100/CSA_VREF pixel
Xpixel_4111 pixel_4111/gring pixel_4111/VDD pixel_4111/GND pixel_4111/VREF pixel_4111/ROW_SEL
+ pixel_4111/NB1 pixel_4111/VBIAS pixel_4111/NB2 pixel_4111/AMP_IN pixel_4111/SF_IB
+ pixel_4111/PIX_OUT pixel_4111/CSA_VREF pixel
Xpixel_4122 pixel_4122/gring pixel_4122/VDD pixel_4122/GND pixel_4122/VREF pixel_4122/ROW_SEL
+ pixel_4122/NB1 pixel_4122/VBIAS pixel_4122/NB2 pixel_4122/AMP_IN pixel_4122/SF_IB
+ pixel_4122/PIX_OUT pixel_4122/CSA_VREF pixel
Xpixel_4133 pixel_4133/gring pixel_4133/VDD pixel_4133/GND pixel_4133/VREF pixel_4133/ROW_SEL
+ pixel_4133/NB1 pixel_4133/VBIAS pixel_4133/NB2 pixel_4133/AMP_IN pixel_4133/SF_IB
+ pixel_4133/PIX_OUT pixel_4133/CSA_VREF pixel
Xpixel_4144 pixel_4144/gring pixel_4144/VDD pixel_4144/GND pixel_4144/VREF pixel_4144/ROW_SEL
+ pixel_4144/NB1 pixel_4144/VBIAS pixel_4144/NB2 pixel_4144/AMP_IN pixel_4144/SF_IB
+ pixel_4144/PIX_OUT pixel_4144/CSA_VREF pixel
Xpixel_172 pixel_172/gring pixel_172/VDD pixel_172/GND pixel_172/VREF pixel_172/ROW_SEL
+ pixel_172/NB1 pixel_172/VBIAS pixel_172/NB2 pixel_172/AMP_IN pixel_172/SF_IB pixel_172/PIX_OUT
+ pixel_172/CSA_VREF pixel
Xpixel_161 pixel_161/gring pixel_161/VDD pixel_161/GND pixel_161/VREF pixel_161/ROW_SEL
+ pixel_161/NB1 pixel_161/VBIAS pixel_161/NB2 pixel_161/AMP_IN pixel_161/SF_IB pixel_161/PIX_OUT
+ pixel_161/CSA_VREF pixel
Xpixel_150 pixel_150/gring pixel_150/VDD pixel_150/GND pixel_150/VREF pixel_150/ROW_SEL
+ pixel_150/NB1 pixel_150/VBIAS pixel_150/NB2 pixel_150/AMP_IN pixel_150/SF_IB pixel_150/PIX_OUT
+ pixel_150/CSA_VREF pixel
Xpixel_3432 pixel_3432/gring pixel_3432/VDD pixel_3432/GND pixel_3432/VREF pixel_3432/ROW_SEL
+ pixel_3432/NB1 pixel_3432/VBIAS pixel_3432/NB2 pixel_3432/AMP_IN pixel_3432/SF_IB
+ pixel_3432/PIX_OUT pixel_3432/CSA_VREF pixel
Xpixel_3421 pixel_3421/gring pixel_3421/VDD pixel_3421/GND pixel_3421/VREF pixel_3421/ROW_SEL
+ pixel_3421/NB1 pixel_3421/VBIAS pixel_3421/NB2 pixel_3421/AMP_IN pixel_3421/SF_IB
+ pixel_3421/PIX_OUT pixel_3421/CSA_VREF pixel
Xpixel_3410 pixel_3410/gring pixel_3410/VDD pixel_3410/GND pixel_3410/VREF pixel_3410/ROW_SEL
+ pixel_3410/NB1 pixel_3410/VBIAS pixel_3410/NB2 pixel_3410/AMP_IN pixel_3410/SF_IB
+ pixel_3410/PIX_OUT pixel_3410/CSA_VREF pixel
Xpixel_4155 pixel_4155/gring pixel_4155/VDD pixel_4155/GND pixel_4155/VREF pixel_4155/ROW_SEL
+ pixel_4155/NB1 pixel_4155/VBIAS pixel_4155/NB2 pixel_4155/AMP_IN pixel_4155/SF_IB
+ pixel_4155/PIX_OUT pixel_4155/CSA_VREF pixel
Xpixel_4166 pixel_4166/gring pixel_4166/VDD pixel_4166/GND pixel_4166/VREF pixel_4166/ROW_SEL
+ pixel_4166/NB1 pixel_4166/VBIAS pixel_4166/NB2 pixel_4166/AMP_IN pixel_4166/SF_IB
+ pixel_4166/PIX_OUT pixel_4166/CSA_VREF pixel
Xpixel_4177 pixel_4177/gring pixel_4177/VDD pixel_4177/GND pixel_4177/VREF pixel_4177/ROW_SEL
+ pixel_4177/NB1 pixel_4177/VBIAS pixel_4177/NB2 pixel_4177/AMP_IN pixel_4177/SF_IB
+ pixel_4177/PIX_OUT pixel_4177/CSA_VREF pixel
Xpixel_194 pixel_194/gring pixel_194/VDD pixel_194/GND pixel_194/VREF pixel_194/ROW_SEL
+ pixel_194/NB1 pixel_194/VBIAS pixel_194/NB2 pixel_194/AMP_IN pixel_194/SF_IB pixel_194/PIX_OUT
+ pixel_194/CSA_VREF pixel
Xpixel_183 pixel_183/gring pixel_183/VDD pixel_183/GND pixel_183/VREF pixel_183/ROW_SEL
+ pixel_183/NB1 pixel_183/VBIAS pixel_183/NB2 pixel_183/AMP_IN pixel_183/SF_IB pixel_183/PIX_OUT
+ pixel_183/CSA_VREF pixel
Xpixel_2731 pixel_2731/gring pixel_2731/VDD pixel_2731/GND pixel_2731/VREF pixel_2731/ROW_SEL
+ pixel_2731/NB1 pixel_2731/VBIAS pixel_2731/NB2 pixel_2731/AMP_IN pixel_2731/SF_IB
+ pixel_2731/PIX_OUT pixel_2731/CSA_VREF pixel
Xpixel_2720 pixel_2720/gring pixel_2720/VDD pixel_2720/GND pixel_2720/VREF pixel_2720/ROW_SEL
+ pixel_2720/NB1 pixel_2720/VBIAS pixel_2720/NB2 pixel_2720/AMP_IN pixel_2720/SF_IB
+ pixel_2720/PIX_OUT pixel_2720/CSA_VREF pixel
Xpixel_3476 pixel_3476/gring pixel_3476/VDD pixel_3476/GND pixel_3476/VREF pixel_3476/ROW_SEL
+ pixel_3476/NB1 pixel_3476/VBIAS pixel_3476/NB2 pixel_3476/AMP_IN pixel_3476/SF_IB
+ pixel_3476/PIX_OUT pixel_3476/CSA_VREF pixel
Xpixel_3465 pixel_3465/gring pixel_3465/VDD pixel_3465/GND pixel_3465/VREF pixel_3465/ROW_SEL
+ pixel_3465/NB1 pixel_3465/VBIAS pixel_3465/NB2 pixel_3465/AMP_IN pixel_3465/SF_IB
+ pixel_3465/PIX_OUT pixel_3465/CSA_VREF pixel
Xpixel_3454 pixel_3454/gring pixel_3454/VDD pixel_3454/GND pixel_3454/VREF pixel_3454/ROW_SEL
+ pixel_3454/NB1 pixel_3454/VBIAS pixel_3454/NB2 pixel_3454/AMP_IN pixel_3454/SF_IB
+ pixel_3454/PIX_OUT pixel_3454/CSA_VREF pixel
Xpixel_3443 pixel_3443/gring pixel_3443/VDD pixel_3443/GND pixel_3443/VREF pixel_3443/ROW_SEL
+ pixel_3443/NB1 pixel_3443/VBIAS pixel_3443/NB2 pixel_3443/AMP_IN pixel_3443/SF_IB
+ pixel_3443/PIX_OUT pixel_3443/CSA_VREF pixel
Xpixel_4188 pixel_4188/gring pixel_4188/VDD pixel_4188/GND pixel_4188/VREF pixel_4188/ROW_SEL
+ pixel_4188/NB1 pixel_4188/VBIAS pixel_4188/NB2 pixel_4188/AMP_IN pixel_4188/SF_IB
+ pixel_4188/PIX_OUT pixel_4188/CSA_VREF pixel
Xpixel_4199 pixel_4199/gring pixel_4199/VDD pixel_4199/GND pixel_4199/VREF pixel_4199/ROW_SEL
+ pixel_4199/NB1 pixel_4199/VBIAS pixel_4199/NB2 pixel_4199/AMP_IN pixel_4199/SF_IB
+ pixel_4199/PIX_OUT pixel_4199/CSA_VREF pixel
Xpixel_2764 pixel_2764/gring pixel_2764/VDD pixel_2764/GND pixel_2764/VREF pixel_2764/ROW_SEL
+ pixel_2764/NB1 pixel_2764/VBIAS pixel_2764/NB2 pixel_2764/AMP_IN pixel_2764/SF_IB
+ pixel_2764/PIX_OUT pixel_2764/CSA_VREF pixel
Xpixel_2753 pixel_2753/gring pixel_2753/VDD pixel_2753/GND pixel_2753/VREF pixel_2753/ROW_SEL
+ pixel_2753/NB1 pixel_2753/VBIAS pixel_2753/NB2 pixel_2753/AMP_IN pixel_2753/SF_IB
+ pixel_2753/PIX_OUT pixel_2753/CSA_VREF pixel
Xpixel_2742 pixel_2742/gring pixel_2742/VDD pixel_2742/GND pixel_2742/VREF pixel_2742/ROW_SEL
+ pixel_2742/NB1 pixel_2742/VBIAS pixel_2742/NB2 pixel_2742/AMP_IN pixel_2742/SF_IB
+ pixel_2742/PIX_OUT pixel_2742/CSA_VREF pixel
Xpixel_3498 pixel_3498/gring pixel_3498/VDD pixel_3498/GND pixel_3498/VREF pixel_3498/ROW_SEL
+ pixel_3498/NB1 pixel_3498/VBIAS pixel_3498/NB2 pixel_3498/AMP_IN pixel_3498/SF_IB
+ pixel_3498/PIX_OUT pixel_3498/CSA_VREF pixel
Xpixel_3487 pixel_3487/gring pixel_3487/VDD pixel_3487/GND pixel_3487/VREF pixel_3487/ROW_SEL
+ pixel_3487/NB1 pixel_3487/VBIAS pixel_3487/NB2 pixel_3487/AMP_IN pixel_3487/SF_IB
+ pixel_3487/PIX_OUT pixel_3487/CSA_VREF pixel
Xpixel_2797 pixel_2797/gring pixel_2797/VDD pixel_2797/GND pixel_2797/VREF pixel_2797/ROW_SEL
+ pixel_2797/NB1 pixel_2797/VBIAS pixel_2797/NB2 pixel_2797/AMP_IN pixel_2797/SF_IB
+ pixel_2797/PIX_OUT pixel_2797/CSA_VREF pixel
Xpixel_2786 pixel_2786/gring pixel_2786/VDD pixel_2786/GND pixel_2786/VREF pixel_2786/ROW_SEL
+ pixel_2786/NB1 pixel_2786/VBIAS pixel_2786/NB2 pixel_2786/AMP_IN pixel_2786/SF_IB
+ pixel_2786/PIX_OUT pixel_2786/CSA_VREF pixel
Xpixel_2775 pixel_2775/gring pixel_2775/VDD pixel_2775/GND pixel_2775/VREF pixel_2775/ROW_SEL
+ pixel_2775/NB1 pixel_2775/VBIAS pixel_2775/NB2 pixel_2775/AMP_IN pixel_2775/SF_IB
+ pixel_2775/PIX_OUT pixel_2775/CSA_VREF pixel
Xpixel_6080 pixel_6080/gring pixel_6080/VDD pixel_6080/GND pixel_6080/VREF pixel_6080/ROW_SEL
+ pixel_6080/NB1 pixel_6080/VBIAS pixel_6080/NB2 pixel_6080/AMP_IN pixel_6080/SF_IB
+ pixel_6080/PIX_OUT pixel_6080/CSA_VREF pixel
Xpixel_6091 pixel_6091/gring pixel_6091/VDD pixel_6091/GND pixel_6091/VREF pixel_6091/ROW_SEL
+ pixel_6091/NB1 pixel_6091/VBIAS pixel_6091/NB2 pixel_6091/AMP_IN pixel_6091/SF_IB
+ pixel_6091/PIX_OUT pixel_6091/CSA_VREF pixel
Xpixel_5390 pixel_5390/gring pixel_5390/VDD pixel_5390/GND pixel_5390/VREF pixel_5390/ROW_SEL
+ pixel_5390/NB1 pixel_5390/VBIAS pixel_5390/NB2 pixel_5390/AMP_IN pixel_5390/SF_IB
+ pixel_5390/PIX_OUT pixel_5390/CSA_VREF pixel
Xpixel_7709 pixel_7709/gring pixel_7709/VDD pixel_7709/GND pixel_7709/VREF pixel_7709/ROW_SEL
+ pixel_7709/NB1 pixel_7709/VBIAS pixel_7709/NB2 pixel_7709/AMP_IN pixel_7709/SF_IB
+ pixel_7709/PIX_OUT pixel_7709/CSA_VREF pixel
Xpixel_2027 pixel_2027/gring pixel_2027/VDD pixel_2027/GND pixel_2027/VREF pixel_2027/ROW_SEL
+ pixel_2027/NB1 pixel_2027/VBIAS pixel_2027/NB2 pixel_2027/AMP_IN pixel_2027/SF_IB
+ pixel_2027/PIX_OUT pixel_2027/CSA_VREF pixel
Xpixel_2016 pixel_2016/gring pixel_2016/VDD pixel_2016/GND pixel_2016/VREF pixel_2016/ROW_SEL
+ pixel_2016/NB1 pixel_2016/VBIAS pixel_2016/NB2 pixel_2016/AMP_IN pixel_2016/SF_IB
+ pixel_2016/PIX_OUT pixel_2016/CSA_VREF pixel
Xpixel_2005 pixel_2005/gring pixel_2005/VDD pixel_2005/GND pixel_2005/VREF pixel_2005/ROW_SEL
+ pixel_2005/NB1 pixel_2005/VBIAS pixel_2005/NB2 pixel_2005/AMP_IN pixel_2005/SF_IB
+ pixel_2005/PIX_OUT pixel_2005/CSA_VREF pixel
Xpixel_1315 pixel_1315/gring pixel_1315/VDD pixel_1315/GND pixel_1315/VREF pixel_1315/ROW_SEL
+ pixel_1315/NB1 pixel_1315/VBIAS pixel_1315/NB2 pixel_1315/AMP_IN pixel_1315/SF_IB
+ pixel_1315/PIX_OUT pixel_1315/CSA_VREF pixel
Xpixel_1304 pixel_1304/gring pixel_1304/VDD pixel_1304/GND pixel_1304/VREF pixel_1304/ROW_SEL
+ pixel_1304/NB1 pixel_1304/VBIAS pixel_1304/NB2 pixel_1304/AMP_IN pixel_1304/SF_IB
+ pixel_1304/PIX_OUT pixel_1304/CSA_VREF pixel
Xpixel_2049 pixel_2049/gring pixel_2049/VDD pixel_2049/GND pixel_2049/VREF pixel_2049/ROW_SEL
+ pixel_2049/NB1 pixel_2049/VBIAS pixel_2049/NB2 pixel_2049/AMP_IN pixel_2049/SF_IB
+ pixel_2049/PIX_OUT pixel_2049/CSA_VREF pixel
Xpixel_2038 pixel_2038/gring pixel_2038/VDD pixel_2038/GND pixel_2038/VREF pixel_2038/ROW_SEL
+ pixel_2038/NB1 pixel_2038/VBIAS pixel_2038/NB2 pixel_2038/AMP_IN pixel_2038/SF_IB
+ pixel_2038/PIX_OUT pixel_2038/CSA_VREF pixel
Xpixel_1348 pixel_1348/gring pixel_1348/VDD pixel_1348/GND pixel_1348/VREF pixel_1348/ROW_SEL
+ pixel_1348/NB1 pixel_1348/VBIAS pixel_1348/NB2 pixel_1348/AMP_IN pixel_1348/SF_IB
+ pixel_1348/PIX_OUT pixel_1348/CSA_VREF pixel
Xpixel_1337 pixel_1337/gring pixel_1337/VDD pixel_1337/GND pixel_1337/VREF pixel_1337/ROW_SEL
+ pixel_1337/NB1 pixel_1337/VBIAS pixel_1337/NB2 pixel_1337/AMP_IN pixel_1337/SF_IB
+ pixel_1337/PIX_OUT pixel_1337/CSA_VREF pixel
Xpixel_1326 pixel_1326/gring pixel_1326/VDD pixel_1326/GND pixel_1326/VREF pixel_1326/ROW_SEL
+ pixel_1326/NB1 pixel_1326/VBIAS pixel_1326/NB2 pixel_1326/AMP_IN pixel_1326/SF_IB
+ pixel_1326/PIX_OUT pixel_1326/CSA_VREF pixel
Xpixel_1359 pixel_1359/gring pixel_1359/VDD pixel_1359/GND pixel_1359/VREF pixel_1359/ROW_SEL
+ pixel_1359/NB1 pixel_1359/VBIAS pixel_1359/NB2 pixel_1359/AMP_IN pixel_1359/SF_IB
+ pixel_1359/PIX_OUT pixel_1359/CSA_VREF pixel
Xpixel_9601 pixel_9601/gring pixel_9601/VDD pixel_9601/GND pixel_9601/VREF pixel_9601/ROW_SEL
+ pixel_9601/NB1 pixel_9601/VBIAS pixel_9601/NB2 pixel_9601/AMP_IN pixel_9601/SF_IB
+ pixel_9601/PIX_OUT pixel_9601/CSA_VREF pixel
Xpixel_9612 pixel_9612/gring pixel_9612/VDD pixel_9612/GND pixel_9612/VREF pixel_9612/ROW_SEL
+ pixel_9612/NB1 pixel_9612/VBIAS pixel_9612/NB2 pixel_9612/AMP_IN pixel_9612/SF_IB
+ pixel_9612/PIX_OUT pixel_9612/CSA_VREF pixel
Xpixel_9623 pixel_9623/gring pixel_9623/VDD pixel_9623/GND pixel_9623/VREF pixel_9623/ROW_SEL
+ pixel_9623/NB1 pixel_9623/VBIAS pixel_9623/NB2 pixel_9623/AMP_IN pixel_9623/SF_IB
+ pixel_9623/PIX_OUT pixel_9623/CSA_VREF pixel
Xpixel_8911 pixel_8911/gring pixel_8911/VDD pixel_8911/GND pixel_8911/VREF pixel_8911/ROW_SEL
+ pixel_8911/NB1 pixel_8911/VBIAS pixel_8911/NB2 pixel_8911/AMP_IN pixel_8911/SF_IB
+ pixel_8911/PIX_OUT pixel_8911/CSA_VREF pixel
Xpixel_8900 pixel_8900/gring pixel_8900/VDD pixel_8900/GND pixel_8900/VREF pixel_8900/ROW_SEL
+ pixel_8900/NB1 pixel_8900/VBIAS pixel_8900/NB2 pixel_8900/AMP_IN pixel_8900/SF_IB
+ pixel_8900/PIX_OUT pixel_8900/CSA_VREF pixel
Xpixel_9634 pixel_9634/gring pixel_9634/VDD pixel_9634/GND pixel_9634/VREF pixel_9634/ROW_SEL
+ pixel_9634/NB1 pixel_9634/VBIAS pixel_9634/NB2 pixel_9634/AMP_IN pixel_9634/SF_IB
+ pixel_9634/PIX_OUT pixel_9634/CSA_VREF pixel
Xpixel_9645 pixel_9645/gring pixel_9645/VDD pixel_9645/GND pixel_9645/VREF pixel_9645/ROW_SEL
+ pixel_9645/NB1 pixel_9645/VBIAS pixel_9645/NB2 pixel_9645/AMP_IN pixel_9645/SF_IB
+ pixel_9645/PIX_OUT pixel_9645/CSA_VREF pixel
Xpixel_9656 pixel_9656/gring pixel_9656/VDD pixel_9656/GND pixel_9656/VREF pixel_9656/ROW_SEL
+ pixel_9656/NB1 pixel_9656/VBIAS pixel_9656/NB2 pixel_9656/AMP_IN pixel_9656/SF_IB
+ pixel_9656/PIX_OUT pixel_9656/CSA_VREF pixel
Xpixel_8955 pixel_8955/gring pixel_8955/VDD pixel_8955/GND pixel_8955/VREF pixel_8955/ROW_SEL
+ pixel_8955/NB1 pixel_8955/VBIAS pixel_8955/NB2 pixel_8955/AMP_IN pixel_8955/SF_IB
+ pixel_8955/PIX_OUT pixel_8955/CSA_VREF pixel
Xpixel_8944 pixel_8944/gring pixel_8944/VDD pixel_8944/GND pixel_8944/VREF pixel_8944/ROW_SEL
+ pixel_8944/NB1 pixel_8944/VBIAS pixel_8944/NB2 pixel_8944/AMP_IN pixel_8944/SF_IB
+ pixel_8944/PIX_OUT pixel_8944/CSA_VREF pixel
Xpixel_8933 pixel_8933/gring pixel_8933/VDD pixel_8933/GND pixel_8933/VREF pixel_8933/ROW_SEL
+ pixel_8933/NB1 pixel_8933/VBIAS pixel_8933/NB2 pixel_8933/AMP_IN pixel_8933/SF_IB
+ pixel_8933/PIX_OUT pixel_8933/CSA_VREF pixel
Xpixel_8922 pixel_8922/gring pixel_8922/VDD pixel_8922/GND pixel_8922/VREF pixel_8922/ROW_SEL
+ pixel_8922/NB1 pixel_8922/VBIAS pixel_8922/NB2 pixel_8922/AMP_IN pixel_8922/SF_IB
+ pixel_8922/PIX_OUT pixel_8922/CSA_VREF pixel
Xpixel_9689 pixel_9689/gring pixel_9689/VDD pixel_9689/GND pixel_9689/VREF pixel_9689/ROW_SEL
+ pixel_9689/NB1 pixel_9689/VBIAS pixel_9689/NB2 pixel_9689/AMP_IN pixel_9689/SF_IB
+ pixel_9689/PIX_OUT pixel_9689/CSA_VREF pixel
Xpixel_9667 pixel_9667/gring pixel_9667/VDD pixel_9667/GND pixel_9667/VREF pixel_9667/ROW_SEL
+ pixel_9667/NB1 pixel_9667/VBIAS pixel_9667/NB2 pixel_9667/AMP_IN pixel_9667/SF_IB
+ pixel_9667/PIX_OUT pixel_9667/CSA_VREF pixel
Xpixel_9678 pixel_9678/gring pixel_9678/VDD pixel_9678/GND pixel_9678/VREF pixel_9678/ROW_SEL
+ pixel_9678/NB1 pixel_9678/VBIAS pixel_9678/NB2 pixel_9678/AMP_IN pixel_9678/SF_IB
+ pixel_9678/PIX_OUT pixel_9678/CSA_VREF pixel
Xpixel_8988 pixel_8988/gring pixel_8988/VDD pixel_8988/GND pixel_8988/VREF pixel_8988/ROW_SEL
+ pixel_8988/NB1 pixel_8988/VBIAS pixel_8988/NB2 pixel_8988/AMP_IN pixel_8988/SF_IB
+ pixel_8988/PIX_OUT pixel_8988/CSA_VREF pixel
Xpixel_8977 pixel_8977/gring pixel_8977/VDD pixel_8977/GND pixel_8977/VREF pixel_8977/ROW_SEL
+ pixel_8977/NB1 pixel_8977/VBIAS pixel_8977/NB2 pixel_8977/AMP_IN pixel_8977/SF_IB
+ pixel_8977/PIX_OUT pixel_8977/CSA_VREF pixel
Xpixel_8966 pixel_8966/gring pixel_8966/VDD pixel_8966/GND pixel_8966/VREF pixel_8966/ROW_SEL
+ pixel_8966/NB1 pixel_8966/VBIAS pixel_8966/NB2 pixel_8966/AMP_IN pixel_8966/SF_IB
+ pixel_8966/PIX_OUT pixel_8966/CSA_VREF pixel
Xpixel_8999 pixel_8999/gring pixel_8999/VDD pixel_8999/GND pixel_8999/VREF pixel_8999/ROW_SEL
+ pixel_8999/NB1 pixel_8999/VBIAS pixel_8999/NB2 pixel_8999/AMP_IN pixel_8999/SF_IB
+ pixel_8999/PIX_OUT pixel_8999/CSA_VREF pixel
Xpixel_3251 pixel_3251/gring pixel_3251/VDD pixel_3251/GND pixel_3251/VREF pixel_3251/ROW_SEL
+ pixel_3251/NB1 pixel_3251/VBIAS pixel_3251/NB2 pixel_3251/AMP_IN pixel_3251/SF_IB
+ pixel_3251/PIX_OUT pixel_3251/CSA_VREF pixel
Xpixel_3240 pixel_3240/gring pixel_3240/VDD pixel_3240/GND pixel_3240/VREF pixel_3240/ROW_SEL
+ pixel_3240/NB1 pixel_3240/VBIAS pixel_3240/NB2 pixel_3240/AMP_IN pixel_3240/SF_IB
+ pixel_3240/PIX_OUT pixel_3240/CSA_VREF pixel
Xpixel_3284 pixel_3284/gring pixel_3284/VDD pixel_3284/GND pixel_3284/VREF pixel_3284/ROW_SEL
+ pixel_3284/NB1 pixel_3284/VBIAS pixel_3284/NB2 pixel_3284/AMP_IN pixel_3284/SF_IB
+ pixel_3284/PIX_OUT pixel_3284/CSA_VREF pixel
Xpixel_3273 pixel_3273/gring pixel_3273/VDD pixel_3273/GND pixel_3273/VREF pixel_3273/ROW_SEL
+ pixel_3273/NB1 pixel_3273/VBIAS pixel_3273/NB2 pixel_3273/AMP_IN pixel_3273/SF_IB
+ pixel_3273/PIX_OUT pixel_3273/CSA_VREF pixel
Xpixel_3262 pixel_3262/gring pixel_3262/VDD pixel_3262/GND pixel_3262/VREF pixel_3262/ROW_SEL
+ pixel_3262/NB1 pixel_3262/VBIAS pixel_3262/NB2 pixel_3262/AMP_IN pixel_3262/SF_IB
+ pixel_3262/PIX_OUT pixel_3262/CSA_VREF pixel
Xpixel_2572 pixel_2572/gring pixel_2572/VDD pixel_2572/GND pixel_2572/VREF pixel_2572/ROW_SEL
+ pixel_2572/NB1 pixel_2572/VBIAS pixel_2572/NB2 pixel_2572/AMP_IN pixel_2572/SF_IB
+ pixel_2572/PIX_OUT pixel_2572/CSA_VREF pixel
Xpixel_2561 pixel_2561/gring pixel_2561/VDD pixel_2561/GND pixel_2561/VREF pixel_2561/ROW_SEL
+ pixel_2561/NB1 pixel_2561/VBIAS pixel_2561/NB2 pixel_2561/AMP_IN pixel_2561/SF_IB
+ pixel_2561/PIX_OUT pixel_2561/CSA_VREF pixel
Xpixel_2550 pixel_2550/gring pixel_2550/VDD pixel_2550/GND pixel_2550/VREF pixel_2550/ROW_SEL
+ pixel_2550/NB1 pixel_2550/VBIAS pixel_2550/NB2 pixel_2550/AMP_IN pixel_2550/SF_IB
+ pixel_2550/PIX_OUT pixel_2550/CSA_VREF pixel
Xpixel_3295 pixel_3295/gring pixel_3295/VDD pixel_3295/GND pixel_3295/VREF pixel_3295/ROW_SEL
+ pixel_3295/NB1 pixel_3295/VBIAS pixel_3295/NB2 pixel_3295/AMP_IN pixel_3295/SF_IB
+ pixel_3295/PIX_OUT pixel_3295/CSA_VREF pixel
Xpixel_1871 pixel_1871/gring pixel_1871/VDD pixel_1871/GND pixel_1871/VREF pixel_1871/ROW_SEL
+ pixel_1871/NB1 pixel_1871/VBIAS pixel_1871/NB2 pixel_1871/AMP_IN pixel_1871/SF_IB
+ pixel_1871/PIX_OUT pixel_1871/CSA_VREF pixel
Xpixel_1860 pixel_1860/gring pixel_1860/VDD pixel_1860/GND pixel_1860/VREF pixel_1860/ROW_SEL
+ pixel_1860/NB1 pixel_1860/VBIAS pixel_1860/NB2 pixel_1860/AMP_IN pixel_1860/SF_IB
+ pixel_1860/PIX_OUT pixel_1860/CSA_VREF pixel
Xpixel_2594 pixel_2594/gring pixel_2594/VDD pixel_2594/GND pixel_2594/VREF pixel_2594/ROW_SEL
+ pixel_2594/NB1 pixel_2594/VBIAS pixel_2594/NB2 pixel_2594/AMP_IN pixel_2594/SF_IB
+ pixel_2594/PIX_OUT pixel_2594/CSA_VREF pixel
Xpixel_2583 pixel_2583/gring pixel_2583/VDD pixel_2583/GND pixel_2583/VREF pixel_2583/ROW_SEL
+ pixel_2583/NB1 pixel_2583/VBIAS pixel_2583/NB2 pixel_2583/AMP_IN pixel_2583/SF_IB
+ pixel_2583/PIX_OUT pixel_2583/CSA_VREF pixel
Xpixel_1893 pixel_1893/gring pixel_1893/VDD pixel_1893/GND pixel_1893/VREF pixel_1893/ROW_SEL
+ pixel_1893/NB1 pixel_1893/VBIAS pixel_1893/NB2 pixel_1893/AMP_IN pixel_1893/SF_IB
+ pixel_1893/PIX_OUT pixel_1893/CSA_VREF pixel
Xpixel_1882 pixel_1882/gring pixel_1882/VDD pixel_1882/GND pixel_1882/VREF pixel_1882/ROW_SEL
+ pixel_1882/NB1 pixel_1882/VBIAS pixel_1882/NB2 pixel_1882/AMP_IN pixel_1882/SF_IB
+ pixel_1882/PIX_OUT pixel_1882/CSA_VREF pixel
Xpixel_919 pixel_919/gring pixel_919/VDD pixel_919/GND pixel_919/VREF pixel_919/ROW_SEL
+ pixel_919/NB1 pixel_919/VBIAS pixel_919/NB2 pixel_919/AMP_IN pixel_919/SF_IB pixel_919/PIX_OUT
+ pixel_919/CSA_VREF pixel
Xpixel_908 pixel_908/gring pixel_908/VDD pixel_908/GND pixel_908/VREF pixel_908/ROW_SEL
+ pixel_908/NB1 pixel_908/VBIAS pixel_908/NB2 pixel_908/AMP_IN pixel_908/SF_IB pixel_908/PIX_OUT
+ pixel_908/CSA_VREF pixel
Xpixel_8207 pixel_8207/gring pixel_8207/VDD pixel_8207/GND pixel_8207/VREF pixel_8207/ROW_SEL
+ pixel_8207/NB1 pixel_8207/VBIAS pixel_8207/NB2 pixel_8207/AMP_IN pixel_8207/SF_IB
+ pixel_8207/PIX_OUT pixel_8207/CSA_VREF pixel
Xpixel_8218 pixel_8218/gring pixel_8218/VDD pixel_8218/GND pixel_8218/VREF pixel_8218/ROW_SEL
+ pixel_8218/NB1 pixel_8218/VBIAS pixel_8218/NB2 pixel_8218/AMP_IN pixel_8218/SF_IB
+ pixel_8218/PIX_OUT pixel_8218/CSA_VREF pixel
Xpixel_8229 pixel_8229/gring pixel_8229/VDD pixel_8229/GND pixel_8229/VREF pixel_8229/ROW_SEL
+ pixel_8229/NB1 pixel_8229/VBIAS pixel_8229/NB2 pixel_8229/AMP_IN pixel_8229/SF_IB
+ pixel_8229/PIX_OUT pixel_8229/CSA_VREF pixel
Xpixel_7506 pixel_7506/gring pixel_7506/VDD pixel_7506/GND pixel_7506/VREF pixel_7506/ROW_SEL
+ pixel_7506/NB1 pixel_7506/VBIAS pixel_7506/NB2 pixel_7506/AMP_IN pixel_7506/SF_IB
+ pixel_7506/PIX_OUT pixel_7506/CSA_VREF pixel
Xpixel_7517 pixel_7517/gring pixel_7517/VDD pixel_7517/GND pixel_7517/VREF pixel_7517/ROW_SEL
+ pixel_7517/NB1 pixel_7517/VBIAS pixel_7517/NB2 pixel_7517/AMP_IN pixel_7517/SF_IB
+ pixel_7517/PIX_OUT pixel_7517/CSA_VREF pixel
Xpixel_7528 pixel_7528/gring pixel_7528/VDD pixel_7528/GND pixel_7528/VREF pixel_7528/ROW_SEL
+ pixel_7528/NB1 pixel_7528/VBIAS pixel_7528/NB2 pixel_7528/AMP_IN pixel_7528/SF_IB
+ pixel_7528/PIX_OUT pixel_7528/CSA_VREF pixel
Xpixel_7539 pixel_7539/gring pixel_7539/VDD pixel_7539/GND pixel_7539/VREF pixel_7539/ROW_SEL
+ pixel_7539/NB1 pixel_7539/VBIAS pixel_7539/NB2 pixel_7539/AMP_IN pixel_7539/SF_IB
+ pixel_7539/PIX_OUT pixel_7539/CSA_VREF pixel
Xpixel_6805 pixel_6805/gring pixel_6805/VDD pixel_6805/GND pixel_6805/VREF pixel_6805/ROW_SEL
+ pixel_6805/NB1 pixel_6805/VBIAS pixel_6805/NB2 pixel_6805/AMP_IN pixel_6805/SF_IB
+ pixel_6805/PIX_OUT pixel_6805/CSA_VREF pixel
Xpixel_6816 pixel_6816/gring pixel_6816/VDD pixel_6816/GND pixel_6816/VREF pixel_6816/ROW_SEL
+ pixel_6816/NB1 pixel_6816/VBIAS pixel_6816/NB2 pixel_6816/AMP_IN pixel_6816/SF_IB
+ pixel_6816/PIX_OUT pixel_6816/CSA_VREF pixel
Xpixel_6827 pixel_6827/gring pixel_6827/VDD pixel_6827/GND pixel_6827/VREF pixel_6827/ROW_SEL
+ pixel_6827/NB1 pixel_6827/VBIAS pixel_6827/NB2 pixel_6827/AMP_IN pixel_6827/SF_IB
+ pixel_6827/PIX_OUT pixel_6827/CSA_VREF pixel
Xpixel_6838 pixel_6838/gring pixel_6838/VDD pixel_6838/GND pixel_6838/VREF pixel_6838/ROW_SEL
+ pixel_6838/NB1 pixel_6838/VBIAS pixel_6838/NB2 pixel_6838/AMP_IN pixel_6838/SF_IB
+ pixel_6838/PIX_OUT pixel_6838/CSA_VREF pixel
Xpixel_6849 pixel_6849/gring pixel_6849/VDD pixel_6849/GND pixel_6849/VREF pixel_6849/ROW_SEL
+ pixel_6849/NB1 pixel_6849/VBIAS pixel_6849/NB2 pixel_6849/AMP_IN pixel_6849/SF_IB
+ pixel_6849/PIX_OUT pixel_6849/CSA_VREF pixel
Xpixel_1123 pixel_1123/gring pixel_1123/VDD pixel_1123/GND pixel_1123/VREF pixel_1123/ROW_SEL
+ pixel_1123/NB1 pixel_1123/VBIAS pixel_1123/NB2 pixel_1123/AMP_IN pixel_1123/SF_IB
+ pixel_1123/PIX_OUT pixel_1123/CSA_VREF pixel
Xpixel_1112 pixel_1112/gring pixel_1112/VDD pixel_1112/GND pixel_1112/VREF pixel_1112/ROW_SEL
+ pixel_1112/NB1 pixel_1112/VBIAS pixel_1112/NB2 pixel_1112/AMP_IN pixel_1112/SF_IB
+ pixel_1112/PIX_OUT pixel_1112/CSA_VREF pixel
Xpixel_1101 pixel_1101/gring pixel_1101/VDD pixel_1101/GND pixel_1101/VREF pixel_1101/ROW_SEL
+ pixel_1101/NB1 pixel_1101/VBIAS pixel_1101/NB2 pixel_1101/AMP_IN pixel_1101/SF_IB
+ pixel_1101/PIX_OUT pixel_1101/CSA_VREF pixel
Xpixel_1156 pixel_1156/gring pixel_1156/VDD pixel_1156/GND pixel_1156/VREF pixel_1156/ROW_SEL
+ pixel_1156/NB1 pixel_1156/VBIAS pixel_1156/NB2 pixel_1156/AMP_IN pixel_1156/SF_IB
+ pixel_1156/PIX_OUT pixel_1156/CSA_VREF pixel
Xpixel_1145 pixel_1145/gring pixel_1145/VDD pixel_1145/GND pixel_1145/VREF pixel_1145/ROW_SEL
+ pixel_1145/NB1 pixel_1145/VBIAS pixel_1145/NB2 pixel_1145/AMP_IN pixel_1145/SF_IB
+ pixel_1145/PIX_OUT pixel_1145/CSA_VREF pixel
Xpixel_1134 pixel_1134/gring pixel_1134/VDD pixel_1134/GND pixel_1134/VREF pixel_1134/ROW_SEL
+ pixel_1134/NB1 pixel_1134/VBIAS pixel_1134/NB2 pixel_1134/AMP_IN pixel_1134/SF_IB
+ pixel_1134/PIX_OUT pixel_1134/CSA_VREF pixel
Xpixel_1189 pixel_1189/gring pixel_1189/VDD pixel_1189/GND pixel_1189/VREF pixel_1189/ROW_SEL
+ pixel_1189/NB1 pixel_1189/VBIAS pixel_1189/NB2 pixel_1189/AMP_IN pixel_1189/SF_IB
+ pixel_1189/PIX_OUT pixel_1189/CSA_VREF pixel
Xpixel_1178 pixel_1178/gring pixel_1178/VDD pixel_1178/GND pixel_1178/VREF pixel_1178/ROW_SEL
+ pixel_1178/NB1 pixel_1178/VBIAS pixel_1178/NB2 pixel_1178/AMP_IN pixel_1178/SF_IB
+ pixel_1178/PIX_OUT pixel_1178/CSA_VREF pixel
Xpixel_1167 pixel_1167/gring pixel_1167/VDD pixel_1167/GND pixel_1167/VREF pixel_1167/ROW_SEL
+ pixel_1167/NB1 pixel_1167/VBIAS pixel_1167/NB2 pixel_1167/AMP_IN pixel_1167/SF_IB
+ pixel_1167/PIX_OUT pixel_1167/CSA_VREF pixel
Xpixel_9431 pixel_9431/gring pixel_9431/VDD pixel_9431/GND pixel_9431/VREF pixel_9431/ROW_SEL
+ pixel_9431/NB1 pixel_9431/VBIAS pixel_9431/NB2 pixel_9431/AMP_IN pixel_9431/SF_IB
+ pixel_9431/PIX_OUT pixel_9431/CSA_VREF pixel
Xpixel_9420 pixel_9420/gring pixel_9420/VDD pixel_9420/GND pixel_9420/VREF pixel_9420/ROW_SEL
+ pixel_9420/NB1 pixel_9420/VBIAS pixel_9420/NB2 pixel_9420/AMP_IN pixel_9420/SF_IB
+ pixel_9420/PIX_OUT pixel_9420/CSA_VREF pixel
Xpixel_8730 pixel_8730/gring pixel_8730/VDD pixel_8730/GND pixel_8730/VREF pixel_8730/ROW_SEL
+ pixel_8730/NB1 pixel_8730/VBIAS pixel_8730/NB2 pixel_8730/AMP_IN pixel_8730/SF_IB
+ pixel_8730/PIX_OUT pixel_8730/CSA_VREF pixel
Xpixel_9464 pixel_9464/gring pixel_9464/VDD pixel_9464/GND pixel_9464/VREF pixel_9464/ROW_SEL
+ pixel_9464/NB1 pixel_9464/VBIAS pixel_9464/NB2 pixel_9464/AMP_IN pixel_9464/SF_IB
+ pixel_9464/PIX_OUT pixel_9464/CSA_VREF pixel
Xpixel_9453 pixel_9453/gring pixel_9453/VDD pixel_9453/GND pixel_9453/VREF pixel_9453/ROW_SEL
+ pixel_9453/NB1 pixel_9453/VBIAS pixel_9453/NB2 pixel_9453/AMP_IN pixel_9453/SF_IB
+ pixel_9453/PIX_OUT pixel_9453/CSA_VREF pixel
Xpixel_9442 pixel_9442/gring pixel_9442/VDD pixel_9442/GND pixel_9442/VREF pixel_9442/ROW_SEL
+ pixel_9442/NB1 pixel_9442/VBIAS pixel_9442/NB2 pixel_9442/AMP_IN pixel_9442/SF_IB
+ pixel_9442/PIX_OUT pixel_9442/CSA_VREF pixel
Xpixel_8763 pixel_8763/gring pixel_8763/VDD pixel_8763/GND pixel_8763/VREF pixel_8763/ROW_SEL
+ pixel_8763/NB1 pixel_8763/VBIAS pixel_8763/NB2 pixel_8763/AMP_IN pixel_8763/SF_IB
+ pixel_8763/PIX_OUT pixel_8763/CSA_VREF pixel
Xpixel_8752 pixel_8752/gring pixel_8752/VDD pixel_8752/GND pixel_8752/VREF pixel_8752/ROW_SEL
+ pixel_8752/NB1 pixel_8752/VBIAS pixel_8752/NB2 pixel_8752/AMP_IN pixel_8752/SF_IB
+ pixel_8752/PIX_OUT pixel_8752/CSA_VREF pixel
Xpixel_8741 pixel_8741/gring pixel_8741/VDD pixel_8741/GND pixel_8741/VREF pixel_8741/ROW_SEL
+ pixel_8741/NB1 pixel_8741/VBIAS pixel_8741/NB2 pixel_8741/AMP_IN pixel_8741/SF_IB
+ pixel_8741/PIX_OUT pixel_8741/CSA_VREF pixel
Xpixel_9497 pixel_9497/gring pixel_9497/VDD pixel_9497/GND pixel_9497/VREF pixel_9497/ROW_SEL
+ pixel_9497/NB1 pixel_9497/VBIAS pixel_9497/NB2 pixel_9497/AMP_IN pixel_9497/SF_IB
+ pixel_9497/PIX_OUT pixel_9497/CSA_VREF pixel
Xpixel_9486 pixel_9486/gring pixel_9486/VDD pixel_9486/GND pixel_9486/VREF pixel_9486/ROW_SEL
+ pixel_9486/NB1 pixel_9486/VBIAS pixel_9486/NB2 pixel_9486/AMP_IN pixel_9486/SF_IB
+ pixel_9486/PIX_OUT pixel_9486/CSA_VREF pixel
Xpixel_9475 pixel_9475/gring pixel_9475/VDD pixel_9475/GND pixel_9475/VREF pixel_9475/ROW_SEL
+ pixel_9475/NB1 pixel_9475/VBIAS pixel_9475/NB2 pixel_9475/AMP_IN pixel_9475/SF_IB
+ pixel_9475/PIX_OUT pixel_9475/CSA_VREF pixel
Xpixel_8796 pixel_8796/gring pixel_8796/VDD pixel_8796/GND pixel_8796/VREF pixel_8796/ROW_SEL
+ pixel_8796/NB1 pixel_8796/VBIAS pixel_8796/NB2 pixel_8796/AMP_IN pixel_8796/SF_IB
+ pixel_8796/PIX_OUT pixel_8796/CSA_VREF pixel
Xpixel_8785 pixel_8785/gring pixel_8785/VDD pixel_8785/GND pixel_8785/VREF pixel_8785/ROW_SEL
+ pixel_8785/NB1 pixel_8785/VBIAS pixel_8785/NB2 pixel_8785/AMP_IN pixel_8785/SF_IB
+ pixel_8785/PIX_OUT pixel_8785/CSA_VREF pixel
Xpixel_8774 pixel_8774/gring pixel_8774/VDD pixel_8774/GND pixel_8774/VREF pixel_8774/ROW_SEL
+ pixel_8774/NB1 pixel_8774/VBIAS pixel_8774/NB2 pixel_8774/AMP_IN pixel_8774/SF_IB
+ pixel_8774/PIX_OUT pixel_8774/CSA_VREF pixel
Xpixel_3092 pixel_3092/gring pixel_3092/VDD pixel_3092/GND pixel_3092/VREF pixel_3092/ROW_SEL
+ pixel_3092/NB1 pixel_3092/VBIAS pixel_3092/NB2 pixel_3092/AMP_IN pixel_3092/SF_IB
+ pixel_3092/PIX_OUT pixel_3092/CSA_VREF pixel
Xpixel_3081 pixel_3081/gring pixel_3081/VDD pixel_3081/GND pixel_3081/VREF pixel_3081/ROW_SEL
+ pixel_3081/NB1 pixel_3081/VBIAS pixel_3081/NB2 pixel_3081/AMP_IN pixel_3081/SF_IB
+ pixel_3081/PIX_OUT pixel_3081/CSA_VREF pixel
Xpixel_3070 pixel_3070/gring pixel_3070/VDD pixel_3070/GND pixel_3070/VREF pixel_3070/ROW_SEL
+ pixel_3070/NB1 pixel_3070/VBIAS pixel_3070/NB2 pixel_3070/AMP_IN pixel_3070/SF_IB
+ pixel_3070/PIX_OUT pixel_3070/CSA_VREF pixel
Xpixel_2391 pixel_2391/gring pixel_2391/VDD pixel_2391/GND pixel_2391/VREF pixel_2391/ROW_SEL
+ pixel_2391/NB1 pixel_2391/VBIAS pixel_2391/NB2 pixel_2391/AMP_IN pixel_2391/SF_IB
+ pixel_2391/PIX_OUT pixel_2391/CSA_VREF pixel
Xpixel_2380 pixel_2380/gring pixel_2380/VDD pixel_2380/GND pixel_2380/VREF pixel_2380/ROW_SEL
+ pixel_2380/NB1 pixel_2380/VBIAS pixel_2380/NB2 pixel_2380/AMP_IN pixel_2380/SF_IB
+ pixel_2380/PIX_OUT pixel_2380/CSA_VREF pixel
Xpixel_1690 pixel_1690/gring pixel_1690/VDD pixel_1690/GND pixel_1690/VREF pixel_1690/ROW_SEL
+ pixel_1690/NB1 pixel_1690/VBIAS pixel_1690/NB2 pixel_1690/AMP_IN pixel_1690/SF_IB
+ pixel_1690/PIX_OUT pixel_1690/CSA_VREF pixel
Xpixel_705 pixel_705/gring pixel_705/VDD pixel_705/GND pixel_705/VREF pixel_705/ROW_SEL
+ pixel_705/NB1 pixel_705/VBIAS pixel_705/NB2 pixel_705/AMP_IN pixel_705/SF_IB pixel_705/PIX_OUT
+ pixel_705/CSA_VREF pixel
Xpixel_738 pixel_738/gring pixel_738/VDD pixel_738/GND pixel_738/VREF pixel_738/ROW_SEL
+ pixel_738/NB1 pixel_738/VBIAS pixel_738/NB2 pixel_738/AMP_IN pixel_738/SF_IB pixel_738/PIX_OUT
+ pixel_738/CSA_VREF pixel
Xpixel_727 pixel_727/gring pixel_727/VDD pixel_727/GND pixel_727/VREF pixel_727/ROW_SEL
+ pixel_727/NB1 pixel_727/VBIAS pixel_727/NB2 pixel_727/AMP_IN pixel_727/SF_IB pixel_727/PIX_OUT
+ pixel_727/CSA_VREF pixel
Xpixel_716 pixel_716/gring pixel_716/VDD pixel_716/GND pixel_716/VREF pixel_716/ROW_SEL
+ pixel_716/NB1 pixel_716/VBIAS pixel_716/NB2 pixel_716/AMP_IN pixel_716/SF_IB pixel_716/PIX_OUT
+ pixel_716/CSA_VREF pixel
Xpixel_749 pixel_749/gring pixel_749/VDD pixel_749/GND pixel_749/VREF pixel_749/ROW_SEL
+ pixel_749/NB1 pixel_749/VBIAS pixel_749/NB2 pixel_749/AMP_IN pixel_749/SF_IB pixel_749/PIX_OUT
+ pixel_749/CSA_VREF pixel
Xpixel_8004 pixel_8004/gring pixel_8004/VDD pixel_8004/GND pixel_8004/VREF pixel_8004/ROW_SEL
+ pixel_8004/NB1 pixel_8004/VBIAS pixel_8004/NB2 pixel_8004/AMP_IN pixel_8004/SF_IB
+ pixel_8004/PIX_OUT pixel_8004/CSA_VREF pixel
Xpixel_8015 pixel_8015/gring pixel_8015/VDD pixel_8015/GND pixel_8015/VREF pixel_8015/ROW_SEL
+ pixel_8015/NB1 pixel_8015/VBIAS pixel_8015/NB2 pixel_8015/AMP_IN pixel_8015/SF_IB
+ pixel_8015/PIX_OUT pixel_8015/CSA_VREF pixel
Xpixel_8026 pixel_8026/gring pixel_8026/VDD pixel_8026/GND pixel_8026/VREF pixel_8026/ROW_SEL
+ pixel_8026/NB1 pixel_8026/VBIAS pixel_8026/NB2 pixel_8026/AMP_IN pixel_8026/SF_IB
+ pixel_8026/PIX_OUT pixel_8026/CSA_VREF pixel
Xpixel_8037 pixel_8037/gring pixel_8037/VDD pixel_8037/GND pixel_8037/VREF pixel_8037/ROW_SEL
+ pixel_8037/NB1 pixel_8037/VBIAS pixel_8037/NB2 pixel_8037/AMP_IN pixel_8037/SF_IB
+ pixel_8037/PIX_OUT pixel_8037/CSA_VREF pixel
Xpixel_8048 pixel_8048/gring pixel_8048/VDD pixel_8048/GND pixel_8048/VREF pixel_8048/ROW_SEL
+ pixel_8048/NB1 pixel_8048/VBIAS pixel_8048/NB2 pixel_8048/AMP_IN pixel_8048/SF_IB
+ pixel_8048/PIX_OUT pixel_8048/CSA_VREF pixel
Xpixel_8059 pixel_8059/gring pixel_8059/VDD pixel_8059/GND pixel_8059/VREF pixel_8059/ROW_SEL
+ pixel_8059/NB1 pixel_8059/VBIAS pixel_8059/NB2 pixel_8059/AMP_IN pixel_8059/SF_IB
+ pixel_8059/PIX_OUT pixel_8059/CSA_VREF pixel
Xpixel_7303 pixel_7303/gring pixel_7303/VDD pixel_7303/GND pixel_7303/VREF pixel_7303/ROW_SEL
+ pixel_7303/NB1 pixel_7303/VBIAS pixel_7303/NB2 pixel_7303/AMP_IN pixel_7303/SF_IB
+ pixel_7303/PIX_OUT pixel_7303/CSA_VREF pixel
Xpixel_7314 pixel_7314/gring pixel_7314/VDD pixel_7314/GND pixel_7314/VREF pixel_7314/ROW_SEL
+ pixel_7314/NB1 pixel_7314/VBIAS pixel_7314/NB2 pixel_7314/AMP_IN pixel_7314/SF_IB
+ pixel_7314/PIX_OUT pixel_7314/CSA_VREF pixel
Xpixel_7325 pixel_7325/gring pixel_7325/VDD pixel_7325/GND pixel_7325/VREF pixel_7325/ROW_SEL
+ pixel_7325/NB1 pixel_7325/VBIAS pixel_7325/NB2 pixel_7325/AMP_IN pixel_7325/SF_IB
+ pixel_7325/PIX_OUT pixel_7325/CSA_VREF pixel
Xpixel_7336 pixel_7336/gring pixel_7336/VDD pixel_7336/GND pixel_7336/VREF pixel_7336/ROW_SEL
+ pixel_7336/NB1 pixel_7336/VBIAS pixel_7336/NB2 pixel_7336/AMP_IN pixel_7336/SF_IB
+ pixel_7336/PIX_OUT pixel_7336/CSA_VREF pixel
Xpixel_7347 pixel_7347/gring pixel_7347/VDD pixel_7347/GND pixel_7347/VREF pixel_7347/ROW_SEL
+ pixel_7347/NB1 pixel_7347/VBIAS pixel_7347/NB2 pixel_7347/AMP_IN pixel_7347/SF_IB
+ pixel_7347/PIX_OUT pixel_7347/CSA_VREF pixel
Xpixel_6602 pixel_6602/gring pixel_6602/VDD pixel_6602/GND pixel_6602/VREF pixel_6602/ROW_SEL
+ pixel_6602/NB1 pixel_6602/VBIAS pixel_6602/NB2 pixel_6602/AMP_IN pixel_6602/SF_IB
+ pixel_6602/PIX_OUT pixel_6602/CSA_VREF pixel
Xpixel_7358 pixel_7358/gring pixel_7358/VDD pixel_7358/GND pixel_7358/VREF pixel_7358/ROW_SEL
+ pixel_7358/NB1 pixel_7358/VBIAS pixel_7358/NB2 pixel_7358/AMP_IN pixel_7358/SF_IB
+ pixel_7358/PIX_OUT pixel_7358/CSA_VREF pixel
Xpixel_7369 pixel_7369/gring pixel_7369/VDD pixel_7369/GND pixel_7369/VREF pixel_7369/ROW_SEL
+ pixel_7369/NB1 pixel_7369/VBIAS pixel_7369/NB2 pixel_7369/AMP_IN pixel_7369/SF_IB
+ pixel_7369/PIX_OUT pixel_7369/CSA_VREF pixel
Xpixel_6613 pixel_6613/gring pixel_6613/VDD pixel_6613/GND pixel_6613/VREF pixel_6613/ROW_SEL
+ pixel_6613/NB1 pixel_6613/VBIAS pixel_6613/NB2 pixel_6613/AMP_IN pixel_6613/SF_IB
+ pixel_6613/PIX_OUT pixel_6613/CSA_VREF pixel
Xpixel_6624 pixel_6624/gring pixel_6624/VDD pixel_6624/GND pixel_6624/VREF pixel_6624/ROW_SEL
+ pixel_6624/NB1 pixel_6624/VBIAS pixel_6624/NB2 pixel_6624/AMP_IN pixel_6624/SF_IB
+ pixel_6624/PIX_OUT pixel_6624/CSA_VREF pixel
Xpixel_6635 pixel_6635/gring pixel_6635/VDD pixel_6635/GND pixel_6635/VREF pixel_6635/ROW_SEL
+ pixel_6635/NB1 pixel_6635/VBIAS pixel_6635/NB2 pixel_6635/AMP_IN pixel_6635/SF_IB
+ pixel_6635/PIX_OUT pixel_6635/CSA_VREF pixel
Xpixel_5901 pixel_5901/gring pixel_5901/VDD pixel_5901/GND pixel_5901/VREF pixel_5901/ROW_SEL
+ pixel_5901/NB1 pixel_5901/VBIAS pixel_5901/NB2 pixel_5901/AMP_IN pixel_5901/SF_IB
+ pixel_5901/PIX_OUT pixel_5901/CSA_VREF pixel
Xpixel_6646 pixel_6646/gring pixel_6646/VDD pixel_6646/GND pixel_6646/VREF pixel_6646/ROW_SEL
+ pixel_6646/NB1 pixel_6646/VBIAS pixel_6646/NB2 pixel_6646/AMP_IN pixel_6646/SF_IB
+ pixel_6646/PIX_OUT pixel_6646/CSA_VREF pixel
Xpixel_6657 pixel_6657/gring pixel_6657/VDD pixel_6657/GND pixel_6657/VREF pixel_6657/ROW_SEL
+ pixel_6657/NB1 pixel_6657/VBIAS pixel_6657/NB2 pixel_6657/AMP_IN pixel_6657/SF_IB
+ pixel_6657/PIX_OUT pixel_6657/CSA_VREF pixel
Xpixel_6668 pixel_6668/gring pixel_6668/VDD pixel_6668/GND pixel_6668/VREF pixel_6668/ROW_SEL
+ pixel_6668/NB1 pixel_6668/VBIAS pixel_6668/NB2 pixel_6668/AMP_IN pixel_6668/SF_IB
+ pixel_6668/PIX_OUT pixel_6668/CSA_VREF pixel
Xpixel_6679 pixel_6679/gring pixel_6679/VDD pixel_6679/GND pixel_6679/VREF pixel_6679/ROW_SEL
+ pixel_6679/NB1 pixel_6679/VBIAS pixel_6679/NB2 pixel_6679/AMP_IN pixel_6679/SF_IB
+ pixel_6679/PIX_OUT pixel_6679/CSA_VREF pixel
Xpixel_5912 pixel_5912/gring pixel_5912/VDD pixel_5912/GND pixel_5912/VREF pixel_5912/ROW_SEL
+ pixel_5912/NB1 pixel_5912/VBIAS pixel_5912/NB2 pixel_5912/AMP_IN pixel_5912/SF_IB
+ pixel_5912/PIX_OUT pixel_5912/CSA_VREF pixel
Xpixel_5923 pixel_5923/gring pixel_5923/VDD pixel_5923/GND pixel_5923/VREF pixel_5923/ROW_SEL
+ pixel_5923/NB1 pixel_5923/VBIAS pixel_5923/NB2 pixel_5923/AMP_IN pixel_5923/SF_IB
+ pixel_5923/PIX_OUT pixel_5923/CSA_VREF pixel
Xpixel_5934 pixel_5934/gring pixel_5934/VDD pixel_5934/GND pixel_5934/VREF pixel_5934/ROW_SEL
+ pixel_5934/NB1 pixel_5934/VBIAS pixel_5934/NB2 pixel_5934/AMP_IN pixel_5934/SF_IB
+ pixel_5934/PIX_OUT pixel_5934/CSA_VREF pixel
Xpixel_5945 pixel_5945/gring pixel_5945/VDD pixel_5945/GND pixel_5945/VREF pixel_5945/ROW_SEL
+ pixel_5945/NB1 pixel_5945/VBIAS pixel_5945/NB2 pixel_5945/AMP_IN pixel_5945/SF_IB
+ pixel_5945/PIX_OUT pixel_5945/CSA_VREF pixel
Xpixel_5956 pixel_5956/gring pixel_5956/VDD pixel_5956/GND pixel_5956/VREF pixel_5956/ROW_SEL
+ pixel_5956/NB1 pixel_5956/VBIAS pixel_5956/NB2 pixel_5956/AMP_IN pixel_5956/SF_IB
+ pixel_5956/PIX_OUT pixel_5956/CSA_VREF pixel
Xpixel_5967 pixel_5967/gring pixel_5967/VDD pixel_5967/GND pixel_5967/VREF pixel_5967/ROW_SEL
+ pixel_5967/NB1 pixel_5967/VBIAS pixel_5967/NB2 pixel_5967/AMP_IN pixel_5967/SF_IB
+ pixel_5967/PIX_OUT pixel_5967/CSA_VREF pixel
Xpixel_5978 pixel_5978/gring pixel_5978/VDD pixel_5978/GND pixel_5978/VREF pixel_5978/ROW_SEL
+ pixel_5978/NB1 pixel_5978/VBIAS pixel_5978/NB2 pixel_5978/AMP_IN pixel_5978/SF_IB
+ pixel_5978/PIX_OUT pixel_5978/CSA_VREF pixel
Xpixel_5989 pixel_5989/gring pixel_5989/VDD pixel_5989/GND pixel_5989/VREF pixel_5989/ROW_SEL
+ pixel_5989/NB1 pixel_5989/VBIAS pixel_5989/NB2 pixel_5989/AMP_IN pixel_5989/SF_IB
+ pixel_5989/PIX_OUT pixel_5989/CSA_VREF pixel
Xpixel_9283 pixel_9283/gring pixel_9283/VDD pixel_9283/GND pixel_9283/VREF pixel_9283/ROW_SEL
+ pixel_9283/NB1 pixel_9283/VBIAS pixel_9283/NB2 pixel_9283/AMP_IN pixel_9283/SF_IB
+ pixel_9283/PIX_OUT pixel_9283/CSA_VREF pixel
Xpixel_9272 pixel_9272/gring pixel_9272/VDD pixel_9272/GND pixel_9272/VREF pixel_9272/ROW_SEL
+ pixel_9272/NB1 pixel_9272/VBIAS pixel_9272/NB2 pixel_9272/AMP_IN pixel_9272/SF_IB
+ pixel_9272/PIX_OUT pixel_9272/CSA_VREF pixel
Xpixel_9261 pixel_9261/gring pixel_9261/VDD pixel_9261/GND pixel_9261/VREF pixel_9261/ROW_SEL
+ pixel_9261/NB1 pixel_9261/VBIAS pixel_9261/NB2 pixel_9261/AMP_IN pixel_9261/SF_IB
+ pixel_9261/PIX_OUT pixel_9261/CSA_VREF pixel
Xpixel_9250 pixel_9250/gring pixel_9250/VDD pixel_9250/GND pixel_9250/VREF pixel_9250/ROW_SEL
+ pixel_9250/NB1 pixel_9250/VBIAS pixel_9250/NB2 pixel_9250/AMP_IN pixel_9250/SF_IB
+ pixel_9250/PIX_OUT pixel_9250/CSA_VREF pixel
Xpixel_8571 pixel_8571/gring pixel_8571/VDD pixel_8571/GND pixel_8571/VREF pixel_8571/ROW_SEL
+ pixel_8571/NB1 pixel_8571/VBIAS pixel_8571/NB2 pixel_8571/AMP_IN pixel_8571/SF_IB
+ pixel_8571/PIX_OUT pixel_8571/CSA_VREF pixel
Xpixel_8560 pixel_8560/gring pixel_8560/VDD pixel_8560/GND pixel_8560/VREF pixel_8560/ROW_SEL
+ pixel_8560/NB1 pixel_8560/VBIAS pixel_8560/NB2 pixel_8560/AMP_IN pixel_8560/SF_IB
+ pixel_8560/PIX_OUT pixel_8560/CSA_VREF pixel
Xpixel_9294 pixel_9294/gring pixel_9294/VDD pixel_9294/GND pixel_9294/VREF pixel_9294/ROW_SEL
+ pixel_9294/NB1 pixel_9294/VBIAS pixel_9294/NB2 pixel_9294/AMP_IN pixel_9294/SF_IB
+ pixel_9294/PIX_OUT pixel_9294/CSA_VREF pixel
Xpixel_8593 pixel_8593/gring pixel_8593/VDD pixel_8593/GND pixel_8593/VREF pixel_8593/ROW_SEL
+ pixel_8593/NB1 pixel_8593/VBIAS pixel_8593/NB2 pixel_8593/AMP_IN pixel_8593/SF_IB
+ pixel_8593/PIX_OUT pixel_8593/CSA_VREF pixel
Xpixel_8582 pixel_8582/gring pixel_8582/VDD pixel_8582/GND pixel_8582/VREF pixel_8582/ROW_SEL
+ pixel_8582/NB1 pixel_8582/VBIAS pixel_8582/NB2 pixel_8582/AMP_IN pixel_8582/SF_IB
+ pixel_8582/PIX_OUT pixel_8582/CSA_VREF pixel
Xpixel_7870 pixel_7870/gring pixel_7870/VDD pixel_7870/GND pixel_7870/VREF pixel_7870/ROW_SEL
+ pixel_7870/NB1 pixel_7870/VBIAS pixel_7870/NB2 pixel_7870/AMP_IN pixel_7870/SF_IB
+ pixel_7870/PIX_OUT pixel_7870/CSA_VREF pixel
Xpixel_7881 pixel_7881/gring pixel_7881/VDD pixel_7881/GND pixel_7881/VREF pixel_7881/ROW_SEL
+ pixel_7881/NB1 pixel_7881/VBIAS pixel_7881/NB2 pixel_7881/AMP_IN pixel_7881/SF_IB
+ pixel_7881/PIX_OUT pixel_7881/CSA_VREF pixel
Xpixel_7892 pixel_7892/gring pixel_7892/VDD pixel_7892/GND pixel_7892/VREF pixel_7892/ROW_SEL
+ pixel_7892/NB1 pixel_7892/VBIAS pixel_7892/NB2 pixel_7892/AMP_IN pixel_7892/SF_IB
+ pixel_7892/PIX_OUT pixel_7892/CSA_VREF pixel
Xpixel_5208 pixel_5208/gring pixel_5208/VDD pixel_5208/GND pixel_5208/VREF pixel_5208/ROW_SEL
+ pixel_5208/NB1 pixel_5208/VBIAS pixel_5208/NB2 pixel_5208/AMP_IN pixel_5208/SF_IB
+ pixel_5208/PIX_OUT pixel_5208/CSA_VREF pixel
Xpixel_5219 pixel_5219/gring pixel_5219/VDD pixel_5219/GND pixel_5219/VREF pixel_5219/ROW_SEL
+ pixel_5219/NB1 pixel_5219/VBIAS pixel_5219/NB2 pixel_5219/AMP_IN pixel_5219/SF_IB
+ pixel_5219/PIX_OUT pixel_5219/CSA_VREF pixel
Xpixel_513 pixel_513/gring pixel_513/VDD pixel_513/GND pixel_513/VREF pixel_513/ROW_SEL
+ pixel_513/NB1 pixel_513/VBIAS pixel_513/NB2 pixel_513/AMP_IN pixel_513/SF_IB pixel_513/PIX_OUT
+ pixel_513/CSA_VREF pixel
Xpixel_502 pixel_502/gring pixel_502/VDD pixel_502/GND pixel_502/VREF pixel_502/ROW_SEL
+ pixel_502/NB1 pixel_502/VBIAS pixel_502/NB2 pixel_502/AMP_IN pixel_502/SF_IB pixel_502/PIX_OUT
+ pixel_502/CSA_VREF pixel
Xpixel_4507 pixel_4507/gring pixel_4507/VDD pixel_4507/GND pixel_4507/VREF pixel_4507/ROW_SEL
+ pixel_4507/NB1 pixel_4507/VBIAS pixel_4507/NB2 pixel_4507/AMP_IN pixel_4507/SF_IB
+ pixel_4507/PIX_OUT pixel_4507/CSA_VREF pixel
Xpixel_4518 pixel_4518/gring pixel_4518/VDD pixel_4518/GND pixel_4518/VREF pixel_4518/ROW_SEL
+ pixel_4518/NB1 pixel_4518/VBIAS pixel_4518/NB2 pixel_4518/AMP_IN pixel_4518/SF_IB
+ pixel_4518/PIX_OUT pixel_4518/CSA_VREF pixel
Xpixel_557 pixel_557/gring pixel_557/VDD pixel_557/GND pixel_557/VREF pixel_557/ROW_SEL
+ pixel_557/NB1 pixel_557/VBIAS pixel_557/NB2 pixel_557/AMP_IN pixel_557/SF_IB pixel_557/PIX_OUT
+ pixel_557/CSA_VREF pixel
Xpixel_546 pixel_546/gring pixel_546/VDD pixel_546/GND pixel_546/VREF pixel_546/ROW_SEL
+ pixel_546/NB1 pixel_546/VBIAS pixel_546/NB2 pixel_546/AMP_IN pixel_546/SF_IB pixel_546/PIX_OUT
+ pixel_546/CSA_VREF pixel
Xpixel_535 pixel_535/gring pixel_535/VDD pixel_535/GND pixel_535/VREF pixel_535/ROW_SEL
+ pixel_535/NB1 pixel_535/VBIAS pixel_535/NB2 pixel_535/AMP_IN pixel_535/SF_IB pixel_535/PIX_OUT
+ pixel_535/CSA_VREF pixel
Xpixel_524 pixel_524/gring pixel_524/VDD pixel_524/GND pixel_524/VREF pixel_524/ROW_SEL
+ pixel_524/NB1 pixel_524/VBIAS pixel_524/NB2 pixel_524/AMP_IN pixel_524/SF_IB pixel_524/PIX_OUT
+ pixel_524/CSA_VREF pixel
Xpixel_4529 pixel_4529/gring pixel_4529/VDD pixel_4529/GND pixel_4529/VREF pixel_4529/ROW_SEL
+ pixel_4529/NB1 pixel_4529/VBIAS pixel_4529/NB2 pixel_4529/AMP_IN pixel_4529/SF_IB
+ pixel_4529/PIX_OUT pixel_4529/CSA_VREF pixel
Xpixel_3806 pixel_3806/gring pixel_3806/VDD pixel_3806/GND pixel_3806/VREF pixel_3806/ROW_SEL
+ pixel_3806/NB1 pixel_3806/VBIAS pixel_3806/NB2 pixel_3806/AMP_IN pixel_3806/SF_IB
+ pixel_3806/PIX_OUT pixel_3806/CSA_VREF pixel
Xpixel_579 pixel_579/gring pixel_579/VDD pixel_579/GND pixel_579/VREF pixel_579/ROW_SEL
+ pixel_579/NB1 pixel_579/VBIAS pixel_579/NB2 pixel_579/AMP_IN pixel_579/SF_IB pixel_579/PIX_OUT
+ pixel_579/CSA_VREF pixel
Xpixel_568 pixel_568/gring pixel_568/VDD pixel_568/GND pixel_568/VREF pixel_568/ROW_SEL
+ pixel_568/NB1 pixel_568/VBIAS pixel_568/NB2 pixel_568/AMP_IN pixel_568/SF_IB pixel_568/PIX_OUT
+ pixel_568/CSA_VREF pixel
Xpixel_3817 pixel_3817/gring pixel_3817/VDD pixel_3817/GND pixel_3817/VREF pixel_3817/ROW_SEL
+ pixel_3817/NB1 pixel_3817/VBIAS pixel_3817/NB2 pixel_3817/AMP_IN pixel_3817/SF_IB
+ pixel_3817/PIX_OUT pixel_3817/CSA_VREF pixel
Xpixel_3828 pixel_3828/gring pixel_3828/VDD pixel_3828/GND pixel_3828/VREF pixel_3828/ROW_SEL
+ pixel_3828/NB1 pixel_3828/VBIAS pixel_3828/NB2 pixel_3828/AMP_IN pixel_3828/SF_IB
+ pixel_3828/PIX_OUT pixel_3828/CSA_VREF pixel
Xpixel_3839 pixel_3839/gring pixel_3839/VDD pixel_3839/GND pixel_3839/VREF pixel_3839/ROW_SEL
+ pixel_3839/NB1 pixel_3839/VBIAS pixel_3839/NB2 pixel_3839/AMP_IN pixel_3839/SF_IB
+ pixel_3839/PIX_OUT pixel_3839/CSA_VREF pixel
Xpixel_7100 pixel_7100/gring pixel_7100/VDD pixel_7100/GND pixel_7100/VREF pixel_7100/ROW_SEL
+ pixel_7100/NB1 pixel_7100/VBIAS pixel_7100/NB2 pixel_7100/AMP_IN pixel_7100/SF_IB
+ pixel_7100/PIX_OUT pixel_7100/CSA_VREF pixel
Xpixel_7111 pixel_7111/gring pixel_7111/VDD pixel_7111/GND pixel_7111/VREF pixel_7111/ROW_SEL
+ pixel_7111/NB1 pixel_7111/VBIAS pixel_7111/NB2 pixel_7111/AMP_IN pixel_7111/SF_IB
+ pixel_7111/PIX_OUT pixel_7111/CSA_VREF pixel
Xpixel_7122 pixel_7122/gring pixel_7122/VDD pixel_7122/GND pixel_7122/VREF pixel_7122/ROW_SEL
+ pixel_7122/NB1 pixel_7122/VBIAS pixel_7122/NB2 pixel_7122/AMP_IN pixel_7122/SF_IB
+ pixel_7122/PIX_OUT pixel_7122/CSA_VREF pixel
Xpixel_7133 pixel_7133/gring pixel_7133/VDD pixel_7133/GND pixel_7133/VREF pixel_7133/ROW_SEL
+ pixel_7133/NB1 pixel_7133/VBIAS pixel_7133/NB2 pixel_7133/AMP_IN pixel_7133/SF_IB
+ pixel_7133/PIX_OUT pixel_7133/CSA_VREF pixel
Xpixel_7144 pixel_7144/gring pixel_7144/VDD pixel_7144/GND pixel_7144/VREF pixel_7144/ROW_SEL
+ pixel_7144/NB1 pixel_7144/VBIAS pixel_7144/NB2 pixel_7144/AMP_IN pixel_7144/SF_IB
+ pixel_7144/PIX_OUT pixel_7144/CSA_VREF pixel
Xpixel_7155 pixel_7155/gring pixel_7155/VDD pixel_7155/GND pixel_7155/VREF pixel_7155/ROW_SEL
+ pixel_7155/NB1 pixel_7155/VBIAS pixel_7155/NB2 pixel_7155/AMP_IN pixel_7155/SF_IB
+ pixel_7155/PIX_OUT pixel_7155/CSA_VREF pixel
Xpixel_6410 pixel_6410/gring pixel_6410/VDD pixel_6410/GND pixel_6410/VREF pixel_6410/ROW_SEL
+ pixel_6410/NB1 pixel_6410/VBIAS pixel_6410/NB2 pixel_6410/AMP_IN pixel_6410/SF_IB
+ pixel_6410/PIX_OUT pixel_6410/CSA_VREF pixel
Xpixel_7166 pixel_7166/gring pixel_7166/VDD pixel_7166/GND pixel_7166/VREF pixel_7166/ROW_SEL
+ pixel_7166/NB1 pixel_7166/VBIAS pixel_7166/NB2 pixel_7166/AMP_IN pixel_7166/SF_IB
+ pixel_7166/PIX_OUT pixel_7166/CSA_VREF pixel
Xpixel_7177 pixel_7177/gring pixel_7177/VDD pixel_7177/GND pixel_7177/VREF pixel_7177/ROW_SEL
+ pixel_7177/NB1 pixel_7177/VBIAS pixel_7177/NB2 pixel_7177/AMP_IN pixel_7177/SF_IB
+ pixel_7177/PIX_OUT pixel_7177/CSA_VREF pixel
Xpixel_7188 pixel_7188/gring pixel_7188/VDD pixel_7188/GND pixel_7188/VREF pixel_7188/ROW_SEL
+ pixel_7188/NB1 pixel_7188/VBIAS pixel_7188/NB2 pixel_7188/AMP_IN pixel_7188/SF_IB
+ pixel_7188/PIX_OUT pixel_7188/CSA_VREF pixel
Xpixel_7199 pixel_7199/gring pixel_7199/VDD pixel_7199/GND pixel_7199/VREF pixel_7199/ROW_SEL
+ pixel_7199/NB1 pixel_7199/VBIAS pixel_7199/NB2 pixel_7199/AMP_IN pixel_7199/SF_IB
+ pixel_7199/PIX_OUT pixel_7199/CSA_VREF pixel
Xpixel_6421 pixel_6421/gring pixel_6421/VDD pixel_6421/GND pixel_6421/VREF pixel_6421/ROW_SEL
+ pixel_6421/NB1 pixel_6421/VBIAS pixel_6421/NB2 pixel_6421/AMP_IN pixel_6421/SF_IB
+ pixel_6421/PIX_OUT pixel_6421/CSA_VREF pixel
Xpixel_6432 pixel_6432/gring pixel_6432/VDD pixel_6432/GND pixel_6432/VREF pixel_6432/ROW_SEL
+ pixel_6432/NB1 pixel_6432/VBIAS pixel_6432/NB2 pixel_6432/AMP_IN pixel_6432/SF_IB
+ pixel_6432/PIX_OUT pixel_6432/CSA_VREF pixel
Xpixel_6443 pixel_6443/gring pixel_6443/VDD pixel_6443/GND pixel_6443/VREF pixel_6443/ROW_SEL
+ pixel_6443/NB1 pixel_6443/VBIAS pixel_6443/NB2 pixel_6443/AMP_IN pixel_6443/SF_IB
+ pixel_6443/PIX_OUT pixel_6443/CSA_VREF pixel
Xpixel_6454 pixel_6454/gring pixel_6454/VDD pixel_6454/GND pixel_6454/VREF pixel_6454/ROW_SEL
+ pixel_6454/NB1 pixel_6454/VBIAS pixel_6454/NB2 pixel_6454/AMP_IN pixel_6454/SF_IB
+ pixel_6454/PIX_OUT pixel_6454/CSA_VREF pixel
Xpixel_6465 pixel_6465/gring pixel_6465/VDD pixel_6465/GND pixel_6465/VREF pixel_6465/ROW_SEL
+ pixel_6465/NB1 pixel_6465/VBIAS pixel_6465/NB2 pixel_6465/AMP_IN pixel_6465/SF_IB
+ pixel_6465/PIX_OUT pixel_6465/CSA_VREF pixel
Xpixel_6476 pixel_6476/gring pixel_6476/VDD pixel_6476/GND pixel_6476/VREF pixel_6476/ROW_SEL
+ pixel_6476/NB1 pixel_6476/VBIAS pixel_6476/NB2 pixel_6476/AMP_IN pixel_6476/SF_IB
+ pixel_6476/PIX_OUT pixel_6476/CSA_VREF pixel
Xpixel_6487 pixel_6487/gring pixel_6487/VDD pixel_6487/GND pixel_6487/VREF pixel_6487/ROW_SEL
+ pixel_6487/NB1 pixel_6487/VBIAS pixel_6487/NB2 pixel_6487/AMP_IN pixel_6487/SF_IB
+ pixel_6487/PIX_OUT pixel_6487/CSA_VREF pixel
Xpixel_5720 pixel_5720/gring pixel_5720/VDD pixel_5720/GND pixel_5720/VREF pixel_5720/ROW_SEL
+ pixel_5720/NB1 pixel_5720/VBIAS pixel_5720/NB2 pixel_5720/AMP_IN pixel_5720/SF_IB
+ pixel_5720/PIX_OUT pixel_5720/CSA_VREF pixel
Xpixel_5731 pixel_5731/gring pixel_5731/VDD pixel_5731/GND pixel_5731/VREF pixel_5731/ROW_SEL
+ pixel_5731/NB1 pixel_5731/VBIAS pixel_5731/NB2 pixel_5731/AMP_IN pixel_5731/SF_IB
+ pixel_5731/PIX_OUT pixel_5731/CSA_VREF pixel
Xpixel_5742 pixel_5742/gring pixel_5742/VDD pixel_5742/GND pixel_5742/VREF pixel_5742/ROW_SEL
+ pixel_5742/NB1 pixel_5742/VBIAS pixel_5742/NB2 pixel_5742/AMP_IN pixel_5742/SF_IB
+ pixel_5742/PIX_OUT pixel_5742/CSA_VREF pixel
Xpixel_6498 pixel_6498/gring pixel_6498/VDD pixel_6498/GND pixel_6498/VREF pixel_6498/ROW_SEL
+ pixel_6498/NB1 pixel_6498/VBIAS pixel_6498/NB2 pixel_6498/AMP_IN pixel_6498/SF_IB
+ pixel_6498/PIX_OUT pixel_6498/CSA_VREF pixel
Xpixel_5753 pixel_5753/gring pixel_5753/VDD pixel_5753/GND pixel_5753/VREF pixel_5753/ROW_SEL
+ pixel_5753/NB1 pixel_5753/VBIAS pixel_5753/NB2 pixel_5753/AMP_IN pixel_5753/SF_IB
+ pixel_5753/PIX_OUT pixel_5753/CSA_VREF pixel
Xpixel_5764 pixel_5764/gring pixel_5764/VDD pixel_5764/GND pixel_5764/VREF pixel_5764/ROW_SEL
+ pixel_5764/NB1 pixel_5764/VBIAS pixel_5764/NB2 pixel_5764/AMP_IN pixel_5764/SF_IB
+ pixel_5764/PIX_OUT pixel_5764/CSA_VREF pixel
Xpixel_5775 pixel_5775/gring pixel_5775/VDD pixel_5775/GND pixel_5775/VREF pixel_5775/ROW_SEL
+ pixel_5775/NB1 pixel_5775/VBIAS pixel_5775/NB2 pixel_5775/AMP_IN pixel_5775/SF_IB
+ pixel_5775/PIX_OUT pixel_5775/CSA_VREF pixel
Xpixel_5786 pixel_5786/gring pixel_5786/VDD pixel_5786/GND pixel_5786/VREF pixel_5786/ROW_SEL
+ pixel_5786/NB1 pixel_5786/VBIAS pixel_5786/NB2 pixel_5786/AMP_IN pixel_5786/SF_IB
+ pixel_5786/PIX_OUT pixel_5786/CSA_VREF pixel
Xpixel_5797 pixel_5797/gring pixel_5797/VDD pixel_5797/GND pixel_5797/VREF pixel_5797/ROW_SEL
+ pixel_5797/NB1 pixel_5797/VBIAS pixel_5797/NB2 pixel_5797/AMP_IN pixel_5797/SF_IB
+ pixel_5797/PIX_OUT pixel_5797/CSA_VREF pixel
Xpixel_9091 pixel_9091/gring pixel_9091/VDD pixel_9091/GND pixel_9091/VREF pixel_9091/ROW_SEL
+ pixel_9091/NB1 pixel_9091/VBIAS pixel_9091/NB2 pixel_9091/AMP_IN pixel_9091/SF_IB
+ pixel_9091/PIX_OUT pixel_9091/CSA_VREF pixel
Xpixel_9080 pixel_9080/gring pixel_9080/VDD pixel_9080/GND pixel_9080/VREF pixel_9080/ROW_SEL
+ pixel_9080/NB1 pixel_9080/VBIAS pixel_9080/NB2 pixel_9080/AMP_IN pixel_9080/SF_IB
+ pixel_9080/PIX_OUT pixel_9080/CSA_VREF pixel
Xpixel_8390 pixel_8390/gring pixel_8390/VDD pixel_8390/GND pixel_8390/VREF pixel_8390/ROW_SEL
+ pixel_8390/NB1 pixel_8390/VBIAS pixel_8390/NB2 pixel_8390/AMP_IN pixel_8390/SF_IB
+ pixel_8390/PIX_OUT pixel_8390/CSA_VREF pixel
Xpixel_91 pixel_91/gring pixel_91/VDD pixel_91/GND pixel_91/VREF pixel_91/ROW_SEL
+ pixel_91/NB1 pixel_91/VBIAS pixel_91/NB2 pixel_91/AMP_IN pixel_91/SF_IB pixel_91/PIX_OUT
+ pixel_91/CSA_VREF pixel
Xpixel_80 pixel_80/gring pixel_80/VDD pixel_80/GND pixel_80/VREF pixel_80/ROW_SEL
+ pixel_80/NB1 pixel_80/VBIAS pixel_80/NB2 pixel_80/AMP_IN pixel_80/SF_IB pixel_80/PIX_OUT
+ pixel_80/CSA_VREF pixel
Xpixel_5005 pixel_5005/gring pixel_5005/VDD pixel_5005/GND pixel_5005/VREF pixel_5005/ROW_SEL
+ pixel_5005/NB1 pixel_5005/VBIAS pixel_5005/NB2 pixel_5005/AMP_IN pixel_5005/SF_IB
+ pixel_5005/PIX_OUT pixel_5005/CSA_VREF pixel
Xpixel_5016 pixel_5016/gring pixel_5016/VDD pixel_5016/GND pixel_5016/VREF pixel_5016/ROW_SEL
+ pixel_5016/NB1 pixel_5016/VBIAS pixel_5016/NB2 pixel_5016/AMP_IN pixel_5016/SF_IB
+ pixel_5016/PIX_OUT pixel_5016/CSA_VREF pixel
Xpixel_5027 pixel_5027/gring pixel_5027/VDD pixel_5027/GND pixel_5027/VREF pixel_5027/ROW_SEL
+ pixel_5027/NB1 pixel_5027/VBIAS pixel_5027/NB2 pixel_5027/AMP_IN pixel_5027/SF_IB
+ pixel_5027/PIX_OUT pixel_5027/CSA_VREF pixel
Xpixel_5038 pixel_5038/gring pixel_5038/VDD pixel_5038/GND pixel_5038/VREF pixel_5038/ROW_SEL
+ pixel_5038/NB1 pixel_5038/VBIAS pixel_5038/NB2 pixel_5038/AMP_IN pixel_5038/SF_IB
+ pixel_5038/PIX_OUT pixel_5038/CSA_VREF pixel
Xpixel_321 pixel_321/gring pixel_321/VDD pixel_321/GND pixel_321/VREF pixel_321/ROW_SEL
+ pixel_321/NB1 pixel_321/VBIAS pixel_321/NB2 pixel_321/AMP_IN pixel_321/SF_IB pixel_321/PIX_OUT
+ pixel_321/CSA_VREF pixel
Xpixel_310 pixel_310/gring pixel_310/VDD pixel_310/GND pixel_310/VREF pixel_310/ROW_SEL
+ pixel_310/NB1 pixel_310/VBIAS pixel_310/NB2 pixel_310/AMP_IN pixel_310/SF_IB pixel_310/PIX_OUT
+ pixel_310/CSA_VREF pixel
Xpixel_5049 pixel_5049/gring pixel_5049/VDD pixel_5049/GND pixel_5049/VREF pixel_5049/ROW_SEL
+ pixel_5049/NB1 pixel_5049/VBIAS pixel_5049/NB2 pixel_5049/AMP_IN pixel_5049/SF_IB
+ pixel_5049/PIX_OUT pixel_5049/CSA_VREF pixel
Xpixel_4304 pixel_4304/gring pixel_4304/VDD pixel_4304/GND pixel_4304/VREF pixel_4304/ROW_SEL
+ pixel_4304/NB1 pixel_4304/VBIAS pixel_4304/NB2 pixel_4304/AMP_IN pixel_4304/SF_IB
+ pixel_4304/PIX_OUT pixel_4304/CSA_VREF pixel
Xpixel_4315 pixel_4315/gring pixel_4315/VDD pixel_4315/GND pixel_4315/VREF pixel_4315/ROW_SEL
+ pixel_4315/NB1 pixel_4315/VBIAS pixel_4315/NB2 pixel_4315/AMP_IN pixel_4315/SF_IB
+ pixel_4315/PIX_OUT pixel_4315/CSA_VREF pixel
Xpixel_4326 pixel_4326/gring pixel_4326/VDD pixel_4326/GND pixel_4326/VREF pixel_4326/ROW_SEL
+ pixel_4326/NB1 pixel_4326/VBIAS pixel_4326/NB2 pixel_4326/AMP_IN pixel_4326/SF_IB
+ pixel_4326/PIX_OUT pixel_4326/CSA_VREF pixel
Xpixel_365 pixel_365/gring pixel_365/VDD pixel_365/GND pixel_365/VREF pixel_365/ROW_SEL
+ pixel_365/NB1 pixel_365/VBIAS pixel_365/NB2 pixel_365/AMP_IN pixel_365/SF_IB pixel_365/PIX_OUT
+ pixel_365/CSA_VREF pixel
Xpixel_354 pixel_354/gring pixel_354/VDD pixel_354/GND pixel_354/VREF pixel_354/ROW_SEL
+ pixel_354/NB1 pixel_354/VBIAS pixel_354/NB2 pixel_354/AMP_IN pixel_354/SF_IB pixel_354/PIX_OUT
+ pixel_354/CSA_VREF pixel
Xpixel_343 pixel_343/gring pixel_343/VDD pixel_343/GND pixel_343/VREF pixel_343/ROW_SEL
+ pixel_343/NB1 pixel_343/VBIAS pixel_343/NB2 pixel_343/AMP_IN pixel_343/SF_IB pixel_343/PIX_OUT
+ pixel_343/CSA_VREF pixel
Xpixel_332 pixel_332/gring pixel_332/VDD pixel_332/GND pixel_332/VREF pixel_332/ROW_SEL
+ pixel_332/NB1 pixel_332/VBIAS pixel_332/NB2 pixel_332/AMP_IN pixel_332/SF_IB pixel_332/PIX_OUT
+ pixel_332/CSA_VREF pixel
Xpixel_3625 pixel_3625/gring pixel_3625/VDD pixel_3625/GND pixel_3625/VREF pixel_3625/ROW_SEL
+ pixel_3625/NB1 pixel_3625/VBIAS pixel_3625/NB2 pixel_3625/AMP_IN pixel_3625/SF_IB
+ pixel_3625/PIX_OUT pixel_3625/CSA_VREF pixel
Xpixel_3614 pixel_3614/gring pixel_3614/VDD pixel_3614/GND pixel_3614/VREF pixel_3614/ROW_SEL
+ pixel_3614/NB1 pixel_3614/VBIAS pixel_3614/NB2 pixel_3614/AMP_IN pixel_3614/SF_IB
+ pixel_3614/PIX_OUT pixel_3614/CSA_VREF pixel
Xpixel_3603 pixel_3603/gring pixel_3603/VDD pixel_3603/GND pixel_3603/VREF pixel_3603/ROW_SEL
+ pixel_3603/NB1 pixel_3603/VBIAS pixel_3603/NB2 pixel_3603/AMP_IN pixel_3603/SF_IB
+ pixel_3603/PIX_OUT pixel_3603/CSA_VREF pixel
Xpixel_4337 pixel_4337/gring pixel_4337/VDD pixel_4337/GND pixel_4337/VREF pixel_4337/ROW_SEL
+ pixel_4337/NB1 pixel_4337/VBIAS pixel_4337/NB2 pixel_4337/AMP_IN pixel_4337/SF_IB
+ pixel_4337/PIX_OUT pixel_4337/CSA_VREF pixel
Xpixel_4348 pixel_4348/gring pixel_4348/VDD pixel_4348/GND pixel_4348/VREF pixel_4348/ROW_SEL
+ pixel_4348/NB1 pixel_4348/VBIAS pixel_4348/NB2 pixel_4348/AMP_IN pixel_4348/SF_IB
+ pixel_4348/PIX_OUT pixel_4348/CSA_VREF pixel
Xpixel_4359 pixel_4359/gring pixel_4359/VDD pixel_4359/GND pixel_4359/VREF pixel_4359/ROW_SEL
+ pixel_4359/NB1 pixel_4359/VBIAS pixel_4359/NB2 pixel_4359/AMP_IN pixel_4359/SF_IB
+ pixel_4359/PIX_OUT pixel_4359/CSA_VREF pixel
Xpixel_398 pixel_398/gring pixel_398/VDD pixel_398/GND pixel_398/VREF pixel_398/ROW_SEL
+ pixel_398/NB1 pixel_398/VBIAS pixel_398/NB2 pixel_398/AMP_IN pixel_398/SF_IB pixel_398/PIX_OUT
+ pixel_398/CSA_VREF pixel
Xpixel_387 pixel_387/gring pixel_387/VDD pixel_387/GND pixel_387/VREF pixel_387/ROW_SEL
+ pixel_387/NB1 pixel_387/VBIAS pixel_387/NB2 pixel_387/AMP_IN pixel_387/SF_IB pixel_387/PIX_OUT
+ pixel_387/CSA_VREF pixel
Xpixel_376 pixel_376/gring pixel_376/VDD pixel_376/GND pixel_376/VREF pixel_376/ROW_SEL
+ pixel_376/NB1 pixel_376/VBIAS pixel_376/NB2 pixel_376/AMP_IN pixel_376/SF_IB pixel_376/PIX_OUT
+ pixel_376/CSA_VREF pixel
Xpixel_2913 pixel_2913/gring pixel_2913/VDD pixel_2913/GND pixel_2913/VREF pixel_2913/ROW_SEL
+ pixel_2913/NB1 pixel_2913/VBIAS pixel_2913/NB2 pixel_2913/AMP_IN pixel_2913/SF_IB
+ pixel_2913/PIX_OUT pixel_2913/CSA_VREF pixel
Xpixel_2902 pixel_2902/gring pixel_2902/VDD pixel_2902/GND pixel_2902/VREF pixel_2902/ROW_SEL
+ pixel_2902/NB1 pixel_2902/VBIAS pixel_2902/NB2 pixel_2902/AMP_IN pixel_2902/SF_IB
+ pixel_2902/PIX_OUT pixel_2902/CSA_VREF pixel
Xpixel_3658 pixel_3658/gring pixel_3658/VDD pixel_3658/GND pixel_3658/VREF pixel_3658/ROW_SEL
+ pixel_3658/NB1 pixel_3658/VBIAS pixel_3658/NB2 pixel_3658/AMP_IN pixel_3658/SF_IB
+ pixel_3658/PIX_OUT pixel_3658/CSA_VREF pixel
Xpixel_3647 pixel_3647/gring pixel_3647/VDD pixel_3647/GND pixel_3647/VREF pixel_3647/ROW_SEL
+ pixel_3647/NB1 pixel_3647/VBIAS pixel_3647/NB2 pixel_3647/AMP_IN pixel_3647/SF_IB
+ pixel_3647/PIX_OUT pixel_3647/CSA_VREF pixel
Xpixel_3636 pixel_3636/gring pixel_3636/VDD pixel_3636/GND pixel_3636/VREF pixel_3636/ROW_SEL
+ pixel_3636/NB1 pixel_3636/VBIAS pixel_3636/NB2 pixel_3636/AMP_IN pixel_3636/SF_IB
+ pixel_3636/PIX_OUT pixel_3636/CSA_VREF pixel
Xpixel_2946 pixel_2946/gring pixel_2946/VDD pixel_2946/GND pixel_2946/VREF pixel_2946/ROW_SEL
+ pixel_2946/NB1 pixel_2946/VBIAS pixel_2946/NB2 pixel_2946/AMP_IN pixel_2946/SF_IB
+ pixel_2946/PIX_OUT pixel_2946/CSA_VREF pixel
Xpixel_2935 pixel_2935/gring pixel_2935/VDD pixel_2935/GND pixel_2935/VREF pixel_2935/ROW_SEL
+ pixel_2935/NB1 pixel_2935/VBIAS pixel_2935/NB2 pixel_2935/AMP_IN pixel_2935/SF_IB
+ pixel_2935/PIX_OUT pixel_2935/CSA_VREF pixel
Xpixel_2924 pixel_2924/gring pixel_2924/VDD pixel_2924/GND pixel_2924/VREF pixel_2924/ROW_SEL
+ pixel_2924/NB1 pixel_2924/VBIAS pixel_2924/NB2 pixel_2924/AMP_IN pixel_2924/SF_IB
+ pixel_2924/PIX_OUT pixel_2924/CSA_VREF pixel
Xpixel_3669 pixel_3669/gring pixel_3669/VDD pixel_3669/GND pixel_3669/VREF pixel_3669/ROW_SEL
+ pixel_3669/NB1 pixel_3669/VBIAS pixel_3669/NB2 pixel_3669/AMP_IN pixel_3669/SF_IB
+ pixel_3669/PIX_OUT pixel_3669/CSA_VREF pixel
Xpixel_2979 pixel_2979/gring pixel_2979/VDD pixel_2979/GND pixel_2979/VREF pixel_2979/ROW_SEL
+ pixel_2979/NB1 pixel_2979/VBIAS pixel_2979/NB2 pixel_2979/AMP_IN pixel_2979/SF_IB
+ pixel_2979/PIX_OUT pixel_2979/CSA_VREF pixel
Xpixel_2968 pixel_2968/gring pixel_2968/VDD pixel_2968/GND pixel_2968/VREF pixel_2968/ROW_SEL
+ pixel_2968/NB1 pixel_2968/VBIAS pixel_2968/NB2 pixel_2968/AMP_IN pixel_2968/SF_IB
+ pixel_2968/PIX_OUT pixel_2968/CSA_VREF pixel
Xpixel_2957 pixel_2957/gring pixel_2957/VDD pixel_2957/GND pixel_2957/VREF pixel_2957/ROW_SEL
+ pixel_2957/NB1 pixel_2957/VBIAS pixel_2957/NB2 pixel_2957/AMP_IN pixel_2957/SF_IB
+ pixel_2957/PIX_OUT pixel_2957/CSA_VREF pixel
Xpixel_6240 pixel_6240/gring pixel_6240/VDD pixel_6240/GND pixel_6240/VREF pixel_6240/ROW_SEL
+ pixel_6240/NB1 pixel_6240/VBIAS pixel_6240/NB2 pixel_6240/AMP_IN pixel_6240/SF_IB
+ pixel_6240/PIX_OUT pixel_6240/CSA_VREF pixel
Xpixel_6251 pixel_6251/gring pixel_6251/VDD pixel_6251/GND pixel_6251/VREF pixel_6251/ROW_SEL
+ pixel_6251/NB1 pixel_6251/VBIAS pixel_6251/NB2 pixel_6251/AMP_IN pixel_6251/SF_IB
+ pixel_6251/PIX_OUT pixel_6251/CSA_VREF pixel
Xpixel_6262 pixel_6262/gring pixel_6262/VDD pixel_6262/GND pixel_6262/VREF pixel_6262/ROW_SEL
+ pixel_6262/NB1 pixel_6262/VBIAS pixel_6262/NB2 pixel_6262/AMP_IN pixel_6262/SF_IB
+ pixel_6262/PIX_OUT pixel_6262/CSA_VREF pixel
Xpixel_6273 pixel_6273/gring pixel_6273/VDD pixel_6273/GND pixel_6273/VREF pixel_6273/ROW_SEL
+ pixel_6273/NB1 pixel_6273/VBIAS pixel_6273/NB2 pixel_6273/AMP_IN pixel_6273/SF_IB
+ pixel_6273/PIX_OUT pixel_6273/CSA_VREF pixel
Xpixel_6284 pixel_6284/gring pixel_6284/VDD pixel_6284/GND pixel_6284/VREF pixel_6284/ROW_SEL
+ pixel_6284/NB1 pixel_6284/VBIAS pixel_6284/NB2 pixel_6284/AMP_IN pixel_6284/SF_IB
+ pixel_6284/PIX_OUT pixel_6284/CSA_VREF pixel
Xpixel_6295 pixel_6295/gring pixel_6295/VDD pixel_6295/GND pixel_6295/VREF pixel_6295/ROW_SEL
+ pixel_6295/NB1 pixel_6295/VBIAS pixel_6295/NB2 pixel_6295/AMP_IN pixel_6295/SF_IB
+ pixel_6295/PIX_OUT pixel_6295/CSA_VREF pixel
Xpixel_5550 pixel_5550/gring pixel_5550/VDD pixel_5550/GND pixel_5550/VREF pixel_5550/ROW_SEL
+ pixel_5550/NB1 pixel_5550/VBIAS pixel_5550/NB2 pixel_5550/AMP_IN pixel_5550/SF_IB
+ pixel_5550/PIX_OUT pixel_5550/CSA_VREF pixel
Xpixel_5561 pixel_5561/gring pixel_5561/VDD pixel_5561/GND pixel_5561/VREF pixel_5561/ROW_SEL
+ pixel_5561/NB1 pixel_5561/VBIAS pixel_5561/NB2 pixel_5561/AMP_IN pixel_5561/SF_IB
+ pixel_5561/PIX_OUT pixel_5561/CSA_VREF pixel
Xpixel_5572 pixel_5572/gring pixel_5572/VDD pixel_5572/GND pixel_5572/VREF pixel_5572/ROW_SEL
+ pixel_5572/NB1 pixel_5572/VBIAS pixel_5572/NB2 pixel_5572/AMP_IN pixel_5572/SF_IB
+ pixel_5572/PIX_OUT pixel_5572/CSA_VREF pixel
Xpixel_5583 pixel_5583/gring pixel_5583/VDD pixel_5583/GND pixel_5583/VREF pixel_5583/ROW_SEL
+ pixel_5583/NB1 pixel_5583/VBIAS pixel_5583/NB2 pixel_5583/AMP_IN pixel_5583/SF_IB
+ pixel_5583/PIX_OUT pixel_5583/CSA_VREF pixel
Xpixel_5594 pixel_5594/gring pixel_5594/VDD pixel_5594/GND pixel_5594/VREF pixel_5594/ROW_SEL
+ pixel_5594/NB1 pixel_5594/VBIAS pixel_5594/NB2 pixel_5594/AMP_IN pixel_5594/SF_IB
+ pixel_5594/PIX_OUT pixel_5594/CSA_VREF pixel
Xpixel_4860 pixel_4860/gring pixel_4860/VDD pixel_4860/GND pixel_4860/VREF pixel_4860/ROW_SEL
+ pixel_4860/NB1 pixel_4860/VBIAS pixel_4860/NB2 pixel_4860/AMP_IN pixel_4860/SF_IB
+ pixel_4860/PIX_OUT pixel_4860/CSA_VREF pixel
Xpixel_4871 pixel_4871/gring pixel_4871/VDD pixel_4871/GND pixel_4871/VREF pixel_4871/ROW_SEL
+ pixel_4871/NB1 pixel_4871/VBIAS pixel_4871/NB2 pixel_4871/AMP_IN pixel_4871/SF_IB
+ pixel_4871/PIX_OUT pixel_4871/CSA_VREF pixel
Xpixel_4882 pixel_4882/gring pixel_4882/VDD pixel_4882/GND pixel_4882/VREF pixel_4882/ROW_SEL
+ pixel_4882/NB1 pixel_4882/VBIAS pixel_4882/NB2 pixel_4882/AMP_IN pixel_4882/SF_IB
+ pixel_4882/PIX_OUT pixel_4882/CSA_VREF pixel
Xpixel_4893 pixel_4893/gring pixel_4893/VDD pixel_4893/GND pixel_4893/VREF pixel_4893/ROW_SEL
+ pixel_4893/NB1 pixel_4893/VBIAS pixel_4893/NB2 pixel_4893/AMP_IN pixel_4893/SF_IB
+ pixel_4893/PIX_OUT pixel_4893/CSA_VREF pixel
Xpixel_2209 pixel_2209/gring pixel_2209/VDD pixel_2209/GND pixel_2209/VREF pixel_2209/ROW_SEL
+ pixel_2209/NB1 pixel_2209/VBIAS pixel_2209/NB2 pixel_2209/AMP_IN pixel_2209/SF_IB
+ pixel_2209/PIX_OUT pixel_2209/CSA_VREF pixel
Xpixel_1519 pixel_1519/gring pixel_1519/VDD pixel_1519/GND pixel_1519/VREF pixel_1519/ROW_SEL
+ pixel_1519/NB1 pixel_1519/VBIAS pixel_1519/NB2 pixel_1519/AMP_IN pixel_1519/SF_IB
+ pixel_1519/PIX_OUT pixel_1519/CSA_VREF pixel
Xpixel_1508 pixel_1508/gring pixel_1508/VDD pixel_1508/GND pixel_1508/VREF pixel_1508/ROW_SEL
+ pixel_1508/NB1 pixel_1508/VBIAS pixel_1508/NB2 pixel_1508/AMP_IN pixel_1508/SF_IB
+ pixel_1508/PIX_OUT pixel_1508/CSA_VREF pixel
Xpixel_9805 pixel_9805/gring pixel_9805/VDD pixel_9805/GND pixel_9805/VREF pixel_9805/ROW_SEL
+ pixel_9805/NB1 pixel_9805/VBIAS pixel_9805/NB2 pixel_9805/AMP_IN pixel_9805/SF_IB
+ pixel_9805/PIX_OUT pixel_9805/CSA_VREF pixel
Xpixel_9838 pixel_9838/gring pixel_9838/VDD pixel_9838/GND pixel_9838/VREF pixel_9838/ROW_SEL
+ pixel_9838/NB1 pixel_9838/VBIAS pixel_9838/NB2 pixel_9838/AMP_IN pixel_9838/SF_IB
+ pixel_9838/PIX_OUT pixel_9838/CSA_VREF pixel
Xpixel_9827 pixel_9827/gring pixel_9827/VDD pixel_9827/GND pixel_9827/VREF pixel_9827/ROW_SEL
+ pixel_9827/NB1 pixel_9827/VBIAS pixel_9827/NB2 pixel_9827/AMP_IN pixel_9827/SF_IB
+ pixel_9827/PIX_OUT pixel_9827/CSA_VREF pixel
Xpixel_9816 pixel_9816/gring pixel_9816/VDD pixel_9816/GND pixel_9816/VREF pixel_9816/ROW_SEL
+ pixel_9816/NB1 pixel_9816/VBIAS pixel_9816/NB2 pixel_9816/AMP_IN pixel_9816/SF_IB
+ pixel_9816/PIX_OUT pixel_9816/CSA_VREF pixel
Xpixel_9849 pixel_9849/gring pixel_9849/VDD pixel_9849/GND pixel_9849/VREF pixel_9849/ROW_SEL
+ pixel_9849/NB1 pixel_9849/VBIAS pixel_9849/NB2 pixel_9849/AMP_IN pixel_9849/SF_IB
+ pixel_9849/PIX_OUT pixel_9849/CSA_VREF pixel
Xpixel_4101 pixel_4101/gring pixel_4101/VDD pixel_4101/GND pixel_4101/VREF pixel_4101/ROW_SEL
+ pixel_4101/NB1 pixel_4101/VBIAS pixel_4101/NB2 pixel_4101/AMP_IN pixel_4101/SF_IB
+ pixel_4101/PIX_OUT pixel_4101/CSA_VREF pixel
Xpixel_140 pixel_140/gring pixel_140/VDD pixel_140/GND pixel_140/VREF pixel_140/ROW_SEL
+ pixel_140/NB1 pixel_140/VBIAS pixel_140/NB2 pixel_140/AMP_IN pixel_140/SF_IB pixel_140/PIX_OUT
+ pixel_140/CSA_VREF pixel
Xpixel_3400 pixel_3400/gring pixel_3400/VDD pixel_3400/GND pixel_3400/VREF pixel_3400/ROW_SEL
+ pixel_3400/NB1 pixel_3400/VBIAS pixel_3400/NB2 pixel_3400/AMP_IN pixel_3400/SF_IB
+ pixel_3400/PIX_OUT pixel_3400/CSA_VREF pixel
Xpixel_4112 pixel_4112/gring pixel_4112/VDD pixel_4112/GND pixel_4112/VREF pixel_4112/ROW_SEL
+ pixel_4112/NB1 pixel_4112/VBIAS pixel_4112/NB2 pixel_4112/AMP_IN pixel_4112/SF_IB
+ pixel_4112/PIX_OUT pixel_4112/CSA_VREF pixel
Xpixel_4123 pixel_4123/gring pixel_4123/VDD pixel_4123/GND pixel_4123/VREF pixel_4123/ROW_SEL
+ pixel_4123/NB1 pixel_4123/VBIAS pixel_4123/NB2 pixel_4123/AMP_IN pixel_4123/SF_IB
+ pixel_4123/PIX_OUT pixel_4123/CSA_VREF pixel
Xpixel_4134 pixel_4134/gring pixel_4134/VDD pixel_4134/GND pixel_4134/VREF pixel_4134/ROW_SEL
+ pixel_4134/NB1 pixel_4134/VBIAS pixel_4134/NB2 pixel_4134/AMP_IN pixel_4134/SF_IB
+ pixel_4134/PIX_OUT pixel_4134/CSA_VREF pixel
Xpixel_173 pixel_173/gring pixel_173/VDD pixel_173/GND pixel_173/VREF pixel_173/ROW_SEL
+ pixel_173/NB1 pixel_173/VBIAS pixel_173/NB2 pixel_173/AMP_IN pixel_173/SF_IB pixel_173/PIX_OUT
+ pixel_173/CSA_VREF pixel
Xpixel_162 pixel_162/gring pixel_162/VDD pixel_162/GND pixel_162/VREF pixel_162/ROW_SEL
+ pixel_162/NB1 pixel_162/VBIAS pixel_162/NB2 pixel_162/AMP_IN pixel_162/SF_IB pixel_162/PIX_OUT
+ pixel_162/CSA_VREF pixel
Xpixel_151 pixel_151/gring pixel_151/VDD pixel_151/GND pixel_151/VREF pixel_151/ROW_SEL
+ pixel_151/NB1 pixel_151/VBIAS pixel_151/NB2 pixel_151/AMP_IN pixel_151/SF_IB pixel_151/PIX_OUT
+ pixel_151/CSA_VREF pixel
Xpixel_3433 pixel_3433/gring pixel_3433/VDD pixel_3433/GND pixel_3433/VREF pixel_3433/ROW_SEL
+ pixel_3433/NB1 pixel_3433/VBIAS pixel_3433/NB2 pixel_3433/AMP_IN pixel_3433/SF_IB
+ pixel_3433/PIX_OUT pixel_3433/CSA_VREF pixel
Xpixel_3422 pixel_3422/gring pixel_3422/VDD pixel_3422/GND pixel_3422/VREF pixel_3422/ROW_SEL
+ pixel_3422/NB1 pixel_3422/VBIAS pixel_3422/NB2 pixel_3422/AMP_IN pixel_3422/SF_IB
+ pixel_3422/PIX_OUT pixel_3422/CSA_VREF pixel
Xpixel_3411 pixel_3411/gring pixel_3411/VDD pixel_3411/GND pixel_3411/VREF pixel_3411/ROW_SEL
+ pixel_3411/NB1 pixel_3411/VBIAS pixel_3411/NB2 pixel_3411/AMP_IN pixel_3411/SF_IB
+ pixel_3411/PIX_OUT pixel_3411/CSA_VREF pixel
Xpixel_4145 pixel_4145/gring pixel_4145/VDD pixel_4145/GND pixel_4145/VREF pixel_4145/ROW_SEL
+ pixel_4145/NB1 pixel_4145/VBIAS pixel_4145/NB2 pixel_4145/AMP_IN pixel_4145/SF_IB
+ pixel_4145/PIX_OUT pixel_4145/CSA_VREF pixel
Xpixel_4156 pixel_4156/gring pixel_4156/VDD pixel_4156/GND pixel_4156/VREF pixel_4156/ROW_SEL
+ pixel_4156/NB1 pixel_4156/VBIAS pixel_4156/NB2 pixel_4156/AMP_IN pixel_4156/SF_IB
+ pixel_4156/PIX_OUT pixel_4156/CSA_VREF pixel
Xpixel_4167 pixel_4167/gring pixel_4167/VDD pixel_4167/GND pixel_4167/VREF pixel_4167/ROW_SEL
+ pixel_4167/NB1 pixel_4167/VBIAS pixel_4167/NB2 pixel_4167/AMP_IN pixel_4167/SF_IB
+ pixel_4167/PIX_OUT pixel_4167/CSA_VREF pixel
Xpixel_4178 pixel_4178/gring pixel_4178/VDD pixel_4178/GND pixel_4178/VREF pixel_4178/ROW_SEL
+ pixel_4178/NB1 pixel_4178/VBIAS pixel_4178/NB2 pixel_4178/AMP_IN pixel_4178/SF_IB
+ pixel_4178/PIX_OUT pixel_4178/CSA_VREF pixel
Xpixel_195 pixel_195/gring pixel_195/VDD pixel_195/GND pixel_195/VREF pixel_195/ROW_SEL
+ pixel_195/NB1 pixel_195/VBIAS pixel_195/NB2 pixel_195/AMP_IN pixel_195/SF_IB pixel_195/PIX_OUT
+ pixel_195/CSA_VREF pixel
Xpixel_184 pixel_184/gring pixel_184/VDD pixel_184/GND pixel_184/VREF pixel_184/ROW_SEL
+ pixel_184/NB1 pixel_184/VBIAS pixel_184/NB2 pixel_184/AMP_IN pixel_184/SF_IB pixel_184/PIX_OUT
+ pixel_184/CSA_VREF pixel
Xpixel_2721 pixel_2721/gring pixel_2721/VDD pixel_2721/GND pixel_2721/VREF pixel_2721/ROW_SEL
+ pixel_2721/NB1 pixel_2721/VBIAS pixel_2721/NB2 pixel_2721/AMP_IN pixel_2721/SF_IB
+ pixel_2721/PIX_OUT pixel_2721/CSA_VREF pixel
Xpixel_2710 pixel_2710/gring pixel_2710/VDD pixel_2710/GND pixel_2710/VREF pixel_2710/ROW_SEL
+ pixel_2710/NB1 pixel_2710/VBIAS pixel_2710/NB2 pixel_2710/AMP_IN pixel_2710/SF_IB
+ pixel_2710/PIX_OUT pixel_2710/CSA_VREF pixel
Xpixel_3466 pixel_3466/gring pixel_3466/VDD pixel_3466/GND pixel_3466/VREF pixel_3466/ROW_SEL
+ pixel_3466/NB1 pixel_3466/VBIAS pixel_3466/NB2 pixel_3466/AMP_IN pixel_3466/SF_IB
+ pixel_3466/PIX_OUT pixel_3466/CSA_VREF pixel
Xpixel_3455 pixel_3455/gring pixel_3455/VDD pixel_3455/GND pixel_3455/VREF pixel_3455/ROW_SEL
+ pixel_3455/NB1 pixel_3455/VBIAS pixel_3455/NB2 pixel_3455/AMP_IN pixel_3455/SF_IB
+ pixel_3455/PIX_OUT pixel_3455/CSA_VREF pixel
Xpixel_3444 pixel_3444/gring pixel_3444/VDD pixel_3444/GND pixel_3444/VREF pixel_3444/ROW_SEL
+ pixel_3444/NB1 pixel_3444/VBIAS pixel_3444/NB2 pixel_3444/AMP_IN pixel_3444/SF_IB
+ pixel_3444/PIX_OUT pixel_3444/CSA_VREF pixel
Xpixel_4189 pixel_4189/gring pixel_4189/VDD pixel_4189/GND pixel_4189/VREF pixel_4189/ROW_SEL
+ pixel_4189/NB1 pixel_4189/VBIAS pixel_4189/NB2 pixel_4189/AMP_IN pixel_4189/SF_IB
+ pixel_4189/PIX_OUT pixel_4189/CSA_VREF pixel
Xpixel_2765 pixel_2765/gring pixel_2765/VDD pixel_2765/GND pixel_2765/VREF pixel_2765/ROW_SEL
+ pixel_2765/NB1 pixel_2765/VBIAS pixel_2765/NB2 pixel_2765/AMP_IN pixel_2765/SF_IB
+ pixel_2765/PIX_OUT pixel_2765/CSA_VREF pixel
Xpixel_2754 pixel_2754/gring pixel_2754/VDD pixel_2754/GND pixel_2754/VREF pixel_2754/ROW_SEL
+ pixel_2754/NB1 pixel_2754/VBIAS pixel_2754/NB2 pixel_2754/AMP_IN pixel_2754/SF_IB
+ pixel_2754/PIX_OUT pixel_2754/CSA_VREF pixel
Xpixel_2743 pixel_2743/gring pixel_2743/VDD pixel_2743/GND pixel_2743/VREF pixel_2743/ROW_SEL
+ pixel_2743/NB1 pixel_2743/VBIAS pixel_2743/NB2 pixel_2743/AMP_IN pixel_2743/SF_IB
+ pixel_2743/PIX_OUT pixel_2743/CSA_VREF pixel
Xpixel_2732 pixel_2732/gring pixel_2732/VDD pixel_2732/GND pixel_2732/VREF pixel_2732/ROW_SEL
+ pixel_2732/NB1 pixel_2732/VBIAS pixel_2732/NB2 pixel_2732/AMP_IN pixel_2732/SF_IB
+ pixel_2732/PIX_OUT pixel_2732/CSA_VREF pixel
Xpixel_3499 pixel_3499/gring pixel_3499/VDD pixel_3499/GND pixel_3499/VREF pixel_3499/ROW_SEL
+ pixel_3499/NB1 pixel_3499/VBIAS pixel_3499/NB2 pixel_3499/AMP_IN pixel_3499/SF_IB
+ pixel_3499/PIX_OUT pixel_3499/CSA_VREF pixel
Xpixel_3488 pixel_3488/gring pixel_3488/VDD pixel_3488/GND pixel_3488/VREF pixel_3488/ROW_SEL
+ pixel_3488/NB1 pixel_3488/VBIAS pixel_3488/NB2 pixel_3488/AMP_IN pixel_3488/SF_IB
+ pixel_3488/PIX_OUT pixel_3488/CSA_VREF pixel
Xpixel_3477 pixel_3477/gring pixel_3477/VDD pixel_3477/GND pixel_3477/VREF pixel_3477/ROW_SEL
+ pixel_3477/NB1 pixel_3477/VBIAS pixel_3477/NB2 pixel_3477/AMP_IN pixel_3477/SF_IB
+ pixel_3477/PIX_OUT pixel_3477/CSA_VREF pixel
Xpixel_2798 pixel_2798/gring pixel_2798/VDD pixel_2798/GND pixel_2798/VREF pixel_2798/ROW_SEL
+ pixel_2798/NB1 pixel_2798/VBIAS pixel_2798/NB2 pixel_2798/AMP_IN pixel_2798/SF_IB
+ pixel_2798/PIX_OUT pixel_2798/CSA_VREF pixel
Xpixel_2787 pixel_2787/gring pixel_2787/VDD pixel_2787/GND pixel_2787/VREF pixel_2787/ROW_SEL
+ pixel_2787/NB1 pixel_2787/VBIAS pixel_2787/NB2 pixel_2787/AMP_IN pixel_2787/SF_IB
+ pixel_2787/PIX_OUT pixel_2787/CSA_VREF pixel
Xpixel_2776 pixel_2776/gring pixel_2776/VDD pixel_2776/GND pixel_2776/VREF pixel_2776/ROW_SEL
+ pixel_2776/NB1 pixel_2776/VBIAS pixel_2776/NB2 pixel_2776/AMP_IN pixel_2776/SF_IB
+ pixel_2776/PIX_OUT pixel_2776/CSA_VREF pixel
Xpixel_6070 pixel_6070/gring pixel_6070/VDD pixel_6070/GND pixel_6070/VREF pixel_6070/ROW_SEL
+ pixel_6070/NB1 pixel_6070/VBIAS pixel_6070/NB2 pixel_6070/AMP_IN pixel_6070/SF_IB
+ pixel_6070/PIX_OUT pixel_6070/CSA_VREF pixel
Xpixel_6081 pixel_6081/gring pixel_6081/VDD pixel_6081/GND pixel_6081/VREF pixel_6081/ROW_SEL
+ pixel_6081/NB1 pixel_6081/VBIAS pixel_6081/NB2 pixel_6081/AMP_IN pixel_6081/SF_IB
+ pixel_6081/PIX_OUT pixel_6081/CSA_VREF pixel
Xpixel_6092 pixel_6092/gring pixel_6092/VDD pixel_6092/GND pixel_6092/VREF pixel_6092/ROW_SEL
+ pixel_6092/NB1 pixel_6092/VBIAS pixel_6092/NB2 pixel_6092/AMP_IN pixel_6092/SF_IB
+ pixel_6092/PIX_OUT pixel_6092/CSA_VREF pixel
Xpixel_5380 pixel_5380/gring pixel_5380/VDD pixel_5380/GND pixel_5380/VREF pixel_5380/ROW_SEL
+ pixel_5380/NB1 pixel_5380/VBIAS pixel_5380/NB2 pixel_5380/AMP_IN pixel_5380/SF_IB
+ pixel_5380/PIX_OUT pixel_5380/CSA_VREF pixel
Xpixel_5391 pixel_5391/gring pixel_5391/VDD pixel_5391/GND pixel_5391/VREF pixel_5391/ROW_SEL
+ pixel_5391/NB1 pixel_5391/VBIAS pixel_5391/NB2 pixel_5391/AMP_IN pixel_5391/SF_IB
+ pixel_5391/PIX_OUT pixel_5391/CSA_VREF pixel
Xpixel_4690 pixel_4690/gring pixel_4690/VDD pixel_4690/GND pixel_4690/VREF pixel_4690/ROW_SEL
+ pixel_4690/NB1 pixel_4690/VBIAS pixel_4690/NB2 pixel_4690/AMP_IN pixel_4690/SF_IB
+ pixel_4690/PIX_OUT pixel_4690/CSA_VREF pixel
Xpixel_2017 pixel_2017/gring pixel_2017/VDD pixel_2017/GND pixel_2017/VREF pixel_2017/ROW_SEL
+ pixel_2017/NB1 pixel_2017/VBIAS pixel_2017/NB2 pixel_2017/AMP_IN pixel_2017/SF_IB
+ pixel_2017/PIX_OUT pixel_2017/CSA_VREF pixel
Xpixel_2006 pixel_2006/gring pixel_2006/VDD pixel_2006/GND pixel_2006/VREF pixel_2006/ROW_SEL
+ pixel_2006/NB1 pixel_2006/VBIAS pixel_2006/NB2 pixel_2006/AMP_IN pixel_2006/SF_IB
+ pixel_2006/PIX_OUT pixel_2006/CSA_VREF pixel
Xpixel_1305 pixel_1305/gring pixel_1305/VDD pixel_1305/GND pixel_1305/VREF pixel_1305/ROW_SEL
+ pixel_1305/NB1 pixel_1305/VBIAS pixel_1305/NB2 pixel_1305/AMP_IN pixel_1305/SF_IB
+ pixel_1305/PIX_OUT pixel_1305/CSA_VREF pixel
Xpixel_2039 pixel_2039/gring pixel_2039/VDD pixel_2039/GND pixel_2039/VREF pixel_2039/ROW_SEL
+ pixel_2039/NB1 pixel_2039/VBIAS pixel_2039/NB2 pixel_2039/AMP_IN pixel_2039/SF_IB
+ pixel_2039/PIX_OUT pixel_2039/CSA_VREF pixel
Xpixel_2028 pixel_2028/gring pixel_2028/VDD pixel_2028/GND pixel_2028/VREF pixel_2028/ROW_SEL
+ pixel_2028/NB1 pixel_2028/VBIAS pixel_2028/NB2 pixel_2028/AMP_IN pixel_2028/SF_IB
+ pixel_2028/PIX_OUT pixel_2028/CSA_VREF pixel
Xpixel_1349 pixel_1349/gring pixel_1349/VDD pixel_1349/GND pixel_1349/VREF pixel_1349/ROW_SEL
+ pixel_1349/NB1 pixel_1349/VBIAS pixel_1349/NB2 pixel_1349/AMP_IN pixel_1349/SF_IB
+ pixel_1349/PIX_OUT pixel_1349/CSA_VREF pixel
Xpixel_1338 pixel_1338/gring pixel_1338/VDD pixel_1338/GND pixel_1338/VREF pixel_1338/ROW_SEL
+ pixel_1338/NB1 pixel_1338/VBIAS pixel_1338/NB2 pixel_1338/AMP_IN pixel_1338/SF_IB
+ pixel_1338/PIX_OUT pixel_1338/CSA_VREF pixel
Xpixel_1327 pixel_1327/gring pixel_1327/VDD pixel_1327/GND pixel_1327/VREF pixel_1327/ROW_SEL
+ pixel_1327/NB1 pixel_1327/VBIAS pixel_1327/NB2 pixel_1327/AMP_IN pixel_1327/SF_IB
+ pixel_1327/PIX_OUT pixel_1327/CSA_VREF pixel
Xpixel_1316 pixel_1316/gring pixel_1316/VDD pixel_1316/GND pixel_1316/VREF pixel_1316/ROW_SEL
+ pixel_1316/NB1 pixel_1316/VBIAS pixel_1316/NB2 pixel_1316/AMP_IN pixel_1316/SF_IB
+ pixel_1316/PIX_OUT pixel_1316/CSA_VREF pixel
Xpixel_9602 pixel_9602/gring pixel_9602/VDD pixel_9602/GND pixel_9602/VREF pixel_9602/ROW_SEL
+ pixel_9602/NB1 pixel_9602/VBIAS pixel_9602/NB2 pixel_9602/AMP_IN pixel_9602/SF_IB
+ pixel_9602/PIX_OUT pixel_9602/CSA_VREF pixel
Xpixel_9613 pixel_9613/gring pixel_9613/VDD pixel_9613/GND pixel_9613/VREF pixel_9613/ROW_SEL
+ pixel_9613/NB1 pixel_9613/VBIAS pixel_9613/NB2 pixel_9613/AMP_IN pixel_9613/SF_IB
+ pixel_9613/PIX_OUT pixel_9613/CSA_VREF pixel
Xpixel_8912 pixel_8912/gring pixel_8912/VDD pixel_8912/GND pixel_8912/VREF pixel_8912/ROW_SEL
+ pixel_8912/NB1 pixel_8912/VBIAS pixel_8912/NB2 pixel_8912/AMP_IN pixel_8912/SF_IB
+ pixel_8912/PIX_OUT pixel_8912/CSA_VREF pixel
Xpixel_8901 pixel_8901/gring pixel_8901/VDD pixel_8901/GND pixel_8901/VREF pixel_8901/ROW_SEL
+ pixel_8901/NB1 pixel_8901/VBIAS pixel_8901/NB2 pixel_8901/AMP_IN pixel_8901/SF_IB
+ pixel_8901/PIX_OUT pixel_8901/CSA_VREF pixel
Xpixel_9624 pixel_9624/gring pixel_9624/VDD pixel_9624/GND pixel_9624/VREF pixel_9624/ROW_SEL
+ pixel_9624/NB1 pixel_9624/VBIAS pixel_9624/NB2 pixel_9624/AMP_IN pixel_9624/SF_IB
+ pixel_9624/PIX_OUT pixel_9624/CSA_VREF pixel
Xpixel_9635 pixel_9635/gring pixel_9635/VDD pixel_9635/GND pixel_9635/VREF pixel_9635/ROW_SEL
+ pixel_9635/NB1 pixel_9635/VBIAS pixel_9635/NB2 pixel_9635/AMP_IN pixel_9635/SF_IB
+ pixel_9635/PIX_OUT pixel_9635/CSA_VREF pixel
Xpixel_9646 pixel_9646/gring pixel_9646/VDD pixel_9646/GND pixel_9646/VREF pixel_9646/ROW_SEL
+ pixel_9646/NB1 pixel_9646/VBIAS pixel_9646/NB2 pixel_9646/AMP_IN pixel_9646/SF_IB
+ pixel_9646/PIX_OUT pixel_9646/CSA_VREF pixel
Xpixel_9657 pixel_9657/gring pixel_9657/VDD pixel_9657/GND pixel_9657/VREF pixel_9657/ROW_SEL
+ pixel_9657/NB1 pixel_9657/VBIAS pixel_9657/NB2 pixel_9657/AMP_IN pixel_9657/SF_IB
+ pixel_9657/PIX_OUT pixel_9657/CSA_VREF pixel
Xpixel_8945 pixel_8945/gring pixel_8945/VDD pixel_8945/GND pixel_8945/VREF pixel_8945/ROW_SEL
+ pixel_8945/NB1 pixel_8945/VBIAS pixel_8945/NB2 pixel_8945/AMP_IN pixel_8945/SF_IB
+ pixel_8945/PIX_OUT pixel_8945/CSA_VREF pixel
Xpixel_8934 pixel_8934/gring pixel_8934/VDD pixel_8934/GND pixel_8934/VREF pixel_8934/ROW_SEL
+ pixel_8934/NB1 pixel_8934/VBIAS pixel_8934/NB2 pixel_8934/AMP_IN pixel_8934/SF_IB
+ pixel_8934/PIX_OUT pixel_8934/CSA_VREF pixel
Xpixel_8923 pixel_8923/gring pixel_8923/VDD pixel_8923/GND pixel_8923/VREF pixel_8923/ROW_SEL
+ pixel_8923/NB1 pixel_8923/VBIAS pixel_8923/NB2 pixel_8923/AMP_IN pixel_8923/SF_IB
+ pixel_8923/PIX_OUT pixel_8923/CSA_VREF pixel
Xpixel_9668 pixel_9668/gring pixel_9668/VDD pixel_9668/GND pixel_9668/VREF pixel_9668/ROW_SEL
+ pixel_9668/NB1 pixel_9668/VBIAS pixel_9668/NB2 pixel_9668/AMP_IN pixel_9668/SF_IB
+ pixel_9668/PIX_OUT pixel_9668/CSA_VREF pixel
Xpixel_9679 pixel_9679/gring pixel_9679/VDD pixel_9679/GND pixel_9679/VREF pixel_9679/ROW_SEL
+ pixel_9679/NB1 pixel_9679/VBIAS pixel_9679/NB2 pixel_9679/AMP_IN pixel_9679/SF_IB
+ pixel_9679/PIX_OUT pixel_9679/CSA_VREF pixel
Xpixel_8978 pixel_8978/gring pixel_8978/VDD pixel_8978/GND pixel_8978/VREF pixel_8978/ROW_SEL
+ pixel_8978/NB1 pixel_8978/VBIAS pixel_8978/NB2 pixel_8978/AMP_IN pixel_8978/SF_IB
+ pixel_8978/PIX_OUT pixel_8978/CSA_VREF pixel
Xpixel_8967 pixel_8967/gring pixel_8967/VDD pixel_8967/GND pixel_8967/VREF pixel_8967/ROW_SEL
+ pixel_8967/NB1 pixel_8967/VBIAS pixel_8967/NB2 pixel_8967/AMP_IN pixel_8967/SF_IB
+ pixel_8967/PIX_OUT pixel_8967/CSA_VREF pixel
Xpixel_8956 pixel_8956/gring pixel_8956/VDD pixel_8956/GND pixel_8956/VREF pixel_8956/ROW_SEL
+ pixel_8956/NB1 pixel_8956/VBIAS pixel_8956/NB2 pixel_8956/AMP_IN pixel_8956/SF_IB
+ pixel_8956/PIX_OUT pixel_8956/CSA_VREF pixel
Xpixel_8989 pixel_8989/gring pixel_8989/VDD pixel_8989/GND pixel_8989/VREF pixel_8989/ROW_SEL
+ pixel_8989/NB1 pixel_8989/VBIAS pixel_8989/NB2 pixel_8989/AMP_IN pixel_8989/SF_IB
+ pixel_8989/PIX_OUT pixel_8989/CSA_VREF pixel
Xpixel_3241 pixel_3241/gring pixel_3241/VDD pixel_3241/GND pixel_3241/VREF pixel_3241/ROW_SEL
+ pixel_3241/NB1 pixel_3241/VBIAS pixel_3241/NB2 pixel_3241/AMP_IN pixel_3241/SF_IB
+ pixel_3241/PIX_OUT pixel_3241/CSA_VREF pixel
Xpixel_3230 pixel_3230/gring pixel_3230/VDD pixel_3230/GND pixel_3230/VREF pixel_3230/ROW_SEL
+ pixel_3230/NB1 pixel_3230/VBIAS pixel_3230/NB2 pixel_3230/AMP_IN pixel_3230/SF_IB
+ pixel_3230/PIX_OUT pixel_3230/CSA_VREF pixel
Xpixel_2540 pixel_2540/gring pixel_2540/VDD pixel_2540/GND pixel_2540/VREF pixel_2540/ROW_SEL
+ pixel_2540/NB1 pixel_2540/VBIAS pixel_2540/NB2 pixel_2540/AMP_IN pixel_2540/SF_IB
+ pixel_2540/PIX_OUT pixel_2540/CSA_VREF pixel
Xpixel_3274 pixel_3274/gring pixel_3274/VDD pixel_3274/GND pixel_3274/VREF pixel_3274/ROW_SEL
+ pixel_3274/NB1 pixel_3274/VBIAS pixel_3274/NB2 pixel_3274/AMP_IN pixel_3274/SF_IB
+ pixel_3274/PIX_OUT pixel_3274/CSA_VREF pixel
Xpixel_3263 pixel_3263/gring pixel_3263/VDD pixel_3263/GND pixel_3263/VREF pixel_3263/ROW_SEL
+ pixel_3263/NB1 pixel_3263/VBIAS pixel_3263/NB2 pixel_3263/AMP_IN pixel_3263/SF_IB
+ pixel_3263/PIX_OUT pixel_3263/CSA_VREF pixel
Xpixel_3252 pixel_3252/gring pixel_3252/VDD pixel_3252/GND pixel_3252/VREF pixel_3252/ROW_SEL
+ pixel_3252/NB1 pixel_3252/VBIAS pixel_3252/NB2 pixel_3252/AMP_IN pixel_3252/SF_IB
+ pixel_3252/PIX_OUT pixel_3252/CSA_VREF pixel
Xpixel_2573 pixel_2573/gring pixel_2573/VDD pixel_2573/GND pixel_2573/VREF pixel_2573/ROW_SEL
+ pixel_2573/NB1 pixel_2573/VBIAS pixel_2573/NB2 pixel_2573/AMP_IN pixel_2573/SF_IB
+ pixel_2573/PIX_OUT pixel_2573/CSA_VREF pixel
Xpixel_2562 pixel_2562/gring pixel_2562/VDD pixel_2562/GND pixel_2562/VREF pixel_2562/ROW_SEL
+ pixel_2562/NB1 pixel_2562/VBIAS pixel_2562/NB2 pixel_2562/AMP_IN pixel_2562/SF_IB
+ pixel_2562/PIX_OUT pixel_2562/CSA_VREF pixel
Xpixel_2551 pixel_2551/gring pixel_2551/VDD pixel_2551/GND pixel_2551/VREF pixel_2551/ROW_SEL
+ pixel_2551/NB1 pixel_2551/VBIAS pixel_2551/NB2 pixel_2551/AMP_IN pixel_2551/SF_IB
+ pixel_2551/PIX_OUT pixel_2551/CSA_VREF pixel
Xpixel_3296 pixel_3296/gring pixel_3296/VDD pixel_3296/GND pixel_3296/VREF pixel_3296/ROW_SEL
+ pixel_3296/NB1 pixel_3296/VBIAS pixel_3296/NB2 pixel_3296/AMP_IN pixel_3296/SF_IB
+ pixel_3296/PIX_OUT pixel_3296/CSA_VREF pixel
Xpixel_3285 pixel_3285/gring pixel_3285/VDD pixel_3285/GND pixel_3285/VREF pixel_3285/ROW_SEL
+ pixel_3285/NB1 pixel_3285/VBIAS pixel_3285/NB2 pixel_3285/AMP_IN pixel_3285/SF_IB
+ pixel_3285/PIX_OUT pixel_3285/CSA_VREF pixel
Xpixel_1861 pixel_1861/gring pixel_1861/VDD pixel_1861/GND pixel_1861/VREF pixel_1861/ROW_SEL
+ pixel_1861/NB1 pixel_1861/VBIAS pixel_1861/NB2 pixel_1861/AMP_IN pixel_1861/SF_IB
+ pixel_1861/PIX_OUT pixel_1861/CSA_VREF pixel
Xpixel_1850 pixel_1850/gring pixel_1850/VDD pixel_1850/GND pixel_1850/VREF pixel_1850/ROW_SEL
+ pixel_1850/NB1 pixel_1850/VBIAS pixel_1850/NB2 pixel_1850/AMP_IN pixel_1850/SF_IB
+ pixel_1850/PIX_OUT pixel_1850/CSA_VREF pixel
Xpixel_2595 pixel_2595/gring pixel_2595/VDD pixel_2595/GND pixel_2595/VREF pixel_2595/ROW_SEL
+ pixel_2595/NB1 pixel_2595/VBIAS pixel_2595/NB2 pixel_2595/AMP_IN pixel_2595/SF_IB
+ pixel_2595/PIX_OUT pixel_2595/CSA_VREF pixel
Xpixel_2584 pixel_2584/gring pixel_2584/VDD pixel_2584/GND pixel_2584/VREF pixel_2584/ROW_SEL
+ pixel_2584/NB1 pixel_2584/VBIAS pixel_2584/NB2 pixel_2584/AMP_IN pixel_2584/SF_IB
+ pixel_2584/PIX_OUT pixel_2584/CSA_VREF pixel
Xpixel_1894 pixel_1894/gring pixel_1894/VDD pixel_1894/GND pixel_1894/VREF pixel_1894/ROW_SEL
+ pixel_1894/NB1 pixel_1894/VBIAS pixel_1894/NB2 pixel_1894/AMP_IN pixel_1894/SF_IB
+ pixel_1894/PIX_OUT pixel_1894/CSA_VREF pixel
Xpixel_1883 pixel_1883/gring pixel_1883/VDD pixel_1883/GND pixel_1883/VREF pixel_1883/ROW_SEL
+ pixel_1883/NB1 pixel_1883/VBIAS pixel_1883/NB2 pixel_1883/AMP_IN pixel_1883/SF_IB
+ pixel_1883/PIX_OUT pixel_1883/CSA_VREF pixel
Xpixel_1872 pixel_1872/gring pixel_1872/VDD pixel_1872/GND pixel_1872/VREF pixel_1872/ROW_SEL
+ pixel_1872/NB1 pixel_1872/VBIAS pixel_1872/NB2 pixel_1872/AMP_IN pixel_1872/SF_IB
+ pixel_1872/PIX_OUT pixel_1872/CSA_VREF pixel
Xpixel_909 pixel_909/gring pixel_909/VDD pixel_909/GND pixel_909/VREF pixel_909/ROW_SEL
+ pixel_909/NB1 pixel_909/VBIAS pixel_909/NB2 pixel_909/AMP_IN pixel_909/SF_IB pixel_909/PIX_OUT
+ pixel_909/CSA_VREF pixel
Xpixel_8208 pixel_8208/gring pixel_8208/VDD pixel_8208/GND pixel_8208/VREF pixel_8208/ROW_SEL
+ pixel_8208/NB1 pixel_8208/VBIAS pixel_8208/NB2 pixel_8208/AMP_IN pixel_8208/SF_IB
+ pixel_8208/PIX_OUT pixel_8208/CSA_VREF pixel
Xpixel_8219 pixel_8219/gring pixel_8219/VDD pixel_8219/GND pixel_8219/VREF pixel_8219/ROW_SEL
+ pixel_8219/NB1 pixel_8219/VBIAS pixel_8219/NB2 pixel_8219/AMP_IN pixel_8219/SF_IB
+ pixel_8219/PIX_OUT pixel_8219/CSA_VREF pixel
Xpixel_7507 pixel_7507/gring pixel_7507/VDD pixel_7507/GND pixel_7507/VREF pixel_7507/ROW_SEL
+ pixel_7507/NB1 pixel_7507/VBIAS pixel_7507/NB2 pixel_7507/AMP_IN pixel_7507/SF_IB
+ pixel_7507/PIX_OUT pixel_7507/CSA_VREF pixel
Xpixel_7518 pixel_7518/gring pixel_7518/VDD pixel_7518/GND pixel_7518/VREF pixel_7518/ROW_SEL
+ pixel_7518/NB1 pixel_7518/VBIAS pixel_7518/NB2 pixel_7518/AMP_IN pixel_7518/SF_IB
+ pixel_7518/PIX_OUT pixel_7518/CSA_VREF pixel
Xpixel_7529 pixel_7529/gring pixel_7529/VDD pixel_7529/GND pixel_7529/VREF pixel_7529/ROW_SEL
+ pixel_7529/NB1 pixel_7529/VBIAS pixel_7529/NB2 pixel_7529/AMP_IN pixel_7529/SF_IB
+ pixel_7529/PIX_OUT pixel_7529/CSA_VREF pixel
Xpixel_6806 pixel_6806/gring pixel_6806/VDD pixel_6806/GND pixel_6806/VREF pixel_6806/ROW_SEL
+ pixel_6806/NB1 pixel_6806/VBIAS pixel_6806/NB2 pixel_6806/AMP_IN pixel_6806/SF_IB
+ pixel_6806/PIX_OUT pixel_6806/CSA_VREF pixel
Xpixel_6817 pixel_6817/gring pixel_6817/VDD pixel_6817/GND pixel_6817/VREF pixel_6817/ROW_SEL
+ pixel_6817/NB1 pixel_6817/VBIAS pixel_6817/NB2 pixel_6817/AMP_IN pixel_6817/SF_IB
+ pixel_6817/PIX_OUT pixel_6817/CSA_VREF pixel
Xpixel_6828 pixel_6828/gring pixel_6828/VDD pixel_6828/GND pixel_6828/VREF pixel_6828/ROW_SEL
+ pixel_6828/NB1 pixel_6828/VBIAS pixel_6828/NB2 pixel_6828/AMP_IN pixel_6828/SF_IB
+ pixel_6828/PIX_OUT pixel_6828/CSA_VREF pixel
Xpixel_6839 pixel_6839/gring pixel_6839/VDD pixel_6839/GND pixel_6839/VREF pixel_6839/ROW_SEL
+ pixel_6839/NB1 pixel_6839/VBIAS pixel_6839/NB2 pixel_6839/AMP_IN pixel_6839/SF_IB
+ pixel_6839/PIX_OUT pixel_6839/CSA_VREF pixel
Xpixel_1124 pixel_1124/gring pixel_1124/VDD pixel_1124/GND pixel_1124/VREF pixel_1124/ROW_SEL
+ pixel_1124/NB1 pixel_1124/VBIAS pixel_1124/NB2 pixel_1124/AMP_IN pixel_1124/SF_IB
+ pixel_1124/PIX_OUT pixel_1124/CSA_VREF pixel
Xpixel_1113 pixel_1113/gring pixel_1113/VDD pixel_1113/GND pixel_1113/VREF pixel_1113/ROW_SEL
+ pixel_1113/NB1 pixel_1113/VBIAS pixel_1113/NB2 pixel_1113/AMP_IN pixel_1113/SF_IB
+ pixel_1113/PIX_OUT pixel_1113/CSA_VREF pixel
Xpixel_1102 pixel_1102/gring pixel_1102/VDD pixel_1102/GND pixel_1102/VREF pixel_1102/ROW_SEL
+ pixel_1102/NB1 pixel_1102/VBIAS pixel_1102/NB2 pixel_1102/AMP_IN pixel_1102/SF_IB
+ pixel_1102/PIX_OUT pixel_1102/CSA_VREF pixel
Xpixel_1157 pixel_1157/gring pixel_1157/VDD pixel_1157/GND pixel_1157/VREF pixel_1157/ROW_SEL
+ pixel_1157/NB1 pixel_1157/VBIAS pixel_1157/NB2 pixel_1157/AMP_IN pixel_1157/SF_IB
+ pixel_1157/PIX_OUT pixel_1157/CSA_VREF pixel
Xpixel_1146 pixel_1146/gring pixel_1146/VDD pixel_1146/GND pixel_1146/VREF pixel_1146/ROW_SEL
+ pixel_1146/NB1 pixel_1146/VBIAS pixel_1146/NB2 pixel_1146/AMP_IN pixel_1146/SF_IB
+ pixel_1146/PIX_OUT pixel_1146/CSA_VREF pixel
Xpixel_1135 pixel_1135/gring pixel_1135/VDD pixel_1135/GND pixel_1135/VREF pixel_1135/ROW_SEL
+ pixel_1135/NB1 pixel_1135/VBIAS pixel_1135/NB2 pixel_1135/AMP_IN pixel_1135/SF_IB
+ pixel_1135/PIX_OUT pixel_1135/CSA_VREF pixel
Xpixel_1179 pixel_1179/gring pixel_1179/VDD pixel_1179/GND pixel_1179/VREF pixel_1179/ROW_SEL
+ pixel_1179/NB1 pixel_1179/VBIAS pixel_1179/NB2 pixel_1179/AMP_IN pixel_1179/SF_IB
+ pixel_1179/PIX_OUT pixel_1179/CSA_VREF pixel
Xpixel_1168 pixel_1168/gring pixel_1168/VDD pixel_1168/GND pixel_1168/VREF pixel_1168/ROW_SEL
+ pixel_1168/NB1 pixel_1168/VBIAS pixel_1168/NB2 pixel_1168/AMP_IN pixel_1168/SF_IB
+ pixel_1168/PIX_OUT pixel_1168/CSA_VREF pixel
Xpixel_9432 pixel_9432/gring pixel_9432/VDD pixel_9432/GND pixel_9432/VREF pixel_9432/ROW_SEL
+ pixel_9432/NB1 pixel_9432/VBIAS pixel_9432/NB2 pixel_9432/AMP_IN pixel_9432/SF_IB
+ pixel_9432/PIX_OUT pixel_9432/CSA_VREF pixel
Xpixel_9421 pixel_9421/gring pixel_9421/VDD pixel_9421/GND pixel_9421/VREF pixel_9421/ROW_SEL
+ pixel_9421/NB1 pixel_9421/VBIAS pixel_9421/NB2 pixel_9421/AMP_IN pixel_9421/SF_IB
+ pixel_9421/PIX_OUT pixel_9421/CSA_VREF pixel
Xpixel_9410 pixel_9410/gring pixel_9410/VDD pixel_9410/GND pixel_9410/VREF pixel_9410/ROW_SEL
+ pixel_9410/NB1 pixel_9410/VBIAS pixel_9410/NB2 pixel_9410/AMP_IN pixel_9410/SF_IB
+ pixel_9410/PIX_OUT pixel_9410/CSA_VREF pixel
Xpixel_8720 pixel_8720/gring pixel_8720/VDD pixel_8720/GND pixel_8720/VREF pixel_8720/ROW_SEL
+ pixel_8720/NB1 pixel_8720/VBIAS pixel_8720/NB2 pixel_8720/AMP_IN pixel_8720/SF_IB
+ pixel_8720/PIX_OUT pixel_8720/CSA_VREF pixel
Xpixel_9465 pixel_9465/gring pixel_9465/VDD pixel_9465/GND pixel_9465/VREF pixel_9465/ROW_SEL
+ pixel_9465/NB1 pixel_9465/VBIAS pixel_9465/NB2 pixel_9465/AMP_IN pixel_9465/SF_IB
+ pixel_9465/PIX_OUT pixel_9465/CSA_VREF pixel
Xpixel_9454 pixel_9454/gring pixel_9454/VDD pixel_9454/GND pixel_9454/VREF pixel_9454/ROW_SEL
+ pixel_9454/NB1 pixel_9454/VBIAS pixel_9454/NB2 pixel_9454/AMP_IN pixel_9454/SF_IB
+ pixel_9454/PIX_OUT pixel_9454/CSA_VREF pixel
Xpixel_9443 pixel_9443/gring pixel_9443/VDD pixel_9443/GND pixel_9443/VREF pixel_9443/ROW_SEL
+ pixel_9443/NB1 pixel_9443/VBIAS pixel_9443/NB2 pixel_9443/AMP_IN pixel_9443/SF_IB
+ pixel_9443/PIX_OUT pixel_9443/CSA_VREF pixel
Xpixel_8753 pixel_8753/gring pixel_8753/VDD pixel_8753/GND pixel_8753/VREF pixel_8753/ROW_SEL
+ pixel_8753/NB1 pixel_8753/VBIAS pixel_8753/NB2 pixel_8753/AMP_IN pixel_8753/SF_IB
+ pixel_8753/PIX_OUT pixel_8753/CSA_VREF pixel
Xpixel_8742 pixel_8742/gring pixel_8742/VDD pixel_8742/GND pixel_8742/VREF pixel_8742/ROW_SEL
+ pixel_8742/NB1 pixel_8742/VBIAS pixel_8742/NB2 pixel_8742/AMP_IN pixel_8742/SF_IB
+ pixel_8742/PIX_OUT pixel_8742/CSA_VREF pixel
Xpixel_8731 pixel_8731/gring pixel_8731/VDD pixel_8731/GND pixel_8731/VREF pixel_8731/ROW_SEL
+ pixel_8731/NB1 pixel_8731/VBIAS pixel_8731/NB2 pixel_8731/AMP_IN pixel_8731/SF_IB
+ pixel_8731/PIX_OUT pixel_8731/CSA_VREF pixel
Xpixel_9498 pixel_9498/gring pixel_9498/VDD pixel_9498/GND pixel_9498/VREF pixel_9498/ROW_SEL
+ pixel_9498/NB1 pixel_9498/VBIAS pixel_9498/NB2 pixel_9498/AMP_IN pixel_9498/SF_IB
+ pixel_9498/PIX_OUT pixel_9498/CSA_VREF pixel
Xpixel_9487 pixel_9487/gring pixel_9487/VDD pixel_9487/GND pixel_9487/VREF pixel_9487/ROW_SEL
+ pixel_9487/NB1 pixel_9487/VBIAS pixel_9487/NB2 pixel_9487/AMP_IN pixel_9487/SF_IB
+ pixel_9487/PIX_OUT pixel_9487/CSA_VREF pixel
Xpixel_9476 pixel_9476/gring pixel_9476/VDD pixel_9476/GND pixel_9476/VREF pixel_9476/ROW_SEL
+ pixel_9476/NB1 pixel_9476/VBIAS pixel_9476/NB2 pixel_9476/AMP_IN pixel_9476/SF_IB
+ pixel_9476/PIX_OUT pixel_9476/CSA_VREF pixel
Xpixel_8797 pixel_8797/gring pixel_8797/VDD pixel_8797/GND pixel_8797/VREF pixel_8797/ROW_SEL
+ pixel_8797/NB1 pixel_8797/VBIAS pixel_8797/NB2 pixel_8797/AMP_IN pixel_8797/SF_IB
+ pixel_8797/PIX_OUT pixel_8797/CSA_VREF pixel
Xpixel_8786 pixel_8786/gring pixel_8786/VDD pixel_8786/GND pixel_8786/VREF pixel_8786/ROW_SEL
+ pixel_8786/NB1 pixel_8786/VBIAS pixel_8786/NB2 pixel_8786/AMP_IN pixel_8786/SF_IB
+ pixel_8786/PIX_OUT pixel_8786/CSA_VREF pixel
Xpixel_8775 pixel_8775/gring pixel_8775/VDD pixel_8775/GND pixel_8775/VREF pixel_8775/ROW_SEL
+ pixel_8775/NB1 pixel_8775/VBIAS pixel_8775/NB2 pixel_8775/AMP_IN pixel_8775/SF_IB
+ pixel_8775/PIX_OUT pixel_8775/CSA_VREF pixel
Xpixel_8764 pixel_8764/gring pixel_8764/VDD pixel_8764/GND pixel_8764/VREF pixel_8764/ROW_SEL
+ pixel_8764/NB1 pixel_8764/VBIAS pixel_8764/NB2 pixel_8764/AMP_IN pixel_8764/SF_IB
+ pixel_8764/PIX_OUT pixel_8764/CSA_VREF pixel
Xpixel_3093 pixel_3093/gring pixel_3093/VDD pixel_3093/GND pixel_3093/VREF pixel_3093/ROW_SEL
+ pixel_3093/NB1 pixel_3093/VBIAS pixel_3093/NB2 pixel_3093/AMP_IN pixel_3093/SF_IB
+ pixel_3093/PIX_OUT pixel_3093/CSA_VREF pixel
Xpixel_3082 pixel_3082/gring pixel_3082/VDD pixel_3082/GND pixel_3082/VREF pixel_3082/ROW_SEL
+ pixel_3082/NB1 pixel_3082/VBIAS pixel_3082/NB2 pixel_3082/AMP_IN pixel_3082/SF_IB
+ pixel_3082/PIX_OUT pixel_3082/CSA_VREF pixel
Xpixel_3071 pixel_3071/gring pixel_3071/VDD pixel_3071/GND pixel_3071/VREF pixel_3071/ROW_SEL
+ pixel_3071/NB1 pixel_3071/VBIAS pixel_3071/NB2 pixel_3071/AMP_IN pixel_3071/SF_IB
+ pixel_3071/PIX_OUT pixel_3071/CSA_VREF pixel
Xpixel_3060 pixel_3060/gring pixel_3060/VDD pixel_3060/GND pixel_3060/VREF pixel_3060/ROW_SEL
+ pixel_3060/NB1 pixel_3060/VBIAS pixel_3060/NB2 pixel_3060/AMP_IN pixel_3060/SF_IB
+ pixel_3060/PIX_OUT pixel_3060/CSA_VREF pixel
Xpixel_2381 pixel_2381/gring pixel_2381/VDD pixel_2381/GND pixel_2381/VREF pixel_2381/ROW_SEL
+ pixel_2381/NB1 pixel_2381/VBIAS pixel_2381/NB2 pixel_2381/AMP_IN pixel_2381/SF_IB
+ pixel_2381/PIX_OUT pixel_2381/CSA_VREF pixel
Xpixel_2370 pixel_2370/gring pixel_2370/VDD pixel_2370/GND pixel_2370/VREF pixel_2370/ROW_SEL
+ pixel_2370/NB1 pixel_2370/VBIAS pixel_2370/NB2 pixel_2370/AMP_IN pixel_2370/SF_IB
+ pixel_2370/PIX_OUT pixel_2370/CSA_VREF pixel
Xpixel_2392 pixel_2392/gring pixel_2392/VDD pixel_2392/GND pixel_2392/VREF pixel_2392/ROW_SEL
+ pixel_2392/NB1 pixel_2392/VBIAS pixel_2392/NB2 pixel_2392/AMP_IN pixel_2392/SF_IB
+ pixel_2392/PIX_OUT pixel_2392/CSA_VREF pixel
Xpixel_1691 pixel_1691/gring pixel_1691/VDD pixel_1691/GND pixel_1691/VREF pixel_1691/ROW_SEL
+ pixel_1691/NB1 pixel_1691/VBIAS pixel_1691/NB2 pixel_1691/AMP_IN pixel_1691/SF_IB
+ pixel_1691/PIX_OUT pixel_1691/CSA_VREF pixel
Xpixel_1680 pixel_1680/gring pixel_1680/VDD pixel_1680/GND pixel_1680/VREF pixel_1680/ROW_SEL
+ pixel_1680/NB1 pixel_1680/VBIAS pixel_1680/NB2 pixel_1680/AMP_IN pixel_1680/SF_IB
+ pixel_1680/PIX_OUT pixel_1680/CSA_VREF pixel
Xpixel_706 pixel_706/gring pixel_706/VDD pixel_706/GND pixel_706/VREF pixel_706/ROW_SEL
+ pixel_706/NB1 pixel_706/VBIAS pixel_706/NB2 pixel_706/AMP_IN pixel_706/SF_IB pixel_706/PIX_OUT
+ pixel_706/CSA_VREF pixel
Xpixel_739 pixel_739/gring pixel_739/VDD pixel_739/GND pixel_739/VREF pixel_739/ROW_SEL
+ pixel_739/NB1 pixel_739/VBIAS pixel_739/NB2 pixel_739/AMP_IN pixel_739/SF_IB pixel_739/PIX_OUT
+ pixel_739/CSA_VREF pixel
Xpixel_728 pixel_728/gring pixel_728/VDD pixel_728/GND pixel_728/VREF pixel_728/ROW_SEL
+ pixel_728/NB1 pixel_728/VBIAS pixel_728/NB2 pixel_728/AMP_IN pixel_728/SF_IB pixel_728/PIX_OUT
+ pixel_728/CSA_VREF pixel
Xpixel_717 pixel_717/gring pixel_717/VDD pixel_717/GND pixel_717/VREF pixel_717/ROW_SEL
+ pixel_717/NB1 pixel_717/VBIAS pixel_717/NB2 pixel_717/AMP_IN pixel_717/SF_IB pixel_717/PIX_OUT
+ pixel_717/CSA_VREF pixel
Xpixel_8005 pixel_8005/gring pixel_8005/VDD pixel_8005/GND pixel_8005/VREF pixel_8005/ROW_SEL
+ pixel_8005/NB1 pixel_8005/VBIAS pixel_8005/NB2 pixel_8005/AMP_IN pixel_8005/SF_IB
+ pixel_8005/PIX_OUT pixel_8005/CSA_VREF pixel
Xpixel_8016 pixel_8016/gring pixel_8016/VDD pixel_8016/GND pixel_8016/VREF pixel_8016/ROW_SEL
+ pixel_8016/NB1 pixel_8016/VBIAS pixel_8016/NB2 pixel_8016/AMP_IN pixel_8016/SF_IB
+ pixel_8016/PIX_OUT pixel_8016/CSA_VREF pixel
Xpixel_8027 pixel_8027/gring pixel_8027/VDD pixel_8027/GND pixel_8027/VREF pixel_8027/ROW_SEL
+ pixel_8027/NB1 pixel_8027/VBIAS pixel_8027/NB2 pixel_8027/AMP_IN pixel_8027/SF_IB
+ pixel_8027/PIX_OUT pixel_8027/CSA_VREF pixel
Xpixel_8038 pixel_8038/gring pixel_8038/VDD pixel_8038/GND pixel_8038/VREF pixel_8038/ROW_SEL
+ pixel_8038/NB1 pixel_8038/VBIAS pixel_8038/NB2 pixel_8038/AMP_IN pixel_8038/SF_IB
+ pixel_8038/PIX_OUT pixel_8038/CSA_VREF pixel
Xpixel_8049 pixel_8049/gring pixel_8049/VDD pixel_8049/GND pixel_8049/VREF pixel_8049/ROW_SEL
+ pixel_8049/NB1 pixel_8049/VBIAS pixel_8049/NB2 pixel_8049/AMP_IN pixel_8049/SF_IB
+ pixel_8049/PIX_OUT pixel_8049/CSA_VREF pixel
Xpixel_7304 pixel_7304/gring pixel_7304/VDD pixel_7304/GND pixel_7304/VREF pixel_7304/ROW_SEL
+ pixel_7304/NB1 pixel_7304/VBIAS pixel_7304/NB2 pixel_7304/AMP_IN pixel_7304/SF_IB
+ pixel_7304/PIX_OUT pixel_7304/CSA_VREF pixel
Xpixel_7315 pixel_7315/gring pixel_7315/VDD pixel_7315/GND pixel_7315/VREF pixel_7315/ROW_SEL
+ pixel_7315/NB1 pixel_7315/VBIAS pixel_7315/NB2 pixel_7315/AMP_IN pixel_7315/SF_IB
+ pixel_7315/PIX_OUT pixel_7315/CSA_VREF pixel
Xpixel_7326 pixel_7326/gring pixel_7326/VDD pixel_7326/GND pixel_7326/VREF pixel_7326/ROW_SEL
+ pixel_7326/NB1 pixel_7326/VBIAS pixel_7326/NB2 pixel_7326/AMP_IN pixel_7326/SF_IB
+ pixel_7326/PIX_OUT pixel_7326/CSA_VREF pixel
Xpixel_7337 pixel_7337/gring pixel_7337/VDD pixel_7337/GND pixel_7337/VREF pixel_7337/ROW_SEL
+ pixel_7337/NB1 pixel_7337/VBIAS pixel_7337/NB2 pixel_7337/AMP_IN pixel_7337/SF_IB
+ pixel_7337/PIX_OUT pixel_7337/CSA_VREF pixel
Xpixel_7348 pixel_7348/gring pixel_7348/VDD pixel_7348/GND pixel_7348/VREF pixel_7348/ROW_SEL
+ pixel_7348/NB1 pixel_7348/VBIAS pixel_7348/NB2 pixel_7348/AMP_IN pixel_7348/SF_IB
+ pixel_7348/PIX_OUT pixel_7348/CSA_VREF pixel
Xpixel_6603 pixel_6603/gring pixel_6603/VDD pixel_6603/GND pixel_6603/VREF pixel_6603/ROW_SEL
+ pixel_6603/NB1 pixel_6603/VBIAS pixel_6603/NB2 pixel_6603/AMP_IN pixel_6603/SF_IB
+ pixel_6603/PIX_OUT pixel_6603/CSA_VREF pixel
Xpixel_7359 pixel_7359/gring pixel_7359/VDD pixel_7359/GND pixel_7359/VREF pixel_7359/ROW_SEL
+ pixel_7359/NB1 pixel_7359/VBIAS pixel_7359/NB2 pixel_7359/AMP_IN pixel_7359/SF_IB
+ pixel_7359/PIX_OUT pixel_7359/CSA_VREF pixel
Xpixel_6614 pixel_6614/gring pixel_6614/VDD pixel_6614/GND pixel_6614/VREF pixel_6614/ROW_SEL
+ pixel_6614/NB1 pixel_6614/VBIAS pixel_6614/NB2 pixel_6614/AMP_IN pixel_6614/SF_IB
+ pixel_6614/PIX_OUT pixel_6614/CSA_VREF pixel
Xpixel_6625 pixel_6625/gring pixel_6625/VDD pixel_6625/GND pixel_6625/VREF pixel_6625/ROW_SEL
+ pixel_6625/NB1 pixel_6625/VBIAS pixel_6625/NB2 pixel_6625/AMP_IN pixel_6625/SF_IB
+ pixel_6625/PIX_OUT pixel_6625/CSA_VREF pixel
Xpixel_6636 pixel_6636/gring pixel_6636/VDD pixel_6636/GND pixel_6636/VREF pixel_6636/ROW_SEL
+ pixel_6636/NB1 pixel_6636/VBIAS pixel_6636/NB2 pixel_6636/AMP_IN pixel_6636/SF_IB
+ pixel_6636/PIX_OUT pixel_6636/CSA_VREF pixel
Xpixel_6647 pixel_6647/gring pixel_6647/VDD pixel_6647/GND pixel_6647/VREF pixel_6647/ROW_SEL
+ pixel_6647/NB1 pixel_6647/VBIAS pixel_6647/NB2 pixel_6647/AMP_IN pixel_6647/SF_IB
+ pixel_6647/PIX_OUT pixel_6647/CSA_VREF pixel
Xpixel_6658 pixel_6658/gring pixel_6658/VDD pixel_6658/GND pixel_6658/VREF pixel_6658/ROW_SEL
+ pixel_6658/NB1 pixel_6658/VBIAS pixel_6658/NB2 pixel_6658/AMP_IN pixel_6658/SF_IB
+ pixel_6658/PIX_OUT pixel_6658/CSA_VREF pixel
Xpixel_6669 pixel_6669/gring pixel_6669/VDD pixel_6669/GND pixel_6669/VREF pixel_6669/ROW_SEL
+ pixel_6669/NB1 pixel_6669/VBIAS pixel_6669/NB2 pixel_6669/AMP_IN pixel_6669/SF_IB
+ pixel_6669/PIX_OUT pixel_6669/CSA_VREF pixel
Xpixel_5902 pixel_5902/gring pixel_5902/VDD pixel_5902/GND pixel_5902/VREF pixel_5902/ROW_SEL
+ pixel_5902/NB1 pixel_5902/VBIAS pixel_5902/NB2 pixel_5902/AMP_IN pixel_5902/SF_IB
+ pixel_5902/PIX_OUT pixel_5902/CSA_VREF pixel
Xpixel_5913 pixel_5913/gring pixel_5913/VDD pixel_5913/GND pixel_5913/VREF pixel_5913/ROW_SEL
+ pixel_5913/NB1 pixel_5913/VBIAS pixel_5913/NB2 pixel_5913/AMP_IN pixel_5913/SF_IB
+ pixel_5913/PIX_OUT pixel_5913/CSA_VREF pixel
Xpixel_5924 pixel_5924/gring pixel_5924/VDD pixel_5924/GND pixel_5924/VREF pixel_5924/ROW_SEL
+ pixel_5924/NB1 pixel_5924/VBIAS pixel_5924/NB2 pixel_5924/AMP_IN pixel_5924/SF_IB
+ pixel_5924/PIX_OUT pixel_5924/CSA_VREF pixel
Xpixel_5935 pixel_5935/gring pixel_5935/VDD pixel_5935/GND pixel_5935/VREF pixel_5935/ROW_SEL
+ pixel_5935/NB1 pixel_5935/VBIAS pixel_5935/NB2 pixel_5935/AMP_IN pixel_5935/SF_IB
+ pixel_5935/PIX_OUT pixel_5935/CSA_VREF pixel
Xpixel_5946 pixel_5946/gring pixel_5946/VDD pixel_5946/GND pixel_5946/VREF pixel_5946/ROW_SEL
+ pixel_5946/NB1 pixel_5946/VBIAS pixel_5946/NB2 pixel_5946/AMP_IN pixel_5946/SF_IB
+ pixel_5946/PIX_OUT pixel_5946/CSA_VREF pixel
Xpixel_5957 pixel_5957/gring pixel_5957/VDD pixel_5957/GND pixel_5957/VREF pixel_5957/ROW_SEL
+ pixel_5957/NB1 pixel_5957/VBIAS pixel_5957/NB2 pixel_5957/AMP_IN pixel_5957/SF_IB
+ pixel_5957/PIX_OUT pixel_5957/CSA_VREF pixel
Xpixel_5968 pixel_5968/gring pixel_5968/VDD pixel_5968/GND pixel_5968/VREF pixel_5968/ROW_SEL
+ pixel_5968/NB1 pixel_5968/VBIAS pixel_5968/NB2 pixel_5968/AMP_IN pixel_5968/SF_IB
+ pixel_5968/PIX_OUT pixel_5968/CSA_VREF pixel
Xpixel_5979 pixel_5979/gring pixel_5979/VDD pixel_5979/GND pixel_5979/VREF pixel_5979/ROW_SEL
+ pixel_5979/NB1 pixel_5979/VBIAS pixel_5979/NB2 pixel_5979/AMP_IN pixel_5979/SF_IB
+ pixel_5979/PIX_OUT pixel_5979/CSA_VREF pixel
Xpixel_9240 pixel_9240/gring pixel_9240/VDD pixel_9240/GND pixel_9240/VREF pixel_9240/ROW_SEL
+ pixel_9240/NB1 pixel_9240/VBIAS pixel_9240/NB2 pixel_9240/AMP_IN pixel_9240/SF_IB
+ pixel_9240/PIX_OUT pixel_9240/CSA_VREF pixel
X0 PIX_OUT83 COL_SEL[83] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X1 PIX_OUT79 COL_SEL[79] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X2 PIX_OUT75 COL_SEL[75] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X3 PIX_OUT71 COL_SEL[71] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X4 PIX_OUT67 COL_SEL[67] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X5 PIX_OUT26 COL_SEL[26] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X6 PIX_OUT64 COL_SEL[64] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X7 PIX_OUT22 COL_SEL[22] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X8 PIX_OUT18 COL_SEL[18] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X9 PIX_OUT60 COL_SEL[60] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X10 PIX_OUT14 COL_SEL[14] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X11 PIX_OUT10 COL_SEL[10] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X12 PIX_OUT86 COL_SEL[86] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X13 PIX_OUT82 COL_SEL[82] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X14 PIX_OUT78 COL_SEL[78] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X15 PIX_OUT74 COL_SEL[74] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X16 PIX_OUT70 COL_SEL[70] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X17 PIX_OUT33 COL_SEL[33] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X18 PIX_OUT29 COL_SEL[29] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X19 PIX_OUT25 COL_SEL[25] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X20 PIX_OUT21 COL_SEL[21] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X21 PIX_OUT17 COL_SEL[17] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X22 PIX_OUT93 COL_SEL[93] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X23 PIX_OUT89 COL_SEL[89] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X24 PIX_OUT85 COL_SEL[85] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X25 PIX_OUT81 COL_SEL[81] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X26 PIX_OUT77 COL_SEL[77] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X27 PIX_OUT36 COL_SEL[36] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X28 PIX_OUT32 COL_SEL[32] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X29 PIX_OUT28 COL_SEL[28] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X30 PIX_OUT24 COL_SEL[24] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X31 PIX_OUT20 COL_SEL[20] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X32 PIX_OUT3 COL_SEL[3] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X33 PIX_OUT96 COL_SEL[96] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X34 PIX_OUT92 COL_SEL[92] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X35 PIX_OUT88 COL_SEL[88] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X36 PIX_OUT84 COL_SEL[84] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X37 PIX_OUT80 COL_SEL[80] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X38 PIX_OUT43 COL_SEL[43] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X39 PIX_OUT0 COL_SEL[0] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X40 PIX_OUT39 COL_SEL[39] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X41 PIX_OUT35 COL_SEL[35] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X42 PIX_OUT31 COL_SEL[31] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X43 PIX_OUT27 COL_SEL[27] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X44 PIX_OUT2 COL_SEL[2] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X45 PIX_OUT99 COL_SEL[99] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X46 PIX_OUT95 COL_SEL[95] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X47 PIX_OUT91 COL_SEL[91] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X48 PIX_OUT87 COL_SEL[87] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X49 PIX_OUT46 COL_SEL[46] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X50 PIX_OUT42 COL_SEL[42] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X51 PIX_OUT38 COL_SEL[38] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X52 PIX_OUT34 COL_SEL[34] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X53 PIX_OUT30 COL_SEL[30] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X54 PIX_OUT1 COL_SEL[1] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X55 PIX_OUT98 COL_SEL[98] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X56 PIX_OUT94 COL_SEL[94] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X57 PIX_OUT90 COL_SEL[90] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X58 PIX_OUT53 COL_SEL[53] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X59 PIX_OUT49 COL_SEL[49] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X60 PIX_OUT45 COL_SEL[45] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X61 PIX_OUT41 COL_SEL[41] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X62 PIX_OUT37 COL_SEL[37] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X63 PIX_OUT97 COL_SEL[97] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X64 PIX_OUT56 COL_SEL[56] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X65 PIX_OUT52 COL_SEL[52] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X66 PIX_OUT6 COL_SEL[6] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X67 PIX_OUT48 COL_SEL[48] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X68 PIX_OUT44 COL_SEL[44] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X69 PIX_OUT40 COL_SEL[40] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X70 PIX_OUT63 COL_SEL[63] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X71 PIX_OUT59 COL_SEL[59] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X72 PIX_OUT55 COL_SEL[55] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X73 PIX_OUT13 COL_SEL[13] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X74 PIX_OUT9 COL_SEL[9] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X75 PIX_OUT51 COL_SEL[51] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X76 PIX_OUT5 COL_SEL[5] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X77 PIX_OUT47 COL_SEL[47] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X78 PIX_OUT73 COL_SEL[73] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X79 PIX_OUT69 COL_SEL[69] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X80 PIX_OUT66 COL_SEL[66] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X81 PIX_OUT62 COL_SEL[62] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X82 PIX_OUT16 COL_SEL[16] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X83 PIX_OUT12 COL_SEL[12] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X84 PIX_OUT58 COL_SEL[58] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X85 PIX_OUT54 COL_SEL[54] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X86 PIX_OUT8 COL_SEL[8] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X87 PIX_OUT50 COL_SEL[50] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X88 PIX_OUT4 COL_SEL[4] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X89 PIX_OUT76 COL_SEL[76] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X90 PIX_OUT72 COL_SEL[72] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X91 PIX_OUT68 COL_SEL[68] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X92 PIX_OUT23 COL_SEL[23] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X93 PIX_OUT19 COL_SEL[19] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X94 PIX_OUT65 COL_SEL[65] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X95 PIX_OUT61 COL_SEL[61] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X96 PIX_OUT15 COL_SEL[15] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X97 PIX_OUT11 COL_SEL[11] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X98 PIX_OUT57 COL_SEL[57] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X99 PIX_OUT7 COL_SEL[7] ARRAY_OUT VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
.ends

