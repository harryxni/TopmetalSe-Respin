magic
tech sky130A
magscale 1 2
timestamp 1758232856
<< metal1 >>
rect 338026 591829 338426 591848
rect 333731 591539 338103 591829
rect 338026 591485 338103 591539
rect 338393 591485 338426 591829
rect 338026 591478 338426 591485
rect 257406 590510 257726 590516
rect 287844 590510 288164 590516
rect 257726 590190 287844 590510
rect 257406 590184 257726 590190
rect 287844 590184 288164 590190
rect 307105 590319 307275 590325
rect 307275 590149 307822 590319
rect 307105 590143 307275 590149
rect 338103 588877 338393 591478
rect 338097 588587 338103 588877
rect 338393 588587 338399 588877
rect 338103 588035 338393 588587
rect 338103 587739 338393 587745
rect 255190 510813 258688 510819
rect 148121 506934 255190 510813
rect 257054 507309 258688 507315
rect 148121 443358 151619 506934
rect 255190 506928 257054 506934
rect 306098 473946 310898 473952
rect 290828 473346 291354 473400
rect 288563 472816 288569 473346
rect 289099 473072 290878 473346
rect 291278 473072 291354 473346
rect 289099 473034 291354 473072
rect 289099 472816 291278 473034
rect 290878 469740 291518 472036
rect 296870 471945 306098 473946
rect 296158 471575 297401 471945
rect 297771 471575 306098 471945
rect 290872 469712 291546 469740
rect 290872 469346 290878 469712
rect 290872 469072 291278 469346
rect 291518 469072 291546 469712
rect 296870 469146 306098 471575
rect 306098 469140 310898 469146
rect 290872 469050 291546 469072
rect 149102 437806 149422 443358
rect 149096 437486 149102 437806
rect 149422 437486 149428 437806
rect 149102 435938 149422 437486
rect 8362 261315 8493 261350
rect 8362 261245 8387 261315
rect 8457 261245 10882 261315
rect 8362 261225 8493 261245
rect 495812 140997 496688 141003
rect 488766 140867 489382 140873
rect 489382 140251 493474 140867
rect 494090 140251 495812 140867
rect 488766 140245 489382 140251
rect 496688 140121 501754 140997
rect 502630 140121 502636 140997
rect 495812 140115 496688 140121
rect 461961 139194 462131 139200
rect 462131 139024 462371 139194
rect 461961 139018 462131 139024
<< via1 >>
rect 338103 591485 338393 591829
rect 257406 590190 257726 590510
rect 287844 590190 288164 590510
rect 307105 590149 307275 590319
rect 338103 588587 338393 588877
rect 338103 587745 338393 588035
rect 255190 507315 258688 510813
rect 255190 506934 257054 507315
rect 288569 472816 289099 473346
rect 290878 473072 291278 473346
rect 297401 471575 297771 471945
rect 290878 469346 291518 469712
rect 291278 469072 291518 469346
rect 306098 469146 310898 473946
rect 149102 437486 149422 437806
rect 8387 261245 8457 261315
rect 488766 140251 489382 140867
rect 493474 140251 494090 140867
rect 495812 140121 496688 140997
rect 501754 140121 502630 140997
rect 461961 139024 462131 139194
<< metal2 >>
rect 306258 599752 344106 600184
rect 274222 595025 276722 595030
rect 274218 592535 274227 595025
rect 276717 593088 276726 595025
rect 306439 593349 306509 599752
rect 289209 593279 306509 593349
rect 307105 594295 308461 594465
rect 308631 594295 308640 594465
rect 275898 592535 276506 592538
rect 276717 592535 279366 593088
rect 274222 592520 279366 592535
rect 288821 592520 289156 592524
rect 274222 592515 289161 592520
rect 274222 592180 288821 592515
rect 289156 592180 289161 592515
rect 298334 592459 298404 593279
rect 274222 592175 289161 592180
rect 274222 590588 279366 592175
rect 288821 592171 289156 592175
rect 288674 591491 289634 591502
rect 291314 591491 291424 592202
rect 288674 591381 291424 591491
rect 257406 590510 257726 590519
rect 287849 590510 288159 590514
rect 257400 590190 257406 590510
rect 257726 590190 257732 590510
rect 287838 590190 287844 590510
rect 288164 590190 288170 590510
rect 257406 590181 257726 590190
rect 287849 590186 288159 590190
rect 288674 588421 289634 591381
rect 307105 590319 307275 594295
rect 338026 591829 338426 591848
rect 338026 591485 338103 591829
rect 338393 591485 338426 591829
rect 338026 591478 338426 591485
rect 338103 591331 338393 591478
rect 338103 590744 338393 591041
rect 338103 590655 338108 590744
rect 338388 590655 338393 590744
rect 338099 590365 338103 590554
rect 338393 590365 338397 590554
rect 270797 587584 270806 588421
rect 271643 587584 289634 588421
rect 291314 587871 291404 590312
rect 307099 590149 307105 590319
rect 307275 590149 307281 590319
rect 338099 590274 338108 590365
rect 338388 590274 338397 590365
rect 338103 588877 338393 590274
rect 338103 588035 338393 588587
rect 288674 587574 289634 587584
rect 289849 587781 291404 587871
rect 234629 587111 234719 587120
rect 289849 587111 289939 587781
rect 338097 587745 338103 588035
rect 338393 587745 338399 588035
rect 234719 587021 289939 587111
rect 234629 587012 234719 587021
rect 236793 586799 236883 586808
rect 291983 586799 292073 587312
rect 236883 586709 292073 586799
rect 338103 586744 338393 587745
rect 236793 586700 236883 586709
rect 338099 586655 338108 586744
rect 338388 586655 338397 586744
rect 338099 586464 338103 586655
rect 338393 586464 338397 586655
rect 338103 586356 338393 586365
rect 240447 584312 240537 584321
rect 240537 584222 292101 584312
rect 240447 584213 240537 584222
rect 306322 583870 308492 584118
rect 265881 578736 265890 579201
rect 266355 579114 286811 579201
rect 266355 578822 286432 579114
rect 286724 578822 286811 579114
rect 266355 578736 286811 578822
rect 243956 571852 244176 571861
rect 291821 571852 292031 571856
rect 244176 571847 292036 571852
rect 244176 571637 291821 571847
rect 292031 571637 292036 571847
rect 244176 571632 292036 571637
rect 243956 571623 244176 571632
rect 291821 571628 292031 571632
rect 291888 570930 292326 571124
rect 247634 570925 292326 570930
rect 247634 570715 291977 570925
rect 292187 570715 292326 570925
rect 247634 570710 292326 570715
rect 249200 570363 249420 570710
rect 291888 570506 292326 570710
rect 249200 570274 249279 570363
rect 249381 570274 249420 570363
rect 249200 570045 249420 570054
rect 292245 568142 292455 568146
rect 229961 567922 229970 568142
rect 230190 568137 292460 568142
rect 230190 567927 292245 568137
rect 292455 567927 292460 568137
rect 230190 567922 292460 567927
rect 292245 567918 292455 567922
rect 255190 532282 258688 532287
rect 255186 528794 255195 532282
rect 258683 528794 258692 532282
rect 255190 528682 258688 528794
rect 257054 526818 258688 528682
rect 255190 510813 258688 526818
rect 255184 506934 255190 510813
rect 258688 507315 258694 510813
rect 257054 506934 257060 507315
rect 293564 478336 293674 583267
rect 306322 581858 306570 583870
rect 303290 581610 306570 581858
rect 308191 579849 308912 580019
rect 308191 575685 308361 579849
rect 332634 575685 332643 575847
rect 308191 575515 332643 575685
rect 332634 575353 332643 575515
rect 333137 575353 333146 575847
rect 343674 486512 344106 599752
rect 347632 585517 347792 585521
rect 461812 585517 461821 585645
rect 347627 585512 461821 585517
rect 347627 585352 347632 585512
rect 347792 585352 461821 585512
rect 347627 585347 461821 585352
rect 347632 585343 347792 585347
rect 461812 585219 461821 585347
rect 462247 585219 462256 585645
rect 371804 575847 372288 575851
rect 371799 575842 444605 575847
rect 371799 575358 371804 575842
rect 372288 575358 444605 575842
rect 371799 575353 444605 575358
rect 445099 575353 445333 575847
rect 371804 575349 372288 575353
rect 343674 485880 344106 486080
rect 415673 478336 416703 478340
rect 152395 477296 152404 478336
rect 153444 478331 416708 478336
rect 153444 477925 415673 478331
rect 153444 477735 291713 477925
rect 291903 477735 415673 477925
rect 153444 477301 415673 477735
rect 416703 477301 416708 478331
rect 153444 477296 416708 477301
rect 415673 477292 416703 477296
rect 343674 475891 344106 475896
rect 343670 475469 343679 475891
rect 344101 475469 344110 475891
rect 343674 475103 344106 475469
rect 153674 475079 422144 475103
rect 431840 475079 432768 475083
rect 153674 475074 432773 475079
rect 153674 474979 431840 475074
rect 153674 474789 292223 474979
rect 292413 474789 431840 474979
rect 153674 474666 431840 474789
rect 153737 472745 154377 474666
rect 343674 474096 344106 474666
rect 417287 474146 431840 474666
rect 432768 474146 432773 475074
rect 417287 474141 432773 474146
rect 431840 474137 432768 474141
rect 309343 473946 314133 473950
rect 288569 473346 289099 473352
rect 290852 473346 291308 473386
rect 288560 472816 288569 473346
rect 289099 472816 289108 473346
rect 290852 473072 290878 473346
rect 291278 473072 291308 473346
rect 290852 473050 291308 473072
rect 288569 472810 289099 472816
rect 153733 472115 153742 472745
rect 154372 472115 154381 472745
rect 153737 472110 154377 472115
rect 290878 469712 291518 469718
rect 290869 469072 290878 469712
rect 291518 469072 291527 469712
rect 290878 469066 291518 469072
rect 294388 464776 294498 472185
rect 296388 471302 296498 472203
rect 297401 471945 297771 471951
rect 297392 471575 297401 471945
rect 297771 471575 297780 471945
rect 297401 471569 297771 471575
rect 296388 471185 301718 471302
rect 296392 468802 301718 471185
rect 306092 469146 306098 473946
rect 310898 473941 314138 473946
rect 314133 469151 314138 473941
rect 310898 469146 314138 469151
rect 309343 469142 314133 469146
rect 299218 467044 301718 468802
rect 466781 467044 469271 467048
rect 299218 467039 469276 467044
rect 294170 459648 296431 464776
rect 299218 464549 466781 467039
rect 469271 464549 469276 467039
rect 299218 464544 469276 464549
rect 466781 464540 469271 464544
rect 453211 459648 455701 459652
rect 294050 459643 455706 459648
rect 294050 457153 453211 459643
rect 455701 457153 455706 459643
rect 294050 457148 455706 457153
rect 453211 457144 455701 457148
rect 151524 442682 151761 442691
rect 150755 442559 151009 442568
rect 150755 441805 151009 442305
rect 150827 441143 150937 441805
rect 151524 440952 151761 442445
rect 140131 439680 140241 439689
rect 140241 439570 141469 439680
rect 140131 439561 140241 439570
rect 454910 438538 455220 438542
rect 454905 438533 515380 438538
rect 454905 438223 454910 438533
rect 455220 438223 515380 438533
rect 454905 438218 515380 438223
rect 515700 438218 515709 438538
rect 454910 438214 455220 438218
rect 149102 437806 149422 437812
rect 149102 437229 149422 437486
rect 149098 436919 149107 437229
rect 149417 436919 149426 437229
rect 149102 436914 149422 436919
rect 149102 436485 149422 436496
rect 149098 436175 149107 436485
rect 149417 436175 149426 436485
rect 149102 436164 149422 436175
rect 454910 435538 455220 435542
rect 454905 435533 515380 435538
rect 454905 435223 454910 435533
rect 455220 435223 515380 435533
rect 454905 435218 515380 435223
rect 515700 435218 515709 435538
rect 454910 435214 455220 435218
rect 454910 432538 455220 432542
rect 454905 432533 515380 432538
rect 454905 432223 454910 432533
rect 455220 432223 515380 432533
rect 454905 432218 515380 432223
rect 515700 432218 515709 432538
rect 454910 432214 455220 432218
rect 454910 429538 455220 429542
rect 454905 429533 515380 429538
rect 454905 429223 454910 429533
rect 455220 429223 515380 429533
rect 454905 429218 515380 429223
rect 515700 429218 515709 429538
rect 454910 429214 455220 429218
rect 454910 426538 455220 426542
rect 454905 426533 515380 426538
rect 454905 426223 454910 426533
rect 455220 426223 515380 426533
rect 454905 426218 515380 426223
rect 515700 426218 515709 426538
rect 454910 426214 455220 426218
rect 454910 423538 455220 423542
rect 454905 423533 515380 423538
rect 454905 423223 454910 423533
rect 455220 423223 515380 423533
rect 454905 423218 515380 423223
rect 515700 423218 515709 423538
rect 454910 423214 455220 423218
rect 454910 420538 455220 420542
rect 454905 420533 515380 420538
rect 454905 420223 454910 420533
rect 455220 420223 515380 420533
rect 454905 420218 515380 420223
rect 515700 420218 515709 420538
rect 454910 420214 455220 420218
rect 454910 417538 455220 417542
rect 454905 417533 515380 417538
rect 454905 417223 454910 417533
rect 455220 417223 515380 417533
rect 454905 417218 515380 417223
rect 515700 417218 515709 417538
rect 454910 417214 455220 417218
rect 454910 414538 455220 414542
rect 454905 414533 515380 414538
rect 454905 414223 454910 414533
rect 455220 414223 515380 414533
rect 454905 414218 515380 414223
rect 515700 414218 515709 414538
rect 454910 414214 455220 414218
rect 454910 411538 455220 411542
rect 454905 411533 515380 411538
rect 454905 411223 454910 411533
rect 455220 411223 515380 411533
rect 454905 411218 515380 411223
rect 515700 411218 515709 411538
rect 454910 411214 455220 411218
rect 454910 408538 455220 408542
rect 454905 408533 515380 408538
rect 454905 408223 454910 408533
rect 455220 408223 515380 408533
rect 454905 408218 515380 408223
rect 515700 408218 515709 408538
rect 454910 408214 455220 408218
rect 454910 405538 455220 405542
rect 454905 405533 515380 405538
rect 454905 405223 454910 405533
rect 455220 405223 515380 405533
rect 454905 405218 515380 405223
rect 515700 405218 515709 405538
rect 454910 405214 455220 405218
rect 454910 402538 455220 402542
rect 454905 402533 515380 402538
rect 454905 402223 454910 402533
rect 455220 402223 515380 402533
rect 454905 402218 515380 402223
rect 515700 402218 515709 402538
rect 454910 402214 455220 402218
rect 454910 399538 455220 399542
rect 454905 399533 515380 399538
rect 454905 399223 454910 399533
rect 455220 399223 515380 399533
rect 454905 399218 515380 399223
rect 515700 399218 515709 399538
rect 454910 399214 455220 399218
rect 454910 396538 455220 396542
rect 454905 396533 515380 396538
rect 454905 396223 454910 396533
rect 455220 396223 515380 396533
rect 454905 396218 515380 396223
rect 515700 396218 515709 396538
rect 454910 396214 455220 396218
rect 454910 393538 455220 393542
rect 454905 393533 515380 393538
rect 454905 393223 454910 393533
rect 455220 393223 515380 393533
rect 454905 393218 515380 393223
rect 515700 393218 515709 393538
rect 454910 393214 455220 393218
rect 454910 390538 455220 390542
rect 454905 390533 515380 390538
rect 454905 390223 454910 390533
rect 455220 390223 515380 390533
rect 454905 390218 515380 390223
rect 515700 390218 515709 390538
rect 454910 390214 455220 390218
rect 454910 387538 455220 387542
rect 454905 387533 515380 387538
rect 454905 387223 454910 387533
rect 455220 387223 515380 387533
rect 454905 387218 515380 387223
rect 515700 387218 515709 387538
rect 454910 387214 455220 387218
rect 454910 384538 455220 384542
rect 454905 384533 515380 384538
rect 454905 384223 454910 384533
rect 455220 384223 515380 384533
rect 454905 384218 515380 384223
rect 515700 384218 515709 384538
rect 454910 384214 455220 384218
rect 454910 381538 455220 381542
rect 454905 381533 515380 381538
rect 454905 381223 454910 381533
rect 455220 381223 515380 381533
rect 454905 381218 515380 381223
rect 515700 381218 515709 381538
rect 454910 381214 455220 381218
rect 454910 378538 455220 378542
rect 454905 378533 515380 378538
rect 454905 378223 454910 378533
rect 455220 378223 515380 378533
rect 454905 378218 515380 378223
rect 515700 378218 515709 378538
rect 454910 378214 455220 378218
rect 454910 375538 455220 375542
rect 454905 375533 515380 375538
rect 454905 375223 454910 375533
rect 455220 375223 515380 375533
rect 454905 375218 515380 375223
rect 515700 375218 515709 375538
rect 454910 375214 455220 375218
rect 454910 372538 455220 372542
rect 454905 372533 515380 372538
rect 454905 372223 454910 372533
rect 455220 372223 515380 372533
rect 454905 372218 515380 372223
rect 515700 372218 515709 372538
rect 454910 372214 455220 372218
rect 454910 369538 455220 369542
rect 454905 369533 515380 369538
rect 454905 369223 454910 369533
rect 455220 369223 515380 369533
rect 454905 369218 515380 369223
rect 515700 369218 515709 369538
rect 454910 369214 455220 369218
rect 454910 366538 455220 366542
rect 454905 366533 515380 366538
rect 454905 366223 454910 366533
rect 455220 366223 515380 366533
rect 454905 366218 515380 366223
rect 515700 366218 515709 366538
rect 454910 366214 455220 366218
rect 454910 363538 455220 363542
rect 454905 363533 515380 363538
rect 454905 363223 454910 363533
rect 455220 363223 515380 363533
rect 454905 363218 515380 363223
rect 515700 363218 515709 363538
rect 454910 363214 455220 363218
rect 454910 360538 455220 360542
rect 454905 360533 515380 360538
rect 454905 360223 454910 360533
rect 455220 360223 515380 360533
rect 454905 360218 515380 360223
rect 515700 360218 515709 360538
rect 454910 360214 455220 360218
rect 454910 357538 455220 357542
rect 454905 357533 515380 357538
rect 454905 357223 454910 357533
rect 455220 357223 515380 357533
rect 454905 357218 515380 357223
rect 515700 357218 515709 357538
rect 454910 357214 455220 357218
rect 454910 354538 455220 354542
rect 454905 354533 515380 354538
rect 454905 354223 454910 354533
rect 455220 354223 515380 354533
rect 454905 354218 515380 354223
rect 515700 354218 515709 354538
rect 454910 354214 455220 354218
rect 454910 351538 455220 351542
rect 454905 351533 515380 351538
rect 454905 351223 454910 351533
rect 455220 351223 515380 351533
rect 454905 351218 515380 351223
rect 515700 351218 515709 351538
rect 454910 351214 455220 351218
rect 454910 348538 455220 348542
rect 454905 348533 515380 348538
rect 454905 348223 454910 348533
rect 455220 348223 515380 348533
rect 454905 348218 515380 348223
rect 515700 348218 515709 348538
rect 454910 348214 455220 348218
rect 454910 345538 455220 345542
rect 454905 345533 515380 345538
rect 454905 345223 454910 345533
rect 455220 345223 515380 345533
rect 454905 345218 515380 345223
rect 515700 345218 515709 345538
rect 454910 345214 455220 345218
rect 454910 342538 455220 342542
rect 454905 342533 515380 342538
rect 454905 342223 454910 342533
rect 455220 342223 515380 342533
rect 454905 342218 515380 342223
rect 515700 342218 515709 342538
rect 454910 342214 455220 342218
rect 454910 339538 455220 339542
rect 454905 339533 515380 339538
rect 454905 339223 454910 339533
rect 455220 339223 515380 339533
rect 454905 339218 515380 339223
rect 515700 339218 515709 339538
rect 454910 339214 455220 339218
rect 5660 336789 5772 336794
rect 5656 336687 5665 336789
rect 5767 336687 5776 336789
rect 5660 327595 5772 336687
rect 454910 336538 455220 336542
rect 454905 336533 515380 336538
rect 454905 336223 454910 336533
rect 455220 336223 515380 336533
rect 454905 336218 515380 336223
rect 515700 336218 515709 336538
rect 454910 336214 455220 336218
rect 454910 333538 455220 333542
rect 454905 333533 515380 333538
rect 454905 333223 454910 333533
rect 455220 333223 515380 333533
rect 454905 333218 515380 333223
rect 515700 333218 515709 333538
rect 454910 333214 455220 333218
rect 454910 330538 455220 330542
rect 454905 330533 515380 330538
rect 454905 330223 454910 330533
rect 455220 330223 515380 330533
rect 454905 330218 515380 330223
rect 515700 330218 515709 330538
rect 454910 330214 455220 330218
rect 454910 327538 455220 327542
rect 5660 327474 5772 327483
rect 454905 327533 515380 327538
rect 454905 327223 454910 327533
rect 455220 327223 515380 327533
rect 454905 327218 515380 327223
rect 515700 327218 515709 327538
rect 454910 327214 455220 327218
rect 454910 324538 455220 324542
rect 454905 324533 515380 324538
rect 454905 324223 454910 324533
rect 455220 324223 515380 324533
rect 454905 324218 515380 324223
rect 515700 324218 515709 324538
rect 454910 324214 455220 324218
rect 454910 321538 455220 321542
rect 454905 321533 515380 321538
rect 454905 321223 454910 321533
rect 455220 321223 515380 321533
rect 454905 321218 515380 321223
rect 515700 321218 515709 321538
rect 454910 321214 455220 321218
rect 454910 318538 455220 318542
rect 454905 318533 515380 318538
rect 454905 318223 454910 318533
rect 455220 318223 515380 318533
rect 454905 318218 515380 318223
rect 515700 318218 515709 318538
rect 454910 318214 455220 318218
rect 454910 315538 455220 315542
rect 454905 315533 515380 315538
rect 454905 315223 454910 315533
rect 455220 315223 515380 315533
rect 454905 315218 515380 315223
rect 515700 315218 515709 315538
rect 454910 315214 455220 315218
rect 454910 312538 455220 312542
rect 454905 312533 515380 312538
rect 454905 312223 454910 312533
rect 455220 312223 515380 312533
rect 454905 312218 515380 312223
rect 515700 312218 515709 312538
rect 454910 312214 455220 312218
rect 454910 309538 455220 309542
rect 454905 309533 515380 309538
rect 454905 309223 454910 309533
rect 455220 309223 515380 309533
rect 454905 309218 515380 309223
rect 515700 309218 515709 309538
rect 454910 309214 455220 309218
rect 454910 306538 455220 306542
rect 454905 306533 515380 306538
rect 454905 306223 454910 306533
rect 455220 306223 515380 306533
rect 454905 306218 515380 306223
rect 515700 306218 515709 306538
rect 454910 306214 455220 306218
rect 454910 303538 455220 303542
rect 454905 303533 515380 303538
rect 454905 303223 454910 303533
rect 455220 303223 515380 303533
rect 454905 303218 515380 303223
rect 515700 303218 515709 303538
rect 454910 303214 455220 303218
rect 454910 300538 455220 300542
rect 454905 300533 515380 300538
rect 454905 300223 454910 300533
rect 455220 300223 515380 300533
rect 454905 300218 515380 300223
rect 515700 300218 515709 300538
rect 454910 300214 455220 300218
rect 454910 297538 455220 297542
rect 454905 297533 515380 297538
rect 454905 297223 454910 297533
rect 455220 297223 515380 297533
rect 454905 297218 515380 297223
rect 515700 297218 515709 297538
rect 454910 297214 455220 297218
rect 454910 294538 455220 294542
rect 454905 294533 515380 294538
rect 454905 294223 454910 294533
rect 455220 294223 515380 294533
rect 454905 294218 515380 294223
rect 515700 294218 515709 294538
rect 454910 294214 455220 294218
rect 454910 291538 455220 291542
rect 454905 291533 515380 291538
rect 454905 291223 454910 291533
rect 455220 291223 515380 291533
rect 454905 291218 515380 291223
rect 515700 291218 515709 291538
rect 454910 291214 455220 291218
rect 454910 288538 455220 288542
rect 454905 288533 515380 288538
rect 454905 288223 454910 288533
rect 455220 288223 515380 288533
rect 454905 288218 515380 288223
rect 515700 288218 515709 288538
rect 454910 288214 455220 288218
rect 454910 285538 455220 285542
rect 454905 285533 515380 285538
rect 454905 285223 454910 285533
rect 455220 285223 515380 285533
rect 454905 285218 515380 285223
rect 515700 285218 515709 285538
rect 454910 285214 455220 285218
rect 454910 282538 455220 282542
rect 454905 282533 515380 282538
rect 454905 282223 454910 282533
rect 455220 282223 515380 282533
rect 454905 282218 515380 282223
rect 515700 282218 515709 282538
rect 454910 282214 455220 282218
rect 454910 279538 455220 279542
rect 454905 279533 515380 279538
rect 454905 279223 454910 279533
rect 455220 279223 515380 279533
rect 454905 279218 515380 279223
rect 515700 279218 515709 279538
rect 454910 279214 455220 279218
rect 454910 276538 455220 276542
rect 454905 276533 515380 276538
rect 454905 276223 454910 276533
rect 455220 276223 515380 276533
rect 454905 276218 515380 276223
rect 515700 276218 515709 276538
rect 454910 276214 455220 276218
rect 454910 273538 455220 273542
rect 454905 273533 515380 273538
rect 454905 273223 454910 273533
rect 455220 273223 515380 273533
rect 454905 273218 515380 273223
rect 515700 273218 515709 273538
rect 454910 273214 455220 273218
rect 454910 270538 455220 270542
rect 454905 270533 515380 270538
rect 454905 270223 454910 270533
rect 455220 270223 515380 270533
rect 454905 270218 515380 270223
rect 515700 270218 515709 270538
rect 454910 270214 455220 270218
rect 454910 267538 455220 267542
rect 454905 267533 515380 267538
rect 454905 267223 454910 267533
rect 455220 267223 515380 267533
rect 454905 267218 515380 267223
rect 515700 267218 515709 267538
rect 454910 267214 455220 267218
rect 454910 264538 455220 264542
rect 454905 264533 515380 264538
rect 454905 264223 454910 264533
rect 455220 264223 515380 264533
rect 454905 264218 515380 264223
rect 515700 264218 515709 264538
rect 454910 264214 455220 264218
rect 454910 261538 455220 261542
rect 454905 261533 515380 261538
rect 8362 261315 8493 261350
rect 8362 261245 8387 261315
rect 8457 261245 8493 261315
rect 8362 261225 8493 261245
rect 454905 261223 454910 261533
rect 455220 261223 515380 261533
rect 454905 261218 515380 261223
rect 515700 261218 515709 261538
rect 454910 261214 455220 261218
rect 454910 258538 455220 258542
rect 454905 258533 515380 258538
rect 454905 258223 454910 258533
rect 455220 258223 515380 258533
rect 454905 258218 515380 258223
rect 515700 258218 515709 258538
rect 454910 258214 455220 258218
rect 454910 255538 455220 255542
rect 454905 255533 515380 255538
rect 454905 255223 454910 255533
rect 455220 255223 515380 255533
rect 454905 255218 515380 255223
rect 515700 255218 515709 255538
rect 454910 255214 455220 255218
rect 454910 252538 455220 252542
rect 454905 252533 515380 252538
rect 454905 252223 454910 252533
rect 455220 252223 515380 252533
rect 454905 252218 515380 252223
rect 515700 252218 515709 252538
rect 454910 252214 455220 252218
rect 454910 249538 455220 249542
rect 454905 249533 515380 249538
rect 454905 249223 454910 249533
rect 455220 249223 515380 249533
rect 454905 249218 515380 249223
rect 515700 249218 515709 249538
rect 454910 249214 455220 249218
rect 454910 246538 455220 246542
rect 454905 246533 515380 246538
rect 454905 246223 454910 246533
rect 455220 246223 515380 246533
rect 454905 246218 515380 246223
rect 515700 246218 515709 246538
rect 454910 246214 455220 246218
rect 454910 243538 455220 243542
rect 454905 243533 515380 243538
rect 454905 243223 454910 243533
rect 455220 243223 515380 243533
rect 454905 243218 515380 243223
rect 515700 243218 515709 243538
rect 454910 243214 455220 243218
rect 454910 240538 455220 240542
rect 454905 240533 515380 240538
rect 454905 240223 454910 240533
rect 455220 240223 515380 240533
rect 454905 240218 515380 240223
rect 515700 240218 515709 240538
rect 454910 240214 455220 240218
rect 454910 237538 455220 237542
rect 454905 237533 515380 237538
rect 454905 237223 454910 237533
rect 455220 237223 515380 237533
rect 454905 237218 515380 237223
rect 515700 237218 515709 237538
rect 454910 237214 455220 237218
rect 454910 234538 455220 234542
rect 454905 234533 515380 234538
rect 454905 234223 454910 234533
rect 455220 234223 515380 234533
rect 454905 234218 515380 234223
rect 515700 234218 515709 234538
rect 454910 234214 455220 234218
rect 454910 231538 455220 231542
rect 454905 231533 515380 231538
rect 454905 231223 454910 231533
rect 455220 231223 515380 231533
rect 454905 231218 515380 231223
rect 515700 231218 515709 231538
rect 454910 231214 455220 231218
rect 454910 228538 455220 228542
rect 454905 228533 515380 228538
rect 454905 228223 454910 228533
rect 455220 228223 515380 228533
rect 454905 228218 515380 228223
rect 515700 228218 515709 228538
rect 454910 228214 455220 228218
rect 454910 225538 455220 225542
rect 454905 225533 515380 225538
rect 454905 225223 454910 225533
rect 455220 225223 515380 225533
rect 454905 225218 515380 225223
rect 515700 225218 515709 225538
rect 454910 225214 455220 225218
rect 454910 222538 455220 222542
rect 454905 222533 515380 222538
rect 454905 222223 454910 222533
rect 455220 222223 515380 222533
rect 454905 222218 515380 222223
rect 515700 222218 515709 222538
rect 454910 222214 455220 222218
rect 454910 219538 455220 219542
rect 454905 219533 515380 219538
rect 454905 219223 454910 219533
rect 455220 219223 515380 219533
rect 454905 219218 515380 219223
rect 515700 219218 515709 219538
rect 454910 219214 455220 219218
rect 454910 216538 455220 216542
rect 454905 216533 515380 216538
rect 454905 216223 454910 216533
rect 455220 216223 515380 216533
rect 454905 216218 515380 216223
rect 515700 216218 515709 216538
rect 454910 216214 455220 216218
rect 454910 213538 455220 213542
rect 454905 213533 515380 213538
rect 454905 213223 454910 213533
rect 455220 213223 515380 213533
rect 454905 213218 515380 213223
rect 515700 213218 515709 213538
rect 454910 213214 455220 213218
rect 454910 210538 455220 210542
rect 454905 210533 515380 210538
rect 454905 210223 454910 210533
rect 455220 210223 515380 210533
rect 454905 210218 515380 210223
rect 515700 210218 515709 210538
rect 454910 210214 455220 210218
rect 454910 207538 455220 207542
rect 454905 207533 515380 207538
rect 454905 207223 454910 207533
rect 455220 207223 515380 207533
rect 454905 207218 515380 207223
rect 515700 207218 515709 207538
rect 454910 207214 455220 207218
rect 454910 204538 455220 204542
rect 454905 204533 515380 204538
rect 454905 204223 454910 204533
rect 455220 204223 515380 204533
rect 454905 204218 515380 204223
rect 515700 204218 515709 204538
rect 454910 204214 455220 204218
rect 454910 201538 455220 201542
rect 454905 201533 515380 201538
rect 454905 201223 454910 201533
rect 455220 201223 515380 201533
rect 454905 201218 515380 201223
rect 515700 201218 515709 201538
rect 454910 201214 455220 201218
rect 454910 198538 455220 198542
rect 454905 198533 515380 198538
rect 454905 198223 454910 198533
rect 455220 198223 515380 198533
rect 454905 198218 515380 198223
rect 515700 198218 515709 198538
rect 454910 198214 455220 198218
rect 454910 195538 455220 195542
rect 454905 195533 515380 195538
rect 454905 195223 454910 195533
rect 455220 195223 515380 195533
rect 454905 195218 515380 195223
rect 515700 195218 515709 195538
rect 454910 195214 455220 195218
rect 454910 192538 455220 192542
rect 454905 192533 515380 192538
rect 454905 192223 454910 192533
rect 455220 192223 515380 192533
rect 454905 192218 515380 192223
rect 515700 192218 515709 192538
rect 454910 192214 455220 192218
rect 9016 191337 9126 191346
rect 9126 191227 10882 191337
rect 9016 191218 9126 191227
rect 454910 189538 455220 189542
rect 454905 189533 515380 189538
rect 454905 189223 454910 189533
rect 455220 189223 515380 189533
rect 454905 189218 515380 189223
rect 515700 189218 515709 189538
rect 454910 189214 455220 189218
rect 454910 186538 455220 186542
rect 454905 186533 515380 186538
rect 454905 186223 454910 186533
rect 455220 186223 515380 186533
rect 454905 186218 515380 186223
rect 515700 186218 515709 186538
rect 454910 186214 455220 186218
rect 454910 183538 455220 183542
rect 454905 183533 515380 183538
rect 454905 183223 454910 183533
rect 455220 183223 515380 183533
rect 454905 183218 515380 183223
rect 515700 183218 515709 183538
rect 454910 183214 455220 183218
rect 454910 180538 455220 180542
rect 454905 180533 515380 180538
rect 454905 180223 454910 180533
rect 455220 180223 515380 180533
rect 454905 180218 515380 180223
rect 515700 180218 515709 180538
rect 454910 180214 455220 180218
rect 454910 177538 455220 177542
rect 454905 177533 515380 177538
rect 454905 177223 454910 177533
rect 455220 177223 515380 177533
rect 454905 177218 515380 177223
rect 515700 177218 515709 177538
rect 454910 177214 455220 177218
rect 454910 174538 455220 174542
rect 454905 174533 515380 174538
rect 454905 174223 454910 174533
rect 455220 174223 515380 174533
rect 454905 174218 515380 174223
rect 515700 174218 515709 174538
rect 454910 174214 455220 174218
rect 454910 171538 455220 171542
rect 454905 171533 515380 171538
rect 454905 171223 454910 171533
rect 455220 171223 515380 171533
rect 454905 171218 515380 171223
rect 515700 171218 515709 171538
rect 454910 171214 455220 171218
rect 454910 168538 455220 168542
rect 454905 168533 515380 168538
rect 454905 168223 454910 168533
rect 455220 168223 515380 168533
rect 454905 168218 515380 168223
rect 515700 168218 515709 168538
rect 454910 168214 455220 168218
rect 454910 165538 455220 165542
rect 454905 165533 515380 165538
rect 454905 165223 454910 165533
rect 455220 165223 515380 165533
rect 454905 165218 515380 165223
rect 515700 165218 515709 165538
rect 454910 165214 455220 165218
rect 454910 162538 455220 162542
rect 454905 162533 515380 162538
rect 454905 162223 454910 162533
rect 455220 162223 515380 162533
rect 454905 162218 515380 162223
rect 515700 162218 515709 162538
rect 454910 162214 455220 162218
rect 454910 159538 455220 159542
rect 454905 159533 515380 159538
rect 454905 159223 454910 159533
rect 455220 159223 515380 159533
rect 454905 159218 515380 159223
rect 515700 159218 515709 159538
rect 454910 159214 455220 159218
rect 454910 156538 455220 156542
rect 454905 156533 515380 156538
rect 454905 156223 454910 156533
rect 455220 156223 515380 156533
rect 454905 156218 515380 156223
rect 515700 156218 515709 156538
rect 454910 156214 455220 156218
rect 454910 153538 455220 153542
rect 454905 153533 515380 153538
rect 454905 153223 454910 153533
rect 455220 153223 515380 153533
rect 454905 153218 515380 153223
rect 515700 153218 515709 153538
rect 454910 153214 455220 153218
rect 454910 150538 455220 150542
rect 454905 150533 515380 150538
rect 454905 150223 454910 150533
rect 455220 150223 515380 150533
rect 454905 150218 515380 150223
rect 515700 150218 515709 150538
rect 454910 150214 455220 150218
rect 501754 140997 502630 141003
rect 493474 140867 494090 140873
rect 495806 140867 495812 140997
rect 488760 140251 488766 140867
rect 489382 140251 493474 140867
rect 494090 140251 495812 140867
rect 493474 140245 494090 140251
rect 495806 140121 495812 140251
rect 496688 140121 501754 140997
rect 502630 140121 503862 140997
rect 501754 140115 502630 140121
rect 461961 139833 462131 139842
rect 461961 139194 462131 139663
rect 461955 139024 461961 139194
rect 462131 139024 462137 139194
rect 126336 133775 127424 133780
rect 126332 132697 126341 133775
rect 127419 132697 127428 133775
rect 456062 133482 463212 133662
rect 462900 132745 463148 133482
rect 126336 129154 127424 132697
rect 144651 129154 145729 129158
rect 127424 129149 146798 129154
rect 127424 128071 144651 129149
rect 145729 128071 146798 129149
rect 460671 128894 460841 128903
rect 460841 128724 463461 128894
rect 460671 128715 460841 128724
rect 127424 128066 146798 128071
rect 126336 127220 127424 128066
rect 144651 128062 145729 128066
rect 19138 125184 19258 125193
rect 19138 118686 19258 125064
rect 21326 124954 21446 124963
rect 21326 120178 21446 124834
rect 27250 124898 27370 124907
rect 130318 124898 130428 124902
rect 27370 124893 130433 124898
rect 27370 124783 130318 124893
rect 130428 124783 130433 124893
rect 27370 124778 130433 124783
rect 27250 124769 27370 124778
rect 130318 124774 130428 124778
rect 24558 123672 24678 123681
rect 24678 123552 124366 123672
rect 24558 123543 24678 123552
rect 124246 120770 124366 123552
rect 134262 120770 134372 120774
rect 124246 120765 134377 120770
rect 124246 120655 134262 120765
rect 134372 120655 134377 120765
rect 124246 120650 134377 120655
rect 134262 120646 134372 120650
rect 138342 120178 138452 120182
rect 21326 120173 138457 120178
rect 21326 120063 138342 120173
rect 138452 120063 138457 120173
rect 21326 120058 138457 120063
rect 138342 120054 138452 120058
rect 142286 118686 142396 118690
rect 19138 118681 142401 118686
rect 19138 118571 142286 118681
rect 142396 118571 142401 118681
rect 19138 118566 142401 118571
rect 142286 118562 142396 118566
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 274227 592538 276717 595025
rect 308461 594295 308631 594465
rect 274227 592535 275898 592538
rect 276506 592535 276717 592538
rect 288821 592180 289156 592515
rect 257406 590190 257726 590510
rect 287849 590195 288159 590505
rect 338103 591485 338393 591775
rect 338103 591041 338393 591331
rect 338108 590655 338388 590744
rect 338103 590365 338393 590655
rect 270806 587584 271643 588421
rect 338108 590274 338388 590365
rect 234629 587021 234719 587111
rect 236793 586709 236883 586799
rect 338108 586655 338388 586744
rect 338103 586365 338393 586655
rect 240447 584222 240537 584312
rect 265890 578736 266355 579201
rect 286432 578822 286724 579114
rect 243956 571632 244176 571852
rect 291821 571637 292031 571847
rect 291977 570715 292187 570925
rect 249279 570274 249381 570363
rect 249200 570054 249420 570274
rect 229970 567922 230190 568142
rect 292245 567927 292455 568137
rect 255195 528794 258683 532282
rect 255190 526818 257054 528682
rect 332643 575353 333137 575847
rect 347632 585352 347792 585512
rect 461821 585219 462247 585645
rect 371804 575358 372288 575842
rect 444605 575353 445099 575847
rect 343674 486080 344106 486512
rect 152404 477296 153444 478336
rect 291713 477735 291903 477925
rect 415673 477301 416703 478331
rect 343679 475469 344101 475891
rect 292223 474789 292413 474979
rect 431840 474146 432768 475074
rect 288569 472816 289099 473346
rect 153742 472115 154372 472745
rect 290878 469346 291518 469712
rect 290878 469072 291278 469346
rect 291278 469072 291518 469346
rect 297401 471575 297771 471945
rect 309343 469151 310898 473941
rect 310898 469151 314133 473941
rect 466781 464549 469271 467039
rect 453211 457153 455701 459643
rect 150755 442305 151009 442559
rect 151524 442445 151761 442682
rect 140131 439570 140241 439680
rect 454910 438223 455220 438533
rect 515380 438218 515700 438538
rect 149107 436919 149417 437229
rect 149107 436175 149417 436485
rect 454910 435223 455220 435533
rect 515380 435218 515700 435538
rect 454910 432223 455220 432533
rect 515380 432218 515700 432538
rect 454910 429223 455220 429533
rect 515380 429218 515700 429538
rect 454910 426223 455220 426533
rect 515380 426218 515700 426538
rect 454910 423223 455220 423533
rect 515380 423218 515700 423538
rect 454910 420223 455220 420533
rect 515380 420218 515700 420538
rect 454910 417223 455220 417533
rect 515380 417218 515700 417538
rect 454910 414223 455220 414533
rect 515380 414218 515700 414538
rect 454910 411223 455220 411533
rect 515380 411218 515700 411538
rect 454910 408223 455220 408533
rect 515380 408218 515700 408538
rect 454910 405223 455220 405533
rect 515380 405218 515700 405538
rect 454910 402223 455220 402533
rect 515380 402218 515700 402538
rect 454910 399223 455220 399533
rect 515380 399218 515700 399538
rect 454910 396223 455220 396533
rect 515380 396218 515700 396538
rect 454910 393223 455220 393533
rect 515380 393218 515700 393538
rect 454910 390223 455220 390533
rect 515380 390218 515700 390538
rect 454910 387223 455220 387533
rect 515380 387218 515700 387538
rect 454910 384223 455220 384533
rect 515380 384218 515700 384538
rect 454910 381223 455220 381533
rect 515380 381218 515700 381538
rect 454910 378223 455220 378533
rect 515380 378218 515700 378538
rect 454910 375223 455220 375533
rect 515380 375218 515700 375538
rect 454910 372223 455220 372533
rect 515380 372218 515700 372538
rect 454910 369223 455220 369533
rect 515380 369218 515700 369538
rect 454910 366223 455220 366533
rect 515380 366218 515700 366538
rect 454910 363223 455220 363533
rect 515380 363218 515700 363538
rect 454910 360223 455220 360533
rect 515380 360218 515700 360538
rect 454910 357223 455220 357533
rect 515380 357218 515700 357538
rect 454910 354223 455220 354533
rect 515380 354218 515700 354538
rect 454910 351223 455220 351533
rect 515380 351218 515700 351538
rect 454910 348223 455220 348533
rect 515380 348218 515700 348538
rect 454910 345223 455220 345533
rect 515380 345218 515700 345538
rect 454910 342223 455220 342533
rect 515380 342218 515700 342538
rect 454910 339223 455220 339533
rect 515380 339218 515700 339538
rect 5665 336687 5767 336789
rect 454910 336223 455220 336533
rect 515380 336218 515700 336538
rect 454910 333223 455220 333533
rect 515380 333218 515700 333538
rect 454910 330223 455220 330533
rect 515380 330218 515700 330538
rect 5660 327483 5772 327595
rect 454910 327223 455220 327533
rect 515380 327218 515700 327538
rect 454910 324223 455220 324533
rect 515380 324218 515700 324538
rect 454910 321223 455220 321533
rect 515380 321218 515700 321538
rect 454910 318223 455220 318533
rect 515380 318218 515700 318538
rect 454910 315223 455220 315533
rect 515380 315218 515700 315538
rect 454910 312223 455220 312533
rect 515380 312218 515700 312538
rect 454910 309223 455220 309533
rect 515380 309218 515700 309538
rect 454910 306223 455220 306533
rect 515380 306218 515700 306538
rect 454910 303223 455220 303533
rect 515380 303218 515700 303538
rect 454910 300223 455220 300533
rect 515380 300218 515700 300538
rect 454910 297223 455220 297533
rect 515380 297218 515700 297538
rect 454910 294223 455220 294533
rect 515380 294218 515700 294538
rect 454910 291223 455220 291533
rect 515380 291218 515700 291538
rect 454910 288223 455220 288533
rect 515380 288218 515700 288538
rect 454910 285223 455220 285533
rect 515380 285218 515700 285538
rect 454910 282223 455220 282533
rect 515380 282218 515700 282538
rect 454910 279223 455220 279533
rect 515380 279218 515700 279538
rect 454910 276223 455220 276533
rect 515380 276218 515700 276538
rect 454910 273223 455220 273533
rect 515380 273218 515700 273538
rect 454910 270223 455220 270533
rect 515380 270218 515700 270538
rect 454910 267223 455220 267533
rect 515380 267218 515700 267538
rect 454910 264223 455220 264533
rect 515380 264218 515700 264538
rect 8387 261245 8457 261315
rect 454910 261223 455220 261533
rect 515380 261218 515700 261538
rect 454910 258223 455220 258533
rect 515380 258218 515700 258538
rect 454910 255223 455220 255533
rect 515380 255218 515700 255538
rect 454910 252223 455220 252533
rect 515380 252218 515700 252538
rect 454910 249223 455220 249533
rect 515380 249218 515700 249538
rect 454910 246223 455220 246533
rect 515380 246218 515700 246538
rect 454910 243223 455220 243533
rect 515380 243218 515700 243538
rect 454910 240223 455220 240533
rect 515380 240218 515700 240538
rect 454910 237223 455220 237533
rect 515380 237218 515700 237538
rect 454910 234223 455220 234533
rect 515380 234218 515700 234538
rect 454910 231223 455220 231533
rect 515380 231218 515700 231538
rect 454910 228223 455220 228533
rect 515380 228218 515700 228538
rect 454910 225223 455220 225533
rect 515380 225218 515700 225538
rect 454910 222223 455220 222533
rect 515380 222218 515700 222538
rect 454910 219223 455220 219533
rect 515380 219218 515700 219538
rect 454910 216223 455220 216533
rect 515380 216218 515700 216538
rect 454910 213223 455220 213533
rect 515380 213218 515700 213538
rect 454910 210223 455220 210533
rect 515380 210218 515700 210538
rect 454910 207223 455220 207533
rect 515380 207218 515700 207538
rect 454910 204223 455220 204533
rect 515380 204218 515700 204538
rect 454910 201223 455220 201533
rect 515380 201218 515700 201538
rect 454910 198223 455220 198533
rect 515380 198218 515700 198538
rect 454910 195223 455220 195533
rect 515380 195218 515700 195538
rect 454910 192223 455220 192533
rect 515380 192218 515700 192538
rect 9016 191227 9126 191337
rect 454910 189223 455220 189533
rect 515380 189218 515700 189538
rect 454910 186223 455220 186533
rect 515380 186218 515700 186538
rect 454910 183223 455220 183533
rect 515380 183218 515700 183538
rect 454910 180223 455220 180533
rect 515380 180218 515700 180538
rect 454910 177223 455220 177533
rect 515380 177218 515700 177538
rect 454910 174223 455220 174533
rect 515380 174218 515700 174538
rect 454910 171223 455220 171533
rect 515380 171218 515700 171538
rect 454910 168223 455220 168533
rect 515380 168218 515700 168538
rect 454910 165223 455220 165533
rect 515380 165218 515700 165538
rect 454910 162223 455220 162533
rect 515380 162218 515700 162538
rect 454910 159223 455220 159533
rect 515380 159218 515700 159538
rect 454910 156223 455220 156533
rect 515380 156218 515700 156538
rect 454910 153223 455220 153533
rect 515380 153218 515700 153538
rect 454910 150223 455220 150533
rect 515380 150218 515700 150538
rect 501754 140121 502630 140997
rect 461961 139663 462131 139833
rect 126341 132697 127419 133775
rect 126336 128066 127424 129154
rect 144651 128071 145729 129149
rect 460671 128724 460841 128894
rect 19138 125064 19258 125184
rect 21326 124834 21446 124954
rect 27250 124778 27370 124898
rect 130318 124783 130428 124893
rect 24558 123552 24678 123672
rect 134262 120655 134372 120765
rect 138342 120063 138452 120173
rect 142286 118571 142396 118681
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703390 418394 704800
rect 413394 703190 427730 703390
rect 413394 702300 418394 703190
rect 18694 696582 21194 702300
rect 18694 694082 66444 696582
rect 18694 693414 21194 694082
rect -800 682742 1700 685242
rect 63944 684066 66444 694082
rect 68940 690186 71440 702300
rect 122330 696788 124830 702300
rect 122330 696678 126146 696788
rect 122330 696013 124830 696678
rect 126036 696013 126146 696678
rect 122330 693513 173102 696013
rect 126036 690672 126146 693513
rect 68940 687686 168136 690186
rect -800 680242 61598 682742
rect 63944 681566 158432 684066
rect 59098 676618 61598 680242
rect 59098 674118 150778 676618
rect 6330 658270 8830 672796
rect 6330 655770 12018 658270
rect -800 643842 5110 648642
rect 148278 645006 150778 674118
rect 155932 650340 158432 681566
rect 165636 662826 168136 687686
rect 170602 669306 173102 693513
rect 177230 680264 179730 702300
rect 228438 698529 229478 698530
rect 228433 697491 228439 698529
rect 229477 697491 229483 698529
rect 331191 698285 332129 698286
rect 228438 686814 229478 697491
rect 331186 697349 331192 698285
rect 332128 697349 332134 698285
rect 228438 685774 316158 686814
rect 177230 677764 284582 680264
rect 170602 666806 276722 669306
rect 165636 660326 272166 662826
rect 155932 647840 265150 650340
rect 148278 642506 258688 645006
rect -800 633842 5110 638642
rect 256188 590510 258688 642506
rect 256188 590190 257406 590510
rect 257726 590190 258688 590510
rect 234624 587111 234724 587116
rect 234624 587021 234629 587111
rect 234719 587021 234724 587111
rect 234624 587016 234724 587021
rect 229965 568142 230195 568147
rect 229965 567922 229970 568142
rect 230190 567922 230195 568142
rect 229965 567917 230195 567922
rect -800 561902 1660 564242
rect -800 559442 1754 561902
rect -800 551902 1660 554242
rect -800 549442 1754 551902
rect 80622 533334 80734 533362
rect 229970 533334 230190 567917
rect 75398 533114 230190 533334
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 891 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect 1366 464931 1478 465323
rect 80622 464931 80734 533114
rect 234629 528757 234719 587016
rect 236788 586799 236888 586804
rect 236788 586709 236793 586799
rect 236883 586709 236888 586799
rect 236788 586704 236888 586709
rect 84431 528667 234719 528757
rect 1366 464874 80766 464931
rect -800 464819 80766 464874
rect -800 464762 1478 464819
rect -800 463580 480 463692
rect -800 462398 702 462510
rect 817 462376 1034 462476
rect 1134 462376 1140 462476
rect -800 425086 803 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 27458 421652
rect -800 420358 591 420470
rect 604 419288 690 419310
rect -800 419276 690 419288
rect -800 419176 717 419276
rect 817 419176 1034 419276
rect 1134 419176 1140 419276
rect -800 381864 979 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect 5660 379054 5772 419818
rect 1356 378430 1468 378793
rect -800 378318 1468 378430
rect 1356 377248 1468 378318
rect 24558 377248 24678 377756
rect -800 377136 824 377248
rect 1285 377136 24682 377248
rect 604 376076 690 376110
rect 604 376066 717 376076
rect -800 375976 717 376066
rect 817 375976 1034 376076
rect 1134 375976 1140 376076
rect -800 375954 690 375976
rect -800 338642 480 338754
rect -800 337460 480 337572
rect 5660 336789 5772 376032
rect 5660 336687 5665 336789
rect 5767 336687 5772 336789
rect 5660 336682 5772 336687
rect -800 336278 480 336390
rect 21326 335208 21446 335228
rect -800 335096 21476 335208
rect -800 333914 480 334026
rect -800 332810 654 332844
rect -800 332776 690 332810
rect -800 332732 717 332776
rect 542 332676 717 332732
rect 817 332676 1034 332776
rect 1134 332676 1140 332776
rect 542 332632 690 332676
rect 578 332608 690 332632
rect 5655 327595 5777 327600
rect 5655 327483 5660 327595
rect 5772 327483 5777 327595
rect 5655 327478 5777 327483
rect -800 295420 680 295532
rect -800 294238 480 294350
rect 5660 293381 5772 327478
rect 5660 293263 5772 293269
rect -800 293056 480 293168
rect 3192 291986 3304 292104
rect -800 291874 3840 291986
rect 3694 290804 3806 291874
rect -800 290692 1908 290804
rect 3672 290692 9839 290804
rect -800 289610 654 289622
rect -800 289576 690 289610
rect -800 289510 717 289576
rect 604 289498 717 289510
rect 660 289476 717 289498
rect 817 289476 1034 289576
rect 1134 289476 1140 289576
rect 9727 289082 9839 290692
rect 19138 289082 19258 291172
rect 9482 288962 19286 289082
rect 9727 288921 9839 288962
rect 8362 261320 8493 261350
rect 8362 261250 8382 261320
rect 8462 261250 8493 261320
rect 8362 261245 8387 261250
rect 8457 261245 8493 261250
rect 8362 261225 8493 261245
rect 19138 253335 19258 288962
rect 21326 253341 21446 335096
rect 24558 260523 24678 377136
rect 24553 260405 24559 260523
rect 24677 260405 24683 260523
rect 24558 260404 24678 260405
rect 27250 258973 27370 421540
rect 27245 258855 27251 258973
rect 27369 258855 27375 258973
rect 27250 258854 27370 258855
rect 19133 253217 19139 253335
rect 19257 253217 19263 253335
rect 21321 253223 21327 253341
rect 21445 253223 21451 253341
rect 21326 253222 21446 253223
rect 19138 253216 19258 253217
rect 5661 253173 5771 253178
rect 5660 253172 10882 253173
rect 5660 253062 5661 253172
rect 5771 253062 10882 253172
rect 5660 253061 10882 253062
rect 5661 253056 5771 253061
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect 84431 248964 84521 528667
rect 236793 525413 236883 586704
rect 240442 584312 240542 584317
rect 240442 584222 240447 584312
rect 240537 584222 240542 584312
rect 240442 584217 240542 584222
rect 90569 525323 236883 525413
rect -800 248852 84746 248964
rect 84431 248166 84521 248852
rect -800 247670 480 247782
rect 19138 247348 19258 247668
rect 604 246600 690 246610
rect -800 246576 690 246600
rect -800 246488 717 246576
rect 588 246476 717 246488
rect 817 246476 1034 246576
rect 1134 246476 1140 246576
rect 588 246407 690 246476
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 10674 191537 10784 191543
rect 10784 191427 10882 191537
rect 10674 191421 10784 191427
rect 9011 191342 9131 191348
rect 9011 191227 9016 191232
rect 9126 191227 9131 191232
rect 9011 191222 9131 191227
rect 2175 177688 3090 177800
rect -800 172888 3090 177688
rect 2175 167688 3090 172888
rect -800 162888 3090 167688
rect 19138 125189 19258 247228
rect 21326 247552 21446 247558
rect 19133 125184 19263 125189
rect 19133 125064 19138 125184
rect 19258 125064 19263 125184
rect 19133 125059 19263 125064
rect 21326 124959 21446 247432
rect 24558 245562 24678 245568
rect 21321 124954 21451 124959
rect -800 124776 480 124888
rect 21321 124834 21326 124954
rect 21446 124834 21451 124954
rect 21321 124829 21451 124834
rect -800 123594 480 123706
rect 24558 123677 24678 245442
rect 27250 244826 27370 244832
rect 27250 124903 27370 244706
rect 27245 124898 27375 124903
rect 27245 124778 27250 124898
rect 27370 124778 27375 124898
rect 27245 124773 27375 124778
rect 24553 123672 24683 123677
rect 24553 123552 24558 123672
rect 24678 123552 24683 123672
rect 24553 123547 24683 123552
rect -800 122412 480 122524
rect 90569 121342 90659 525323
rect 240447 524479 240537 584217
rect 256188 578600 258688 590190
rect 243951 571852 244181 571857
rect 243951 571632 243956 571852
rect 244176 571632 244181 571852
rect 243951 571627 244181 571632
rect -800 121230 90659 121342
rect -800 120048 480 120160
rect 604 118984 690 119010
rect 445 118978 690 118984
rect -800 118976 690 118978
rect -800 118876 717 118976
rect 817 118876 1034 118976
rect 1134 118876 1140 118976
rect -800 118866 480 118876
rect 90569 113839 90659 121230
rect 96745 524389 240537 524479
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect 96745 78120 96835 524389
rect 243956 520756 244176 571627
rect 249200 570363 249420 570892
rect 249200 570279 249279 570363
rect 249195 570274 249279 570279
rect 249381 570279 249420 570363
rect 249381 570274 249425 570279
rect 249195 570054 249200 570274
rect 249420 570054 249425 570274
rect 249195 570049 249425 570054
rect 249200 569732 249420 570049
rect 102724 520536 244176 520756
rect -800 78008 96840 78120
rect -800 76826 480 76938
rect 604 75776 690 75810
rect 604 75756 717 75776
rect -800 75676 717 75756
rect 817 75676 1034 75776
rect 1134 75676 1140 75776
rect -800 75644 662 75676
rect 96745 71505 96835 78008
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect 102724 34898 102944 520536
rect 249274 518820 249386 569732
rect 255190 532282 258688 578600
rect 255190 528794 255195 532282
rect 258683 528794 258688 532282
rect 255190 528789 258688 528794
rect 262650 579201 265150 647840
rect 269666 588421 272166 660326
rect 269406 587584 270806 588421
rect 271643 587584 272166 588421
rect 269666 587380 272166 587584
rect 265885 579201 266360 579206
rect 262650 578736 265890 579201
rect 266355 578736 266360 579201
rect 255190 528687 257054 528789
rect 255185 528682 257059 528687
rect 255185 526818 255190 528682
rect 257054 526818 257059 528682
rect 255185 526813 257059 526818
rect -800 34786 102944 34898
rect 102724 34178 102944 34786
rect 110138 518708 249386 518820
rect -800 33604 480 33716
rect 604 32534 690 32577
rect -800 32422 690 32534
rect 604 32376 690 32422
rect 604 32298 717 32376
rect 660 32276 717 32298
rect 817 32276 1034 32376
rect 1134 32276 1140 32376
rect -800 16910 480 17022
rect 110138 16048 110250 518708
rect 262650 500548 265150 578736
rect 265885 578731 266360 578736
rect 137358 498048 265150 500548
rect 137784 441645 139433 498048
rect 269658 496755 272166 587380
rect 125868 439996 139433 441645
rect 139873 496322 272166 496755
rect 274222 595025 276722 666806
rect 274222 592535 274227 595025
rect 275898 592535 276506 592538
rect 276717 592535 276722 595025
rect 139873 496129 272158 496322
rect 125868 133775 127897 439996
rect 139873 439680 140499 496129
rect 269658 496118 272158 496129
rect 274222 494642 276722 592535
rect 282082 581021 284582 677764
rect 315118 608532 316158 685774
rect 331191 627679 332129 697349
rect 415894 693150 418394 702300
rect 427530 693150 427730 703190
rect 465394 702300 470394 704800
rect 415894 690650 456486 693150
rect 427530 688862 427730 690650
rect 331191 626741 432773 627679
rect 315118 607492 416708 608532
rect 308456 594465 308636 594470
rect 308456 594295 308461 594465
rect 308631 594295 347797 594465
rect 308456 594290 308636 594295
rect 288816 592515 289161 592520
rect 288816 592402 288821 592515
rect 288522 592292 288821 592402
rect 288816 592180 288821 592292
rect 289156 592402 289161 592515
rect 289696 592402 289804 592407
rect 289156 592401 289805 592402
rect 289156 592293 289696 592401
rect 289804 592293 289805 592401
rect 289156 592292 289805 592293
rect 289156 592180 289161 592292
rect 289696 592287 289804 592292
rect 288816 592175 289161 592180
rect 338103 592197 338393 592203
rect 338103 591780 338393 591907
rect 338098 591775 338398 591780
rect 338098 591485 338103 591775
rect 338393 591485 338398 591775
rect 338098 591480 338398 591485
rect 338103 591336 338393 591480
rect 338098 591331 338398 591336
rect 338098 591041 338103 591331
rect 338393 591041 338398 591331
rect 338098 591036 338398 591041
rect 338103 590776 338393 591036
rect 337998 590744 338462 590776
rect 337998 590655 338108 590744
rect 338388 590655 338462 590744
rect 287845 590510 288163 590515
rect 287844 590509 288164 590510
rect 287844 590191 287845 590509
rect 288163 590191 288164 590509
rect 287844 590190 288164 590191
rect 337998 590365 338103 590655
rect 338393 590365 338462 590655
rect 337998 590274 338108 590365
rect 338388 590274 338462 590365
rect 287845 590185 288163 590190
rect 337998 590046 338462 590274
rect 338103 586744 338393 590046
rect 338103 586660 338108 586744
rect 338098 586655 338108 586660
rect 338388 586660 338393 586744
rect 338388 586655 338398 586660
rect 338098 586365 338103 586655
rect 338393 586365 338398 586655
rect 338098 586360 338398 586365
rect 347627 585512 347797 594295
rect 347627 585352 347632 585512
rect 347792 585352 347797 585512
rect 347627 585347 347797 585352
rect 293114 581021 293204 584901
rect 282082 580719 293310 581021
rect 282082 576984 284582 580719
rect 293114 579712 293204 580719
rect 289792 579119 290092 579124
rect 286427 579118 290093 579119
rect 286427 579114 289792 579118
rect 286427 578822 286432 579114
rect 286724 578822 289792 579114
rect 286427 578818 289792 578822
rect 290092 578818 290093 579118
rect 286427 578817 290093 578818
rect 289792 578812 290092 578817
rect 308982 578275 309667 578281
rect 308982 577584 309667 577590
rect 282082 574484 291184 576984
rect 332638 575847 333142 575852
rect 332638 575353 332643 575847
rect 333137 575842 372293 575847
rect 333137 575358 371804 575842
rect 372288 575358 372293 575842
rect 333137 575353 372293 575358
rect 332638 575348 333142 575353
rect 141510 493746 276986 494642
rect 141510 441759 142406 493746
rect 274222 493676 276722 493746
rect 288684 490736 291184 574484
rect 291817 571852 292035 571857
rect 291816 571851 292036 571852
rect 291816 571633 291817 571851
rect 292035 571633 292036 571851
rect 291816 571632 292036 571633
rect 291817 571627 292035 571632
rect 291888 570929 292326 571124
rect 291888 570711 291973 570929
rect 292191 570711 292326 570929
rect 291888 570506 292326 570711
rect 292241 568142 292459 568147
rect 292240 568141 292460 568142
rect 292240 567923 292241 568141
rect 292459 567923 292460 568141
rect 292240 567922 292460 567923
rect 292241 567917 292459 567922
rect 148059 489641 291184 490736
rect 141510 441500 141829 441759
rect 142088 441500 142406 441759
rect 141510 440950 142406 441500
rect 148349 441443 148864 489641
rect 150248 478336 151288 484306
rect 152399 478336 153449 478341
rect 149648 477296 152404 478336
rect 153444 477296 153449 478336
rect 150248 442824 151288 477296
rect 152399 477291 153449 477296
rect 288684 473608 291184 489641
rect 343669 486512 344111 486517
rect 343669 486080 343674 486512
rect 344106 486080 344111 486512
rect 343669 486075 344111 486080
rect 291708 477925 291908 477930
rect 291708 477735 291713 477925
rect 291903 477735 291908 477925
rect 153737 472745 154377 473120
rect 288558 472811 288564 473351
rect 289094 473346 289104 473351
rect 289099 472816 289104 473346
rect 289718 473208 290319 473608
rect 289094 472811 289104 472816
rect 153737 472115 153742 472745
rect 154372 472115 154377 472745
rect 150755 442564 151009 442824
rect 151519 442682 151766 442687
rect 153737 442682 154377 472115
rect 289973 471179 290063 473208
rect 291708 472920 291908 477735
rect 343674 475891 344106 486075
rect 415668 478331 416708 607492
rect 415668 477301 415673 478331
rect 416703 477301 416708 478331
rect 415668 477296 416708 477301
rect 343674 475469 343679 475891
rect 344101 475469 344106 475891
rect 343674 475464 344106 475469
rect 431835 475074 432773 626741
rect 444600 575847 445104 575852
rect 453206 575847 455706 690650
rect 461816 585645 462252 585650
rect 466776 585645 469276 702300
rect 510594 698160 515394 704800
rect 520594 698160 525394 704800
rect 566594 702300 571594 704800
rect 566594 690142 571476 702300
rect 554148 689282 571476 690142
rect 547286 669777 548114 669782
rect 561083 669777 561913 689282
rect 566594 674025 571476 689282
rect 574600 682984 582176 683000
rect 574600 682800 584800 682984
rect 574440 682402 584800 682800
rect 574440 678818 575238 682402
rect 582000 678818 584800 682402
rect 574440 678370 584800 678818
rect 582300 677984 584800 678370
rect 547285 669776 561913 669777
rect 547285 668948 547286 669776
rect 548114 668948 561913 669776
rect 566588 669143 566594 674025
rect 571476 669143 571482 674025
rect 547285 668947 561913 668948
rect 547286 668942 548114 668947
rect 534064 644852 543338 645740
rect 534064 639522 535706 644852
rect 541456 644584 543338 644852
rect 541456 639784 584800 644584
rect 541456 639522 543338 639784
rect 534064 639002 543338 639522
rect 534308 634678 543582 635078
rect 534308 629610 536566 634678
rect 541812 634584 543582 634678
rect 541812 629784 584800 634584
rect 541812 629610 543582 629784
rect 534308 628340 543582 629610
rect 577935 629044 578045 629784
rect 577922 629014 578088 629044
rect 577922 628906 577936 629014
rect 578044 628906 578088 629014
rect 577922 628894 578088 628906
rect 577935 625014 578045 628894
rect 577930 624906 577936 625014
rect 578044 624906 578050 625014
rect 577935 624905 578045 624906
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 461816 585219 461821 585645
rect 462247 585219 469276 585645
rect 461816 585214 462252 585219
rect 444600 575353 444605 575847
rect 445099 575353 455706 575847
rect 444600 575348 445104 575353
rect 292218 474979 292418 474984
rect 292218 474789 292223 474979
rect 292413 474789 292418 474979
rect 292218 472964 292418 474789
rect 431835 474146 431840 475074
rect 432768 474146 432773 475074
rect 431835 474141 432773 474146
rect 314131 473946 318929 473951
rect 309338 473945 318930 473946
rect 309338 473941 314131 473945
rect 291188 471179 291278 472125
rect 297396 471945 297406 471950
rect 297396 471575 297401 471945
rect 297396 471570 297406 471575
rect 297776 471570 297782 471950
rect 289973 471089 291278 471179
rect 290873 469712 290883 469717
rect 290873 469072 290878 469712
rect 290873 469067 290883 469072
rect 291523 469067 291529 469717
rect 309338 469151 309343 473941
rect 309338 469147 314131 469151
rect 318929 469147 318930 473945
rect 309338 469146 318930 469147
rect 314131 469141 318929 469146
rect 453206 462143 455706 575353
rect 466776 467039 469276 585219
rect 583520 584744 584800 584856
rect 581085 583562 584800 583674
rect 582340 555352 584800 555362
rect 581085 554285 584800 555352
rect 578987 550570 584800 554285
rect 582340 550562 584800 550570
rect 581085 544277 584800 545362
rect 578987 540562 584800 544277
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 534554 494140 584800 494252
rect 466776 464549 466781 467039
rect 469271 464549 469276 467039
rect 453206 459643 461052 462143
rect 453206 457153 453211 459643
rect 455701 457153 455706 459643
rect 453206 457148 455706 457153
rect 150750 442559 151014 442564
rect 150750 442305 150755 442559
rect 151009 442305 151014 442559
rect 151519 442445 151524 442682
rect 151761 442445 154377 442682
rect 151519 442440 151766 442445
rect 150750 442300 151014 442305
rect 153737 442243 154377 442445
rect 148349 441353 150467 441443
rect 148349 441141 148864 441353
rect 139873 439570 140131 439680
rect 140241 439570 140499 439680
rect 139873 439312 140499 439570
rect 454906 438538 455224 438543
rect 454905 438537 455225 438538
rect 454905 438219 454906 438537
rect 455224 438219 455225 438537
rect 454905 438218 455225 438219
rect 454906 438213 455224 438218
rect 149102 437233 149422 437234
rect 149097 436915 149103 437233
rect 149421 436915 149427 437233
rect 149102 436914 149422 436915
rect 149102 436489 149422 436490
rect 149097 436171 149103 436489
rect 149421 436171 149427 436489
rect 149102 436170 149422 436171
rect 454906 435538 455224 435543
rect 454905 435537 455225 435538
rect 454905 435219 454906 435537
rect 455224 435219 455225 435537
rect 454905 435218 455225 435219
rect 454906 435213 455224 435218
rect 454906 432538 455224 432543
rect 454905 432537 455225 432538
rect 454905 432219 454906 432537
rect 455224 432219 455225 432537
rect 454905 432218 455225 432219
rect 454906 432213 455224 432218
rect 454906 429538 455224 429543
rect 454905 429537 455225 429538
rect 454905 429219 454906 429537
rect 455224 429219 455225 429537
rect 454905 429218 455225 429219
rect 454906 429213 455224 429218
rect 454906 426538 455224 426543
rect 454905 426537 455225 426538
rect 454905 426219 454906 426537
rect 455224 426219 455225 426537
rect 454905 426218 455225 426219
rect 454906 426213 455224 426218
rect 454906 423538 455224 423543
rect 454905 423537 455225 423538
rect 454905 423219 454906 423537
rect 455224 423219 455225 423537
rect 454905 423218 455225 423219
rect 454906 423213 455224 423218
rect 454906 420538 455224 420543
rect 454905 420537 455225 420538
rect 454905 420219 454906 420537
rect 455224 420219 455225 420537
rect 454905 420218 455225 420219
rect 454906 420213 455224 420218
rect 454906 417538 455224 417543
rect 454905 417537 455225 417538
rect 454905 417219 454906 417537
rect 455224 417219 455225 417537
rect 454905 417218 455225 417219
rect 454906 417213 455224 417218
rect 454906 414538 455224 414543
rect 454905 414537 455225 414538
rect 454905 414219 454906 414537
rect 455224 414219 455225 414537
rect 454905 414218 455225 414219
rect 454906 414213 455224 414218
rect 454906 411538 455224 411543
rect 454905 411537 455225 411538
rect 454905 411219 454906 411537
rect 455224 411219 455225 411537
rect 454905 411218 455225 411219
rect 454906 411213 455224 411218
rect 454906 408538 455224 408543
rect 454905 408537 455225 408538
rect 454905 408219 454906 408537
rect 455224 408219 455225 408537
rect 454905 408218 455225 408219
rect 454906 408213 455224 408218
rect 454906 405538 455224 405543
rect 454905 405537 455225 405538
rect 454905 405219 454906 405537
rect 455224 405219 455225 405537
rect 454905 405218 455225 405219
rect 454906 405213 455224 405218
rect 454906 402538 455224 402543
rect 454905 402537 455225 402538
rect 454905 402219 454906 402537
rect 455224 402219 455225 402537
rect 454905 402218 455225 402219
rect 454906 402213 455224 402218
rect 454906 399538 455224 399543
rect 454905 399537 455225 399538
rect 454905 399219 454906 399537
rect 455224 399219 455225 399537
rect 454905 399218 455225 399219
rect 454906 399213 455224 399218
rect 454906 396538 455224 396543
rect 454905 396537 455225 396538
rect 454905 396219 454906 396537
rect 455224 396219 455225 396537
rect 454905 396218 455225 396219
rect 454906 396213 455224 396218
rect 454906 393538 455224 393543
rect 454905 393537 455225 393538
rect 454905 393219 454906 393537
rect 455224 393219 455225 393537
rect 454905 393218 455225 393219
rect 454906 393213 455224 393218
rect 454906 390538 455224 390543
rect 454905 390537 455225 390538
rect 454905 390219 454906 390537
rect 455224 390219 455225 390537
rect 454905 390218 455225 390219
rect 454906 390213 455224 390218
rect 454906 387538 455224 387543
rect 454905 387537 455225 387538
rect 454905 387219 454906 387537
rect 455224 387219 455225 387537
rect 454905 387218 455225 387219
rect 454906 387213 455224 387218
rect 454906 384538 455224 384543
rect 454905 384537 455225 384538
rect 454905 384219 454906 384537
rect 455224 384219 455225 384537
rect 454905 384218 455225 384219
rect 454906 384213 455224 384218
rect 454906 381538 455224 381543
rect 454905 381537 455225 381538
rect 454905 381219 454906 381537
rect 455224 381219 455225 381537
rect 454905 381218 455225 381219
rect 454906 381213 455224 381218
rect 454906 378538 455224 378543
rect 454905 378537 455225 378538
rect 454905 378219 454906 378537
rect 455224 378219 455225 378537
rect 454905 378218 455225 378219
rect 454906 378213 455224 378218
rect 454906 375538 455224 375543
rect 454905 375537 455225 375538
rect 454905 375219 454906 375537
rect 455224 375219 455225 375537
rect 454905 375218 455225 375219
rect 454906 375213 455224 375218
rect 454906 372538 455224 372543
rect 454905 372537 455225 372538
rect 454905 372219 454906 372537
rect 455224 372219 455225 372537
rect 454905 372218 455225 372219
rect 454906 372213 455224 372218
rect 454906 369538 455224 369543
rect 454905 369537 455225 369538
rect 454905 369219 454906 369537
rect 455224 369219 455225 369537
rect 454905 369218 455225 369219
rect 454906 369213 455224 369218
rect 454906 366538 455224 366543
rect 454905 366537 455225 366538
rect 454905 366219 454906 366537
rect 455224 366219 455225 366537
rect 454905 366218 455225 366219
rect 454906 366213 455224 366218
rect 454906 363538 455224 363543
rect 454905 363537 455225 363538
rect 454905 363219 454906 363537
rect 455224 363219 455225 363537
rect 454905 363218 455225 363219
rect 454906 363213 455224 363218
rect 454906 360538 455224 360543
rect 454905 360537 455225 360538
rect 454905 360219 454906 360537
rect 455224 360219 455225 360537
rect 454905 360218 455225 360219
rect 454906 360213 455224 360218
rect 454906 357538 455224 357543
rect 454905 357537 455225 357538
rect 454905 357219 454906 357537
rect 455224 357219 455225 357537
rect 454905 357218 455225 357219
rect 454906 357213 455224 357218
rect 454906 354538 455224 354543
rect 454905 354537 455225 354538
rect 454905 354219 454906 354537
rect 455224 354219 455225 354537
rect 454905 354218 455225 354219
rect 454906 354213 455224 354218
rect 454906 351538 455224 351543
rect 454905 351537 455225 351538
rect 454905 351219 454906 351537
rect 455224 351219 455225 351537
rect 454905 351218 455225 351219
rect 454906 351213 455224 351218
rect 454906 348538 455224 348543
rect 454905 348537 455225 348538
rect 454905 348219 454906 348537
rect 455224 348219 455225 348537
rect 454905 348218 455225 348219
rect 454906 348213 455224 348218
rect 454906 345538 455224 345543
rect 454905 345537 455225 345538
rect 454905 345219 454906 345537
rect 455224 345219 455225 345537
rect 454905 345218 455225 345219
rect 454906 345213 455224 345218
rect 454906 342538 455224 342543
rect 454905 342537 455225 342538
rect 454905 342219 454906 342537
rect 455224 342219 455225 342537
rect 454905 342218 455225 342219
rect 454906 342213 455224 342218
rect 454906 339538 455224 339543
rect 454905 339537 455225 339538
rect 454905 339219 454906 339537
rect 455224 339219 455225 339537
rect 454905 339218 455225 339219
rect 454906 339213 455224 339218
rect 454906 336538 455224 336543
rect 454905 336537 455225 336538
rect 454905 336219 454906 336537
rect 455224 336219 455225 336537
rect 454905 336218 455225 336219
rect 454906 336213 455224 336218
rect 454906 333538 455224 333543
rect 454905 333537 455225 333538
rect 454905 333219 454906 333537
rect 455224 333219 455225 333537
rect 454905 333218 455225 333219
rect 454906 333213 455224 333218
rect 454906 330538 455224 330543
rect 454905 330537 455225 330538
rect 454905 330219 454906 330537
rect 455224 330219 455225 330537
rect 454905 330218 455225 330219
rect 454906 330213 455224 330218
rect 454906 327538 455224 327543
rect 454905 327537 455225 327538
rect 454905 327219 454906 327537
rect 455224 327219 455225 327537
rect 454905 327218 455225 327219
rect 454906 327213 455224 327218
rect 454906 324538 455224 324543
rect 454905 324537 455225 324538
rect 454905 324219 454906 324537
rect 455224 324219 455225 324537
rect 454905 324218 455225 324219
rect 454906 324213 455224 324218
rect 454906 321538 455224 321543
rect 454905 321537 455225 321538
rect 454905 321219 454906 321537
rect 455224 321219 455225 321537
rect 454905 321218 455225 321219
rect 454906 321213 455224 321218
rect 454906 318538 455224 318543
rect 454905 318537 455225 318538
rect 454905 318219 454906 318537
rect 455224 318219 455225 318537
rect 454905 318218 455225 318219
rect 454906 318213 455224 318218
rect 454906 315538 455224 315543
rect 454905 315537 455225 315538
rect 454905 315219 454906 315537
rect 455224 315219 455225 315537
rect 454905 315218 455225 315219
rect 454906 315213 455224 315218
rect 454906 312538 455224 312543
rect 454905 312537 455225 312538
rect 454905 312219 454906 312537
rect 455224 312219 455225 312537
rect 454905 312218 455225 312219
rect 454906 312213 455224 312218
rect 454906 309538 455224 309543
rect 454905 309537 455225 309538
rect 454905 309219 454906 309537
rect 455224 309219 455225 309537
rect 454905 309218 455225 309219
rect 454906 309213 455224 309218
rect 454906 306538 455224 306543
rect 454905 306537 455225 306538
rect 454905 306219 454906 306537
rect 455224 306219 455225 306537
rect 454905 306218 455225 306219
rect 454906 306213 455224 306218
rect 454906 303538 455224 303543
rect 454905 303537 455225 303538
rect 454905 303219 454906 303537
rect 455224 303219 455225 303537
rect 454905 303218 455225 303219
rect 454906 303213 455224 303218
rect 454906 300538 455224 300543
rect 454905 300537 455225 300538
rect 454905 300219 454906 300537
rect 455224 300219 455225 300537
rect 454905 300218 455225 300219
rect 454906 300213 455224 300218
rect 454906 297538 455224 297543
rect 454905 297537 455225 297538
rect 454905 297219 454906 297537
rect 455224 297219 455225 297537
rect 454905 297218 455225 297219
rect 454906 297213 455224 297218
rect 454906 294538 455224 294543
rect 454905 294537 455225 294538
rect 454905 294219 454906 294537
rect 455224 294219 455225 294537
rect 454905 294218 455225 294219
rect 454906 294213 455224 294218
rect 454906 291538 455224 291543
rect 454905 291537 455225 291538
rect 454905 291219 454906 291537
rect 455224 291219 455225 291537
rect 454905 291218 455225 291219
rect 454906 291213 455224 291218
rect 454906 288538 455224 288543
rect 454905 288537 455225 288538
rect 454905 288219 454906 288537
rect 455224 288219 455225 288537
rect 454905 288218 455225 288219
rect 454906 288213 455224 288218
rect 454906 285538 455224 285543
rect 454905 285537 455225 285538
rect 454905 285219 454906 285537
rect 455224 285219 455225 285537
rect 454905 285218 455225 285219
rect 454906 285213 455224 285218
rect 454906 282538 455224 282543
rect 454905 282537 455225 282538
rect 454905 282219 454906 282537
rect 455224 282219 455225 282537
rect 454905 282218 455225 282219
rect 454906 282213 455224 282218
rect 454906 279538 455224 279543
rect 454905 279537 455225 279538
rect 454905 279219 454906 279537
rect 455224 279219 455225 279537
rect 454905 279218 455225 279219
rect 454906 279213 455224 279218
rect 454906 276538 455224 276543
rect 454905 276537 455225 276538
rect 454905 276219 454906 276537
rect 455224 276219 455225 276537
rect 454905 276218 455225 276219
rect 454906 276213 455224 276218
rect 454906 273538 455224 273543
rect 454905 273537 455225 273538
rect 454905 273219 454906 273537
rect 455224 273219 455225 273537
rect 454905 273218 455225 273219
rect 454906 273213 455224 273218
rect 454906 270538 455224 270543
rect 454905 270537 455225 270538
rect 454905 270219 454906 270537
rect 455224 270219 455225 270537
rect 454905 270218 455225 270219
rect 454906 270213 455224 270218
rect 454906 267538 455224 267543
rect 454905 267537 455225 267538
rect 454905 267219 454906 267537
rect 455224 267219 455225 267537
rect 454905 267218 455225 267219
rect 454906 267213 455224 267218
rect 454906 264538 455224 264543
rect 454905 264537 455225 264538
rect 454905 264219 454906 264537
rect 455224 264219 455225 264537
rect 454905 264218 455225 264219
rect 454906 264213 455224 264218
rect 454906 261538 455224 261543
rect 454905 261537 455225 261538
rect 454905 261219 454906 261537
rect 455224 261219 455225 261537
rect 454905 261218 455225 261219
rect 454906 261213 455224 261218
rect 454906 258538 455224 258543
rect 454905 258537 455225 258538
rect 454905 258219 454906 258537
rect 455224 258219 455225 258537
rect 454905 258218 455225 258219
rect 454906 258213 455224 258218
rect 454906 255538 455224 255543
rect 454905 255537 455225 255538
rect 454905 255219 454906 255537
rect 455224 255219 455225 255537
rect 454905 255218 455225 255219
rect 454906 255213 455224 255218
rect 454906 252538 455224 252543
rect 454905 252537 455225 252538
rect 454905 252219 454906 252537
rect 455224 252219 455225 252537
rect 454905 252218 455225 252219
rect 454906 252213 455224 252218
rect 454906 249538 455224 249543
rect 454905 249537 455225 249538
rect 454905 249219 454906 249537
rect 455224 249219 455225 249537
rect 454905 249218 455225 249219
rect 454906 249213 455224 249218
rect 454906 246538 455224 246543
rect 454905 246537 455225 246538
rect 454905 246219 454906 246537
rect 455224 246219 455225 246537
rect 454905 246218 455225 246219
rect 454906 246213 455224 246218
rect 454906 243538 455224 243543
rect 454905 243537 455225 243538
rect 454905 243219 454906 243537
rect 455224 243219 455225 243537
rect 454905 243218 455225 243219
rect 454906 243213 455224 243218
rect 454906 240538 455224 240543
rect 454905 240537 455225 240538
rect 454905 240219 454906 240537
rect 455224 240219 455225 240537
rect 454905 240218 455225 240219
rect 454906 240213 455224 240218
rect 454906 237538 455224 237543
rect 454905 237537 455225 237538
rect 454905 237219 454906 237537
rect 455224 237219 455225 237537
rect 454905 237218 455225 237219
rect 454906 237213 455224 237218
rect 454906 234538 455224 234543
rect 454905 234537 455225 234538
rect 454905 234219 454906 234537
rect 455224 234219 455225 234537
rect 454905 234218 455225 234219
rect 454906 234213 455224 234218
rect 454906 231538 455224 231543
rect 454905 231537 455225 231538
rect 454905 231219 454906 231537
rect 455224 231219 455225 231537
rect 454905 231218 455225 231219
rect 454906 231213 455224 231218
rect 454906 228538 455224 228543
rect 454905 228537 455225 228538
rect 454905 228219 454906 228537
rect 455224 228219 455225 228537
rect 454905 228218 455225 228219
rect 454906 228213 455224 228218
rect 454906 225538 455224 225543
rect 454905 225537 455225 225538
rect 454905 225219 454906 225537
rect 455224 225219 455225 225537
rect 454905 225218 455225 225219
rect 454906 225213 455224 225218
rect 454906 222538 455224 222543
rect 454905 222537 455225 222538
rect 454905 222219 454906 222537
rect 455224 222219 455225 222537
rect 454905 222218 455225 222219
rect 454906 222213 455224 222218
rect 454906 219538 455224 219543
rect 454905 219537 455225 219538
rect 454905 219219 454906 219537
rect 455224 219219 455225 219537
rect 454905 219218 455225 219219
rect 454906 219213 455224 219218
rect 454906 216538 455224 216543
rect 454905 216537 455225 216538
rect 454905 216219 454906 216537
rect 455224 216219 455225 216537
rect 454905 216218 455225 216219
rect 454906 216213 455224 216218
rect 454906 213538 455224 213543
rect 454905 213537 455225 213538
rect 454905 213219 454906 213537
rect 455224 213219 455225 213537
rect 454905 213218 455225 213219
rect 454906 213213 455224 213218
rect 454906 210538 455224 210543
rect 454905 210537 455225 210538
rect 454905 210219 454906 210537
rect 455224 210219 455225 210537
rect 454905 210218 455225 210219
rect 454906 210213 455224 210218
rect 454906 207538 455224 207543
rect 454905 207537 455225 207538
rect 454905 207219 454906 207537
rect 455224 207219 455225 207537
rect 454905 207218 455225 207219
rect 454906 207213 455224 207218
rect 454906 204538 455224 204543
rect 454905 204537 455225 204538
rect 454905 204219 454906 204537
rect 455224 204219 455225 204537
rect 454905 204218 455225 204219
rect 454906 204213 455224 204218
rect 454906 201538 455224 201543
rect 454905 201537 455225 201538
rect 454905 201219 454906 201537
rect 455224 201219 455225 201537
rect 454905 201218 455225 201219
rect 454906 201213 455224 201218
rect 454906 198538 455224 198543
rect 454905 198537 455225 198538
rect 454905 198219 454906 198537
rect 455224 198219 455225 198537
rect 454905 198218 455225 198219
rect 454906 198213 455224 198218
rect 454906 195538 455224 195543
rect 454905 195537 455225 195538
rect 454905 195219 454906 195537
rect 455224 195219 455225 195537
rect 454905 195218 455225 195219
rect 454906 195213 455224 195218
rect 454906 192538 455224 192543
rect 454905 192537 455225 192538
rect 454905 192219 454906 192537
rect 455224 192219 455225 192537
rect 454905 192218 455225 192219
rect 454906 192213 455224 192218
rect 454906 189538 455224 189543
rect 454905 189537 455225 189538
rect 454905 189219 454906 189537
rect 455224 189219 455225 189537
rect 454905 189218 455225 189219
rect 454906 189213 455224 189218
rect 454906 186538 455224 186543
rect 454905 186537 455225 186538
rect 454905 186219 454906 186537
rect 455224 186219 455225 186537
rect 454905 186218 455225 186219
rect 454906 186213 455224 186218
rect 454906 183538 455224 183543
rect 454905 183537 455225 183538
rect 454905 183219 454906 183537
rect 455224 183219 455225 183537
rect 454905 183218 455225 183219
rect 454906 183213 455224 183218
rect 454906 180538 455224 180543
rect 454905 180537 455225 180538
rect 454905 180219 454906 180537
rect 455224 180219 455225 180537
rect 454905 180218 455225 180219
rect 454906 180213 455224 180218
rect 454906 177538 455224 177543
rect 454905 177537 455225 177538
rect 454905 177219 454906 177537
rect 455224 177219 455225 177537
rect 454905 177218 455225 177219
rect 454906 177213 455224 177218
rect 454906 174538 455224 174543
rect 454905 174537 455225 174538
rect 454905 174219 454906 174537
rect 455224 174219 455225 174537
rect 454905 174218 455225 174219
rect 454906 174213 455224 174218
rect 454906 171538 455224 171543
rect 454905 171537 455225 171538
rect 454905 171219 454906 171537
rect 455224 171219 455225 171537
rect 454905 171218 455225 171219
rect 454906 171213 455224 171218
rect 454906 168538 455224 168543
rect 454905 168537 455225 168538
rect 454905 168219 454906 168537
rect 455224 168219 455225 168537
rect 454905 168218 455225 168219
rect 454906 168213 455224 168218
rect 454906 165538 455224 165543
rect 454905 165537 455225 165538
rect 454905 165219 454906 165537
rect 455224 165219 455225 165537
rect 454905 165218 455225 165219
rect 454906 165213 455224 165218
rect 454906 162538 455224 162543
rect 454905 162537 455225 162538
rect 454905 162219 454906 162537
rect 455224 162219 455225 162537
rect 454905 162218 455225 162219
rect 454906 162213 455224 162218
rect 454906 159538 455224 159543
rect 454905 159537 455225 159538
rect 454905 159219 454906 159537
rect 455224 159219 455225 159537
rect 454905 159218 455225 159219
rect 454906 159213 455224 159218
rect 454906 156538 455224 156543
rect 454905 156537 455225 156538
rect 454905 156219 454906 156537
rect 455224 156219 455225 156537
rect 454905 156218 455225 156219
rect 454906 156213 455224 156218
rect 454906 153538 455224 153543
rect 454905 153537 455225 153538
rect 454905 153219 454906 153537
rect 455224 153219 455225 153537
rect 454905 153218 455225 153219
rect 454906 153213 455224 153218
rect 454906 150538 455224 150543
rect 454905 150537 455225 150538
rect 454905 150219 454906 150537
rect 455224 150219 455225 150537
rect 454905 150218 455225 150219
rect 454906 150213 455224 150218
rect 125868 132697 126341 133775
rect 127419 132697 127897 133775
rect 125868 129154 127897 132697
rect 125868 128636 126336 129154
rect 126331 128066 126336 128636
rect 127424 128636 127897 129154
rect 127424 128066 127429 128636
rect 126331 128061 127429 128066
rect 130313 124893 130433 131530
rect 130313 124783 130318 124893
rect 130428 124783 130433 124893
rect 130313 124778 130433 124783
rect 134257 120765 134377 131548
rect 134257 120655 134262 120765
rect 134372 120655 134377 120765
rect 134257 120650 134377 120655
rect 138337 120173 138457 131448
rect 138337 120063 138342 120173
rect 138452 120063 138457 120173
rect 138337 120058 138457 120063
rect 142281 118681 142401 131424
rect 144647 129154 145733 129159
rect 144646 129153 145734 129154
rect 144646 128067 144647 129153
rect 145733 128067 145734 129153
rect 460671 128899 460841 459643
rect 466776 459040 469276 464549
rect 461524 456540 469276 459040
rect 461823 139833 462269 456540
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 534554 449718 584800 449830
rect 515375 438538 515385 438543
rect 515375 438218 515380 438538
rect 515375 438213 515385 438218
rect 515705 438213 515711 438543
rect 515375 435538 515385 435543
rect 515375 435218 515380 435538
rect 515375 435213 515385 435218
rect 515705 435213 515711 435543
rect 515375 432538 515385 432543
rect 515375 432218 515380 432538
rect 515375 432213 515385 432218
rect 515705 432213 515711 432543
rect 515375 429538 515385 429543
rect 515375 429218 515380 429538
rect 515375 429213 515385 429218
rect 515705 429213 515711 429543
rect 515375 426538 515385 426543
rect 515375 426218 515380 426538
rect 515375 426213 515385 426218
rect 515705 426213 515711 426543
rect 515375 423538 515385 423543
rect 515375 423218 515380 423538
rect 515375 423213 515385 423218
rect 515705 423213 515711 423543
rect 515375 420538 515385 420543
rect 515375 420218 515380 420538
rect 515375 420213 515385 420218
rect 515705 420213 515711 420543
rect 515375 417538 515385 417543
rect 515375 417218 515380 417538
rect 515375 417213 515385 417218
rect 515705 417213 515711 417543
rect 515375 414538 515385 414543
rect 515375 414218 515380 414538
rect 515375 414213 515385 414218
rect 515705 414213 515711 414543
rect 515375 411538 515385 411543
rect 515375 411218 515380 411538
rect 515375 411213 515385 411218
rect 515705 411213 515711 411543
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 515375 408538 515385 408543
rect 515375 408218 515380 408538
rect 515375 408213 515385 408218
rect 515705 408213 515711 408543
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 515375 405538 515385 405543
rect 515375 405218 515380 405538
rect 515375 405213 515385 405218
rect 515705 405213 515711 405543
rect 583520 405296 584800 405408
rect 515375 402538 515385 402543
rect 515375 402218 515380 402538
rect 515375 402213 515385 402218
rect 515705 402213 515711 402543
rect 515375 399538 515385 399543
rect 515375 399218 515380 399538
rect 515375 399213 515385 399218
rect 515705 399213 515711 399543
rect 515375 396538 515385 396543
rect 515375 396218 515380 396538
rect 515375 396213 515385 396218
rect 515705 396213 515711 396543
rect 515375 393538 515385 393543
rect 515375 393218 515380 393538
rect 515375 393213 515385 393218
rect 515705 393213 515711 393543
rect 515375 390538 515385 390543
rect 515375 390218 515380 390538
rect 515375 390213 515385 390218
rect 515705 390213 515711 390543
rect 515375 387538 515385 387543
rect 515375 387218 515380 387538
rect 515375 387213 515385 387218
rect 515705 387213 515711 387543
rect 515375 384538 515385 384543
rect 515375 384218 515380 384538
rect 515375 384213 515385 384218
rect 515705 384213 515711 384543
rect 515375 381538 515385 381543
rect 515375 381218 515380 381538
rect 515375 381213 515385 381218
rect 515705 381213 515711 381543
rect 515375 378538 515385 378543
rect 515375 378218 515380 378538
rect 515375 378213 515385 378218
rect 515705 378213 515711 378543
rect 515375 375538 515385 375543
rect 515375 375218 515380 375538
rect 515375 375213 515385 375218
rect 515705 375213 515711 375543
rect 515375 372538 515385 372543
rect 515375 372218 515380 372538
rect 515375 372213 515385 372218
rect 515705 372213 515711 372543
rect 515375 369538 515385 369543
rect 515375 369218 515380 369538
rect 515375 369213 515385 369218
rect 515705 369213 515711 369543
rect 582538 368886 582656 368894
rect 582538 368786 582546 368886
rect 582646 368786 582656 368886
rect 582538 368778 582656 368786
rect 515375 366538 515385 366543
rect 515375 366218 515380 366538
rect 515375 366213 515385 366218
rect 515705 366213 515711 366543
rect 582476 364801 582546 364886
rect 582482 364786 582546 364801
rect 582646 364786 582787 364886
rect 582918 364784 584800 364896
rect 583520 363602 584800 363714
rect 515375 363538 515385 363543
rect 515375 363218 515380 363538
rect 515375 363213 515385 363218
rect 515705 363213 515711 363543
rect 534554 362420 584800 362532
rect 515375 360538 515385 360543
rect 515375 360218 515380 360538
rect 515375 360213 515385 360218
rect 515705 360213 515711 360543
rect 515375 357538 515385 357543
rect 515375 357218 515380 357538
rect 515375 357213 515385 357218
rect 515705 357213 515711 357543
rect 515375 354538 515385 354543
rect 515375 354218 515380 354538
rect 515375 354213 515385 354218
rect 515705 354213 515711 354543
rect 515375 351538 515385 351543
rect 515375 351218 515380 351538
rect 515375 351213 515385 351218
rect 515705 351213 515711 351543
rect 515375 348538 515385 348543
rect 515375 348218 515380 348538
rect 515375 348213 515385 348218
rect 515705 348213 515711 348543
rect 515375 345538 515385 345543
rect 515375 345218 515380 345538
rect 515375 345213 515385 345218
rect 515705 345213 515711 345543
rect 515375 342538 515385 342543
rect 515375 342218 515380 342538
rect 515375 342213 515385 342218
rect 515705 342213 515711 342543
rect 515375 339538 515385 339543
rect 515375 339218 515380 339538
rect 515375 339213 515385 339218
rect 515705 339213 515711 339543
rect 515375 336538 515385 336543
rect 515375 336218 515380 336538
rect 515375 336213 515385 336218
rect 515705 336213 515711 336543
rect 515375 333538 515385 333543
rect 515375 333218 515380 333538
rect 515375 333213 515385 333218
rect 515705 333213 515711 333543
rect 515375 330538 515385 330543
rect 515375 330218 515380 330538
rect 515375 330213 515385 330218
rect 515705 330213 515711 330543
rect 515375 327538 515385 327543
rect 515375 327218 515380 327538
rect 515375 327213 515385 327218
rect 515705 327213 515711 327543
rect 515375 324538 515385 324543
rect 515375 324218 515380 324538
rect 515375 324213 515385 324218
rect 515705 324213 515711 324543
rect 515375 321538 515385 321543
rect 515375 321218 515380 321538
rect 515375 321213 515385 321218
rect 515705 321213 515711 321543
rect 515375 318538 515385 318543
rect 515375 318218 515380 318538
rect 515375 318213 515385 318218
rect 515705 318213 515711 318543
rect 515375 315538 515385 315543
rect 515375 315218 515380 315538
rect 515375 315213 515385 315218
rect 515705 315213 515711 315543
rect 515375 312538 515385 312543
rect 515375 312218 515380 312538
rect 515375 312213 515385 312218
rect 515705 312213 515711 312543
rect 515375 309538 515385 309543
rect 515375 309218 515380 309538
rect 515375 309213 515385 309218
rect 515705 309213 515711 309543
rect 515375 306538 515385 306543
rect 515375 306218 515380 306538
rect 515375 306213 515385 306218
rect 515705 306213 515711 306543
rect 515375 303538 515385 303543
rect 515375 303218 515380 303538
rect 515375 303213 515385 303218
rect 515705 303213 515711 303543
rect 515375 300538 515385 300543
rect 515375 300218 515380 300538
rect 515375 300213 515385 300218
rect 515705 300213 515711 300543
rect 515375 297538 515385 297543
rect 515375 297218 515380 297538
rect 515375 297213 515385 297218
rect 515705 297213 515711 297543
rect 515375 294538 515385 294543
rect 515375 294218 515380 294538
rect 515375 294213 515385 294218
rect 515705 294213 515711 294543
rect 515375 291538 515385 291543
rect 515375 291218 515380 291538
rect 515375 291213 515385 291218
rect 515705 291213 515711 291543
rect 515375 288538 515385 288543
rect 515375 288218 515380 288538
rect 515375 288213 515385 288218
rect 515705 288213 515711 288543
rect 515375 285538 515385 285543
rect 515375 285218 515380 285538
rect 515375 285213 515385 285218
rect 515705 285213 515711 285543
rect 515375 282538 515385 282543
rect 515375 282218 515380 282538
rect 515375 282213 515385 282218
rect 515705 282213 515711 282543
rect 515375 279538 515385 279543
rect 515375 279218 515380 279538
rect 515375 279213 515385 279218
rect 515705 279213 515711 279543
rect 515375 276538 515385 276543
rect 515375 276218 515380 276538
rect 515375 276213 515385 276218
rect 515705 276213 515711 276543
rect 515375 273538 515385 273543
rect 515375 273218 515380 273538
rect 515375 273213 515385 273218
rect 515705 273213 515711 273543
rect 515375 270538 515385 270543
rect 515375 270218 515380 270538
rect 515375 270213 515385 270218
rect 515705 270213 515711 270543
rect 515375 267538 515385 267543
rect 515375 267218 515380 267538
rect 515375 267213 515385 267218
rect 515705 267213 515711 267543
rect 515375 264538 515385 264543
rect 515375 264218 515380 264538
rect 515375 264213 515385 264218
rect 515705 264213 515711 264543
rect 515375 261538 515385 261543
rect 515375 261218 515380 261538
rect 515375 261213 515385 261218
rect 515705 261213 515711 261543
rect 515375 258538 515385 258543
rect 515375 258218 515380 258538
rect 515375 258213 515385 258218
rect 515705 258213 515711 258543
rect 515375 255538 515385 255543
rect 515375 255218 515380 255538
rect 515375 255213 515385 255218
rect 515705 255213 515711 255543
rect 515375 252538 515385 252543
rect 515375 252218 515380 252538
rect 515375 252213 515385 252218
rect 515705 252213 515711 252543
rect 515375 249538 515385 249543
rect 515375 249218 515380 249538
rect 515375 249213 515385 249218
rect 515705 249213 515711 249543
rect 515375 246538 515385 246543
rect 515375 246218 515380 246538
rect 515375 246213 515385 246218
rect 515705 246213 515711 246543
rect 515375 243538 515385 243543
rect 515375 243218 515380 243538
rect 515375 243213 515385 243218
rect 515705 243213 515711 243543
rect 515375 240538 515385 240543
rect 515375 240218 515380 240538
rect 515375 240213 515385 240218
rect 515705 240213 515711 240543
rect 515375 237538 515385 237543
rect 515375 237218 515380 237538
rect 515375 237213 515385 237218
rect 515705 237213 515711 237543
rect 515375 234538 515385 234543
rect 515375 234218 515380 234538
rect 515375 234213 515385 234218
rect 515705 234213 515711 234543
rect 515375 231538 515385 231543
rect 515375 231218 515380 231538
rect 515375 231213 515385 231218
rect 515705 231213 515711 231543
rect 515375 228538 515385 228543
rect 515375 228218 515380 228538
rect 515375 228213 515385 228218
rect 515705 228213 515711 228543
rect 515375 225538 515385 225543
rect 515375 225218 515380 225538
rect 515375 225213 515385 225218
rect 515705 225213 515711 225543
rect 515375 222538 515385 222543
rect 515375 222218 515380 222538
rect 515375 222213 515385 222218
rect 515705 222213 515711 222543
rect 515375 219538 515385 219543
rect 515375 219218 515380 219538
rect 515375 219213 515385 219218
rect 515705 219213 515711 219543
rect 515375 216538 515385 216543
rect 515375 216218 515380 216538
rect 515375 216213 515385 216218
rect 515705 216213 515711 216543
rect 515375 213538 515385 213543
rect 515375 213218 515380 213538
rect 515375 213213 515385 213218
rect 515705 213213 515711 213543
rect 515375 210538 515385 210543
rect 515375 210218 515380 210538
rect 515375 210213 515385 210218
rect 515705 210213 515711 210543
rect 515375 207538 515385 207543
rect 515375 207218 515380 207538
rect 515375 207213 515385 207218
rect 515705 207213 515711 207543
rect 515375 204538 515385 204543
rect 515375 204218 515380 204538
rect 515375 204213 515385 204218
rect 515705 204213 515711 204543
rect 515375 201538 515385 201543
rect 515375 201218 515380 201538
rect 515375 201213 515385 201218
rect 515705 201213 515711 201543
rect 515375 198538 515385 198543
rect 515375 198218 515380 198538
rect 515375 198213 515385 198218
rect 515705 198213 515711 198543
rect 515375 195538 515385 195543
rect 515375 195218 515380 195538
rect 515375 195213 515385 195218
rect 515705 195213 515711 195543
rect 515375 192538 515385 192543
rect 515375 192218 515380 192538
rect 515375 192213 515385 192218
rect 515705 192213 515711 192543
rect 515375 189538 515385 189543
rect 515375 189218 515380 189538
rect 515375 189213 515385 189218
rect 515705 189213 515711 189543
rect 515375 186538 515385 186543
rect 515375 186218 515380 186538
rect 515375 186213 515385 186218
rect 515705 186213 515711 186543
rect 515375 183538 515385 183543
rect 515375 183218 515380 183538
rect 515375 183213 515385 183218
rect 515705 183213 515711 183543
rect 515375 180538 515385 180543
rect 515375 180218 515380 180538
rect 515375 180213 515385 180218
rect 515705 180213 515711 180543
rect 515375 177538 515385 177543
rect 515375 177218 515380 177538
rect 515375 177213 515385 177218
rect 515705 177213 515711 177543
rect 515375 174538 515385 174543
rect 515375 174218 515380 174538
rect 515375 174213 515385 174218
rect 515705 174213 515711 174543
rect 515375 171538 515385 171543
rect 515375 171218 515380 171538
rect 515375 171213 515385 171218
rect 515705 171213 515711 171543
rect 515375 168538 515385 168543
rect 515375 168218 515380 168538
rect 515375 168213 515385 168218
rect 515705 168213 515711 168543
rect 515375 165538 515385 165543
rect 515375 165218 515380 165538
rect 515375 165213 515385 165218
rect 515705 165213 515711 165543
rect 515375 162538 515385 162543
rect 515375 162218 515380 162538
rect 515375 162213 515385 162218
rect 515705 162213 515711 162543
rect 515375 159538 515385 159543
rect 515375 159218 515380 159538
rect 515375 159213 515385 159218
rect 515705 159213 515711 159543
rect 515375 156538 515385 156543
rect 515375 156218 515380 156538
rect 515375 156213 515385 156218
rect 515705 156213 515711 156543
rect 515375 153538 515385 153543
rect 515375 153218 515380 153538
rect 515375 153213 515385 153218
rect 515705 153213 515711 153543
rect 515375 150538 515385 150543
rect 515375 150218 515380 150538
rect 515375 150213 515385 150218
rect 515705 150213 515711 150543
rect 503116 141266 504528 141271
rect 499369 139852 499375 141266
rect 500789 141265 504529 141266
rect 500789 140997 503116 141265
rect 500789 140121 501754 140997
rect 502630 140121 503116 140997
rect 500789 139853 503116 140121
rect 504528 140997 504529 141265
rect 504528 140121 505628 140997
rect 506504 140121 506510 140997
rect 504528 139853 504529 140121
rect 500789 139852 504529 139853
rect 503116 139847 504528 139852
rect 461823 139663 461961 139833
rect 462131 139663 462269 139833
rect 461823 139525 462269 139663
rect 460666 128894 460846 128899
rect 456132 128660 458042 128780
rect 460666 128724 460671 128894
rect 460841 128724 460846 128894
rect 460666 128719 460846 128724
rect 144646 128066 145734 128067
rect 144647 128061 145733 128066
rect 457922 126066 458042 128660
rect 463525 126465 463531 127150
rect 464216 126465 464222 127150
rect 534554 126066 534666 362420
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583093 358874 584800 358986
rect 542712 344507 542832 344508
rect 542640 344387 570754 344507
rect 457922 125946 534814 126066
rect 542712 124836 542832 344387
rect 570634 317310 570754 344387
rect 582536 323646 582660 323652
rect 582536 323546 582546 323646
rect 582646 323546 582660 323646
rect 582536 323540 582660 323546
rect 583138 319656 584800 319674
rect 582918 319646 584800 319656
rect 582476 319561 582546 319646
rect 582482 319546 582546 319561
rect 582646 319546 582787 319646
rect 582887 319562 584800 319646
rect 582887 319546 583364 319562
rect 582918 319544 583364 319546
rect 583520 318380 584800 318492
rect 570463 317198 584800 317310
rect 570634 316193 570754 317198
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 581256 313652 584800 313764
rect 582536 279246 582654 279250
rect 582536 279146 582546 279246
rect 582646 279146 582654 279246
rect 582536 279140 582654 279146
rect 456202 124716 542832 124836
rect 544022 276244 580683 276364
rect 544022 120756 544142 276244
rect 580563 272888 580683 276244
rect 582918 275252 583364 275256
rect 582918 275246 584800 275252
rect 582476 275161 582546 275246
rect 582482 275146 582546 275161
rect 582646 275146 582787 275246
rect 582887 275146 584800 275246
rect 582918 275144 584800 275146
rect 583156 275140 584800 275144
rect 583520 273958 584800 274070
rect 580563 272776 584800 272888
rect 580563 272105 580683 272776
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 582310 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 578645 198242 579069 198298
rect 552812 196966 579468 198242
rect 552812 196230 554140 196966
rect 550944 191768 554140 196230
rect 578296 196230 579468 196966
rect 578296 191768 584800 196230
rect 550944 191430 584800 191768
rect 552812 190928 579468 191430
rect 553276 187154 558076 190928
rect 551320 186340 579660 187154
rect 551320 186230 553050 186340
rect 550944 181430 553050 186230
rect 551320 181150 553050 181430
rect 576862 186230 579660 186340
rect 576862 181430 584800 186230
rect 576862 181150 579660 181430
rect 551320 180540 579660 181150
rect 553276 164626 558076 180540
rect 552718 164209 558786 164626
rect 552718 159411 553277 164209
rect 558075 159411 558786 164209
rect 552718 158880 558786 159411
rect 582340 149347 584800 151630
rect 576060 146887 584800 149347
rect 582340 146830 584800 146887
rect 582340 139290 584800 141630
rect 576060 136830 584800 139290
rect 456280 120636 544278 120756
rect 544022 120620 544142 120636
rect 461464 119798 571679 119918
rect 142281 118571 142286 118681
rect 142396 118571 142401 118681
rect 142281 118566 142401 118571
rect 461620 116812 461740 119798
rect 456242 116692 461740 116812
rect 571559 92866 571679 119798
rect 582532 99246 582656 99252
rect 582532 99146 582546 99246
rect 582646 99146 582656 99246
rect 582532 99138 582656 99146
rect 582918 95246 583364 95256
rect 582476 95161 582546 95246
rect 582482 95146 582546 95161
rect 582646 95146 582787 95246
rect 582887 95230 583364 95246
rect 582887 95146 584800 95230
rect 582918 95144 584800 95146
rect 583184 95118 584800 95144
rect 583520 93936 584800 94048
rect 570398 92754 584800 92866
rect 571559 89505 571679 92754
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 583520 16910 584800 17022
rect 10662 15936 110250 16048
rect -800 15728 480 15840
rect -800 14546 480 14658
rect 10662 13476 10774 15936
rect 583520 15728 584800 15840
rect 583520 14546 584800 14658
rect -800 13364 10882 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11010 674 11112
rect -800 11000 690 11010
rect 583520 11000 584800 11112
rect 562 10976 690 11000
rect 562 10876 717 10976
rect 817 10876 1034 10976
rect 1134 10876 1140 10976
rect 562 10868 674 10876
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 1849 8748
rect 583520 8636 584800 8748
rect -800 7454 584 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 354 4020
rect 466 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 717 419176 817 419276
rect 717 375976 817 376076
rect 717 332676 817 332776
rect 717 289476 817 289576
rect 717 246476 817 246576
rect 717 118876 817 118976
rect 717 75676 817 75776
rect 717 32276 817 32376
rect 582787 319546 582887 319646
rect 582787 275146 582887 275246
rect 582787 95146 582887 95246
rect 717 10876 817 10976
<< via3 >>
rect 228439 697491 229477 698529
rect 331192 697349 332128 698285
rect 1034 462376 1134 462476
rect 1034 419176 1134 419276
rect 1034 375976 1134 376076
rect 1034 332676 1134 332776
rect 5660 293269 5772 293381
rect 1034 289476 1134 289576
rect 8382 261315 8462 261320
rect 8382 261250 8387 261315
rect 8387 261250 8457 261315
rect 8457 261250 8462 261315
rect 24559 260405 24677 260523
rect 27251 258855 27369 258973
rect 19139 253217 19257 253335
rect 21327 253223 21445 253341
rect 5661 253062 5771 253172
rect 19138 247228 19258 247348
rect 1034 246476 1134 246576
rect 10674 191427 10784 191537
rect 9011 191337 9131 191342
rect 9011 191232 9016 191337
rect 9016 191232 9126 191337
rect 9126 191232 9131 191337
rect 21326 247432 21446 247552
rect 24558 245442 24678 245562
rect 27250 244706 27370 244826
rect 1034 118876 1134 118976
rect 1034 75676 1134 75776
rect 1034 32276 1134 32376
rect 289696 592293 289804 592401
rect 338103 591907 338393 592197
rect 287845 590505 288163 590509
rect 287845 590195 287849 590505
rect 287849 590195 288159 590505
rect 288159 590195 288163 590505
rect 287845 590191 288163 590195
rect 289792 578818 290092 579118
rect 308982 577590 309667 578275
rect 291817 571847 292035 571851
rect 291817 571637 291821 571847
rect 291821 571637 292031 571847
rect 292031 571637 292035 571847
rect 291817 571633 292035 571637
rect 291973 570925 292191 570929
rect 291973 570715 291977 570925
rect 291977 570715 292187 570925
rect 292187 570715 292191 570925
rect 291973 570711 292191 570715
rect 292241 568137 292459 568141
rect 292241 567927 292245 568137
rect 292245 567927 292455 568137
rect 292455 567927 292459 568137
rect 292241 567923 292459 567927
rect 141829 441500 142088 441759
rect 288564 473346 289094 473351
rect 288564 472816 288569 473346
rect 288569 472816 289094 473346
rect 288564 472811 289094 472816
rect 575238 678818 582000 682402
rect 547286 668948 548114 669776
rect 566594 669143 571476 674025
rect 535706 639522 541456 644852
rect 536566 629610 541812 634678
rect 577936 628906 578044 629014
rect 577936 624906 578044 625014
rect 314131 473941 318929 473945
rect 297406 471945 297776 471950
rect 297406 471575 297771 471945
rect 297771 471575 297776 471945
rect 297406 471570 297776 471575
rect 290883 469712 291523 469717
rect 290883 469072 291518 469712
rect 291518 469072 291523 469712
rect 290883 469067 291523 469072
rect 314131 469151 314133 473941
rect 314133 469151 318929 473941
rect 314131 469147 318929 469151
rect 454906 438533 455224 438537
rect 454906 438223 454910 438533
rect 454910 438223 455220 438533
rect 455220 438223 455224 438533
rect 454906 438219 455224 438223
rect 149103 437229 149421 437233
rect 149103 436919 149107 437229
rect 149107 436919 149417 437229
rect 149417 436919 149421 437229
rect 149103 436915 149421 436919
rect 149103 436485 149421 436489
rect 149103 436175 149107 436485
rect 149107 436175 149417 436485
rect 149417 436175 149421 436485
rect 149103 436171 149421 436175
rect 454906 435533 455224 435537
rect 454906 435223 454910 435533
rect 454910 435223 455220 435533
rect 455220 435223 455224 435533
rect 454906 435219 455224 435223
rect 454906 432533 455224 432537
rect 454906 432223 454910 432533
rect 454910 432223 455220 432533
rect 455220 432223 455224 432533
rect 454906 432219 455224 432223
rect 454906 429533 455224 429537
rect 454906 429223 454910 429533
rect 454910 429223 455220 429533
rect 455220 429223 455224 429533
rect 454906 429219 455224 429223
rect 454906 426533 455224 426537
rect 454906 426223 454910 426533
rect 454910 426223 455220 426533
rect 455220 426223 455224 426533
rect 454906 426219 455224 426223
rect 454906 423533 455224 423537
rect 454906 423223 454910 423533
rect 454910 423223 455220 423533
rect 455220 423223 455224 423533
rect 454906 423219 455224 423223
rect 454906 420533 455224 420537
rect 454906 420223 454910 420533
rect 454910 420223 455220 420533
rect 455220 420223 455224 420533
rect 454906 420219 455224 420223
rect 454906 417533 455224 417537
rect 454906 417223 454910 417533
rect 454910 417223 455220 417533
rect 455220 417223 455224 417533
rect 454906 417219 455224 417223
rect 454906 414533 455224 414537
rect 454906 414223 454910 414533
rect 454910 414223 455220 414533
rect 455220 414223 455224 414533
rect 454906 414219 455224 414223
rect 454906 411533 455224 411537
rect 454906 411223 454910 411533
rect 454910 411223 455220 411533
rect 455220 411223 455224 411533
rect 454906 411219 455224 411223
rect 454906 408533 455224 408537
rect 454906 408223 454910 408533
rect 454910 408223 455220 408533
rect 455220 408223 455224 408533
rect 454906 408219 455224 408223
rect 454906 405533 455224 405537
rect 454906 405223 454910 405533
rect 454910 405223 455220 405533
rect 455220 405223 455224 405533
rect 454906 405219 455224 405223
rect 454906 402533 455224 402537
rect 454906 402223 454910 402533
rect 454910 402223 455220 402533
rect 455220 402223 455224 402533
rect 454906 402219 455224 402223
rect 454906 399533 455224 399537
rect 454906 399223 454910 399533
rect 454910 399223 455220 399533
rect 455220 399223 455224 399533
rect 454906 399219 455224 399223
rect 454906 396533 455224 396537
rect 454906 396223 454910 396533
rect 454910 396223 455220 396533
rect 455220 396223 455224 396533
rect 454906 396219 455224 396223
rect 454906 393533 455224 393537
rect 454906 393223 454910 393533
rect 454910 393223 455220 393533
rect 455220 393223 455224 393533
rect 454906 393219 455224 393223
rect 454906 390533 455224 390537
rect 454906 390223 454910 390533
rect 454910 390223 455220 390533
rect 455220 390223 455224 390533
rect 454906 390219 455224 390223
rect 454906 387533 455224 387537
rect 454906 387223 454910 387533
rect 454910 387223 455220 387533
rect 455220 387223 455224 387533
rect 454906 387219 455224 387223
rect 454906 384533 455224 384537
rect 454906 384223 454910 384533
rect 454910 384223 455220 384533
rect 455220 384223 455224 384533
rect 454906 384219 455224 384223
rect 454906 381533 455224 381537
rect 454906 381223 454910 381533
rect 454910 381223 455220 381533
rect 455220 381223 455224 381533
rect 454906 381219 455224 381223
rect 454906 378533 455224 378537
rect 454906 378223 454910 378533
rect 454910 378223 455220 378533
rect 455220 378223 455224 378533
rect 454906 378219 455224 378223
rect 454906 375533 455224 375537
rect 454906 375223 454910 375533
rect 454910 375223 455220 375533
rect 455220 375223 455224 375533
rect 454906 375219 455224 375223
rect 454906 372533 455224 372537
rect 454906 372223 454910 372533
rect 454910 372223 455220 372533
rect 455220 372223 455224 372533
rect 454906 372219 455224 372223
rect 454906 369533 455224 369537
rect 454906 369223 454910 369533
rect 454910 369223 455220 369533
rect 455220 369223 455224 369533
rect 454906 369219 455224 369223
rect 454906 366533 455224 366537
rect 454906 366223 454910 366533
rect 454910 366223 455220 366533
rect 455220 366223 455224 366533
rect 454906 366219 455224 366223
rect 454906 363533 455224 363537
rect 454906 363223 454910 363533
rect 454910 363223 455220 363533
rect 455220 363223 455224 363533
rect 454906 363219 455224 363223
rect 454906 360533 455224 360537
rect 454906 360223 454910 360533
rect 454910 360223 455220 360533
rect 455220 360223 455224 360533
rect 454906 360219 455224 360223
rect 454906 357533 455224 357537
rect 454906 357223 454910 357533
rect 454910 357223 455220 357533
rect 455220 357223 455224 357533
rect 454906 357219 455224 357223
rect 454906 354533 455224 354537
rect 454906 354223 454910 354533
rect 454910 354223 455220 354533
rect 455220 354223 455224 354533
rect 454906 354219 455224 354223
rect 454906 351533 455224 351537
rect 454906 351223 454910 351533
rect 454910 351223 455220 351533
rect 455220 351223 455224 351533
rect 454906 351219 455224 351223
rect 454906 348533 455224 348537
rect 454906 348223 454910 348533
rect 454910 348223 455220 348533
rect 455220 348223 455224 348533
rect 454906 348219 455224 348223
rect 454906 345533 455224 345537
rect 454906 345223 454910 345533
rect 454910 345223 455220 345533
rect 455220 345223 455224 345533
rect 454906 345219 455224 345223
rect 454906 342533 455224 342537
rect 454906 342223 454910 342533
rect 454910 342223 455220 342533
rect 455220 342223 455224 342533
rect 454906 342219 455224 342223
rect 454906 339533 455224 339537
rect 454906 339223 454910 339533
rect 454910 339223 455220 339533
rect 455220 339223 455224 339533
rect 454906 339219 455224 339223
rect 454906 336533 455224 336537
rect 454906 336223 454910 336533
rect 454910 336223 455220 336533
rect 455220 336223 455224 336533
rect 454906 336219 455224 336223
rect 454906 333533 455224 333537
rect 454906 333223 454910 333533
rect 454910 333223 455220 333533
rect 455220 333223 455224 333533
rect 454906 333219 455224 333223
rect 454906 330533 455224 330537
rect 454906 330223 454910 330533
rect 454910 330223 455220 330533
rect 455220 330223 455224 330533
rect 454906 330219 455224 330223
rect 454906 327533 455224 327537
rect 454906 327223 454910 327533
rect 454910 327223 455220 327533
rect 455220 327223 455224 327533
rect 454906 327219 455224 327223
rect 454906 324533 455224 324537
rect 454906 324223 454910 324533
rect 454910 324223 455220 324533
rect 455220 324223 455224 324533
rect 454906 324219 455224 324223
rect 454906 321533 455224 321537
rect 454906 321223 454910 321533
rect 454910 321223 455220 321533
rect 455220 321223 455224 321533
rect 454906 321219 455224 321223
rect 454906 318533 455224 318537
rect 454906 318223 454910 318533
rect 454910 318223 455220 318533
rect 455220 318223 455224 318533
rect 454906 318219 455224 318223
rect 454906 315533 455224 315537
rect 454906 315223 454910 315533
rect 454910 315223 455220 315533
rect 455220 315223 455224 315533
rect 454906 315219 455224 315223
rect 454906 312533 455224 312537
rect 454906 312223 454910 312533
rect 454910 312223 455220 312533
rect 455220 312223 455224 312533
rect 454906 312219 455224 312223
rect 454906 309533 455224 309537
rect 454906 309223 454910 309533
rect 454910 309223 455220 309533
rect 455220 309223 455224 309533
rect 454906 309219 455224 309223
rect 454906 306533 455224 306537
rect 454906 306223 454910 306533
rect 454910 306223 455220 306533
rect 455220 306223 455224 306533
rect 454906 306219 455224 306223
rect 454906 303533 455224 303537
rect 454906 303223 454910 303533
rect 454910 303223 455220 303533
rect 455220 303223 455224 303533
rect 454906 303219 455224 303223
rect 454906 300533 455224 300537
rect 454906 300223 454910 300533
rect 454910 300223 455220 300533
rect 455220 300223 455224 300533
rect 454906 300219 455224 300223
rect 454906 297533 455224 297537
rect 454906 297223 454910 297533
rect 454910 297223 455220 297533
rect 455220 297223 455224 297533
rect 454906 297219 455224 297223
rect 454906 294533 455224 294537
rect 454906 294223 454910 294533
rect 454910 294223 455220 294533
rect 455220 294223 455224 294533
rect 454906 294219 455224 294223
rect 454906 291533 455224 291537
rect 454906 291223 454910 291533
rect 454910 291223 455220 291533
rect 455220 291223 455224 291533
rect 454906 291219 455224 291223
rect 454906 288533 455224 288537
rect 454906 288223 454910 288533
rect 454910 288223 455220 288533
rect 455220 288223 455224 288533
rect 454906 288219 455224 288223
rect 454906 285533 455224 285537
rect 454906 285223 454910 285533
rect 454910 285223 455220 285533
rect 455220 285223 455224 285533
rect 454906 285219 455224 285223
rect 454906 282533 455224 282537
rect 454906 282223 454910 282533
rect 454910 282223 455220 282533
rect 455220 282223 455224 282533
rect 454906 282219 455224 282223
rect 454906 279533 455224 279537
rect 454906 279223 454910 279533
rect 454910 279223 455220 279533
rect 455220 279223 455224 279533
rect 454906 279219 455224 279223
rect 454906 276533 455224 276537
rect 454906 276223 454910 276533
rect 454910 276223 455220 276533
rect 455220 276223 455224 276533
rect 454906 276219 455224 276223
rect 454906 273533 455224 273537
rect 454906 273223 454910 273533
rect 454910 273223 455220 273533
rect 455220 273223 455224 273533
rect 454906 273219 455224 273223
rect 454906 270533 455224 270537
rect 454906 270223 454910 270533
rect 454910 270223 455220 270533
rect 455220 270223 455224 270533
rect 454906 270219 455224 270223
rect 454906 267533 455224 267537
rect 454906 267223 454910 267533
rect 454910 267223 455220 267533
rect 455220 267223 455224 267533
rect 454906 267219 455224 267223
rect 454906 264533 455224 264537
rect 454906 264223 454910 264533
rect 454910 264223 455220 264533
rect 455220 264223 455224 264533
rect 454906 264219 455224 264223
rect 454906 261533 455224 261537
rect 454906 261223 454910 261533
rect 454910 261223 455220 261533
rect 455220 261223 455224 261533
rect 454906 261219 455224 261223
rect 454906 258533 455224 258537
rect 454906 258223 454910 258533
rect 454910 258223 455220 258533
rect 455220 258223 455224 258533
rect 454906 258219 455224 258223
rect 454906 255533 455224 255537
rect 454906 255223 454910 255533
rect 454910 255223 455220 255533
rect 455220 255223 455224 255533
rect 454906 255219 455224 255223
rect 454906 252533 455224 252537
rect 454906 252223 454910 252533
rect 454910 252223 455220 252533
rect 455220 252223 455224 252533
rect 454906 252219 455224 252223
rect 454906 249533 455224 249537
rect 454906 249223 454910 249533
rect 454910 249223 455220 249533
rect 455220 249223 455224 249533
rect 454906 249219 455224 249223
rect 454906 246533 455224 246537
rect 454906 246223 454910 246533
rect 454910 246223 455220 246533
rect 455220 246223 455224 246533
rect 454906 246219 455224 246223
rect 454906 243533 455224 243537
rect 454906 243223 454910 243533
rect 454910 243223 455220 243533
rect 455220 243223 455224 243533
rect 454906 243219 455224 243223
rect 454906 240533 455224 240537
rect 454906 240223 454910 240533
rect 454910 240223 455220 240533
rect 455220 240223 455224 240533
rect 454906 240219 455224 240223
rect 454906 237533 455224 237537
rect 454906 237223 454910 237533
rect 454910 237223 455220 237533
rect 455220 237223 455224 237533
rect 454906 237219 455224 237223
rect 454906 234533 455224 234537
rect 454906 234223 454910 234533
rect 454910 234223 455220 234533
rect 455220 234223 455224 234533
rect 454906 234219 455224 234223
rect 454906 231533 455224 231537
rect 454906 231223 454910 231533
rect 454910 231223 455220 231533
rect 455220 231223 455224 231533
rect 454906 231219 455224 231223
rect 454906 228533 455224 228537
rect 454906 228223 454910 228533
rect 454910 228223 455220 228533
rect 455220 228223 455224 228533
rect 454906 228219 455224 228223
rect 454906 225533 455224 225537
rect 454906 225223 454910 225533
rect 454910 225223 455220 225533
rect 455220 225223 455224 225533
rect 454906 225219 455224 225223
rect 454906 222533 455224 222537
rect 454906 222223 454910 222533
rect 454910 222223 455220 222533
rect 455220 222223 455224 222533
rect 454906 222219 455224 222223
rect 454906 219533 455224 219537
rect 454906 219223 454910 219533
rect 454910 219223 455220 219533
rect 455220 219223 455224 219533
rect 454906 219219 455224 219223
rect 454906 216533 455224 216537
rect 454906 216223 454910 216533
rect 454910 216223 455220 216533
rect 455220 216223 455224 216533
rect 454906 216219 455224 216223
rect 454906 213533 455224 213537
rect 454906 213223 454910 213533
rect 454910 213223 455220 213533
rect 455220 213223 455224 213533
rect 454906 213219 455224 213223
rect 454906 210533 455224 210537
rect 454906 210223 454910 210533
rect 454910 210223 455220 210533
rect 455220 210223 455224 210533
rect 454906 210219 455224 210223
rect 454906 207533 455224 207537
rect 454906 207223 454910 207533
rect 454910 207223 455220 207533
rect 455220 207223 455224 207533
rect 454906 207219 455224 207223
rect 454906 204533 455224 204537
rect 454906 204223 454910 204533
rect 454910 204223 455220 204533
rect 455220 204223 455224 204533
rect 454906 204219 455224 204223
rect 454906 201533 455224 201537
rect 454906 201223 454910 201533
rect 454910 201223 455220 201533
rect 455220 201223 455224 201533
rect 454906 201219 455224 201223
rect 454906 198533 455224 198537
rect 454906 198223 454910 198533
rect 454910 198223 455220 198533
rect 455220 198223 455224 198533
rect 454906 198219 455224 198223
rect 454906 195533 455224 195537
rect 454906 195223 454910 195533
rect 454910 195223 455220 195533
rect 455220 195223 455224 195533
rect 454906 195219 455224 195223
rect 454906 192533 455224 192537
rect 454906 192223 454910 192533
rect 454910 192223 455220 192533
rect 455220 192223 455224 192533
rect 454906 192219 455224 192223
rect 454906 189533 455224 189537
rect 454906 189223 454910 189533
rect 454910 189223 455220 189533
rect 455220 189223 455224 189533
rect 454906 189219 455224 189223
rect 454906 186533 455224 186537
rect 454906 186223 454910 186533
rect 454910 186223 455220 186533
rect 455220 186223 455224 186533
rect 454906 186219 455224 186223
rect 454906 183533 455224 183537
rect 454906 183223 454910 183533
rect 454910 183223 455220 183533
rect 455220 183223 455224 183533
rect 454906 183219 455224 183223
rect 454906 180533 455224 180537
rect 454906 180223 454910 180533
rect 454910 180223 455220 180533
rect 455220 180223 455224 180533
rect 454906 180219 455224 180223
rect 454906 177533 455224 177537
rect 454906 177223 454910 177533
rect 454910 177223 455220 177533
rect 455220 177223 455224 177533
rect 454906 177219 455224 177223
rect 454906 174533 455224 174537
rect 454906 174223 454910 174533
rect 454910 174223 455220 174533
rect 455220 174223 455224 174533
rect 454906 174219 455224 174223
rect 454906 171533 455224 171537
rect 454906 171223 454910 171533
rect 454910 171223 455220 171533
rect 455220 171223 455224 171533
rect 454906 171219 455224 171223
rect 454906 168533 455224 168537
rect 454906 168223 454910 168533
rect 454910 168223 455220 168533
rect 455220 168223 455224 168533
rect 454906 168219 455224 168223
rect 454906 165533 455224 165537
rect 454906 165223 454910 165533
rect 454910 165223 455220 165533
rect 455220 165223 455224 165533
rect 454906 165219 455224 165223
rect 454906 162533 455224 162537
rect 454906 162223 454910 162533
rect 454910 162223 455220 162533
rect 455220 162223 455224 162533
rect 454906 162219 455224 162223
rect 454906 159533 455224 159537
rect 454906 159223 454910 159533
rect 454910 159223 455220 159533
rect 455220 159223 455224 159533
rect 454906 159219 455224 159223
rect 454906 156533 455224 156537
rect 454906 156223 454910 156533
rect 454910 156223 455220 156533
rect 455220 156223 455224 156533
rect 454906 156219 455224 156223
rect 454906 153533 455224 153537
rect 454906 153223 454910 153533
rect 454910 153223 455220 153533
rect 455220 153223 455224 153533
rect 454906 153219 455224 153223
rect 454906 150533 455224 150537
rect 454906 150223 454910 150533
rect 454910 150223 455220 150533
rect 455220 150223 455224 150533
rect 454906 150219 455224 150223
rect 144647 129149 145733 129153
rect 144647 128071 144651 129149
rect 144651 128071 145729 129149
rect 145729 128071 145733 129149
rect 144647 128067 145733 128071
rect 515385 438538 515705 438543
rect 515385 438218 515700 438538
rect 515700 438218 515705 438538
rect 515385 438213 515705 438218
rect 515385 435538 515705 435543
rect 515385 435218 515700 435538
rect 515700 435218 515705 435538
rect 515385 435213 515705 435218
rect 515385 432538 515705 432543
rect 515385 432218 515700 432538
rect 515700 432218 515705 432538
rect 515385 432213 515705 432218
rect 515385 429538 515705 429543
rect 515385 429218 515700 429538
rect 515700 429218 515705 429538
rect 515385 429213 515705 429218
rect 515385 426538 515705 426543
rect 515385 426218 515700 426538
rect 515700 426218 515705 426538
rect 515385 426213 515705 426218
rect 515385 423538 515705 423543
rect 515385 423218 515700 423538
rect 515700 423218 515705 423538
rect 515385 423213 515705 423218
rect 515385 420538 515705 420543
rect 515385 420218 515700 420538
rect 515700 420218 515705 420538
rect 515385 420213 515705 420218
rect 515385 417538 515705 417543
rect 515385 417218 515700 417538
rect 515700 417218 515705 417538
rect 515385 417213 515705 417218
rect 515385 414538 515705 414543
rect 515385 414218 515700 414538
rect 515700 414218 515705 414538
rect 515385 414213 515705 414218
rect 515385 411538 515705 411543
rect 515385 411218 515700 411538
rect 515700 411218 515705 411538
rect 515385 411213 515705 411218
rect 515385 408538 515705 408543
rect 515385 408218 515700 408538
rect 515700 408218 515705 408538
rect 515385 408213 515705 408218
rect 515385 405538 515705 405543
rect 515385 405218 515700 405538
rect 515700 405218 515705 405538
rect 515385 405213 515705 405218
rect 515385 402538 515705 402543
rect 515385 402218 515700 402538
rect 515700 402218 515705 402538
rect 515385 402213 515705 402218
rect 515385 399538 515705 399543
rect 515385 399218 515700 399538
rect 515700 399218 515705 399538
rect 515385 399213 515705 399218
rect 515385 396538 515705 396543
rect 515385 396218 515700 396538
rect 515700 396218 515705 396538
rect 515385 396213 515705 396218
rect 515385 393538 515705 393543
rect 515385 393218 515700 393538
rect 515700 393218 515705 393538
rect 515385 393213 515705 393218
rect 515385 390538 515705 390543
rect 515385 390218 515700 390538
rect 515700 390218 515705 390538
rect 515385 390213 515705 390218
rect 515385 387538 515705 387543
rect 515385 387218 515700 387538
rect 515700 387218 515705 387538
rect 515385 387213 515705 387218
rect 515385 384538 515705 384543
rect 515385 384218 515700 384538
rect 515700 384218 515705 384538
rect 515385 384213 515705 384218
rect 515385 381538 515705 381543
rect 515385 381218 515700 381538
rect 515700 381218 515705 381538
rect 515385 381213 515705 381218
rect 515385 378538 515705 378543
rect 515385 378218 515700 378538
rect 515700 378218 515705 378538
rect 515385 378213 515705 378218
rect 515385 375538 515705 375543
rect 515385 375218 515700 375538
rect 515700 375218 515705 375538
rect 515385 375213 515705 375218
rect 515385 372538 515705 372543
rect 515385 372218 515700 372538
rect 515700 372218 515705 372538
rect 515385 372213 515705 372218
rect 515385 369538 515705 369543
rect 515385 369218 515700 369538
rect 515700 369218 515705 369538
rect 515385 369213 515705 369218
rect 582546 368786 582646 368886
rect 515385 366538 515705 366543
rect 515385 366218 515700 366538
rect 515700 366218 515705 366538
rect 515385 366213 515705 366218
rect 582546 364786 582646 364886
rect 515385 363538 515705 363543
rect 515385 363218 515700 363538
rect 515700 363218 515705 363538
rect 515385 363213 515705 363218
rect 515385 360538 515705 360543
rect 515385 360218 515700 360538
rect 515700 360218 515705 360538
rect 515385 360213 515705 360218
rect 515385 357538 515705 357543
rect 515385 357218 515700 357538
rect 515700 357218 515705 357538
rect 515385 357213 515705 357218
rect 515385 354538 515705 354543
rect 515385 354218 515700 354538
rect 515700 354218 515705 354538
rect 515385 354213 515705 354218
rect 515385 351538 515705 351543
rect 515385 351218 515700 351538
rect 515700 351218 515705 351538
rect 515385 351213 515705 351218
rect 515385 348538 515705 348543
rect 515385 348218 515700 348538
rect 515700 348218 515705 348538
rect 515385 348213 515705 348218
rect 515385 345538 515705 345543
rect 515385 345218 515700 345538
rect 515700 345218 515705 345538
rect 515385 345213 515705 345218
rect 515385 342538 515705 342543
rect 515385 342218 515700 342538
rect 515700 342218 515705 342538
rect 515385 342213 515705 342218
rect 515385 339538 515705 339543
rect 515385 339218 515700 339538
rect 515700 339218 515705 339538
rect 515385 339213 515705 339218
rect 515385 336538 515705 336543
rect 515385 336218 515700 336538
rect 515700 336218 515705 336538
rect 515385 336213 515705 336218
rect 515385 333538 515705 333543
rect 515385 333218 515700 333538
rect 515700 333218 515705 333538
rect 515385 333213 515705 333218
rect 515385 330538 515705 330543
rect 515385 330218 515700 330538
rect 515700 330218 515705 330538
rect 515385 330213 515705 330218
rect 515385 327538 515705 327543
rect 515385 327218 515700 327538
rect 515700 327218 515705 327538
rect 515385 327213 515705 327218
rect 515385 324538 515705 324543
rect 515385 324218 515700 324538
rect 515700 324218 515705 324538
rect 515385 324213 515705 324218
rect 515385 321538 515705 321543
rect 515385 321218 515700 321538
rect 515700 321218 515705 321538
rect 515385 321213 515705 321218
rect 515385 318538 515705 318543
rect 515385 318218 515700 318538
rect 515700 318218 515705 318538
rect 515385 318213 515705 318218
rect 515385 315538 515705 315543
rect 515385 315218 515700 315538
rect 515700 315218 515705 315538
rect 515385 315213 515705 315218
rect 515385 312538 515705 312543
rect 515385 312218 515700 312538
rect 515700 312218 515705 312538
rect 515385 312213 515705 312218
rect 515385 309538 515705 309543
rect 515385 309218 515700 309538
rect 515700 309218 515705 309538
rect 515385 309213 515705 309218
rect 515385 306538 515705 306543
rect 515385 306218 515700 306538
rect 515700 306218 515705 306538
rect 515385 306213 515705 306218
rect 515385 303538 515705 303543
rect 515385 303218 515700 303538
rect 515700 303218 515705 303538
rect 515385 303213 515705 303218
rect 515385 300538 515705 300543
rect 515385 300218 515700 300538
rect 515700 300218 515705 300538
rect 515385 300213 515705 300218
rect 515385 297538 515705 297543
rect 515385 297218 515700 297538
rect 515700 297218 515705 297538
rect 515385 297213 515705 297218
rect 515385 294538 515705 294543
rect 515385 294218 515700 294538
rect 515700 294218 515705 294538
rect 515385 294213 515705 294218
rect 515385 291538 515705 291543
rect 515385 291218 515700 291538
rect 515700 291218 515705 291538
rect 515385 291213 515705 291218
rect 515385 288538 515705 288543
rect 515385 288218 515700 288538
rect 515700 288218 515705 288538
rect 515385 288213 515705 288218
rect 515385 285538 515705 285543
rect 515385 285218 515700 285538
rect 515700 285218 515705 285538
rect 515385 285213 515705 285218
rect 515385 282538 515705 282543
rect 515385 282218 515700 282538
rect 515700 282218 515705 282538
rect 515385 282213 515705 282218
rect 515385 279538 515705 279543
rect 515385 279218 515700 279538
rect 515700 279218 515705 279538
rect 515385 279213 515705 279218
rect 515385 276538 515705 276543
rect 515385 276218 515700 276538
rect 515700 276218 515705 276538
rect 515385 276213 515705 276218
rect 515385 273538 515705 273543
rect 515385 273218 515700 273538
rect 515700 273218 515705 273538
rect 515385 273213 515705 273218
rect 515385 270538 515705 270543
rect 515385 270218 515700 270538
rect 515700 270218 515705 270538
rect 515385 270213 515705 270218
rect 515385 267538 515705 267543
rect 515385 267218 515700 267538
rect 515700 267218 515705 267538
rect 515385 267213 515705 267218
rect 515385 264538 515705 264543
rect 515385 264218 515700 264538
rect 515700 264218 515705 264538
rect 515385 264213 515705 264218
rect 515385 261538 515705 261543
rect 515385 261218 515700 261538
rect 515700 261218 515705 261538
rect 515385 261213 515705 261218
rect 515385 258538 515705 258543
rect 515385 258218 515700 258538
rect 515700 258218 515705 258538
rect 515385 258213 515705 258218
rect 515385 255538 515705 255543
rect 515385 255218 515700 255538
rect 515700 255218 515705 255538
rect 515385 255213 515705 255218
rect 515385 252538 515705 252543
rect 515385 252218 515700 252538
rect 515700 252218 515705 252538
rect 515385 252213 515705 252218
rect 515385 249538 515705 249543
rect 515385 249218 515700 249538
rect 515700 249218 515705 249538
rect 515385 249213 515705 249218
rect 515385 246538 515705 246543
rect 515385 246218 515700 246538
rect 515700 246218 515705 246538
rect 515385 246213 515705 246218
rect 515385 243538 515705 243543
rect 515385 243218 515700 243538
rect 515700 243218 515705 243538
rect 515385 243213 515705 243218
rect 515385 240538 515705 240543
rect 515385 240218 515700 240538
rect 515700 240218 515705 240538
rect 515385 240213 515705 240218
rect 515385 237538 515705 237543
rect 515385 237218 515700 237538
rect 515700 237218 515705 237538
rect 515385 237213 515705 237218
rect 515385 234538 515705 234543
rect 515385 234218 515700 234538
rect 515700 234218 515705 234538
rect 515385 234213 515705 234218
rect 515385 231538 515705 231543
rect 515385 231218 515700 231538
rect 515700 231218 515705 231538
rect 515385 231213 515705 231218
rect 515385 228538 515705 228543
rect 515385 228218 515700 228538
rect 515700 228218 515705 228538
rect 515385 228213 515705 228218
rect 515385 225538 515705 225543
rect 515385 225218 515700 225538
rect 515700 225218 515705 225538
rect 515385 225213 515705 225218
rect 515385 222538 515705 222543
rect 515385 222218 515700 222538
rect 515700 222218 515705 222538
rect 515385 222213 515705 222218
rect 515385 219538 515705 219543
rect 515385 219218 515700 219538
rect 515700 219218 515705 219538
rect 515385 219213 515705 219218
rect 515385 216538 515705 216543
rect 515385 216218 515700 216538
rect 515700 216218 515705 216538
rect 515385 216213 515705 216218
rect 515385 213538 515705 213543
rect 515385 213218 515700 213538
rect 515700 213218 515705 213538
rect 515385 213213 515705 213218
rect 515385 210538 515705 210543
rect 515385 210218 515700 210538
rect 515700 210218 515705 210538
rect 515385 210213 515705 210218
rect 515385 207538 515705 207543
rect 515385 207218 515700 207538
rect 515700 207218 515705 207538
rect 515385 207213 515705 207218
rect 515385 204538 515705 204543
rect 515385 204218 515700 204538
rect 515700 204218 515705 204538
rect 515385 204213 515705 204218
rect 515385 201538 515705 201543
rect 515385 201218 515700 201538
rect 515700 201218 515705 201538
rect 515385 201213 515705 201218
rect 515385 198538 515705 198543
rect 515385 198218 515700 198538
rect 515700 198218 515705 198538
rect 515385 198213 515705 198218
rect 515385 195538 515705 195543
rect 515385 195218 515700 195538
rect 515700 195218 515705 195538
rect 515385 195213 515705 195218
rect 515385 192538 515705 192543
rect 515385 192218 515700 192538
rect 515700 192218 515705 192538
rect 515385 192213 515705 192218
rect 515385 189538 515705 189543
rect 515385 189218 515700 189538
rect 515700 189218 515705 189538
rect 515385 189213 515705 189218
rect 515385 186538 515705 186543
rect 515385 186218 515700 186538
rect 515700 186218 515705 186538
rect 515385 186213 515705 186218
rect 515385 183538 515705 183543
rect 515385 183218 515700 183538
rect 515700 183218 515705 183538
rect 515385 183213 515705 183218
rect 515385 180538 515705 180543
rect 515385 180218 515700 180538
rect 515700 180218 515705 180538
rect 515385 180213 515705 180218
rect 515385 177538 515705 177543
rect 515385 177218 515700 177538
rect 515700 177218 515705 177538
rect 515385 177213 515705 177218
rect 515385 174538 515705 174543
rect 515385 174218 515700 174538
rect 515700 174218 515705 174538
rect 515385 174213 515705 174218
rect 515385 171538 515705 171543
rect 515385 171218 515700 171538
rect 515700 171218 515705 171538
rect 515385 171213 515705 171218
rect 515385 168538 515705 168543
rect 515385 168218 515700 168538
rect 515700 168218 515705 168538
rect 515385 168213 515705 168218
rect 515385 165538 515705 165543
rect 515385 165218 515700 165538
rect 515700 165218 515705 165538
rect 515385 165213 515705 165218
rect 515385 162538 515705 162543
rect 515385 162218 515700 162538
rect 515700 162218 515705 162538
rect 515385 162213 515705 162218
rect 515385 159538 515705 159543
rect 515385 159218 515700 159538
rect 515700 159218 515705 159538
rect 515385 159213 515705 159218
rect 515385 156538 515705 156543
rect 515385 156218 515700 156538
rect 515700 156218 515705 156538
rect 515385 156213 515705 156218
rect 515385 153538 515705 153543
rect 515385 153218 515700 153538
rect 515700 153218 515705 153538
rect 515385 153213 515705 153218
rect 515385 150538 515705 150543
rect 515385 150218 515700 150538
rect 515700 150218 515705 150538
rect 515385 150213 515705 150218
rect 499375 139852 500789 141266
rect 503116 139853 504528 141265
rect 505628 140121 506504 140997
rect 463531 126465 464216 127150
rect 582546 323546 582646 323646
rect 582546 319546 582646 319646
rect 582546 279146 582646 279246
rect 582546 275146 582646 275246
rect 554140 191768 578296 196966
rect 553050 181150 576862 186340
rect 553277 159411 558075 164209
rect 582546 99146 582646 99246
rect 582546 95146 582646 95246
rect 1034 10876 1134 10976
rect 354 3908 466 4020
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329590 701834 334030 701858
rect 229190 699708 231180 699960
rect 229190 698530 229597 699708
rect 228350 698529 229597 698530
rect 228350 697491 228439 698529
rect 229477 697552 229597 698529
rect 229477 697491 231180 697552
rect 228350 697490 231180 697491
rect 229190 697460 231180 697490
rect 329590 697442 329614 701834
rect 334006 697442 334030 701834
rect 329590 697349 331192 697442
rect 332128 697349 334030 697442
rect 329590 694172 334030 697349
rect 574553 682650 577887 682687
rect 574553 682402 582200 682650
rect 574553 678818 575238 682402
rect 582000 678818 582200 682402
rect 574553 678570 582200 678818
rect 566593 674025 571477 674026
rect 1033 462476 1135 462477
rect 2440 462476 2540 462606
rect 1033 462376 1034 462476
rect 1134 462376 2540 462476
rect 1033 462375 1135 462376
rect 1033 419276 1135 419277
rect 2440 419276 2540 462376
rect 8387 422228 8457 672796
rect 9016 422228 9126 672796
rect 10674 422228 10784 672796
rect 478811 669776 566594 674025
rect 478811 668948 547286 669776
rect 548114 669143 566594 669776
rect 571476 669143 571477 674025
rect 548114 668948 548311 669143
rect 566593 669142 571477 669143
rect 478811 668947 548311 668948
rect 478811 597477 483889 668947
rect 574553 665164 577887 678570
rect 303894 592806 304214 596286
rect 339885 593924 483889 597477
rect 335215 593094 483889 593924
rect 303894 592534 303918 592806
rect 304190 592534 304214 592806
rect 303894 592510 304214 592534
rect 289695 592401 292013 592402
rect 289695 592293 289696 592401
rect 289804 592293 292013 592401
rect 339885 592399 483889 593094
rect 490227 661830 577887 665164
rect 289695 592292 292013 592293
rect 338102 592197 338394 592198
rect 338102 591907 338103 592197
rect 338393 591907 338394 592197
rect 338102 591906 338394 591907
rect 287844 591878 292634 591902
rect 287844 591606 292338 591878
rect 292610 591606 292634 591878
rect 287844 591582 292634 591606
rect 287844 590509 288164 591582
rect 287844 590191 287845 590509
rect 288163 590191 288164 590509
rect 338103 590460 338393 591906
rect 287844 590190 288164 590191
rect 338103 586460 338393 590140
rect 293834 579119 293944 582037
rect 289791 579118 294040 579119
rect 289791 578818 289792 579118
rect 290092 578818 294040 579118
rect 289791 578817 294040 578818
rect 294534 571852 294754 581972
rect 291816 571851 294754 571852
rect 291816 571633 291817 571851
rect 292035 571633 294754 571851
rect 291816 571632 294754 571633
rect 291888 570930 292326 571124
rect 297534 570930 297754 582004
rect 291888 570929 297754 570930
rect 291888 570711 291973 570929
rect 292191 570711 297754 570929
rect 291888 570710 297754 570711
rect 291888 570506 292326 570710
rect 300534 568142 300754 582016
rect 308981 578275 309668 578276
rect 308981 577590 308982 578275
rect 309667 577590 309668 578275
rect 308981 577589 309668 577590
rect 292240 568141 300754 568142
rect 292240 567923 292241 568141
rect 292459 567923 300754 568141
rect 292240 567922 300754 567923
rect 308982 557285 309667 577589
rect 314130 473945 339500 473946
rect 289093 473351 289095 473352
rect 289094 472811 289095 473351
rect 289093 472810 289095 472811
rect 297405 471950 297407 471951
rect 297405 471570 297406 471950
rect 297405 471569 297407 471570
rect 290882 469717 290884 469718
rect 290882 469067 290883 469717
rect 314130 469147 314131 473945
rect 318929 473922 339500 473945
rect 318929 469170 334724 473922
rect 339476 469170 339500 473922
rect 318929 469147 339500 469170
rect 314130 469146 339500 469147
rect 290882 469066 290884 469067
rect 141828 441759 142089 441760
rect 141828 441500 141829 441759
rect 142088 441500 142089 441759
rect 141828 439981 142089 441500
rect 162784 438802 163104 454558
rect 162784 438530 162808 438802
rect 163080 438530 163104 438802
rect 162784 438506 163104 438530
rect 165784 438802 166104 454558
rect 165784 438530 165808 438802
rect 166080 438530 166104 438802
rect 165784 438506 166104 438530
rect 168784 438802 169104 454558
rect 168784 438530 168808 438802
rect 169080 438530 169104 438802
rect 168784 438506 169104 438530
rect 171784 438802 172104 454558
rect 171784 438530 171808 438802
rect 172080 438530 172104 438802
rect 171784 438506 172104 438530
rect 174784 438802 175104 454558
rect 174784 438530 174808 438802
rect 175080 438530 175104 438802
rect 174784 438506 175104 438530
rect 177784 438802 178104 454558
rect 177784 438530 177808 438802
rect 178080 438530 178104 438802
rect 177784 438506 178104 438530
rect 180784 438802 181104 454558
rect 180784 438530 180808 438802
rect 181080 438530 181104 438802
rect 180784 438506 181104 438530
rect 183784 438802 184104 454558
rect 183784 438530 183808 438802
rect 184080 438530 184104 438802
rect 183784 438506 184104 438530
rect 186784 438802 187104 454558
rect 186784 438530 186808 438802
rect 187080 438530 187104 438802
rect 186784 438506 187104 438530
rect 189784 438802 190104 454558
rect 189784 438530 189808 438802
rect 190080 438530 190104 438802
rect 189784 438506 190104 438530
rect 192784 438802 193104 454558
rect 192784 438530 192808 438802
rect 193080 438530 193104 438802
rect 192784 438506 193104 438530
rect 195784 438802 196104 454558
rect 195784 438530 195808 438802
rect 196080 438530 196104 438802
rect 195784 438506 196104 438530
rect 198784 438802 199104 454558
rect 198784 438530 198808 438802
rect 199080 438530 199104 438802
rect 198784 438506 199104 438530
rect 201784 438802 202104 454558
rect 201784 438530 201808 438802
rect 202080 438530 202104 438802
rect 201784 438506 202104 438530
rect 204784 438802 205104 454558
rect 204784 438530 204808 438802
rect 205080 438530 205104 438802
rect 204784 438506 205104 438530
rect 207784 438802 208104 454558
rect 207784 438530 207808 438802
rect 208080 438530 208104 438802
rect 207784 438506 208104 438530
rect 210784 438802 211104 454558
rect 210784 438530 210808 438802
rect 211080 438530 211104 438802
rect 210784 438506 211104 438530
rect 213784 438802 214104 454558
rect 213784 438530 213808 438802
rect 214080 438530 214104 438802
rect 213784 438506 214104 438530
rect 216784 438802 217104 454558
rect 216784 438530 216808 438802
rect 217080 438530 217104 438802
rect 216784 438506 217104 438530
rect 219784 438802 220104 454558
rect 219784 438530 219808 438802
rect 220080 438530 220104 438802
rect 219784 438506 220104 438530
rect 222784 438802 223104 454558
rect 222784 438530 222808 438802
rect 223080 438530 223104 438802
rect 222784 438506 223104 438530
rect 225784 438802 226104 454558
rect 225784 438530 225808 438802
rect 226080 438530 226104 438802
rect 225784 438506 226104 438530
rect 228784 438802 229104 454558
rect 228784 438530 228808 438802
rect 229080 438530 229104 438802
rect 228784 438506 229104 438530
rect 231784 438802 232104 454558
rect 231784 438530 231808 438802
rect 232080 438530 232104 438802
rect 231784 438506 232104 438530
rect 234784 438802 235104 454558
rect 234784 438530 234808 438802
rect 235080 438530 235104 438802
rect 234784 438506 235104 438530
rect 237784 438802 238104 454558
rect 237784 438530 237808 438802
rect 238080 438530 238104 438802
rect 237784 438506 238104 438530
rect 240784 438802 241104 454558
rect 240784 438530 240808 438802
rect 241080 438530 241104 438802
rect 240784 438506 241104 438530
rect 243784 438802 244104 454558
rect 243784 438530 243808 438802
rect 244080 438530 244104 438802
rect 243784 438506 244104 438530
rect 246784 438802 247104 454558
rect 246784 438530 246808 438802
rect 247080 438530 247104 438802
rect 246784 438506 247104 438530
rect 249784 438802 250104 454558
rect 249784 438530 249808 438802
rect 250080 438530 250104 438802
rect 249784 438506 250104 438530
rect 252784 438802 253104 454558
rect 252784 438530 252808 438802
rect 253080 438530 253104 438802
rect 252784 438506 253104 438530
rect 255784 438802 256104 454558
rect 255784 438530 255808 438802
rect 256080 438530 256104 438802
rect 255784 438506 256104 438530
rect 258784 438802 259104 454558
rect 258784 438530 258808 438802
rect 259080 438530 259104 438802
rect 258784 438506 259104 438530
rect 261784 438802 262104 454558
rect 261784 438530 261808 438802
rect 262080 438530 262104 438802
rect 261784 438506 262104 438530
rect 264784 438802 265104 454558
rect 264784 438530 264808 438802
rect 265080 438530 265104 438802
rect 264784 438506 265104 438530
rect 267784 438802 268104 454558
rect 267784 438530 267808 438802
rect 268080 438530 268104 438802
rect 267784 438506 268104 438530
rect 270784 438802 271104 454558
rect 270784 438530 270808 438802
rect 271080 438530 271104 438802
rect 270784 438506 271104 438530
rect 273784 438802 274104 454558
rect 273784 438530 273808 438802
rect 274080 438530 274104 438802
rect 273784 438506 274104 438530
rect 276784 438802 277104 454558
rect 276784 438530 276808 438802
rect 277080 438530 277104 438802
rect 276784 438506 277104 438530
rect 279784 438802 280104 454558
rect 279784 438530 279808 438802
rect 280080 438530 280104 438802
rect 279784 438506 280104 438530
rect 282784 438802 283104 454558
rect 282784 438530 282808 438802
rect 283080 438530 283104 438802
rect 282784 438506 283104 438530
rect 285784 438802 286104 454558
rect 285784 438530 285808 438802
rect 286080 438530 286104 438802
rect 285784 438506 286104 438530
rect 288784 438802 289104 454558
rect 288784 438530 288808 438802
rect 289080 438530 289104 438802
rect 288784 438506 289104 438530
rect 291784 438802 292104 454558
rect 291784 438530 291808 438802
rect 292080 438530 292104 438802
rect 291784 438506 292104 438530
rect 294784 438802 295104 454558
rect 294784 438530 294808 438802
rect 295080 438530 295104 438802
rect 294784 438506 295104 438530
rect 297784 438802 298104 454558
rect 297784 438530 297808 438802
rect 298080 438530 298104 438802
rect 297784 438506 298104 438530
rect 300784 438802 301104 454558
rect 300784 438530 300808 438802
rect 301080 438530 301104 438802
rect 300784 438506 301104 438530
rect 303784 438802 304104 454558
rect 303784 438530 303808 438802
rect 304080 438530 304104 438802
rect 303784 438506 304104 438530
rect 306784 438802 307104 454558
rect 306784 438530 306808 438802
rect 307080 438530 307104 438802
rect 306784 438506 307104 438530
rect 309784 438802 310104 454558
rect 309784 438530 309808 438802
rect 310080 438530 310104 438802
rect 309784 438506 310104 438530
rect 312784 438802 313104 454558
rect 312784 438530 312808 438802
rect 313080 438530 313104 438802
rect 312784 438506 313104 438530
rect 315784 438802 316104 454558
rect 315784 438530 315808 438802
rect 316080 438530 316104 438802
rect 315784 438506 316104 438530
rect 318784 438802 319104 454558
rect 318784 438530 318808 438802
rect 319080 438530 319104 438802
rect 318784 438506 319104 438530
rect 321784 438802 322104 454558
rect 321784 438530 321808 438802
rect 322080 438530 322104 438802
rect 321784 438506 322104 438530
rect 324784 438802 325104 454558
rect 324784 438530 324808 438802
rect 325080 438530 325104 438802
rect 324784 438506 325104 438530
rect 327784 438802 328104 454558
rect 327784 438530 327808 438802
rect 328080 438530 328104 438802
rect 327784 438506 328104 438530
rect 330784 438802 331104 454558
rect 330784 438530 330808 438802
rect 331080 438530 331104 438802
rect 330784 438506 331104 438530
rect 333784 438802 334104 454558
rect 333784 438530 333808 438802
rect 334080 438530 334104 438802
rect 333784 438506 334104 438530
rect 336784 438802 337104 454558
rect 336784 438530 336808 438802
rect 337080 438530 337104 438802
rect 336784 438506 337104 438530
rect 339784 438802 340104 454558
rect 339784 438530 339808 438802
rect 340080 438530 340104 438802
rect 339784 438506 340104 438530
rect 342784 438802 343104 454558
rect 342784 438530 342808 438802
rect 343080 438530 343104 438802
rect 342784 438506 343104 438530
rect 345784 438802 346104 454558
rect 345784 438530 345808 438802
rect 346080 438530 346104 438802
rect 345784 438506 346104 438530
rect 348784 438802 349104 454558
rect 348784 438530 348808 438802
rect 349080 438530 349104 438802
rect 348784 438506 349104 438530
rect 351784 438802 352104 454558
rect 351784 438530 351808 438802
rect 352080 438530 352104 438802
rect 351784 438506 352104 438530
rect 354784 438802 355104 454558
rect 354784 438530 354808 438802
rect 355080 438530 355104 438802
rect 354784 438506 355104 438530
rect 357784 438802 358104 454558
rect 357784 438530 357808 438802
rect 358080 438530 358104 438802
rect 357784 438506 358104 438530
rect 360784 438802 361104 454558
rect 360784 438530 360808 438802
rect 361080 438530 361104 438802
rect 360784 438506 361104 438530
rect 363784 438802 364104 454558
rect 363784 438530 363808 438802
rect 364080 438530 364104 438802
rect 363784 438506 364104 438530
rect 366784 438802 367104 454558
rect 366784 438530 366808 438802
rect 367080 438530 367104 438802
rect 366784 438506 367104 438530
rect 369784 438802 370104 454558
rect 369784 438530 369808 438802
rect 370080 438530 370104 438802
rect 369784 438506 370104 438530
rect 372784 438802 373104 454558
rect 372784 438530 372808 438802
rect 373080 438530 373104 438802
rect 372784 438506 373104 438530
rect 375784 438802 376104 454558
rect 375784 438530 375808 438802
rect 376080 438530 376104 438802
rect 375784 438506 376104 438530
rect 378784 438802 379104 454558
rect 378784 438530 378808 438802
rect 379080 438530 379104 438802
rect 378784 438506 379104 438530
rect 381784 438802 382104 454558
rect 381784 438530 381808 438802
rect 382080 438530 382104 438802
rect 381784 438506 382104 438530
rect 384784 438802 385104 454558
rect 384784 438530 384808 438802
rect 385080 438530 385104 438802
rect 384784 438506 385104 438530
rect 387784 438802 388104 454558
rect 387784 438530 387808 438802
rect 388080 438530 388104 438802
rect 387784 438506 388104 438530
rect 390784 438802 391104 454558
rect 390784 438530 390808 438802
rect 391080 438530 391104 438802
rect 390784 438506 391104 438530
rect 393784 438802 394104 454558
rect 393784 438530 393808 438802
rect 394080 438530 394104 438802
rect 393784 438506 394104 438530
rect 396784 438802 397104 454558
rect 396784 438530 396808 438802
rect 397080 438530 397104 438802
rect 396784 438506 397104 438530
rect 399784 438802 400104 454558
rect 399784 438530 399808 438802
rect 400080 438530 400104 438802
rect 399784 438506 400104 438530
rect 402784 438802 403104 454558
rect 402784 438530 402808 438802
rect 403080 438530 403104 438802
rect 402784 438506 403104 438530
rect 405784 438802 406104 454558
rect 405784 438530 405808 438802
rect 406080 438530 406104 438802
rect 405784 438506 406104 438530
rect 408784 438802 409104 454558
rect 408784 438530 408808 438802
rect 409080 438530 409104 438802
rect 408784 438506 409104 438530
rect 411784 438802 412104 454558
rect 411784 438530 411808 438802
rect 412080 438530 412104 438802
rect 411784 438506 412104 438530
rect 414784 438802 415104 454558
rect 414784 438530 414808 438802
rect 415080 438530 415104 438802
rect 414784 438506 415104 438530
rect 417784 438802 418104 454558
rect 417784 438530 417808 438802
rect 418080 438530 418104 438802
rect 417784 438506 418104 438530
rect 420784 438802 421104 454558
rect 420784 438530 420808 438802
rect 421080 438530 421104 438802
rect 420784 438506 421104 438530
rect 423784 438802 424104 454558
rect 423784 438530 423808 438802
rect 424080 438530 424104 438802
rect 423784 438506 424104 438530
rect 426784 438802 427104 454558
rect 426784 438530 426808 438802
rect 427080 438530 427104 438802
rect 426784 438506 427104 438530
rect 429784 438802 430104 454558
rect 429784 438530 429808 438802
rect 430080 438530 430104 438802
rect 429784 438506 430104 438530
rect 432784 438802 433104 454558
rect 432784 438530 432808 438802
rect 433080 438530 433104 438802
rect 432784 438506 433104 438530
rect 435784 438802 436104 454558
rect 435784 438530 435808 438802
rect 436080 438530 436104 438802
rect 435784 438506 436104 438530
rect 438784 438802 439104 454558
rect 438784 438530 438808 438802
rect 439080 438530 439104 438802
rect 438784 438506 439104 438530
rect 441784 438802 442104 454558
rect 441784 438530 441808 438802
rect 442080 438530 442104 438802
rect 441784 438506 442104 438530
rect 444784 438802 445104 454558
rect 444784 438530 444808 438802
rect 445080 438530 445104 438802
rect 444784 438506 445104 438530
rect 447784 438802 448104 454558
rect 447784 438530 447808 438802
rect 448080 438530 448104 438802
rect 447784 438506 448104 438530
rect 454905 438537 455225 438538
rect 454905 438219 454906 438537
rect 455224 438219 455225 438537
rect 454905 438218 455225 438219
rect 149102 437233 149422 437234
rect 149102 436915 149103 437233
rect 149421 436915 149422 437233
rect 149102 436914 149422 436915
rect 149102 436489 149422 436490
rect 149102 436171 149103 436489
rect 149421 436171 149422 436489
rect 149102 436170 149422 436171
rect 120572 436088 129377 436112
rect 120572 435816 129081 436088
rect 129353 435816 129377 436088
rect 120572 435792 129377 435816
rect 454905 435537 455225 435538
rect 454905 435219 454906 435537
rect 455224 435219 455225 435537
rect 454905 435218 455225 435219
rect 454905 432537 455225 432538
rect 454905 432219 454906 432537
rect 455224 432219 455225 432537
rect 454905 432218 455225 432219
rect 120572 432088 129377 432112
rect 120572 431816 129081 432088
rect 129353 431816 129377 432088
rect 120572 431792 129377 431816
rect 454905 429537 455225 429538
rect 454905 429219 454906 429537
rect 455224 429219 455225 429537
rect 454905 429218 455225 429219
rect 120572 428088 129377 428112
rect 120572 427816 129081 428088
rect 129353 427816 129377 428088
rect 120572 427792 129377 427816
rect 454905 426537 455225 426538
rect 454905 426219 454906 426537
rect 455224 426219 455225 426537
rect 454905 426218 455225 426219
rect 120572 424088 129377 424112
rect 120572 423816 129081 424088
rect 129353 423816 129377 424088
rect 120572 423792 129377 423816
rect 454905 423537 455225 423538
rect 454905 423219 454906 423537
rect 455224 423219 455225 423537
rect 454905 423218 455225 423219
rect 454905 420537 455225 420538
rect 454905 420219 454906 420537
rect 455224 420219 455225 420537
rect 454905 420218 455225 420219
rect 1033 419176 1034 419276
rect 1134 419176 2540 419276
rect 1033 419175 1135 419176
rect 1033 376076 1135 376077
rect 2440 376076 2540 419176
rect 8387 379054 8457 419818
rect 9016 379054 9126 419818
rect 10674 379054 10784 419818
rect 120572 420088 129377 420112
rect 120572 419816 129081 420088
rect 129353 419816 129377 420088
rect 120572 419792 129377 419816
rect 454905 417537 455225 417538
rect 454905 417219 454906 417537
rect 455224 417219 455225 417537
rect 454905 417218 455225 417219
rect 120572 416088 129377 416112
rect 120572 415816 129081 416088
rect 129353 415816 129377 416088
rect 120572 415792 129377 415816
rect 454905 414537 455225 414538
rect 454905 414219 454906 414537
rect 455224 414219 455225 414537
rect 454905 414218 455225 414219
rect 120572 412088 129377 412112
rect 120572 411816 129081 412088
rect 129353 411816 129377 412088
rect 120572 411792 129377 411816
rect 454905 411537 455225 411538
rect 454905 411219 454906 411537
rect 455224 411219 455225 411537
rect 454905 411218 455225 411219
rect 454905 408537 455225 408538
rect 454905 408219 454906 408537
rect 455224 408219 455225 408537
rect 454905 408218 455225 408219
rect 120572 408088 129377 408112
rect 120572 407816 129081 408088
rect 129353 407816 129377 408088
rect 120572 407792 129377 407816
rect 454905 405537 455225 405538
rect 454905 405219 454906 405537
rect 455224 405219 455225 405537
rect 454905 405218 455225 405219
rect 120572 404088 129377 404112
rect 120572 403816 129081 404088
rect 129353 403816 129377 404088
rect 120572 403792 129377 403816
rect 454905 402537 455225 402538
rect 454905 402219 454906 402537
rect 455224 402219 455225 402537
rect 454905 402218 455225 402219
rect 120572 400088 129377 400112
rect 120572 399816 129081 400088
rect 129353 399816 129377 400088
rect 120572 399792 129377 399816
rect 454905 399537 455225 399538
rect 454905 399219 454906 399537
rect 455224 399219 455225 399537
rect 454905 399218 455225 399219
rect 454905 396537 455225 396538
rect 454905 396219 454906 396537
rect 455224 396219 455225 396537
rect 454905 396218 455225 396219
rect 120572 396088 129377 396112
rect 120572 395816 129081 396088
rect 129353 395816 129377 396088
rect 120572 395792 129377 395816
rect 454905 393537 455225 393538
rect 454905 393219 454906 393537
rect 455224 393219 455225 393537
rect 454905 393218 455225 393219
rect 120572 392088 129377 392112
rect 120572 391816 129081 392088
rect 129353 391816 129377 392088
rect 120572 391792 129377 391816
rect 454905 390537 455225 390538
rect 454905 390219 454906 390537
rect 455224 390219 455225 390537
rect 454905 390218 455225 390219
rect 120572 388088 129377 388112
rect 120572 387816 129081 388088
rect 129353 387816 129377 388088
rect 120572 387792 129377 387816
rect 454905 387537 455225 387538
rect 454905 387219 454906 387537
rect 455224 387219 455225 387537
rect 454905 387218 455225 387219
rect 454905 384537 455225 384538
rect 454905 384219 454906 384537
rect 455224 384219 455225 384537
rect 454905 384218 455225 384219
rect 120572 384088 129377 384112
rect 120572 383816 129081 384088
rect 129353 383816 129377 384088
rect 120572 383792 129377 383816
rect 454905 381537 455225 381538
rect 454905 381219 454906 381537
rect 455224 381219 455225 381537
rect 454905 381218 455225 381219
rect 120572 380088 129377 380112
rect 120572 379816 129081 380088
rect 129353 379816 129377 380088
rect 120572 379792 129377 379816
rect 454905 378537 455225 378538
rect 454905 378219 454906 378537
rect 455224 378219 455225 378537
rect 454905 378218 455225 378219
rect 1033 375976 1034 376076
rect 1134 375976 2540 376076
rect 1033 375975 1135 375976
rect 1033 332776 1135 332777
rect 2440 332776 2540 375976
rect 1033 332676 1034 332776
rect 1134 332676 2540 332776
rect 1033 332675 1135 332676
rect 1033 289576 1135 289577
rect 2440 289576 2540 332676
rect 5659 293381 5773 293382
rect 5659 293269 5660 293381
rect 5772 293269 5773 293381
rect 5659 293268 5773 293269
rect 1033 289476 1034 289576
rect 1134 289476 2540 289576
rect 1033 289475 1135 289476
rect 1033 246576 1135 246577
rect 2440 246576 2540 289476
rect 5660 253172 5772 293268
rect 8387 261321 8457 376032
rect 8381 261320 8463 261321
rect 8381 261250 8382 261320
rect 8462 261250 8463 261320
rect 8381 261249 8463 261250
rect 5660 253062 5661 253172
rect 5771 253062 5772 253172
rect 5660 253061 5772 253062
rect 1033 246476 1034 246576
rect 1134 246476 2540 246576
rect 1033 246475 1135 246476
rect 2440 178862 2540 246476
rect 9016 191343 9126 376032
rect 10674 191538 10784 376032
rect 120572 376088 129377 376112
rect 120572 375816 129081 376088
rect 129353 375816 129377 376088
rect 120572 375792 129377 375816
rect 454905 375537 455225 375538
rect 454905 375219 454906 375537
rect 455224 375219 455225 375537
rect 454905 375218 455225 375219
rect 454905 372537 455225 372538
rect 454905 372219 454906 372537
rect 455224 372219 455225 372537
rect 454905 372218 455225 372219
rect 120572 372088 129377 372112
rect 120572 371816 129081 372088
rect 129353 371816 129377 372088
rect 120572 371792 129377 371816
rect 454905 369537 455225 369538
rect 454905 369219 454906 369537
rect 455224 369219 455225 369537
rect 454905 369218 455225 369219
rect 120572 368088 129377 368112
rect 120572 367816 129081 368088
rect 129353 367816 129377 368088
rect 120572 367792 129377 367816
rect 454905 366537 455225 366538
rect 454905 366219 454906 366537
rect 455224 366219 455225 366537
rect 454905 366218 455225 366219
rect 120572 364088 129377 364112
rect 120572 363816 129081 364088
rect 129353 363816 129377 364088
rect 120572 363792 129377 363816
rect 454905 363537 455225 363538
rect 454905 363219 454906 363537
rect 455224 363219 455225 363537
rect 454905 363218 455225 363219
rect 454905 360537 455225 360538
rect 454905 360219 454906 360537
rect 455224 360219 455225 360537
rect 454905 360218 455225 360219
rect 120572 360088 129377 360112
rect 120572 359816 129081 360088
rect 129353 359816 129377 360088
rect 120572 359792 129377 359816
rect 454905 357537 455225 357538
rect 454905 357219 454906 357537
rect 455224 357219 455225 357537
rect 454905 357218 455225 357219
rect 120572 356088 129377 356112
rect 120572 355816 129081 356088
rect 129353 355816 129377 356088
rect 120572 355792 129377 355816
rect 454905 354537 455225 354538
rect 454905 354219 454906 354537
rect 455224 354219 455225 354537
rect 454905 354218 455225 354219
rect 120572 352088 129377 352112
rect 120572 351816 129081 352088
rect 129353 351816 129377 352088
rect 120572 351792 129377 351816
rect 454905 351537 455225 351538
rect 454905 351219 454906 351537
rect 455224 351219 455225 351537
rect 454905 351218 455225 351219
rect 454905 348537 455225 348538
rect 454905 348219 454906 348537
rect 455224 348219 455225 348537
rect 454905 348218 455225 348219
rect 120572 348088 129377 348112
rect 120572 347816 129081 348088
rect 129353 347816 129377 348088
rect 120572 347792 129377 347816
rect 454905 345537 455225 345538
rect 454905 345219 454906 345537
rect 455224 345219 455225 345537
rect 454905 345218 455225 345219
rect 120572 344088 129377 344112
rect 120572 343816 129081 344088
rect 129353 343816 129377 344088
rect 120572 343792 129377 343816
rect 454905 342537 455225 342538
rect 454905 342219 454906 342537
rect 455224 342219 455225 342537
rect 454905 342218 455225 342219
rect 120572 340088 129377 340112
rect 120572 339816 129081 340088
rect 129353 339816 129377 340088
rect 120572 339792 129377 339816
rect 454905 339537 455225 339538
rect 454905 339219 454906 339537
rect 455224 339219 455225 339537
rect 454905 339218 455225 339219
rect 454905 336537 455225 336538
rect 454905 336219 454906 336537
rect 455224 336219 455225 336537
rect 454905 336218 455225 336219
rect 120572 336088 129377 336112
rect 120572 335816 129081 336088
rect 129353 335816 129377 336088
rect 120572 335792 129377 335816
rect 454905 333537 455225 333538
rect 454905 333219 454906 333537
rect 455224 333219 455225 333537
rect 454905 333218 455225 333219
rect 120572 332088 129377 332112
rect 120572 331816 129081 332088
rect 129353 331816 129377 332088
rect 120572 331792 129377 331816
rect 454905 330537 455225 330538
rect 454905 330219 454906 330537
rect 455224 330219 455225 330537
rect 454905 330218 455225 330219
rect 120572 328088 129377 328112
rect 120572 327816 129081 328088
rect 129353 327816 129377 328088
rect 120572 327792 129377 327816
rect 454905 327537 455225 327538
rect 454905 327219 454906 327537
rect 455224 327219 455225 327537
rect 454905 327218 455225 327219
rect 454905 324537 455225 324538
rect 454905 324219 454906 324537
rect 455224 324219 455225 324537
rect 454905 324218 455225 324219
rect 120572 324088 129377 324112
rect 120572 323816 129081 324088
rect 129353 323816 129377 324088
rect 120572 323792 129377 323816
rect 454905 321537 455225 321538
rect 454905 321219 454906 321537
rect 455224 321219 455225 321537
rect 454905 321218 455225 321219
rect 120572 320088 129377 320112
rect 120572 319816 129081 320088
rect 129353 319816 129377 320088
rect 120572 319792 129377 319816
rect 454905 318537 455225 318538
rect 454905 318219 454906 318537
rect 455224 318219 455225 318537
rect 454905 318218 455225 318219
rect 120572 316088 129377 316112
rect 120572 315816 129081 316088
rect 129353 315816 129377 316088
rect 120572 315792 129377 315816
rect 454905 315537 455225 315538
rect 454905 315219 454906 315537
rect 455224 315219 455225 315537
rect 454905 315218 455225 315219
rect 454905 312537 455225 312538
rect 454905 312219 454906 312537
rect 455224 312219 455225 312537
rect 454905 312218 455225 312219
rect 120572 312088 129377 312112
rect 120572 311816 129081 312088
rect 129353 311816 129377 312088
rect 120572 311792 129377 311816
rect 454905 309537 455225 309538
rect 454905 309219 454906 309537
rect 455224 309219 455225 309537
rect 454905 309218 455225 309219
rect 120572 308088 129377 308112
rect 120572 307816 129081 308088
rect 129353 307816 129377 308088
rect 120572 307792 129377 307816
rect 454905 306537 455225 306538
rect 454905 306219 454906 306537
rect 455224 306219 455225 306537
rect 454905 306218 455225 306219
rect 120572 304088 129377 304112
rect 120572 303816 129081 304088
rect 129353 303816 129377 304088
rect 120572 303792 129377 303816
rect 454905 303537 455225 303538
rect 454905 303219 454906 303537
rect 455224 303219 455225 303537
rect 454905 303218 455225 303219
rect 454905 300537 455225 300538
rect 454905 300219 454906 300537
rect 455224 300219 455225 300537
rect 454905 300218 455225 300219
rect 120572 300088 129377 300112
rect 120572 299816 129081 300088
rect 129353 299816 129377 300088
rect 120572 299792 129377 299816
rect 454905 297537 455225 297538
rect 454905 297219 454906 297537
rect 455224 297219 455225 297537
rect 454905 297218 455225 297219
rect 120572 296088 129377 296112
rect 120572 295816 129081 296088
rect 129353 295816 129377 296088
rect 120572 295792 129377 295816
rect 454905 294537 455225 294538
rect 454905 294219 454906 294537
rect 455224 294219 455225 294537
rect 454905 294218 455225 294219
rect 120572 292088 129377 292112
rect 120572 291816 129081 292088
rect 129353 291816 129377 292088
rect 120572 291792 129377 291816
rect 454905 291537 455225 291538
rect 454905 291219 454906 291537
rect 455224 291219 455225 291537
rect 454905 291218 455225 291219
rect 454905 288537 455225 288538
rect 454905 288219 454906 288537
rect 455224 288219 455225 288537
rect 454905 288218 455225 288219
rect 120572 288088 129377 288112
rect 120572 287816 129081 288088
rect 129353 287816 129377 288088
rect 120572 287792 129377 287816
rect 454905 285537 455225 285538
rect 454905 285219 454906 285537
rect 455224 285219 455225 285537
rect 454905 285218 455225 285219
rect 120572 284088 129377 284112
rect 120572 283816 129081 284088
rect 129353 283816 129377 284088
rect 120572 283792 129377 283816
rect 454905 282537 455225 282538
rect 454905 282219 454906 282537
rect 455224 282219 455225 282537
rect 454905 282218 455225 282219
rect 120572 280088 129377 280112
rect 120572 279816 129081 280088
rect 129353 279816 129377 280088
rect 120572 279792 129377 279816
rect 454905 279537 455225 279538
rect 454905 279219 454906 279537
rect 455224 279219 455225 279537
rect 454905 279218 455225 279219
rect 454905 276537 455225 276538
rect 454905 276219 454906 276537
rect 455224 276219 455225 276537
rect 454905 276218 455225 276219
rect 120572 276088 129377 276112
rect 120572 275816 129081 276088
rect 129353 275816 129377 276088
rect 120572 275792 129377 275816
rect 454905 273537 455225 273538
rect 454905 273219 454906 273537
rect 455224 273219 455225 273537
rect 454905 273218 455225 273219
rect 120572 272088 129377 272112
rect 120572 271816 129081 272088
rect 129353 271816 129377 272088
rect 120572 271792 129377 271816
rect 454905 270537 455225 270538
rect 454905 270219 454906 270537
rect 455224 270219 455225 270537
rect 454905 270218 455225 270219
rect 120572 268088 129377 268112
rect 120572 267816 129081 268088
rect 129353 267816 129377 268088
rect 120572 267792 129377 267816
rect 454905 267537 455225 267538
rect 454905 267219 454906 267537
rect 455224 267219 455225 267537
rect 454905 267218 455225 267219
rect 454905 264537 455225 264538
rect 454905 264219 454906 264537
rect 455224 264219 455225 264537
rect 454905 264218 455225 264219
rect 120572 264088 129377 264112
rect 120572 263816 129081 264088
rect 129353 263816 129377 264088
rect 120572 263792 129377 263816
rect 454905 261537 455225 261538
rect 454905 261219 454906 261537
rect 455224 261219 455225 261537
rect 454905 261218 455225 261219
rect 24558 260523 24678 260524
rect 24558 260405 24559 260523
rect 24677 260405 24678 260523
rect 19138 253335 19258 254086
rect 19138 253217 19139 253335
rect 19257 253217 19258 253335
rect 19138 247349 19258 253217
rect 21326 253341 21446 253342
rect 21326 253223 21327 253341
rect 21445 253223 21446 253341
rect 21326 247553 21446 253223
rect 21325 247552 21447 247553
rect 21325 247432 21326 247552
rect 21446 247432 21447 247552
rect 21325 247431 21447 247432
rect 19137 247348 19259 247349
rect 19137 247228 19138 247348
rect 19258 247228 19259 247348
rect 19137 247227 19259 247228
rect 24558 245563 24678 260405
rect 120572 260088 129377 260112
rect 120572 259816 129081 260088
rect 129353 259816 129377 260088
rect 120572 259792 129377 259816
rect 27250 258973 27370 258974
rect 27250 258855 27251 258973
rect 27369 258855 27370 258973
rect 24557 245562 24679 245563
rect 24557 245442 24558 245562
rect 24678 245442 24679 245562
rect 24557 245441 24679 245442
rect 27250 244827 27370 258855
rect 454905 258537 455225 258538
rect 454905 258219 454906 258537
rect 455224 258219 455225 258537
rect 454905 258218 455225 258219
rect 120572 256088 129377 256112
rect 120572 255816 129081 256088
rect 129353 255816 129377 256088
rect 120572 255792 129377 255816
rect 454905 255537 455225 255538
rect 454905 255219 454906 255537
rect 455224 255219 455225 255537
rect 454905 255218 455225 255219
rect 454905 252537 455225 252538
rect 454905 252219 454906 252537
rect 455224 252219 455225 252537
rect 454905 252218 455225 252219
rect 120572 252088 129377 252112
rect 120572 251816 129081 252088
rect 129353 251816 129377 252088
rect 120572 251792 129377 251816
rect 454905 249537 455225 249538
rect 454905 249219 454906 249537
rect 455224 249219 455225 249537
rect 454905 249218 455225 249219
rect 120572 248088 129377 248112
rect 120572 247816 129081 248088
rect 129353 247816 129377 248088
rect 120572 247792 129377 247816
rect 454905 246537 455225 246538
rect 454905 246219 454906 246537
rect 455224 246219 455225 246537
rect 454905 246218 455225 246219
rect 27249 244826 27371 244827
rect 27249 244706 27250 244826
rect 27370 244706 27371 244826
rect 27249 244705 27371 244706
rect 120572 244088 129377 244112
rect 120572 243816 129081 244088
rect 129353 243816 129377 244088
rect 120572 243792 129377 243816
rect 454905 243537 455225 243538
rect 454905 243219 454906 243537
rect 455224 243219 455225 243537
rect 454905 243218 455225 243219
rect 454905 240537 455225 240538
rect 454905 240219 454906 240537
rect 455224 240219 455225 240537
rect 454905 240218 455225 240219
rect 120572 240088 129377 240112
rect 120572 239816 129081 240088
rect 129353 239816 129377 240088
rect 120572 239792 129377 239816
rect 454905 237537 455225 237538
rect 454905 237219 454906 237537
rect 455224 237219 455225 237537
rect 454905 237218 455225 237219
rect 120572 236088 129377 236112
rect 120572 235816 129081 236088
rect 129353 235816 129377 236088
rect 120572 235792 129377 235816
rect 454905 234537 455225 234538
rect 454905 234219 454906 234537
rect 455224 234219 455225 234537
rect 454905 234218 455225 234219
rect 120572 232088 129377 232112
rect 120572 231816 129081 232088
rect 129353 231816 129377 232088
rect 120572 231792 129377 231816
rect 454905 231537 455225 231538
rect 454905 231219 454906 231537
rect 455224 231219 455225 231537
rect 454905 231218 455225 231219
rect 454905 228537 455225 228538
rect 454905 228219 454906 228537
rect 455224 228219 455225 228537
rect 454905 228218 455225 228219
rect 120572 228088 129377 228112
rect 120572 227816 129081 228088
rect 129353 227816 129377 228088
rect 120572 227792 129377 227816
rect 454905 225537 455225 225538
rect 454905 225219 454906 225537
rect 455224 225219 455225 225537
rect 454905 225218 455225 225219
rect 120572 224088 129377 224112
rect 120572 223816 129081 224088
rect 129353 223816 129377 224088
rect 120572 223792 129377 223816
rect 454905 222537 455225 222538
rect 454905 222219 454906 222537
rect 455224 222219 455225 222537
rect 454905 222218 455225 222219
rect 120572 220088 129377 220112
rect 120572 219816 129081 220088
rect 129353 219816 129377 220088
rect 120572 219792 129377 219816
rect 454905 219537 455225 219538
rect 454905 219219 454906 219537
rect 455224 219219 455225 219537
rect 454905 219218 455225 219219
rect 454905 216537 455225 216538
rect 454905 216219 454906 216537
rect 455224 216219 455225 216537
rect 454905 216218 455225 216219
rect 120572 216088 129377 216112
rect 120572 215816 129081 216088
rect 129353 215816 129377 216088
rect 120572 215792 129377 215816
rect 454905 213537 455225 213538
rect 454905 213219 454906 213537
rect 455224 213219 455225 213537
rect 454905 213218 455225 213219
rect 120572 212088 129377 212112
rect 120572 211816 129081 212088
rect 129353 211816 129377 212088
rect 120572 211792 129377 211816
rect 454905 210537 455225 210538
rect 454905 210219 454906 210537
rect 455224 210219 455225 210537
rect 454905 210218 455225 210219
rect 120572 208088 129377 208112
rect 120572 207816 129081 208088
rect 129353 207816 129377 208088
rect 120572 207792 129377 207816
rect 454905 207537 455225 207538
rect 454905 207219 454906 207537
rect 455224 207219 455225 207537
rect 454905 207218 455225 207219
rect 454905 204537 455225 204538
rect 454905 204219 454906 204537
rect 455224 204219 455225 204537
rect 454905 204218 455225 204219
rect 120572 204088 129377 204112
rect 120572 203816 129081 204088
rect 129353 203816 129377 204088
rect 120572 203792 129377 203816
rect 454905 201537 455225 201538
rect 454905 201219 454906 201537
rect 455224 201219 455225 201537
rect 454905 201218 455225 201219
rect 120572 200088 129377 200112
rect 120572 199816 129081 200088
rect 129353 199816 129377 200088
rect 120572 199792 129377 199816
rect 454905 198537 455225 198538
rect 454905 198219 454906 198537
rect 455224 198219 455225 198537
rect 454905 198218 455225 198219
rect 120572 196088 129377 196112
rect 120572 195816 129081 196088
rect 129353 195816 129377 196088
rect 120572 195792 129377 195816
rect 454905 195537 455225 195538
rect 454905 195219 454906 195537
rect 455224 195219 455225 195537
rect 454905 195218 455225 195219
rect 454905 192537 455225 192538
rect 454905 192219 454906 192537
rect 455224 192219 455225 192537
rect 454905 192218 455225 192219
rect 120572 192088 129377 192112
rect 120572 191816 129081 192088
rect 129353 191816 129377 192088
rect 120572 191792 129377 191816
rect 10673 191537 10785 191538
rect 10673 191427 10674 191537
rect 10784 191427 10785 191537
rect 10673 191426 10785 191427
rect 9010 191342 9132 191343
rect 9010 191232 9011 191342
rect 9131 191232 9132 191342
rect 9010 191231 9132 191232
rect 454905 189537 455225 189538
rect 454905 189219 454906 189537
rect 455224 189219 455225 189537
rect 454905 189218 455225 189219
rect 120572 188088 129377 188112
rect 120572 187816 129081 188088
rect 129353 187816 129377 188088
rect 120572 187792 129377 187816
rect 454905 186537 455225 186538
rect 454905 186219 454906 186537
rect 455224 186219 455225 186537
rect 454905 186218 455225 186219
rect 4379 181780 4624 184240
rect 120572 184088 129377 184112
rect 120572 183816 129081 184088
rect 129353 183816 129377 184088
rect 120572 183792 129377 183816
rect 454905 183537 455225 183538
rect 454905 183219 454906 183537
rect 455224 183219 455225 183537
rect 454905 183218 455225 183219
rect 454905 180537 455225 180538
rect 454905 180219 454906 180537
rect 455224 180219 455225 180537
rect 454905 180218 455225 180219
rect 120572 180088 129377 180112
rect 120572 179816 129081 180088
rect 129353 179816 129377 180088
rect 120572 179792 129377 179816
rect 2440 178762 4664 178862
rect 1919 174762 2440 178276
rect 2540 174862 3090 178276
rect 1919 164695 3090 174762
rect 2175 163346 3090 164695
rect 4564 160876 4664 178762
rect 454905 177537 455225 177538
rect 454905 177219 454906 177537
rect 455224 177219 455225 177537
rect 454905 177218 455225 177219
rect 120572 176088 129377 176112
rect 120572 175816 129081 176088
rect 129353 175816 129377 176088
rect 120572 175792 129377 175816
rect 454905 174537 455225 174538
rect 454905 174219 454906 174537
rect 455224 174219 455225 174537
rect 454905 174218 455225 174219
rect 120572 172088 129377 172112
rect 120572 171816 129081 172088
rect 129353 171816 129377 172088
rect 120572 171792 129377 171816
rect 454905 171537 455225 171538
rect 454905 171219 454906 171537
rect 455224 171219 455225 171537
rect 454905 171218 455225 171219
rect 454905 168537 455225 168538
rect 454905 168219 454906 168537
rect 455224 168219 455225 168537
rect 454905 168218 455225 168219
rect 120572 168088 129377 168112
rect 120572 167816 129081 168088
rect 129353 167816 129377 168088
rect 120572 167792 129377 167816
rect 454905 165537 455225 165538
rect 454905 165219 454906 165537
rect 455224 165219 455225 165537
rect 454905 165218 455225 165219
rect 120572 164088 129377 164112
rect 120572 163816 129081 164088
rect 129353 163816 129377 164088
rect 120572 163792 129377 163816
rect 454905 162537 455225 162538
rect 454905 162219 454906 162537
rect 455224 162219 455225 162537
rect 454905 162218 455225 162219
rect 2622 160776 4664 160876
rect 1033 118976 1135 118977
rect 2622 118976 2722 160776
rect 120572 160088 129377 160112
rect 120572 159816 129081 160088
rect 129353 159816 129377 160088
rect 120572 159792 129377 159816
rect 454905 159537 455225 159538
rect 454905 159219 454906 159537
rect 455224 159219 455225 159537
rect 454905 159218 455225 159219
rect 454905 156537 455225 156538
rect 454905 156219 454906 156537
rect 455224 156219 455225 156537
rect 454905 156218 455225 156219
rect 120572 156088 129377 156112
rect 120572 155816 129081 156088
rect 129353 155816 129377 156088
rect 120572 155792 129377 155816
rect 454905 153537 455225 153538
rect 454905 153219 454906 153537
rect 455224 153219 455225 153537
rect 454905 153218 455225 153219
rect 120572 152088 129377 152112
rect 120572 151816 129081 152088
rect 129353 151816 129377 152088
rect 120572 151792 129377 151816
rect 454905 150537 455225 150538
rect 454905 150219 454906 150537
rect 455224 150219 455225 150537
rect 454905 150218 455225 150219
rect 120572 148088 129377 148112
rect 120572 147816 129081 148088
rect 129353 147816 129377 148088
rect 120572 147792 129377 147816
rect 490227 145105 493561 661830
rect 534064 644852 543338 645740
rect 534064 639522 535706 644852
rect 541456 639522 543338 644852
rect 534064 639002 543338 639522
rect 534308 634678 543582 635078
rect 534308 629610 536566 634678
rect 541812 629610 543582 634678
rect 534308 628340 543582 629610
rect 577922 629014 578088 629044
rect 577922 628906 577936 629014
rect 578044 628906 578088 629014
rect 577922 628894 578088 628906
rect 577935 625014 578045 625015
rect 577935 624906 577936 625014
rect 578044 624906 578045 625014
rect 508868 559006 533522 559030
rect 508868 557261 528746 559006
rect 508868 556624 509895 557261
rect 510532 556624 528746 557261
rect 508868 554254 528746 556624
rect 533498 554254 533522 559006
rect 508868 554230 533522 554254
rect 577935 539255 578045 624906
rect 577935 539145 582651 539255
rect 511640 473922 537996 473946
rect 511640 469170 533220 473922
rect 537972 469170 537996 473922
rect 511640 469146 537996 469170
rect 507116 457972 534522 457996
rect 507116 453220 507140 457972
rect 511892 453220 534522 457972
rect 507116 453196 534522 453220
rect 515384 438543 515386 438544
rect 515384 438213 515385 438543
rect 515384 438212 515386 438213
rect 515384 435543 515386 435544
rect 515384 435213 515385 435543
rect 515384 435212 515386 435213
rect 515384 432543 515386 432544
rect 515384 432213 515385 432543
rect 515384 432212 515386 432213
rect 515384 429543 515386 429544
rect 515384 429213 515385 429543
rect 515384 429212 515386 429213
rect 515384 426543 515386 426544
rect 515384 426213 515385 426543
rect 515384 426212 515386 426213
rect 515384 423543 515386 423544
rect 515384 423213 515385 423543
rect 515384 423212 515386 423213
rect 515384 420543 515386 420544
rect 515384 420213 515385 420543
rect 515384 420212 515386 420213
rect 515384 417543 515386 417544
rect 515384 417213 515385 417543
rect 515384 417212 515386 417213
rect 515384 414543 515386 414544
rect 515384 414213 515385 414543
rect 515384 414212 515386 414213
rect 515384 411543 515386 411544
rect 515384 411213 515385 411543
rect 515384 411212 515386 411213
rect 515384 408543 515386 408544
rect 515384 408213 515385 408543
rect 515384 408212 515386 408213
rect 515384 405543 515386 405544
rect 515384 405213 515385 405543
rect 515384 405212 515386 405213
rect 515384 402543 515386 402544
rect 515384 402213 515385 402543
rect 515384 402212 515386 402213
rect 515384 399543 515386 399544
rect 515384 399213 515385 399543
rect 515384 399212 515386 399213
rect 515384 396543 515386 396544
rect 515384 396213 515385 396543
rect 515384 396212 515386 396213
rect 515384 393543 515386 393544
rect 515384 393213 515385 393543
rect 515384 393212 515386 393213
rect 515384 390543 515386 390544
rect 515384 390213 515385 390543
rect 515384 390212 515386 390213
rect 515384 387543 515386 387544
rect 515384 387213 515385 387543
rect 515384 387212 515386 387213
rect 515384 384543 515386 384544
rect 515384 384213 515385 384543
rect 515384 384212 515386 384213
rect 515384 381543 515386 381544
rect 515384 381213 515385 381543
rect 515384 381212 515386 381213
rect 515384 378543 515386 378544
rect 515384 378213 515385 378543
rect 515384 378212 515386 378213
rect 515384 375543 515386 375544
rect 515384 375213 515385 375543
rect 515384 375212 515386 375213
rect 515384 372543 515386 372544
rect 515384 372213 515385 372543
rect 515384 372212 515386 372213
rect 515384 369543 515386 369544
rect 515384 369213 515385 369543
rect 515384 369212 515386 369213
rect 582541 368886 582651 539145
rect 582541 368786 582546 368886
rect 582646 368786 582651 368886
rect 515384 366543 515386 366544
rect 515384 366213 515385 366543
rect 515384 366212 515386 366213
rect 582541 364996 582651 368786
rect 582436 364886 582756 364996
rect 582436 364786 582546 364886
rect 582646 364786 582756 364886
rect 582436 364676 582756 364786
rect 515384 363543 515386 363544
rect 515384 363213 515385 363543
rect 515384 363212 515386 363213
rect 515384 360543 515386 360544
rect 515384 360213 515385 360543
rect 515384 360212 515386 360213
rect 515384 357543 515386 357544
rect 515384 357213 515385 357543
rect 515384 357212 515386 357213
rect 515384 354543 515386 354544
rect 515384 354213 515385 354543
rect 515384 354212 515386 354213
rect 515384 351543 515386 351544
rect 515384 351213 515385 351543
rect 515384 351212 515386 351213
rect 515384 348543 515386 348544
rect 515384 348213 515385 348543
rect 515384 348212 515386 348213
rect 515384 345543 515386 345544
rect 515384 345213 515385 345543
rect 515384 345212 515386 345213
rect 515384 342543 515386 342544
rect 515384 342213 515385 342543
rect 515384 342212 515386 342213
rect 515384 339543 515386 339544
rect 515384 339213 515385 339543
rect 515384 339212 515386 339213
rect 515384 336543 515386 336544
rect 515384 336213 515385 336543
rect 515384 336212 515386 336213
rect 515384 333543 515386 333544
rect 515384 333213 515385 333543
rect 515384 333212 515386 333213
rect 515384 330543 515386 330544
rect 515384 330213 515385 330543
rect 515384 330212 515386 330213
rect 515384 327543 515386 327544
rect 515384 327213 515385 327543
rect 515384 327212 515386 327213
rect 515384 324543 515386 324544
rect 515384 324213 515385 324543
rect 515384 324212 515386 324213
rect 582541 323646 582651 364676
rect 582541 323546 582546 323646
rect 582646 323546 582651 323646
rect 515384 321543 515386 321544
rect 515384 321213 515385 321543
rect 515384 321212 515386 321213
rect 582541 319756 582651 323546
rect 582436 319646 582756 319756
rect 582436 319546 582546 319646
rect 582646 319546 582756 319646
rect 582436 319436 582756 319546
rect 515384 318543 515386 318544
rect 515384 318213 515385 318543
rect 515384 318212 515386 318213
rect 515384 315543 515386 315544
rect 515384 315213 515385 315543
rect 515384 315212 515386 315213
rect 515384 312543 515386 312544
rect 515384 312213 515385 312543
rect 515384 312212 515386 312213
rect 515384 309543 515386 309544
rect 515384 309213 515385 309543
rect 515384 309212 515386 309213
rect 515384 306543 515386 306544
rect 515384 306213 515385 306543
rect 515384 306212 515386 306213
rect 515384 303543 515386 303544
rect 515384 303213 515385 303543
rect 515384 303212 515386 303213
rect 515384 300543 515386 300544
rect 515384 300213 515385 300543
rect 515384 300212 515386 300213
rect 515384 297543 515386 297544
rect 515384 297213 515385 297543
rect 515384 297212 515386 297213
rect 515384 294543 515386 294544
rect 515384 294213 515385 294543
rect 515384 294212 515386 294213
rect 515384 291543 515386 291544
rect 515384 291213 515385 291543
rect 515384 291212 515386 291213
rect 515384 288543 515386 288544
rect 515384 288213 515385 288543
rect 515384 288212 515386 288213
rect 515384 285543 515386 285544
rect 515384 285213 515385 285543
rect 515384 285212 515386 285213
rect 515384 282543 515386 282544
rect 515384 282213 515385 282543
rect 515384 282212 515386 282213
rect 515384 279543 515386 279544
rect 515384 279213 515385 279543
rect 515384 279212 515386 279213
rect 582541 279246 582651 319436
rect 582541 279146 582546 279246
rect 582646 279146 582651 279246
rect 515384 276543 515386 276544
rect 515384 276213 515385 276543
rect 515384 276212 515386 276213
rect 582541 275356 582651 279146
rect 582436 275246 582756 275356
rect 582436 275146 582546 275246
rect 582646 275146 582756 275246
rect 582436 275036 582756 275146
rect 515384 273543 515386 273544
rect 515384 273213 515385 273543
rect 515384 273212 515386 273213
rect 515384 270543 515386 270544
rect 515384 270213 515385 270543
rect 515384 270212 515386 270213
rect 515384 267543 515386 267544
rect 515384 267213 515385 267543
rect 515384 267212 515386 267213
rect 515384 264543 515386 264544
rect 515384 264213 515385 264543
rect 515384 264212 515386 264213
rect 515384 261543 515386 261544
rect 515384 261213 515385 261543
rect 515384 261212 515386 261213
rect 515384 258543 515386 258544
rect 515384 258213 515385 258543
rect 515384 258212 515386 258213
rect 515384 255543 515386 255544
rect 515384 255213 515385 255543
rect 515384 255212 515386 255213
rect 515384 252543 515386 252544
rect 515384 252213 515385 252543
rect 515384 252212 515386 252213
rect 515384 249543 515386 249544
rect 515384 249213 515385 249543
rect 515384 249212 515386 249213
rect 515384 246543 515386 246544
rect 515384 246213 515385 246543
rect 515384 246212 515386 246213
rect 515384 243543 515386 243544
rect 515384 243213 515385 243543
rect 515384 243212 515386 243213
rect 580888 242005 581188 245316
rect 582541 242005 582651 275036
rect 580888 241895 582651 242005
rect 515384 240543 515386 240544
rect 515384 240213 515385 240543
rect 515384 240212 515386 240213
rect 515384 237543 515386 237544
rect 515384 237213 515385 237543
rect 515384 237212 515386 237213
rect 515384 234543 515386 234544
rect 515384 234213 515385 234543
rect 515384 234212 515386 234213
rect 515384 231543 515386 231544
rect 515384 231213 515385 231543
rect 515384 231212 515386 231213
rect 515384 228543 515386 228544
rect 515384 228213 515385 228543
rect 515384 228212 515386 228213
rect 515384 225543 515386 225544
rect 515384 225213 515385 225543
rect 515384 225212 515386 225213
rect 515384 222543 515386 222544
rect 515384 222213 515385 222543
rect 515384 222212 515386 222213
rect 515384 219543 515386 219544
rect 515384 219213 515385 219543
rect 515384 219212 515386 219213
rect 515384 216543 515386 216544
rect 515384 216213 515385 216543
rect 515384 216212 515386 216213
rect 515384 213543 515386 213544
rect 515384 213213 515385 213543
rect 515384 213212 515386 213213
rect 515384 210543 515386 210544
rect 515384 210213 515385 210543
rect 515384 210212 515386 210213
rect 515384 207543 515386 207544
rect 515384 207213 515385 207543
rect 515384 207212 515386 207213
rect 515384 204543 515386 204544
rect 515384 204213 515385 204543
rect 515384 204212 515386 204213
rect 515384 201543 515386 201544
rect 515384 201213 515385 201543
rect 515384 201212 515386 201213
rect 515384 198543 515386 198544
rect 515384 198213 515385 198543
rect 515384 198212 515386 198213
rect 552812 196966 579468 198242
rect 515384 195543 515386 195544
rect 515384 195213 515385 195543
rect 515384 195212 515386 195213
rect 515384 192543 515386 192544
rect 515384 192213 515385 192543
rect 515384 192212 515386 192213
rect 552812 191768 554140 196966
rect 578296 191768 579468 196966
rect 552812 190928 579468 191768
rect 515384 189543 515386 189544
rect 515384 189213 515385 189543
rect 515384 189212 515386 189213
rect 515384 186543 515386 186544
rect 515384 186213 515385 186543
rect 515384 186212 515386 186213
rect 551320 186340 579660 187154
rect 515384 183543 515386 183544
rect 515384 183213 515385 183543
rect 515384 183212 515386 183213
rect 551320 181150 553050 186340
rect 576862 181150 579660 186340
rect 515384 180543 515386 180544
rect 515384 180213 515385 180543
rect 551320 180540 579660 181150
rect 515384 180212 515386 180213
rect 515384 177543 515386 177544
rect 515384 177213 515385 177543
rect 515384 177212 515386 177213
rect 515384 174543 515386 174544
rect 515384 174213 515385 174543
rect 515384 174212 515386 174213
rect 515384 171543 515386 171544
rect 515384 171213 515385 171543
rect 515384 171212 515386 171213
rect 515384 168543 515386 168544
rect 515384 168213 515385 168543
rect 515384 168212 515386 168213
rect 515384 165543 515386 165544
rect 515384 165213 515385 165543
rect 515384 165212 515386 165213
rect 552718 164209 558786 164626
rect 515384 162543 515386 162544
rect 515384 162213 515385 162543
rect 515384 162212 515386 162213
rect 515384 159543 515386 159544
rect 515384 159213 515385 159543
rect 515384 159212 515386 159213
rect 552718 159411 553277 164209
rect 558075 159411 558786 164209
rect 552718 158880 558786 159411
rect 580888 159120 581188 241895
rect 582541 241680 582651 241895
rect 580888 158290 581422 159120
rect 515384 156543 515386 156544
rect 515384 156213 515385 156543
rect 515384 156212 515386 156213
rect 515384 153543 515386 153544
rect 515384 153213 515385 153543
rect 515384 153212 515386 153213
rect 515384 150543 515386 150544
rect 515384 150213 515385 150543
rect 515384 150212 515386 150213
rect 120572 144088 129377 144112
rect 120572 143816 129081 144088
rect 129353 143816 129377 144088
rect 120572 143792 129377 143816
rect 462379 141771 493561 145105
rect 499374 141266 500790 141267
rect 494841 141242 499375 141266
rect 120572 140088 129377 140112
rect 120572 139816 129081 140088
rect 129353 139816 129377 140088
rect 494841 139876 495525 141242
rect 496891 139876 499375 141242
rect 494841 139852 499375 139876
rect 500789 141265 507515 141266
rect 500789 139853 503116 141265
rect 504528 140997 507515 141265
rect 504528 140121 505628 140997
rect 506504 140121 507515 140997
rect 504528 139853 507515 140121
rect 500789 139852 507515 139853
rect 499374 139851 500790 139852
rect 120572 139792 129377 139816
rect 459182 134644 459867 134700
rect 453395 134620 461504 134644
rect 453395 134348 453419 134620
rect 453691 134348 461504 134620
rect 453395 134324 461504 134348
rect 144646 129153 145734 129154
rect 144646 128067 144647 129153
rect 145733 128067 145734 129153
rect 144646 128066 145734 128067
rect 459182 127150 459867 134324
rect 581122 132708 581422 158290
rect 582515 132708 582625 134578
rect 581122 132408 582720 132708
rect 463530 127150 464217 127151
rect 459182 126465 463531 127150
rect 464216 126465 557323 127150
rect 463530 126464 464217 126465
rect 1033 118876 1034 118976
rect 1134 118876 2722 118976
rect 1033 118875 1135 118876
rect 1033 75776 1135 75777
rect 2622 75776 2722 118876
rect 150296 115072 150616 115096
rect 150296 114800 150320 115072
rect 150592 114800 150616 115072
rect 150296 95142 150616 114800
rect 153296 115072 153616 115096
rect 153296 114800 153320 115072
rect 153592 114800 153616 115072
rect 153296 95142 153616 114800
rect 156296 115072 156616 115096
rect 156296 114800 156320 115072
rect 156592 114800 156616 115072
rect 156296 95142 156616 114800
rect 159296 115072 159616 115096
rect 159296 114800 159320 115072
rect 159592 114800 159616 115072
rect 159296 95142 159616 114800
rect 162296 115072 162616 115096
rect 162296 114800 162320 115072
rect 162592 114800 162616 115072
rect 162296 95142 162616 114800
rect 165296 115072 165616 115096
rect 165296 114800 165320 115072
rect 165592 114800 165616 115072
rect 165296 95142 165616 114800
rect 168296 115072 168616 115096
rect 168296 114800 168320 115072
rect 168592 114800 168616 115072
rect 168296 95142 168616 114800
rect 171296 115072 171616 115096
rect 171296 114800 171320 115072
rect 171592 114800 171616 115072
rect 171296 95142 171616 114800
rect 174296 115072 174616 115096
rect 174296 114800 174320 115072
rect 174592 114800 174616 115072
rect 174296 95142 174616 114800
rect 177296 115072 177616 115096
rect 177296 114800 177320 115072
rect 177592 114800 177616 115072
rect 177296 95142 177616 114800
rect 180296 115072 180616 115096
rect 180296 114800 180320 115072
rect 180592 114800 180616 115072
rect 180296 95142 180616 114800
rect 183296 115072 183616 115096
rect 183296 114800 183320 115072
rect 183592 114800 183616 115072
rect 183296 95142 183616 114800
rect 186296 115072 186616 115096
rect 186296 114800 186320 115072
rect 186592 114800 186616 115072
rect 186296 95142 186616 114800
rect 189296 115072 189616 115096
rect 189296 114800 189320 115072
rect 189592 114800 189616 115072
rect 189296 95142 189616 114800
rect 192296 115072 192616 115096
rect 192296 114800 192320 115072
rect 192592 114800 192616 115072
rect 192296 95142 192616 114800
rect 195296 115072 195616 115096
rect 195296 114800 195320 115072
rect 195592 114800 195616 115072
rect 195296 95142 195616 114800
rect 198296 115072 198616 115096
rect 198296 114800 198320 115072
rect 198592 114800 198616 115072
rect 198296 95142 198616 114800
rect 201296 115072 201616 115096
rect 201296 114800 201320 115072
rect 201592 114800 201616 115072
rect 201296 95142 201616 114800
rect 204296 115072 204616 115096
rect 204296 114800 204320 115072
rect 204592 114800 204616 115072
rect 204296 95142 204616 114800
rect 207296 115072 207616 115096
rect 207296 114800 207320 115072
rect 207592 114800 207616 115072
rect 207296 95142 207616 114800
rect 210296 115072 210616 115096
rect 210296 114800 210320 115072
rect 210592 114800 210616 115072
rect 210296 95142 210616 114800
rect 213296 115072 213616 115096
rect 213296 114800 213320 115072
rect 213592 114800 213616 115072
rect 213296 95142 213616 114800
rect 216296 115072 216616 115096
rect 216296 114800 216320 115072
rect 216592 114800 216616 115072
rect 216296 95142 216616 114800
rect 219296 115072 219616 115096
rect 219296 114800 219320 115072
rect 219592 114800 219616 115072
rect 219296 95142 219616 114800
rect 222296 115072 222616 115096
rect 222296 114800 222320 115072
rect 222592 114800 222616 115072
rect 222296 95142 222616 114800
rect 225296 115072 225616 115096
rect 225296 114800 225320 115072
rect 225592 114800 225616 115072
rect 225296 95142 225616 114800
rect 228296 115072 228616 115096
rect 228296 114800 228320 115072
rect 228592 114800 228616 115072
rect 228296 95142 228616 114800
rect 231296 115072 231616 115096
rect 231296 114800 231320 115072
rect 231592 114800 231616 115072
rect 231296 95142 231616 114800
rect 234296 115072 234616 115096
rect 234296 114800 234320 115072
rect 234592 114800 234616 115072
rect 234296 95142 234616 114800
rect 237296 115072 237616 115096
rect 237296 114800 237320 115072
rect 237592 114800 237616 115072
rect 237296 95142 237616 114800
rect 240296 115072 240616 115096
rect 240296 114800 240320 115072
rect 240592 114800 240616 115072
rect 240296 95142 240616 114800
rect 243296 115072 243616 115096
rect 243296 114800 243320 115072
rect 243592 114800 243616 115072
rect 243296 95142 243616 114800
rect 246296 115072 246616 115096
rect 246296 114800 246320 115072
rect 246592 114800 246616 115072
rect 246296 95142 246616 114800
rect 249296 115072 249616 115096
rect 249296 114800 249320 115072
rect 249592 114800 249616 115072
rect 249296 95142 249616 114800
rect 252296 115072 252616 115096
rect 252296 114800 252320 115072
rect 252592 114800 252616 115072
rect 252296 95142 252616 114800
rect 255296 115072 255616 115096
rect 255296 114800 255320 115072
rect 255592 114800 255616 115072
rect 255296 95142 255616 114800
rect 258296 115072 258616 115096
rect 258296 114800 258320 115072
rect 258592 114800 258616 115072
rect 258296 95142 258616 114800
rect 261296 115072 261616 115096
rect 261296 114800 261320 115072
rect 261592 114800 261616 115072
rect 261296 95142 261616 114800
rect 264296 115072 264616 115096
rect 264296 114800 264320 115072
rect 264592 114800 264616 115072
rect 264296 95142 264616 114800
rect 267296 115072 267616 115096
rect 267296 114800 267320 115072
rect 267592 114800 267616 115072
rect 267296 95142 267616 114800
rect 270296 115072 270616 115096
rect 270296 114800 270320 115072
rect 270592 114800 270616 115072
rect 270296 95142 270616 114800
rect 273296 115072 273616 115096
rect 273296 114800 273320 115072
rect 273592 114800 273616 115072
rect 273296 95142 273616 114800
rect 276296 115072 276616 115096
rect 276296 114800 276320 115072
rect 276592 114800 276616 115072
rect 276296 95142 276616 114800
rect 279296 115072 279616 115096
rect 279296 114800 279320 115072
rect 279592 114800 279616 115072
rect 279296 95142 279616 114800
rect 282296 115072 282616 115096
rect 282296 114800 282320 115072
rect 282592 114800 282616 115072
rect 282296 95142 282616 114800
rect 285296 115072 285616 115096
rect 285296 114800 285320 115072
rect 285592 114800 285616 115072
rect 285296 95142 285616 114800
rect 288296 115072 288616 115096
rect 288296 114800 288320 115072
rect 288592 114800 288616 115072
rect 288296 95142 288616 114800
rect 291296 115072 291616 115096
rect 291296 114800 291320 115072
rect 291592 114800 291616 115072
rect 291296 95142 291616 114800
rect 294296 115072 294616 115096
rect 294296 114800 294320 115072
rect 294592 114800 294616 115072
rect 294296 95142 294616 114800
rect 297296 115072 297616 115096
rect 297296 114800 297320 115072
rect 297592 114800 297616 115072
rect 297296 95142 297616 114800
rect 300296 115072 300616 115096
rect 300296 114800 300320 115072
rect 300592 114800 300616 115072
rect 300296 95142 300616 114800
rect 303296 115072 303616 115096
rect 303296 114800 303320 115072
rect 303592 114800 303616 115072
rect 303296 95142 303616 114800
rect 306296 115072 306616 115096
rect 306296 114800 306320 115072
rect 306592 114800 306616 115072
rect 306296 95142 306616 114800
rect 309296 115072 309616 115096
rect 309296 114800 309320 115072
rect 309592 114800 309616 115072
rect 309296 95142 309616 114800
rect 312296 115072 312616 115096
rect 312296 114800 312320 115072
rect 312592 114800 312616 115072
rect 312296 95142 312616 114800
rect 315296 115072 315616 115096
rect 315296 114800 315320 115072
rect 315592 114800 315616 115072
rect 315296 95142 315616 114800
rect 318296 115072 318616 115096
rect 318296 114800 318320 115072
rect 318592 114800 318616 115072
rect 318296 95142 318616 114800
rect 321296 115072 321616 115096
rect 321296 114800 321320 115072
rect 321592 114800 321616 115072
rect 321296 95142 321616 114800
rect 324296 115072 324616 115096
rect 324296 114800 324320 115072
rect 324592 114800 324616 115072
rect 324296 95142 324616 114800
rect 327296 115072 327616 115096
rect 327296 114800 327320 115072
rect 327592 114800 327616 115072
rect 327296 95142 327616 114800
rect 330296 115072 330616 115096
rect 330296 114800 330320 115072
rect 330592 114800 330616 115072
rect 330296 95142 330616 114800
rect 333296 115072 333616 115096
rect 333296 114800 333320 115072
rect 333592 114800 333616 115072
rect 333296 95142 333616 114800
rect 336296 115072 336616 115096
rect 336296 114800 336320 115072
rect 336592 114800 336616 115072
rect 336296 95142 336616 114800
rect 339296 115072 339616 115096
rect 339296 114800 339320 115072
rect 339592 114800 339616 115072
rect 339296 95142 339616 114800
rect 342296 115072 342616 115096
rect 342296 114800 342320 115072
rect 342592 114800 342616 115072
rect 342296 95142 342616 114800
rect 345296 115072 345616 115096
rect 345296 114800 345320 115072
rect 345592 114800 345616 115072
rect 345296 95142 345616 114800
rect 348296 115072 348616 115096
rect 348296 114800 348320 115072
rect 348592 114800 348616 115072
rect 348296 95142 348616 114800
rect 351296 115072 351616 115096
rect 351296 114800 351320 115072
rect 351592 114800 351616 115072
rect 351296 95142 351616 114800
rect 354296 115072 354616 115096
rect 354296 114800 354320 115072
rect 354592 114800 354616 115072
rect 354296 95142 354616 114800
rect 357296 115072 357616 115096
rect 357296 114800 357320 115072
rect 357592 114800 357616 115072
rect 357296 95142 357616 114800
rect 360296 115072 360616 115096
rect 360296 114800 360320 115072
rect 360592 114800 360616 115072
rect 360296 95142 360616 114800
rect 363296 115072 363616 115096
rect 363296 114800 363320 115072
rect 363592 114800 363616 115072
rect 363296 95142 363616 114800
rect 366296 115072 366616 115096
rect 366296 114800 366320 115072
rect 366592 114800 366616 115072
rect 366296 95142 366616 114800
rect 369296 115072 369616 115096
rect 369296 114800 369320 115072
rect 369592 114800 369616 115072
rect 369296 95142 369616 114800
rect 372296 115072 372616 115096
rect 372296 114800 372320 115072
rect 372592 114800 372616 115072
rect 372296 95142 372616 114800
rect 375296 115072 375616 115096
rect 375296 114800 375320 115072
rect 375592 114800 375616 115072
rect 375296 95142 375616 114800
rect 378296 115072 378616 115096
rect 378296 114800 378320 115072
rect 378592 114800 378616 115072
rect 378296 95142 378616 114800
rect 381296 115072 381616 115096
rect 381296 114800 381320 115072
rect 381592 114800 381616 115072
rect 381296 95142 381616 114800
rect 384296 115072 384616 115096
rect 384296 114800 384320 115072
rect 384592 114800 384616 115072
rect 384296 95142 384616 114800
rect 387296 115072 387616 115096
rect 387296 114800 387320 115072
rect 387592 114800 387616 115072
rect 387296 95142 387616 114800
rect 390296 115072 390616 115096
rect 390296 114800 390320 115072
rect 390592 114800 390616 115072
rect 390296 95142 390616 114800
rect 393296 115072 393616 115096
rect 393296 114800 393320 115072
rect 393592 114800 393616 115072
rect 393296 95142 393616 114800
rect 396296 115072 396616 115096
rect 396296 114800 396320 115072
rect 396592 114800 396616 115072
rect 396296 95142 396616 114800
rect 399296 115072 399616 115096
rect 399296 114800 399320 115072
rect 399592 114800 399616 115072
rect 399296 95142 399616 114800
rect 402296 115072 402616 115096
rect 402296 114800 402320 115072
rect 402592 114800 402616 115072
rect 402296 95142 402616 114800
rect 405296 115072 405616 115096
rect 405296 114800 405320 115072
rect 405592 114800 405616 115072
rect 405296 95142 405616 114800
rect 408296 115072 408616 115096
rect 408296 114800 408320 115072
rect 408592 114800 408616 115072
rect 408296 95142 408616 114800
rect 411296 115072 411616 115096
rect 411296 114800 411320 115072
rect 411592 114800 411616 115072
rect 411296 95142 411616 114800
rect 414296 115072 414616 115096
rect 414296 114800 414320 115072
rect 414592 114800 414616 115072
rect 414296 95142 414616 114800
rect 420296 115072 420616 115096
rect 420296 114800 420320 115072
rect 420592 114800 420616 115072
rect 417296 95142 417616 112994
rect 420296 95142 420616 114800
rect 423296 115072 423616 115096
rect 423296 114800 423320 115072
rect 423592 114800 423616 115072
rect 423296 95142 423616 114800
rect 426296 115072 426616 115096
rect 426296 114800 426320 115072
rect 426592 114800 426616 115072
rect 426296 95142 426616 114800
rect 429296 115072 429616 115096
rect 429296 114800 429320 115072
rect 429592 114800 429616 115072
rect 429296 95142 429616 114800
rect 432296 115072 432616 115096
rect 432296 114800 432320 115072
rect 432592 114800 432616 115072
rect 432296 95142 432616 114800
rect 435296 115072 435616 115096
rect 435296 114800 435320 115072
rect 435592 114800 435616 115072
rect 435296 95142 435616 114800
rect 438296 115072 438616 115096
rect 438296 114800 438320 115072
rect 438592 114800 438616 115072
rect 438296 95142 438616 114800
rect 441296 115072 441616 115096
rect 441296 114800 441320 115072
rect 441592 114800 441616 115072
rect 441296 95142 441616 114800
rect 444296 115072 444616 115096
rect 444296 114800 444320 115072
rect 444592 114800 444616 115072
rect 444296 95142 444616 114800
rect 464812 95142 465497 126465
rect 489067 95142 489752 126465
rect 582420 99246 582720 132408
rect 582420 99146 582546 99246
rect 582646 99146 582720 99246
rect 582420 95356 582720 99146
rect 582420 95246 582756 95356
rect 582420 95146 582546 95246
rect 582646 95146 582756 95246
rect 101340 95118 558076 95142
rect 101340 90366 553300 95118
rect 558052 90366 558076 95118
rect 101340 90342 558076 90366
rect 582420 95036 582756 95146
rect 150296 89870 150616 90342
rect 153296 89870 153616 90342
rect 156296 89870 156616 90342
rect 159296 89870 159616 90342
rect 162296 89870 162616 90342
rect 165296 89870 165616 90342
rect 168296 89870 168616 90342
rect 171296 89870 171616 90342
rect 174296 89870 174616 90342
rect 177296 89870 177616 90342
rect 180296 89870 180616 90342
rect 183296 89870 183616 90342
rect 186296 89870 186616 90342
rect 189296 89870 189616 90342
rect 192296 89870 192616 90342
rect 195296 89870 195616 90342
rect 198296 89870 198616 90342
rect 201296 89870 201616 90342
rect 204296 89870 204616 90342
rect 207296 89870 207616 90342
rect 210296 89870 210616 90342
rect 213296 89870 213616 90342
rect 216296 89870 216616 90342
rect 219296 89870 219616 90342
rect 222296 89870 222616 90342
rect 225296 89870 225616 90342
rect 228296 89870 228616 90342
rect 231296 89870 231616 90342
rect 234296 89870 234616 90342
rect 237296 89870 237616 90342
rect 240296 89870 240616 90342
rect 243296 89870 243616 90342
rect 246296 89870 246616 90342
rect 249296 89870 249616 90342
rect 252296 89870 252616 90342
rect 255296 89870 255616 90342
rect 258296 89870 258616 90342
rect 261296 89870 261616 90342
rect 264296 89870 264616 90342
rect 267296 89870 267616 90342
rect 270296 89870 270616 90342
rect 273296 89870 273616 90342
rect 276296 89870 276616 90342
rect 279296 89870 279616 90342
rect 282296 89870 282616 90342
rect 285296 89870 285616 90342
rect 288296 89870 288616 90342
rect 291296 89870 291616 90342
rect 294296 89870 294616 90342
rect 297296 89870 297616 90342
rect 300296 89870 300616 90342
rect 303296 89870 303616 90342
rect 306296 89870 306616 90342
rect 309296 89870 309616 90342
rect 312296 89870 312616 90342
rect 315296 89870 315616 90342
rect 318296 89870 318616 90342
rect 321296 89870 321616 90342
rect 324296 89870 324616 90342
rect 327296 89870 327616 90342
rect 330296 89870 330616 90342
rect 333296 89870 333616 90342
rect 336296 89870 336616 90342
rect 339296 89870 339616 90342
rect 342296 89870 342616 90342
rect 345296 89870 345616 90342
rect 348296 89870 348616 90342
rect 351296 89870 351616 90342
rect 354296 89870 354616 90342
rect 357296 89870 357616 90342
rect 360296 89870 360616 90342
rect 363296 89870 363616 90342
rect 366296 89870 366616 90342
rect 369296 89870 369616 90342
rect 372296 89870 372616 90342
rect 375296 89870 375616 90342
rect 378296 89870 378616 90342
rect 381296 89870 381616 90342
rect 384296 89870 384616 90342
rect 387296 89870 387616 90342
rect 390296 89870 390616 90342
rect 393296 89870 393616 90342
rect 396296 89870 396616 90342
rect 399296 89870 399616 90342
rect 402296 89870 402616 90342
rect 405296 89870 405616 90342
rect 408296 89870 408616 90342
rect 411296 89870 411616 90342
rect 414296 89870 414616 90342
rect 417296 89870 417616 90342
rect 420296 89870 420616 90342
rect 423296 89870 423616 90342
rect 426296 89870 426616 90342
rect 429296 89870 429616 90342
rect 432296 89870 432616 90342
rect 435296 89870 435616 90342
rect 438296 89870 438616 90342
rect 441296 89870 441616 90342
rect 444296 89870 444616 90342
rect 1033 75676 1034 75776
rect 1134 75676 2722 75776
rect 1033 75675 1135 75676
rect 1033 32376 1135 32377
rect 2622 32376 2722 75676
rect 1033 32276 1034 32376
rect 1134 32276 2722 32376
rect 1033 32275 1135 32276
rect 1033 10976 1135 10977
rect 2622 10976 2722 32276
rect 1033 10876 1034 10976
rect 1134 10876 2722 10976
rect 1033 10875 1135 10876
rect 2622 7266 2722 10876
rect 2324 6966 2866 7266
rect 353 4020 467 4021
rect 353 3908 354 4020
rect 466 3908 467 4020
rect 353 3907 467 3908
rect 2324 3730 2624 6966
rect 582420 3730 582720 95036
rect 2324 3430 582720 3730
<< via4 >>
rect 229597 697552 231180 699708
rect 329614 698285 334006 701834
rect 329614 697442 331192 698285
rect 331192 697442 332128 698285
rect 332128 697442 334006 698285
rect 303918 596606 304190 596630
rect 303894 596286 304214 596606
rect 303918 592534 304190 592806
rect 292338 591606 292610 591878
rect 338088 590140 338408 590460
rect 338088 586140 338408 586460
rect 308982 556600 309667 557285
rect 288563 473351 289093 473352
rect 288563 472811 288564 473351
rect 288564 472811 289093 473351
rect 288563 472810 289093 472811
rect 297407 471950 297777 471951
rect 297407 471570 297776 471950
rect 297776 471570 297777 471950
rect 297407 471569 297777 471570
rect 290884 469717 291524 469718
rect 290884 469067 291523 469717
rect 291523 469067 291524 469717
rect 334724 469170 339476 473922
rect 290884 469066 291524 469067
rect 162784 454558 163104 454878
rect 162808 438530 163080 438802
rect 165784 454558 166104 454878
rect 165808 438530 166080 438802
rect 168784 454558 169104 454878
rect 168808 438530 169080 438802
rect 171784 454558 172104 454878
rect 171808 438530 172080 438802
rect 174784 454558 175104 454878
rect 174808 438530 175080 438802
rect 177784 454558 178104 454878
rect 177808 438530 178080 438802
rect 180784 454558 181104 454878
rect 180808 438530 181080 438802
rect 183784 454558 184104 454878
rect 183808 438530 184080 438802
rect 186784 454558 187104 454878
rect 186808 438530 187080 438802
rect 189784 454558 190104 454878
rect 189808 438530 190080 438802
rect 192784 454558 193104 454878
rect 192808 438530 193080 438802
rect 195784 454558 196104 454878
rect 195808 438530 196080 438802
rect 198784 454558 199104 454878
rect 198808 438530 199080 438802
rect 201784 454558 202104 454878
rect 201808 438530 202080 438802
rect 204784 454558 205104 454878
rect 204808 438530 205080 438802
rect 207784 454558 208104 454878
rect 207808 438530 208080 438802
rect 210784 454558 211104 454878
rect 210808 438530 211080 438802
rect 213784 454558 214104 454878
rect 213808 438530 214080 438802
rect 216784 454558 217104 454878
rect 216808 438530 217080 438802
rect 219784 454558 220104 454878
rect 219808 438530 220080 438802
rect 222784 454558 223104 454878
rect 222808 438530 223080 438802
rect 225784 454558 226104 454878
rect 225808 438530 226080 438802
rect 228784 454558 229104 454878
rect 228808 438530 229080 438802
rect 231784 454558 232104 454878
rect 231808 438530 232080 438802
rect 234784 454558 235104 454878
rect 234808 438530 235080 438802
rect 237784 454558 238104 454878
rect 237808 438530 238080 438802
rect 240784 454558 241104 454878
rect 240808 438530 241080 438802
rect 243784 454558 244104 454878
rect 243808 438530 244080 438802
rect 246784 454558 247104 454878
rect 246808 438530 247080 438802
rect 249784 454558 250104 454878
rect 249808 438530 250080 438802
rect 252784 454558 253104 454878
rect 252808 438530 253080 438802
rect 255784 454558 256104 454878
rect 255808 438530 256080 438802
rect 258784 454558 259104 454878
rect 258808 438530 259080 438802
rect 261784 454558 262104 454878
rect 261808 438530 262080 438802
rect 264784 454558 265104 454878
rect 264808 438530 265080 438802
rect 267784 454558 268104 454878
rect 267808 438530 268080 438802
rect 270784 454558 271104 454878
rect 270808 438530 271080 438802
rect 273784 454558 274104 454878
rect 273808 438530 274080 438802
rect 276784 454558 277104 454878
rect 276808 438530 277080 438802
rect 279784 454558 280104 454878
rect 279808 438530 280080 438802
rect 282784 454558 283104 454878
rect 282808 438530 283080 438802
rect 285784 454558 286104 454878
rect 285808 438530 286080 438802
rect 288784 454558 289104 454878
rect 288808 438530 289080 438802
rect 291784 454558 292104 454878
rect 291808 438530 292080 438802
rect 294784 454558 295104 454878
rect 294808 438530 295080 438802
rect 297784 454558 298104 454878
rect 297808 438530 298080 438802
rect 300784 454558 301104 454878
rect 300808 438530 301080 438802
rect 303784 454558 304104 454878
rect 303808 438530 304080 438802
rect 306784 454558 307104 454878
rect 306808 438530 307080 438802
rect 309784 454558 310104 454878
rect 309808 438530 310080 438802
rect 312784 454558 313104 454878
rect 312808 438530 313080 438802
rect 315784 454558 316104 454878
rect 315808 438530 316080 438802
rect 318784 454558 319104 454878
rect 318808 438530 319080 438802
rect 321784 454558 322104 454878
rect 321808 438530 322080 438802
rect 324784 454558 325104 454878
rect 324808 438530 325080 438802
rect 327784 454558 328104 454878
rect 327808 438530 328080 438802
rect 330784 454558 331104 454878
rect 330808 438530 331080 438802
rect 333784 454558 334104 454878
rect 333808 438530 334080 438802
rect 336784 454558 337104 454878
rect 336808 438530 337080 438802
rect 339784 454558 340104 454878
rect 339808 438530 340080 438802
rect 342784 454558 343104 454878
rect 342808 438530 343080 438802
rect 345784 454558 346104 454878
rect 345808 438530 346080 438802
rect 348784 454558 349104 454878
rect 348808 438530 349080 438802
rect 351784 454558 352104 454878
rect 351808 438530 352080 438802
rect 354784 454558 355104 454878
rect 354808 438530 355080 438802
rect 357784 454558 358104 454878
rect 357808 438530 358080 438802
rect 360784 454558 361104 454878
rect 360808 438530 361080 438802
rect 363784 454558 364104 454878
rect 363808 438530 364080 438802
rect 366784 454558 367104 454878
rect 366808 438530 367080 438802
rect 369784 454558 370104 454878
rect 369808 438530 370080 438802
rect 372784 454558 373104 454878
rect 372808 438530 373080 438802
rect 375784 454558 376104 454878
rect 375808 438530 376080 438802
rect 378784 454558 379104 454878
rect 378808 438530 379080 438802
rect 381784 454558 382104 454878
rect 381808 438530 382080 438802
rect 384784 454558 385104 454878
rect 384808 438530 385080 438802
rect 387784 454558 388104 454878
rect 387808 438530 388080 438802
rect 390784 454558 391104 454878
rect 390808 438530 391080 438802
rect 393784 454558 394104 454878
rect 393808 438530 394080 438802
rect 396784 454558 397104 454878
rect 396808 438530 397080 438802
rect 399784 454558 400104 454878
rect 399808 438530 400080 438802
rect 402784 454558 403104 454878
rect 402808 438530 403080 438802
rect 405784 454558 406104 454878
rect 405808 438530 406080 438802
rect 408784 454558 409104 454878
rect 408808 438530 409080 438802
rect 411784 454558 412104 454878
rect 411808 438530 412080 438802
rect 414784 454558 415104 454878
rect 414808 438530 415080 438802
rect 417784 454558 418104 454878
rect 417808 438530 418080 438802
rect 420784 454558 421104 454878
rect 420808 438530 421080 438802
rect 423784 454558 424104 454878
rect 423808 438530 424080 438802
rect 426784 454558 427104 454878
rect 426808 438530 427080 438802
rect 429784 454558 430104 454878
rect 429808 438530 430080 438802
rect 432784 454558 433104 454878
rect 432808 438530 433080 438802
rect 435784 454558 436104 454878
rect 435808 438530 436080 438802
rect 438784 454558 439104 454878
rect 438808 438530 439080 438802
rect 441784 454558 442104 454878
rect 441808 438530 442080 438802
rect 444784 454558 445104 454878
rect 444808 438530 445080 438802
rect 447784 454558 448104 454878
rect 447808 438530 448080 438802
rect 454929 438242 455201 438514
rect 149126 436938 149398 437210
rect 149126 436194 149398 436466
rect 120252 435792 120572 436112
rect 129081 435816 129353 436088
rect 454929 435242 455201 435514
rect 454929 432242 455201 432514
rect 120252 431792 120572 432112
rect 129081 431816 129353 432088
rect 454929 429242 455201 429514
rect 120252 427792 120572 428112
rect 129081 427816 129353 428088
rect 454929 426242 455201 426514
rect 120252 423792 120572 424112
rect 129081 423816 129353 424088
rect 454929 423242 455201 423514
rect 454929 420242 455201 420514
rect 120252 419792 120572 420112
rect 129081 419816 129353 420088
rect 454929 417242 455201 417514
rect 120252 415792 120572 416112
rect 129081 415816 129353 416088
rect 454929 414242 455201 414514
rect 120252 411792 120572 412112
rect 129081 411816 129353 412088
rect 454929 411242 455201 411514
rect 454929 408242 455201 408514
rect 120252 407792 120572 408112
rect 129081 407816 129353 408088
rect 454929 405242 455201 405514
rect 120252 403792 120572 404112
rect 129081 403816 129353 404088
rect 454929 402242 455201 402514
rect 120252 399792 120572 400112
rect 129081 399816 129353 400088
rect 454929 399242 455201 399514
rect 454929 396242 455201 396514
rect 120252 395792 120572 396112
rect 129081 395816 129353 396088
rect 454929 393242 455201 393514
rect 120252 391792 120572 392112
rect 129081 391816 129353 392088
rect 454929 390242 455201 390514
rect 120252 387792 120572 388112
rect 129081 387816 129353 388088
rect 454929 387242 455201 387514
rect 454929 384242 455201 384514
rect 120252 383792 120572 384112
rect 129081 383816 129353 384088
rect 454929 381242 455201 381514
rect 120252 379792 120572 380112
rect 129081 379816 129353 380088
rect 454929 378242 455201 378514
rect 120252 375792 120572 376112
rect 129081 375816 129353 376088
rect 454929 375242 455201 375514
rect 454929 372242 455201 372514
rect 120252 371792 120572 372112
rect 129081 371816 129353 372088
rect 454929 369242 455201 369514
rect 120252 367792 120572 368112
rect 129081 367816 129353 368088
rect 454929 366242 455201 366514
rect 120252 363792 120572 364112
rect 129081 363816 129353 364088
rect 454929 363242 455201 363514
rect 454929 360242 455201 360514
rect 120252 359792 120572 360112
rect 129081 359816 129353 360088
rect 454929 357242 455201 357514
rect 120252 355792 120572 356112
rect 129081 355816 129353 356088
rect 454929 354242 455201 354514
rect 120252 351792 120572 352112
rect 129081 351816 129353 352088
rect 454929 351242 455201 351514
rect 454929 348242 455201 348514
rect 120252 347792 120572 348112
rect 129081 347816 129353 348088
rect 454929 345242 455201 345514
rect 120252 343792 120572 344112
rect 129081 343816 129353 344088
rect 454929 342242 455201 342514
rect 120252 339792 120572 340112
rect 129081 339816 129353 340088
rect 454929 339242 455201 339514
rect 454929 336242 455201 336514
rect 120252 335792 120572 336112
rect 129081 335816 129353 336088
rect 454929 333242 455201 333514
rect 120252 331792 120572 332112
rect 129081 331816 129353 332088
rect 454929 330242 455201 330514
rect 120252 327792 120572 328112
rect 129081 327816 129353 328088
rect 454929 327242 455201 327514
rect 454929 324242 455201 324514
rect 120252 323792 120572 324112
rect 129081 323816 129353 324088
rect 454929 321242 455201 321514
rect 120252 319792 120572 320112
rect 129081 319816 129353 320088
rect 454929 318242 455201 318514
rect 120252 315792 120572 316112
rect 129081 315816 129353 316088
rect 454929 315242 455201 315514
rect 454929 312242 455201 312514
rect 120252 311792 120572 312112
rect 129081 311816 129353 312088
rect 454929 309242 455201 309514
rect 120252 307792 120572 308112
rect 129081 307816 129353 308088
rect 454929 306242 455201 306514
rect 120252 303792 120572 304112
rect 129081 303816 129353 304088
rect 454929 303242 455201 303514
rect 454929 300242 455201 300514
rect 120252 299792 120572 300112
rect 129081 299816 129353 300088
rect 454929 297242 455201 297514
rect 120252 295792 120572 296112
rect 129081 295816 129353 296088
rect 454929 294242 455201 294514
rect 120252 291792 120572 292112
rect 129081 291816 129353 292088
rect 454929 291242 455201 291514
rect 454929 288242 455201 288514
rect 120252 287792 120572 288112
rect 129081 287816 129353 288088
rect 454929 285242 455201 285514
rect 120252 283792 120572 284112
rect 129081 283816 129353 284088
rect 454929 282242 455201 282514
rect 120252 279792 120572 280112
rect 129081 279816 129353 280088
rect 454929 279242 455201 279514
rect 454929 276242 455201 276514
rect 120252 275792 120572 276112
rect 129081 275816 129353 276088
rect 454929 273242 455201 273514
rect 120252 271792 120572 272112
rect 129081 271816 129353 272088
rect 454929 270242 455201 270514
rect 120252 267792 120572 268112
rect 129081 267816 129353 268088
rect 454929 267242 455201 267514
rect 454929 264242 455201 264514
rect 120252 263792 120572 264112
rect 129081 263816 129353 264088
rect 454929 261242 455201 261514
rect 120252 259792 120572 260112
rect 129081 259816 129353 260088
rect 454929 258242 455201 258514
rect 120252 255792 120572 256112
rect 129081 255816 129353 256088
rect 454929 255242 455201 255514
rect 454929 252242 455201 252514
rect 120252 251792 120572 252112
rect 129081 251816 129353 252088
rect 454929 249242 455201 249514
rect 120252 247792 120572 248112
rect 129081 247816 129353 248088
rect 454929 246242 455201 246514
rect 120252 243792 120572 244112
rect 129081 243816 129353 244088
rect 454929 243242 455201 243514
rect 454929 240242 455201 240514
rect 120252 239792 120572 240112
rect 129081 239816 129353 240088
rect 454929 237242 455201 237514
rect 120252 235792 120572 236112
rect 129081 235816 129353 236088
rect 454929 234242 455201 234514
rect 120252 231792 120572 232112
rect 129081 231816 129353 232088
rect 454929 231242 455201 231514
rect 454929 228242 455201 228514
rect 120252 227792 120572 228112
rect 129081 227816 129353 228088
rect 454929 225242 455201 225514
rect 120252 223792 120572 224112
rect 129081 223816 129353 224088
rect 454929 222242 455201 222514
rect 120252 219792 120572 220112
rect 129081 219816 129353 220088
rect 454929 219242 455201 219514
rect 454929 216242 455201 216514
rect 120252 215792 120572 216112
rect 129081 215816 129353 216088
rect 454929 213242 455201 213514
rect 120252 211792 120572 212112
rect 129081 211816 129353 212088
rect 454929 210242 455201 210514
rect 120252 207792 120572 208112
rect 129081 207816 129353 208088
rect 454929 207242 455201 207514
rect 454929 204242 455201 204514
rect 120252 203792 120572 204112
rect 129081 203816 129353 204088
rect 454929 201242 455201 201514
rect 120252 199792 120572 200112
rect 129081 199816 129353 200088
rect 454929 198242 455201 198514
rect 120252 195792 120572 196112
rect 129081 195816 129353 196088
rect 454929 195242 455201 195514
rect 454929 192242 455201 192514
rect 120252 191792 120572 192112
rect 129081 191816 129353 192088
rect 454929 189242 455201 189514
rect 120252 187792 120572 188112
rect 129081 187816 129353 188088
rect 454929 186242 455201 186514
rect 120252 183792 120572 184112
rect 129081 183816 129353 184088
rect 454929 183242 455201 183514
rect 454929 180242 455201 180514
rect 120252 179792 120572 180112
rect 129081 179816 129353 180088
rect 454929 177242 455201 177514
rect 120252 175792 120572 176112
rect 129081 175816 129353 176088
rect 454929 174242 455201 174514
rect 120252 171792 120572 172112
rect 129081 171816 129353 172088
rect 454929 171242 455201 171514
rect 454929 168242 455201 168514
rect 120252 167792 120572 168112
rect 129081 167816 129353 168088
rect 454929 165242 455201 165514
rect 120252 163792 120572 164112
rect 129081 163816 129353 164088
rect 454929 162242 455201 162514
rect 120252 159792 120572 160112
rect 129081 159816 129353 160088
rect 454929 159242 455201 159514
rect 454929 156242 455201 156514
rect 120252 155792 120572 156112
rect 129081 155816 129353 156088
rect 454929 153242 455201 153514
rect 120252 151792 120572 152112
rect 129081 151816 129353 152088
rect 454929 150242 455201 150514
rect 120252 147792 120572 148112
rect 129081 147816 129353 148088
rect 536033 639783 540833 644609
rect 536767 629783 541567 634609
rect 504068 554230 508868 559030
rect 509895 556624 510532 557261
rect 528746 554254 533498 559006
rect 506840 469146 511640 473946
rect 533220 469170 537972 473922
rect 507140 453220 511892 457972
rect 534522 453196 539322 457996
rect 515386 438543 515706 438544
rect 515386 438213 515705 438543
rect 515705 438213 515706 438543
rect 515386 438212 515706 438213
rect 515386 435543 515706 435544
rect 515386 435213 515705 435543
rect 515705 435213 515706 435543
rect 515386 435212 515706 435213
rect 515386 432543 515706 432544
rect 515386 432213 515705 432543
rect 515705 432213 515706 432543
rect 515386 432212 515706 432213
rect 515386 429543 515706 429544
rect 515386 429213 515705 429543
rect 515705 429213 515706 429543
rect 515386 429212 515706 429213
rect 515386 426543 515706 426544
rect 515386 426213 515705 426543
rect 515705 426213 515706 426543
rect 515386 426212 515706 426213
rect 515386 423543 515706 423544
rect 515386 423213 515705 423543
rect 515705 423213 515706 423543
rect 515386 423212 515706 423213
rect 515386 420543 515706 420544
rect 515386 420213 515705 420543
rect 515705 420213 515706 420543
rect 515386 420212 515706 420213
rect 515386 417543 515706 417544
rect 515386 417213 515705 417543
rect 515705 417213 515706 417543
rect 515386 417212 515706 417213
rect 515386 414543 515706 414544
rect 515386 414213 515705 414543
rect 515705 414213 515706 414543
rect 515386 414212 515706 414213
rect 515386 411543 515706 411544
rect 515386 411213 515705 411543
rect 515705 411213 515706 411543
rect 515386 411212 515706 411213
rect 515386 408543 515706 408544
rect 515386 408213 515705 408543
rect 515705 408213 515706 408543
rect 515386 408212 515706 408213
rect 515386 405543 515706 405544
rect 515386 405213 515705 405543
rect 515705 405213 515706 405543
rect 515386 405212 515706 405213
rect 515386 402543 515706 402544
rect 515386 402213 515705 402543
rect 515705 402213 515706 402543
rect 515386 402212 515706 402213
rect 515386 399543 515706 399544
rect 515386 399213 515705 399543
rect 515705 399213 515706 399543
rect 515386 399212 515706 399213
rect 515386 396543 515706 396544
rect 515386 396213 515705 396543
rect 515705 396213 515706 396543
rect 515386 396212 515706 396213
rect 515386 393543 515706 393544
rect 515386 393213 515705 393543
rect 515705 393213 515706 393543
rect 515386 393212 515706 393213
rect 515386 390543 515706 390544
rect 515386 390213 515705 390543
rect 515705 390213 515706 390543
rect 515386 390212 515706 390213
rect 515386 387543 515706 387544
rect 515386 387213 515705 387543
rect 515705 387213 515706 387543
rect 515386 387212 515706 387213
rect 515386 384543 515706 384544
rect 515386 384213 515705 384543
rect 515705 384213 515706 384543
rect 515386 384212 515706 384213
rect 515386 381543 515706 381544
rect 515386 381213 515705 381543
rect 515705 381213 515706 381543
rect 515386 381212 515706 381213
rect 515386 378543 515706 378544
rect 515386 378213 515705 378543
rect 515705 378213 515706 378543
rect 515386 378212 515706 378213
rect 515386 375543 515706 375544
rect 515386 375213 515705 375543
rect 515705 375213 515706 375543
rect 515386 375212 515706 375213
rect 515386 372543 515706 372544
rect 515386 372213 515705 372543
rect 515705 372213 515706 372543
rect 515386 372212 515706 372213
rect 515386 369543 515706 369544
rect 515386 369213 515705 369543
rect 515705 369213 515706 369543
rect 515386 369212 515706 369213
rect 515386 366543 515706 366544
rect 515386 366213 515705 366543
rect 515705 366213 515706 366543
rect 515386 366212 515706 366213
rect 515386 363543 515706 363544
rect 515386 363213 515705 363543
rect 515705 363213 515706 363543
rect 515386 363212 515706 363213
rect 515386 360543 515706 360544
rect 515386 360213 515705 360543
rect 515705 360213 515706 360543
rect 515386 360212 515706 360213
rect 515386 357543 515706 357544
rect 515386 357213 515705 357543
rect 515705 357213 515706 357543
rect 515386 357212 515706 357213
rect 515386 354543 515706 354544
rect 515386 354213 515705 354543
rect 515705 354213 515706 354543
rect 515386 354212 515706 354213
rect 515386 351543 515706 351544
rect 515386 351213 515705 351543
rect 515705 351213 515706 351543
rect 515386 351212 515706 351213
rect 515386 348543 515706 348544
rect 515386 348213 515705 348543
rect 515705 348213 515706 348543
rect 515386 348212 515706 348213
rect 515386 345543 515706 345544
rect 515386 345213 515705 345543
rect 515705 345213 515706 345543
rect 515386 345212 515706 345213
rect 515386 342543 515706 342544
rect 515386 342213 515705 342543
rect 515705 342213 515706 342543
rect 515386 342212 515706 342213
rect 515386 339543 515706 339544
rect 515386 339213 515705 339543
rect 515705 339213 515706 339543
rect 515386 339212 515706 339213
rect 515386 336543 515706 336544
rect 515386 336213 515705 336543
rect 515705 336213 515706 336543
rect 515386 336212 515706 336213
rect 515386 333543 515706 333544
rect 515386 333213 515705 333543
rect 515705 333213 515706 333543
rect 515386 333212 515706 333213
rect 515386 330543 515706 330544
rect 515386 330213 515705 330543
rect 515705 330213 515706 330543
rect 515386 330212 515706 330213
rect 515386 327543 515706 327544
rect 515386 327213 515705 327543
rect 515705 327213 515706 327543
rect 515386 327212 515706 327213
rect 515386 324543 515706 324544
rect 515386 324213 515705 324543
rect 515705 324213 515706 324543
rect 515386 324212 515706 324213
rect 515386 321543 515706 321544
rect 515386 321213 515705 321543
rect 515705 321213 515706 321543
rect 515386 321212 515706 321213
rect 515386 318543 515706 318544
rect 515386 318213 515705 318543
rect 515705 318213 515706 318543
rect 515386 318212 515706 318213
rect 515386 315543 515706 315544
rect 515386 315213 515705 315543
rect 515705 315213 515706 315543
rect 515386 315212 515706 315213
rect 515386 312543 515706 312544
rect 515386 312213 515705 312543
rect 515705 312213 515706 312543
rect 515386 312212 515706 312213
rect 515386 309543 515706 309544
rect 515386 309213 515705 309543
rect 515705 309213 515706 309543
rect 515386 309212 515706 309213
rect 515386 306543 515706 306544
rect 515386 306213 515705 306543
rect 515705 306213 515706 306543
rect 515386 306212 515706 306213
rect 515386 303543 515706 303544
rect 515386 303213 515705 303543
rect 515705 303213 515706 303543
rect 515386 303212 515706 303213
rect 515386 300543 515706 300544
rect 515386 300213 515705 300543
rect 515705 300213 515706 300543
rect 515386 300212 515706 300213
rect 515386 297543 515706 297544
rect 515386 297213 515705 297543
rect 515705 297213 515706 297543
rect 515386 297212 515706 297213
rect 515386 294543 515706 294544
rect 515386 294213 515705 294543
rect 515705 294213 515706 294543
rect 515386 294212 515706 294213
rect 515386 291543 515706 291544
rect 515386 291213 515705 291543
rect 515705 291213 515706 291543
rect 515386 291212 515706 291213
rect 515386 288543 515706 288544
rect 515386 288213 515705 288543
rect 515705 288213 515706 288543
rect 515386 288212 515706 288213
rect 515386 285543 515706 285544
rect 515386 285213 515705 285543
rect 515705 285213 515706 285543
rect 515386 285212 515706 285213
rect 515386 282543 515706 282544
rect 515386 282213 515705 282543
rect 515705 282213 515706 282543
rect 515386 282212 515706 282213
rect 515386 279543 515706 279544
rect 515386 279213 515705 279543
rect 515705 279213 515706 279543
rect 515386 279212 515706 279213
rect 515386 276543 515706 276544
rect 515386 276213 515705 276543
rect 515705 276213 515706 276543
rect 515386 276212 515706 276213
rect 515386 273543 515706 273544
rect 515386 273213 515705 273543
rect 515705 273213 515706 273543
rect 515386 273212 515706 273213
rect 515386 270543 515706 270544
rect 515386 270213 515705 270543
rect 515705 270213 515706 270543
rect 515386 270212 515706 270213
rect 515386 267543 515706 267544
rect 515386 267213 515705 267543
rect 515705 267213 515706 267543
rect 515386 267212 515706 267213
rect 515386 264543 515706 264544
rect 515386 264213 515705 264543
rect 515705 264213 515706 264543
rect 515386 264212 515706 264213
rect 515386 261543 515706 261544
rect 515386 261213 515705 261543
rect 515705 261213 515706 261543
rect 515386 261212 515706 261213
rect 515386 258543 515706 258544
rect 515386 258213 515705 258543
rect 515705 258213 515706 258543
rect 515386 258212 515706 258213
rect 515386 255543 515706 255544
rect 515386 255213 515705 255543
rect 515705 255213 515706 255543
rect 515386 255212 515706 255213
rect 515386 252543 515706 252544
rect 515386 252213 515705 252543
rect 515705 252213 515706 252543
rect 515386 252212 515706 252213
rect 515386 249543 515706 249544
rect 515386 249213 515705 249543
rect 515705 249213 515706 249543
rect 515386 249212 515706 249213
rect 515386 246543 515706 246544
rect 515386 246213 515705 246543
rect 515705 246213 515706 246543
rect 515386 246212 515706 246213
rect 515386 243543 515706 243544
rect 515386 243213 515705 243543
rect 515705 243213 515706 243543
rect 515386 243212 515706 243213
rect 515386 240543 515706 240544
rect 515386 240213 515705 240543
rect 515705 240213 515706 240543
rect 515386 240212 515706 240213
rect 515386 237543 515706 237544
rect 515386 237213 515705 237543
rect 515705 237213 515706 237543
rect 515386 237212 515706 237213
rect 515386 234543 515706 234544
rect 515386 234213 515705 234543
rect 515705 234213 515706 234543
rect 515386 234212 515706 234213
rect 515386 231543 515706 231544
rect 515386 231213 515705 231543
rect 515705 231213 515706 231543
rect 515386 231212 515706 231213
rect 515386 228543 515706 228544
rect 515386 228213 515705 228543
rect 515705 228213 515706 228543
rect 515386 228212 515706 228213
rect 515386 225543 515706 225544
rect 515386 225213 515705 225543
rect 515705 225213 515706 225543
rect 515386 225212 515706 225213
rect 515386 222543 515706 222544
rect 515386 222213 515705 222543
rect 515705 222213 515706 222543
rect 515386 222212 515706 222213
rect 515386 219543 515706 219544
rect 515386 219213 515705 219543
rect 515705 219213 515706 219543
rect 515386 219212 515706 219213
rect 515386 216543 515706 216544
rect 515386 216213 515705 216543
rect 515705 216213 515706 216543
rect 515386 216212 515706 216213
rect 515386 213543 515706 213544
rect 515386 213213 515705 213543
rect 515705 213213 515706 213543
rect 515386 213212 515706 213213
rect 515386 210543 515706 210544
rect 515386 210213 515705 210543
rect 515705 210213 515706 210543
rect 515386 210212 515706 210213
rect 515386 207543 515706 207544
rect 515386 207213 515705 207543
rect 515705 207213 515706 207543
rect 515386 207212 515706 207213
rect 515386 204543 515706 204544
rect 515386 204213 515705 204543
rect 515705 204213 515706 204543
rect 515386 204212 515706 204213
rect 515386 201543 515706 201544
rect 515386 201213 515705 201543
rect 515705 201213 515706 201543
rect 515386 201212 515706 201213
rect 515386 198543 515706 198544
rect 515386 198213 515705 198543
rect 515705 198213 515706 198543
rect 515386 198212 515706 198213
rect 515386 195543 515706 195544
rect 515386 195213 515705 195543
rect 515705 195213 515706 195543
rect 515386 195212 515706 195213
rect 515386 192543 515706 192544
rect 515386 192213 515705 192543
rect 515705 192213 515706 192543
rect 515386 192212 515706 192213
rect 554140 191768 578296 196966
rect 515386 189543 515706 189544
rect 515386 189213 515705 189543
rect 515705 189213 515706 189543
rect 515386 189212 515706 189213
rect 515386 186543 515706 186544
rect 515386 186213 515705 186543
rect 515705 186213 515706 186543
rect 515386 186212 515706 186213
rect 515386 183543 515706 183544
rect 515386 183213 515705 183543
rect 515705 183213 515706 183543
rect 515386 183212 515706 183213
rect 553050 181150 576862 186340
rect 515386 180543 515706 180544
rect 515386 180213 515705 180543
rect 515705 180213 515706 180543
rect 515386 180212 515706 180213
rect 515386 177543 515706 177544
rect 515386 177213 515705 177543
rect 515705 177213 515706 177543
rect 515386 177212 515706 177213
rect 515386 174543 515706 174544
rect 515386 174213 515705 174543
rect 515705 174213 515706 174543
rect 515386 174212 515706 174213
rect 515386 171543 515706 171544
rect 515386 171213 515705 171543
rect 515705 171213 515706 171543
rect 515386 171212 515706 171213
rect 515386 168543 515706 168544
rect 515386 168213 515705 168543
rect 515705 168213 515706 168543
rect 515386 168212 515706 168213
rect 515386 165543 515706 165544
rect 515386 165213 515705 165543
rect 515705 165213 515706 165543
rect 515386 165212 515706 165213
rect 515386 162543 515706 162544
rect 515386 162213 515705 162543
rect 515705 162213 515706 162543
rect 515386 162212 515706 162213
rect 515386 159543 515706 159544
rect 515386 159213 515705 159543
rect 515705 159213 515706 159543
rect 515386 159212 515706 159213
rect 553300 159434 558052 164186
rect 515386 156543 515706 156544
rect 515386 156213 515705 156543
rect 515705 156213 515706 156543
rect 515386 156212 515706 156213
rect 515386 153543 515706 153544
rect 515386 153213 515705 153543
rect 515705 153213 515706 153543
rect 515386 153212 515706 153213
rect 515386 150543 515706 150544
rect 515386 150213 515705 150543
rect 515705 150213 515706 150543
rect 515386 150212 515706 150213
rect 120252 143792 120572 144112
rect 129081 143816 129353 144088
rect 120252 139792 120572 140112
rect 129081 139816 129353 140088
rect 495525 139876 496891 141242
rect 507515 139852 510119 141266
rect 453419 134348 453691 134620
rect 557323 126465 558008 127150
rect 150320 114800 150592 115072
rect 153320 114800 153592 115072
rect 156320 114800 156592 115072
rect 159320 114800 159592 115072
rect 162320 114800 162592 115072
rect 165320 114800 165592 115072
rect 168320 114800 168592 115072
rect 171320 114800 171592 115072
rect 174320 114800 174592 115072
rect 177320 114800 177592 115072
rect 180320 114800 180592 115072
rect 183320 114800 183592 115072
rect 186320 114800 186592 115072
rect 189320 114800 189592 115072
rect 192320 114800 192592 115072
rect 195320 114800 195592 115072
rect 198320 114800 198592 115072
rect 201320 114800 201592 115072
rect 204320 114800 204592 115072
rect 207320 114800 207592 115072
rect 210320 114800 210592 115072
rect 213320 114800 213592 115072
rect 216320 114800 216592 115072
rect 219320 114800 219592 115072
rect 222320 114800 222592 115072
rect 225320 114800 225592 115072
rect 228320 114800 228592 115072
rect 231320 114800 231592 115072
rect 234320 114800 234592 115072
rect 237320 114800 237592 115072
rect 240320 114800 240592 115072
rect 243320 114800 243592 115072
rect 246320 114800 246592 115072
rect 249320 114800 249592 115072
rect 252320 114800 252592 115072
rect 255320 114800 255592 115072
rect 258320 114800 258592 115072
rect 261320 114800 261592 115072
rect 264320 114800 264592 115072
rect 267320 114800 267592 115072
rect 270320 114800 270592 115072
rect 273320 114800 273592 115072
rect 276320 114800 276592 115072
rect 279320 114800 279592 115072
rect 282320 114800 282592 115072
rect 285320 114800 285592 115072
rect 288320 114800 288592 115072
rect 291320 114800 291592 115072
rect 294320 114800 294592 115072
rect 297320 114800 297592 115072
rect 300320 114800 300592 115072
rect 303320 114800 303592 115072
rect 306320 114800 306592 115072
rect 309320 114800 309592 115072
rect 312320 114800 312592 115072
rect 315320 114800 315592 115072
rect 318320 114800 318592 115072
rect 321320 114800 321592 115072
rect 324320 114800 324592 115072
rect 327320 114800 327592 115072
rect 330320 114800 330592 115072
rect 333320 114800 333592 115072
rect 336320 114800 336592 115072
rect 339320 114800 339592 115072
rect 342320 114800 342592 115072
rect 345320 114800 345592 115072
rect 348320 114800 348592 115072
rect 351320 114800 351592 115072
rect 354320 114800 354592 115072
rect 357320 114800 357592 115072
rect 360320 114800 360592 115072
rect 363320 114800 363592 115072
rect 366320 114800 366592 115072
rect 369320 114800 369592 115072
rect 372320 114800 372592 115072
rect 375320 114800 375592 115072
rect 378320 114800 378592 115072
rect 381320 114800 381592 115072
rect 384320 114800 384592 115072
rect 387320 114800 387592 115072
rect 390320 114800 390592 115072
rect 393320 114800 393592 115072
rect 396320 114800 396592 115072
rect 399320 114800 399592 115072
rect 402320 114800 402592 115072
rect 405320 114800 405592 115072
rect 408320 114800 408592 115072
rect 411320 114800 411592 115072
rect 414320 114800 414592 115072
rect 420320 114800 420592 115072
rect 423320 114800 423592 115072
rect 426320 114800 426592 115072
rect 429320 114800 429592 115072
rect 432320 114800 432592 115072
rect 435320 114800 435592 115072
rect 438320 114800 438592 115072
rect 441320 114800 441592 115072
rect 444320 114800 444592 115072
rect 96540 90342 101340 95142
rect 553300 90366 558052 95118
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 229160 699708 231660 702300
rect 229160 697552 229597 699708
rect 231180 697552 231660 699708
rect 229160 697490 231660 697552
rect 329590 701834 334230 702300
rect 329590 697442 329614 701834
rect 334006 700360 334230 701834
rect 334006 697442 334030 700360
rect 329590 697418 334030 697442
rect 518241 644584 520957 646724
rect 534064 644609 543338 645740
rect 534064 644584 536033 644609
rect 518241 639784 536033 644584
rect 209568 634844 210568 635244
rect 208168 634444 210568 634844
rect 207168 634244 210568 634444
rect 206168 633844 210568 634244
rect 205168 633444 210568 633844
rect 518241 634584 520957 639784
rect 534064 639783 536033 639784
rect 540833 639783 543338 644609
rect 534064 639002 543338 639783
rect 534308 634609 543582 635078
rect 534308 634584 536767 634609
rect 203968 633244 210168 633444
rect 202968 632844 209168 633244
rect 201568 632444 208168 632844
rect 200168 632244 207168 632444
rect 199168 631844 206168 632244
rect 197968 631444 204968 631844
rect 196568 631244 203968 631444
rect 195168 630844 202568 631244
rect 193968 630444 201568 630844
rect 90568 630244 91568 630444
rect 192568 630244 200168 630444
rect 90568 629844 92968 630244
rect 191168 629844 199168 630244
rect 90568 629444 94168 629844
rect 189568 629444 197968 629844
rect 518241 629784 536767 634584
rect 90568 629244 95568 629444
rect 188168 629244 196568 629444
rect 91568 628844 96968 629244
rect 186568 628844 195168 629244
rect 92568 628444 98168 628844
rect 184968 628444 193968 628844
rect 93968 628244 99968 628444
rect 183568 628244 192568 628444
rect 94968 627844 101568 628244
rect 181968 627844 190968 628244
rect 96168 627444 103168 627844
rect 163968 627444 164568 627844
rect 179968 627444 189568 627844
rect 97568 627244 105168 627444
rect 162568 627244 165968 627444
rect 178168 627244 187968 627444
rect 98968 626844 107168 627244
rect 161968 626844 166568 627244
rect 176168 626844 186568 627244
rect 100568 626444 109568 626844
rect 161568 626444 166968 626844
rect 174168 626444 184968 626844
rect 101968 626244 111968 626444
rect 160968 626244 167168 626444
rect 172168 626244 183168 626444
rect 103968 625844 114568 626244
rect 160168 625844 167568 626244
rect 169568 625844 181568 626244
rect 105568 625444 117568 625844
rect 143968 625444 147168 625844
rect 159968 625444 179568 625844
rect 107568 625244 120968 625444
rect 143168 625244 147968 625444
rect 159568 625244 177968 625444
rect 109968 624844 124968 625244
rect 142568 624844 148968 625244
rect 159568 624844 175968 625244
rect 111968 624444 129968 624844
rect 142168 624444 149568 624844
rect 155968 624444 173568 624844
rect 114568 624244 137568 624444
rect 141968 624244 171568 624444
rect 117168 623844 168968 624244
rect 120568 623444 167168 623844
rect 123968 623244 166968 623444
rect 128568 622844 165968 623244
rect 134568 622444 153168 622844
rect 158168 622444 164168 622844
rect 141168 622244 151168 622444
rect 141568 621844 151168 622244
rect 141968 621444 151168 621844
rect 158168 622244 163568 622444
rect 158168 621444 163168 622244
rect 142568 621244 151568 621444
rect 145568 620844 151568 621244
rect 145968 620444 151568 620844
rect 146168 619244 151568 620444
rect 157968 621244 163168 621444
rect 157968 619444 162968 621244
rect 146168 616844 151968 619244
rect 145968 615844 151968 616844
rect 145568 614444 151968 615844
rect 145168 613244 151968 614444
rect 144968 612244 151968 613244
rect 144568 611244 151968 612244
rect 144168 609844 151968 611244
rect 143968 609244 151968 609844
rect 157968 617844 163168 619444
rect 157968 616844 163568 617844
rect 157968 615444 163968 616844
rect 157968 614244 164168 615444
rect 157968 613244 164568 614244
rect 157968 612244 164968 613244
rect 157968 610844 165168 612244
rect 157968 609444 165568 610844
rect 143968 608444 151568 609244
rect 143568 606444 151568 608444
rect 157968 607444 165968 609444
rect 157968 606844 166168 607444
rect 143168 603244 151568 606444
rect 158168 604444 166168 606844
rect 143168 597844 151168 603244
rect 158168 602244 166568 604444
rect 158568 599244 166568 602244
rect 158168 598844 166568 599244
rect 143168 595844 151568 597844
rect 158168 597244 166168 598844
rect 157968 596844 166168 597244
rect 156968 596444 166168 596844
rect 155968 596244 166168 596444
rect 303840 596630 304276 596670
rect 303840 596606 303918 596630
rect 304190 596606 304276 596630
rect 303840 596286 303894 596606
rect 304214 596286 340720 596606
rect 303840 596250 304276 596286
rect 155568 595844 166168 596244
rect 126168 595444 128968 595844
rect 123968 595244 130168 595444
rect 122968 594844 131168 595244
rect 121568 594444 131968 594844
rect 143168 594444 151968 595844
rect 154968 595444 166168 595844
rect 154568 595244 166168 595444
rect 154168 594844 166168 595244
rect 153968 594444 166168 594844
rect 120968 594244 132568 594444
rect 143568 594244 151968 594444
rect 120168 593844 132968 594244
rect 119568 593444 133168 593844
rect 118968 593244 133968 593444
rect 143568 593244 152168 594244
rect 153568 593844 166168 594444
rect 304812 594242 307352 594562
rect 153168 593444 166168 593844
rect 118168 592844 134168 593244
rect 117968 592444 134568 592844
rect 143568 592444 152568 593244
rect 153168 592844 165968 593444
rect 152968 592444 165968 592844
rect 303894 592806 304214 592830
rect 303894 592534 303918 592806
rect 304190 592534 304214 592806
rect 303894 592510 304214 592534
rect 117568 592244 134968 592444
rect 143568 592244 165968 592444
rect 117168 591844 124968 592244
rect 129168 591844 135168 592244
rect 116968 591444 123168 591844
rect 130168 591444 135568 591844
rect 143968 591444 165968 592244
rect 292314 591878 292634 591902
rect 292314 591606 292338 591878
rect 292610 591606 292634 591878
rect 292314 591582 292634 591606
rect 116568 591244 122168 591444
rect 130968 591244 135968 591444
rect 116168 590844 121568 591244
rect 131568 590844 136168 591244
rect 116168 590444 120968 590844
rect 131968 590444 136568 590844
rect 143968 590444 165568 591444
rect 337754 590460 340470 596286
rect 115968 590244 120568 590444
rect 132168 590244 136968 590444
rect 115568 589844 120168 590244
rect 132568 589844 137168 590244
rect 115568 589444 119568 589844
rect 132968 589444 137168 589844
rect 144168 589444 165968 590444
rect 337754 590140 338088 590460
rect 338408 590140 340470 590460
rect 115168 589244 119168 589444
rect 133168 589244 137568 589444
rect 115168 588844 118968 589244
rect 133568 588844 137968 589244
rect 144568 588844 166168 589444
rect 114968 588444 118568 588844
rect 133968 588444 138168 588844
rect 144568 588444 166568 588844
rect 337754 588588 340470 590140
rect 518241 588588 520957 629784
rect 534308 629783 536767 629784
rect 541567 629783 543582 634609
rect 534308 628340 543582 629783
rect 114968 588244 118168 588444
rect 134168 588244 138168 588444
rect 144968 588244 166968 588444
rect 114968 587844 117968 588244
rect 134168 587844 138568 588244
rect 114568 587444 117968 587844
rect 134568 587444 138568 587844
rect 145168 587844 167168 588244
rect 145168 587444 167568 587844
rect 114568 587244 117568 587444
rect 134568 587244 138968 587444
rect 145568 587244 167568 587444
rect 114568 586844 117168 587244
rect 114168 586444 117168 586844
rect 134968 586844 138968 587244
rect 145968 586844 167968 587244
rect 114168 586244 116968 586444
rect 134968 586244 139168 586844
rect 146168 586444 167968 586844
rect 146568 586244 167968 586444
rect 337754 586460 520957 588588
rect 114168 585244 116568 586244
rect 135168 585244 139568 586244
rect 146568 585444 167568 586244
rect 337754 586140 338088 586460
rect 338408 586140 520957 586460
rect 337754 585872 520957 586140
rect 146568 585244 167168 585444
rect 114168 584244 116168 585244
rect 114168 583444 115968 584244
rect 135568 583444 139968 585244
rect 146168 584844 167168 585244
rect 146168 584444 166968 584844
rect 146168 584244 166568 584444
rect 146168 583844 162168 584244
rect 162968 583844 165968 584244
rect 114568 582844 115568 583444
rect 135968 579444 139968 583444
rect 145968 583444 162168 583844
rect 145968 582844 162568 583444
rect 145968 581844 162968 582844
rect 145568 580444 163168 581844
rect 145168 579844 163168 580444
rect 135568 578244 139568 579444
rect 145168 578844 163568 579844
rect 144968 578444 163568 578844
rect 135568 577844 139168 578244
rect 135168 576844 139168 577844
rect 144968 577444 163968 578444
rect 134968 575844 138968 576844
rect 144568 575844 163968 577444
rect 134968 575444 138568 575844
rect 134568 574844 138568 575444
rect 144168 575244 163968 575844
rect 134568 573844 138168 574844
rect 144168 574244 163568 575244
rect 134568 573244 137968 573844
rect 134168 572244 137968 573244
rect 144168 573444 163168 574244
rect 144168 572844 162968 573444
rect 134168 570244 137568 572244
rect 143968 571844 162568 572844
rect 143968 571244 162168 571844
rect 143968 570844 161968 571244
rect 144168 570444 161968 570844
rect 134568 569244 137568 570244
rect 143968 570244 161568 570444
rect 143968 569844 161168 570244
rect 143968 569444 160968 569844
rect 134568 568244 137968 569244
rect 134968 567844 137968 568244
rect 143968 568844 160568 569444
rect 143968 568444 160168 568844
rect 143968 567844 159968 568444
rect 134968 567244 138168 567844
rect 143568 567244 159568 567844
rect 135168 566844 138568 567244
rect 135168 566244 138968 566844
rect 143568 566444 159168 567244
rect 135568 565844 139168 566244
rect 135568 565444 139568 565844
rect 135968 565244 140168 565444
rect 143168 565244 158968 566444
rect 136168 564844 140568 565244
rect 142968 564844 158968 565244
rect 136168 564444 141168 564844
rect 142968 564444 159568 564844
rect 136568 564244 141968 564444
rect 142968 564244 159968 564444
rect 136968 563844 160568 564244
rect 137168 563444 160968 563844
rect 137968 563244 161568 563444
rect 138168 562844 162168 563244
rect 138568 562444 162968 562844
rect 139168 562244 163168 562444
rect 139568 561844 163968 562244
rect 139968 561444 164568 561844
rect 140568 561244 164968 561444
rect 140968 560844 165568 561244
rect 140568 560444 166168 560844
rect 140568 560244 166968 560444
rect 140168 559844 167168 560244
rect 140168 559444 167968 559844
rect 139968 559244 168568 559444
rect 139968 558844 168968 559244
rect 290594 559030 290914 582110
rect 304924 559030 305244 580778
rect 504044 559030 508892 559054
rect 139568 558444 169568 558844
rect 139568 558244 169968 558444
rect 139168 557844 170568 558244
rect 139168 557444 170968 557844
rect 138968 557244 171168 557444
rect 283960 557285 504068 559030
rect 138968 556844 171568 557244
rect 138568 556244 149168 556844
rect 149568 556444 171968 556844
rect 283960 556600 308982 557285
rect 309667 556600 504068 557285
rect 150568 556244 172168 556444
rect 138168 555844 148968 556244
rect 151568 555844 172568 556244
rect 137968 555444 148568 555844
rect 152568 555444 172568 555844
rect 137568 555244 148568 555444
rect 154168 555244 172968 555444
rect 137168 554844 148168 555244
rect 155968 554844 172968 555244
rect 136568 554444 148168 554844
rect 157968 554444 173168 554844
rect 130168 554244 147968 554444
rect 159968 554244 173168 554444
rect 126568 553844 147568 554244
rect 161568 553844 173168 554244
rect 283960 554230 504068 556600
rect 508868 557285 508892 559030
rect 508868 557261 510556 557285
rect 508868 556624 509895 557261
rect 510532 556624 510556 557261
rect 508868 556600 510556 556624
rect 508868 554230 508892 556600
rect 504044 554206 508892 554230
rect 124968 553444 147568 553844
rect 162968 553444 173568 553844
rect 123968 553244 147168 553444
rect 163968 553244 173568 553444
rect 123168 552844 147168 553244
rect 164968 552844 173568 553244
rect 122968 552444 146968 552844
rect 165568 552444 173568 552844
rect 122568 551844 146568 552444
rect 165968 552244 173568 552444
rect 165968 551844 173968 552244
rect 122568 551444 146168 551844
rect 122168 551244 145968 551444
rect 122168 550444 145568 551244
rect 122168 550244 145168 550444
rect 166168 550244 173968 551844
rect 122168 549844 144968 550244
rect 122168 549444 144568 549844
rect 166568 549444 173968 550244
rect 122168 549244 144168 549444
rect 122168 548844 143968 549244
rect 122168 548444 143168 548844
rect 122168 548244 142568 548444
rect 166568 548244 174168 549444
rect 122168 547844 142168 548244
rect 122568 547444 141568 547844
rect 122568 547244 139968 547444
rect 122568 545844 128568 547244
rect 130568 546844 137968 547244
rect 132168 546444 134168 546844
rect 166968 546444 174168 548244
rect 122968 544844 128568 545844
rect 122968 544444 128968 544844
rect 167168 544444 174168 546444
rect 123168 544244 128968 544444
rect 123168 543444 129168 544244
rect 123568 543244 129568 543444
rect 123568 542844 129968 543244
rect 167568 542844 174168 544444
rect 179968 544244 183968 544444
rect 178168 543844 184168 544244
rect 176968 543444 184568 543844
rect 175568 543244 184568 543444
rect 174968 542844 184168 543244
rect 123968 542444 130168 542844
rect 167568 542444 184168 542844
rect 123968 542244 130568 542444
rect 167568 542244 183968 542444
rect 124168 541844 130968 542244
rect 167968 541844 183568 542244
rect 124168 541444 131568 541844
rect 167968 541444 183168 541844
rect 124968 541244 131968 541444
rect 167968 541244 182568 541444
rect 125168 540844 132168 541244
rect 167968 540844 181968 541244
rect 126168 540444 132568 540844
rect 167968 540444 180968 540844
rect 127568 540244 132968 540444
rect 168168 540244 180168 540444
rect 128568 539844 133168 540244
rect 168168 539844 179168 540244
rect 128968 539444 133568 539844
rect 168168 539444 178168 539844
rect 129568 539244 133968 539444
rect 168168 539244 177168 539444
rect 129968 538844 133968 539244
rect 168568 538844 176168 539244
rect 130968 538444 134168 538844
rect 168568 538444 175168 538844
rect 131968 538244 134168 538444
rect 168968 538244 174168 538444
rect 132968 537844 134168 538244
rect 169168 537844 173168 538244
rect 169968 537444 171968 537844
rect 518241 489282 520957 585872
rect 528722 559006 552198 559030
rect 528722 554254 528746 559006
rect 533498 554254 558076 559006
rect 528722 554230 558076 554254
rect 284208 486566 520957 489282
rect 284208 473346 286924 486566
rect 506816 473946 511664 473970
rect 296978 473922 506840 473946
rect 288539 473352 289117 473376
rect 288539 473346 288563 473352
rect 284208 472816 288563 473346
rect 284208 471752 286924 472816
rect 288539 472810 288563 472816
rect 289093 472810 289117 473352
rect 288539 472786 289117 472810
rect 296978 471951 334724 473922
rect 296978 471569 297407 471951
rect 297777 471569 334724 471951
rect 290860 469718 291548 469742
rect 290860 469066 290884 469718
rect 291524 469712 291548 469718
rect 296978 469712 334724 471569
rect 291524 469170 334724 469712
rect 339476 469170 506840 473922
rect 291524 469146 506840 469170
rect 511640 469146 511664 473946
rect 291524 469072 302376 469146
rect 506816 469122 511664 469146
rect 291524 469066 291548 469072
rect 290860 469042 291548 469066
rect 96586 457972 511916 457996
rect 96586 454878 507140 457972
rect 96586 454558 162784 454878
rect 163104 454558 165784 454878
rect 166104 454558 168784 454878
rect 169104 454558 171784 454878
rect 172104 454558 174784 454878
rect 175104 454558 177784 454878
rect 178104 454558 180784 454878
rect 181104 454558 183784 454878
rect 184104 454558 186784 454878
rect 187104 454558 189784 454878
rect 190104 454558 192784 454878
rect 193104 454558 195784 454878
rect 196104 454558 198784 454878
rect 199104 454558 201784 454878
rect 202104 454558 204784 454878
rect 205104 454558 207784 454878
rect 208104 454558 210784 454878
rect 211104 454558 213784 454878
rect 214104 454558 216784 454878
rect 217104 454558 219784 454878
rect 220104 454558 222784 454878
rect 223104 454558 225784 454878
rect 226104 454558 228784 454878
rect 229104 454558 231784 454878
rect 232104 454558 234784 454878
rect 235104 454558 237784 454878
rect 238104 454558 240784 454878
rect 241104 454558 243784 454878
rect 244104 454558 246784 454878
rect 247104 454558 249784 454878
rect 250104 454558 252784 454878
rect 253104 454558 255784 454878
rect 256104 454558 258784 454878
rect 259104 454558 261784 454878
rect 262104 454558 264784 454878
rect 265104 454558 267784 454878
rect 268104 454558 270784 454878
rect 271104 454558 273784 454878
rect 274104 454558 276784 454878
rect 277104 454558 279784 454878
rect 280104 454558 282784 454878
rect 283104 454558 285784 454878
rect 286104 454558 288784 454878
rect 289104 454558 291784 454878
rect 292104 454558 294784 454878
rect 295104 454558 297784 454878
rect 298104 454558 300784 454878
rect 301104 454558 303784 454878
rect 304104 454558 306784 454878
rect 307104 454558 309784 454878
rect 310104 454558 312784 454878
rect 313104 454558 315784 454878
rect 316104 454558 318784 454878
rect 319104 454558 321784 454878
rect 322104 454558 324784 454878
rect 325104 454558 327784 454878
rect 328104 454558 330784 454878
rect 331104 454558 333784 454878
rect 334104 454558 336784 454878
rect 337104 454558 339784 454878
rect 340104 454558 342784 454878
rect 343104 454558 345784 454878
rect 346104 454558 348784 454878
rect 349104 454558 351784 454878
rect 352104 454558 354784 454878
rect 355104 454558 357784 454878
rect 358104 454558 360784 454878
rect 361104 454558 363784 454878
rect 364104 454558 366784 454878
rect 367104 454558 369784 454878
rect 370104 454558 372784 454878
rect 373104 454558 375784 454878
rect 376104 454558 378784 454878
rect 379104 454558 381784 454878
rect 382104 454558 384784 454878
rect 385104 454558 387784 454878
rect 388104 454558 390784 454878
rect 391104 454558 393784 454878
rect 394104 454558 396784 454878
rect 397104 454558 399784 454878
rect 400104 454558 402784 454878
rect 403104 454558 405784 454878
rect 406104 454558 408784 454878
rect 409104 454558 411784 454878
rect 412104 454558 414784 454878
rect 415104 454558 417784 454878
rect 418104 454558 420784 454878
rect 421104 454558 423784 454878
rect 424104 454558 426784 454878
rect 427104 454558 429784 454878
rect 430104 454558 432784 454878
rect 433104 454558 435784 454878
rect 436104 454558 438784 454878
rect 439104 454558 441784 454878
rect 442104 454558 444784 454878
rect 445104 454558 447784 454878
rect 448104 454558 507140 454878
rect 96586 453220 507140 454558
rect 511892 453220 511916 457972
rect 96586 453196 511916 453220
rect 96586 95166 101386 453196
rect 518241 446868 520957 486566
rect 553276 473946 558076 554230
rect 533196 473922 558076 473946
rect 533196 469170 533220 473922
rect 537972 469170 558076 473922
rect 533196 469146 558076 469170
rect 534498 457996 539346 458020
rect 553276 457996 558076 469146
rect 534498 453196 534522 457996
rect 539322 453196 558076 457996
rect 534498 453172 539346 453196
rect 118982 444152 520957 446868
rect 118982 436112 121698 444152
rect 162784 438802 163104 438826
rect 162784 438530 162808 438802
rect 163080 438530 163104 438802
rect 162784 438506 163104 438530
rect 165784 438802 166104 438826
rect 165784 438530 165808 438802
rect 166080 438530 166104 438802
rect 165784 438506 166104 438530
rect 168784 438802 169104 438826
rect 168784 438530 168808 438802
rect 169080 438530 169104 438802
rect 168784 438506 169104 438530
rect 171784 438802 172104 438826
rect 171784 438530 171808 438802
rect 172080 438530 172104 438802
rect 171784 438506 172104 438530
rect 174784 438802 175104 438826
rect 174784 438530 174808 438802
rect 175080 438530 175104 438802
rect 174784 438506 175104 438530
rect 177784 438802 178104 438826
rect 177784 438530 177808 438802
rect 178080 438530 178104 438802
rect 177784 438506 178104 438530
rect 180784 438802 181104 438826
rect 180784 438530 180808 438802
rect 181080 438530 181104 438802
rect 180784 438506 181104 438530
rect 183784 438802 184104 438826
rect 183784 438530 183808 438802
rect 184080 438530 184104 438802
rect 183784 438506 184104 438530
rect 186784 438802 187104 438826
rect 186784 438530 186808 438802
rect 187080 438530 187104 438802
rect 186784 438506 187104 438530
rect 189784 438802 190104 438826
rect 189784 438530 189808 438802
rect 190080 438530 190104 438802
rect 189784 438506 190104 438530
rect 192784 438802 193104 438826
rect 192784 438530 192808 438802
rect 193080 438530 193104 438802
rect 192784 438506 193104 438530
rect 195784 438802 196104 438826
rect 195784 438530 195808 438802
rect 196080 438530 196104 438802
rect 195784 438506 196104 438530
rect 198784 438802 199104 438826
rect 198784 438530 198808 438802
rect 199080 438530 199104 438802
rect 198784 438506 199104 438530
rect 201784 438802 202104 438826
rect 201784 438530 201808 438802
rect 202080 438530 202104 438802
rect 201784 438506 202104 438530
rect 204784 438802 205104 438826
rect 204784 438530 204808 438802
rect 205080 438530 205104 438802
rect 204784 438506 205104 438530
rect 207784 438802 208104 438826
rect 207784 438530 207808 438802
rect 208080 438530 208104 438802
rect 207784 438506 208104 438530
rect 210784 438802 211104 438826
rect 210784 438530 210808 438802
rect 211080 438530 211104 438802
rect 210784 438506 211104 438530
rect 213784 438802 214104 438826
rect 213784 438530 213808 438802
rect 214080 438530 214104 438802
rect 213784 438506 214104 438530
rect 216784 438802 217104 438826
rect 216784 438530 216808 438802
rect 217080 438530 217104 438802
rect 216784 438506 217104 438530
rect 219784 438802 220104 438826
rect 219784 438530 219808 438802
rect 220080 438530 220104 438802
rect 219784 438506 220104 438530
rect 222784 438802 223104 438826
rect 222784 438530 222808 438802
rect 223080 438530 223104 438802
rect 222784 438506 223104 438530
rect 225784 438802 226104 438826
rect 225784 438530 225808 438802
rect 226080 438530 226104 438802
rect 225784 438506 226104 438530
rect 228784 438802 229104 438826
rect 228784 438530 228808 438802
rect 229080 438530 229104 438802
rect 228784 438506 229104 438530
rect 231784 438802 232104 438826
rect 231784 438530 231808 438802
rect 232080 438530 232104 438802
rect 231784 438506 232104 438530
rect 234784 438802 235104 438826
rect 234784 438530 234808 438802
rect 235080 438530 235104 438802
rect 234784 438506 235104 438530
rect 237784 438802 238104 438826
rect 237784 438530 237808 438802
rect 238080 438530 238104 438802
rect 237784 438506 238104 438530
rect 240784 438802 241104 438826
rect 240784 438530 240808 438802
rect 241080 438530 241104 438802
rect 240784 438506 241104 438530
rect 243784 438802 244104 438826
rect 243784 438530 243808 438802
rect 244080 438530 244104 438802
rect 243784 438506 244104 438530
rect 246784 438802 247104 438826
rect 246784 438530 246808 438802
rect 247080 438530 247104 438802
rect 246784 438506 247104 438530
rect 249784 438802 250104 438826
rect 249784 438530 249808 438802
rect 250080 438530 250104 438802
rect 249784 438506 250104 438530
rect 252784 438802 253104 438826
rect 252784 438530 252808 438802
rect 253080 438530 253104 438802
rect 252784 438506 253104 438530
rect 255784 438802 256104 438826
rect 255784 438530 255808 438802
rect 256080 438530 256104 438802
rect 255784 438506 256104 438530
rect 258784 438802 259104 438826
rect 258784 438530 258808 438802
rect 259080 438530 259104 438802
rect 258784 438506 259104 438530
rect 261784 438802 262104 438826
rect 261784 438530 261808 438802
rect 262080 438530 262104 438802
rect 261784 438506 262104 438530
rect 264784 438802 265104 438826
rect 264784 438530 264808 438802
rect 265080 438530 265104 438802
rect 264784 438506 265104 438530
rect 267784 438802 268104 438826
rect 267784 438530 267808 438802
rect 268080 438530 268104 438802
rect 267784 438506 268104 438530
rect 270784 438802 271104 438826
rect 270784 438530 270808 438802
rect 271080 438530 271104 438802
rect 270784 438506 271104 438530
rect 273784 438802 274104 438826
rect 273784 438530 273808 438802
rect 274080 438530 274104 438802
rect 273784 438506 274104 438530
rect 276784 438802 277104 438826
rect 276784 438530 276808 438802
rect 277080 438530 277104 438802
rect 276784 438506 277104 438530
rect 279784 438802 280104 438826
rect 279784 438530 279808 438802
rect 280080 438530 280104 438802
rect 279784 438506 280104 438530
rect 282784 438802 283104 438826
rect 282784 438530 282808 438802
rect 283080 438530 283104 438802
rect 282784 438506 283104 438530
rect 285784 438802 286104 438826
rect 285784 438530 285808 438802
rect 286080 438530 286104 438802
rect 285784 438506 286104 438530
rect 288784 438802 289104 438826
rect 288784 438530 288808 438802
rect 289080 438530 289104 438802
rect 288784 438506 289104 438530
rect 291784 438802 292104 438826
rect 291784 438530 291808 438802
rect 292080 438530 292104 438802
rect 291784 438506 292104 438530
rect 294784 438802 295104 438826
rect 294784 438530 294808 438802
rect 295080 438530 295104 438802
rect 294784 438506 295104 438530
rect 297784 438802 298104 438826
rect 297784 438530 297808 438802
rect 298080 438530 298104 438802
rect 297784 438506 298104 438530
rect 300784 438802 301104 438826
rect 300784 438530 300808 438802
rect 301080 438530 301104 438802
rect 300784 438506 301104 438530
rect 303784 438802 304104 438826
rect 303784 438530 303808 438802
rect 304080 438530 304104 438802
rect 303784 438506 304104 438530
rect 306784 438802 307104 438826
rect 306784 438530 306808 438802
rect 307080 438530 307104 438802
rect 306784 438506 307104 438530
rect 309784 438802 310104 438826
rect 309784 438530 309808 438802
rect 310080 438530 310104 438802
rect 309784 438506 310104 438530
rect 312784 438802 313104 438826
rect 312784 438530 312808 438802
rect 313080 438530 313104 438802
rect 312784 438506 313104 438530
rect 315784 438802 316104 438826
rect 315784 438530 315808 438802
rect 316080 438530 316104 438802
rect 315784 438506 316104 438530
rect 318784 438802 319104 438826
rect 318784 438530 318808 438802
rect 319080 438530 319104 438802
rect 318784 438506 319104 438530
rect 321784 438802 322104 438826
rect 321784 438530 321808 438802
rect 322080 438530 322104 438802
rect 321784 438506 322104 438530
rect 324784 438802 325104 438826
rect 324784 438530 324808 438802
rect 325080 438530 325104 438802
rect 324784 438506 325104 438530
rect 327784 438802 328104 438826
rect 327784 438530 327808 438802
rect 328080 438530 328104 438802
rect 327784 438506 328104 438530
rect 330784 438802 331104 438826
rect 330784 438530 330808 438802
rect 331080 438530 331104 438802
rect 330784 438506 331104 438530
rect 333784 438802 334104 438826
rect 333784 438530 333808 438802
rect 334080 438530 334104 438802
rect 333784 438506 334104 438530
rect 336784 438802 337104 438826
rect 336784 438530 336808 438802
rect 337080 438530 337104 438802
rect 336784 438506 337104 438530
rect 339784 438802 340104 438826
rect 339784 438530 339808 438802
rect 340080 438530 340104 438802
rect 339784 438506 340104 438530
rect 342784 438802 343104 438826
rect 342784 438530 342808 438802
rect 343080 438530 343104 438802
rect 342784 438506 343104 438530
rect 345784 438802 346104 438826
rect 345784 438530 345808 438802
rect 346080 438530 346104 438802
rect 345784 438506 346104 438530
rect 348784 438802 349104 438826
rect 348784 438530 348808 438802
rect 349080 438530 349104 438802
rect 348784 438506 349104 438530
rect 351784 438802 352104 438826
rect 351784 438530 351808 438802
rect 352080 438530 352104 438802
rect 351784 438506 352104 438530
rect 354784 438802 355104 438826
rect 354784 438530 354808 438802
rect 355080 438530 355104 438802
rect 354784 438506 355104 438530
rect 357784 438802 358104 438826
rect 357784 438530 357808 438802
rect 358080 438530 358104 438802
rect 357784 438506 358104 438530
rect 360784 438802 361104 438826
rect 360784 438530 360808 438802
rect 361080 438530 361104 438802
rect 360784 438506 361104 438530
rect 363784 438802 364104 438826
rect 363784 438530 363808 438802
rect 364080 438530 364104 438802
rect 363784 438506 364104 438530
rect 366784 438802 367104 438826
rect 366784 438530 366808 438802
rect 367080 438530 367104 438802
rect 366784 438506 367104 438530
rect 369784 438802 370104 438826
rect 369784 438530 369808 438802
rect 370080 438530 370104 438802
rect 369784 438506 370104 438530
rect 372784 438802 373104 438826
rect 372784 438530 372808 438802
rect 373080 438530 373104 438802
rect 372784 438506 373104 438530
rect 375784 438802 376104 438826
rect 375784 438530 375808 438802
rect 376080 438530 376104 438802
rect 375784 438506 376104 438530
rect 378784 438802 379104 438826
rect 378784 438530 378808 438802
rect 379080 438530 379104 438802
rect 378784 438506 379104 438530
rect 381784 438802 382104 438826
rect 381784 438530 381808 438802
rect 382080 438530 382104 438802
rect 381784 438506 382104 438530
rect 384784 438802 385104 438826
rect 384784 438530 384808 438802
rect 385080 438530 385104 438802
rect 384784 438506 385104 438530
rect 387784 438802 388104 438826
rect 387784 438530 387808 438802
rect 388080 438530 388104 438802
rect 387784 438506 388104 438530
rect 390784 438802 391104 438826
rect 390784 438530 390808 438802
rect 391080 438530 391104 438802
rect 390784 438506 391104 438530
rect 393784 438802 394104 438826
rect 393784 438530 393808 438802
rect 394080 438530 394104 438802
rect 393784 438506 394104 438530
rect 396784 438802 397104 438826
rect 396784 438530 396808 438802
rect 397080 438530 397104 438802
rect 396784 438506 397104 438530
rect 399784 438802 400104 438826
rect 399784 438530 399808 438802
rect 400080 438530 400104 438802
rect 399784 438506 400104 438530
rect 402784 438802 403104 438826
rect 402784 438530 402808 438802
rect 403080 438530 403104 438802
rect 402784 438506 403104 438530
rect 405784 438802 406104 438826
rect 405784 438530 405808 438802
rect 406080 438530 406104 438802
rect 405784 438506 406104 438530
rect 408784 438802 409104 438826
rect 408784 438530 408808 438802
rect 409080 438530 409104 438802
rect 408784 438506 409104 438530
rect 411784 438802 412104 438826
rect 411784 438530 411808 438802
rect 412080 438530 412104 438802
rect 411784 438506 412104 438530
rect 414784 438802 415104 438826
rect 414784 438530 414808 438802
rect 415080 438530 415104 438802
rect 414784 438506 415104 438530
rect 417784 438802 418104 438826
rect 417784 438530 417808 438802
rect 418080 438530 418104 438802
rect 417784 438506 418104 438530
rect 420784 438802 421104 438826
rect 420784 438530 420808 438802
rect 421080 438530 421104 438802
rect 420784 438506 421104 438530
rect 423784 438802 424104 438826
rect 423784 438530 423808 438802
rect 424080 438530 424104 438802
rect 423784 438506 424104 438530
rect 426784 438802 427104 438826
rect 426784 438530 426808 438802
rect 427080 438530 427104 438802
rect 426784 438506 427104 438530
rect 429784 438802 430104 438826
rect 429784 438530 429808 438802
rect 430080 438530 430104 438802
rect 429784 438506 430104 438530
rect 432784 438802 433104 438826
rect 432784 438530 432808 438802
rect 433080 438530 433104 438802
rect 432784 438506 433104 438530
rect 435784 438802 436104 438826
rect 435784 438530 435808 438802
rect 436080 438530 436104 438802
rect 435784 438506 436104 438530
rect 438784 438802 439104 438826
rect 438784 438530 438808 438802
rect 439080 438530 439104 438802
rect 438784 438506 439104 438530
rect 441784 438802 442104 438826
rect 441784 438530 441808 438802
rect 442080 438530 442104 438802
rect 441784 438506 442104 438530
rect 444784 438802 445104 438826
rect 444784 438530 444808 438802
rect 445080 438530 445104 438802
rect 444784 438506 445104 438530
rect 447784 438802 448104 438826
rect 447784 438530 447808 438802
rect 448080 438530 448104 438802
rect 515362 438544 515730 438568
rect 447784 438506 448104 438530
rect 454905 438514 455225 438538
rect 454905 438242 454929 438514
rect 455201 438242 455225 438514
rect 454905 438218 455225 438242
rect 515362 438212 515386 438544
rect 515706 438538 515730 438544
rect 518241 438538 520957 444152
rect 515706 438218 520957 438538
rect 515706 438212 515730 438218
rect 515362 438188 515730 438212
rect 149102 437210 149422 437234
rect 149102 436938 149126 437210
rect 149398 436938 149422 437210
rect 149102 436466 149422 436938
rect 149102 436194 149126 436466
rect 149398 436194 149422 436466
rect 118982 435792 120252 436112
rect 120572 435792 121698 436112
rect 129057 436088 129377 436112
rect 129057 435816 129081 436088
rect 129353 435816 129377 436088
rect 129057 435792 129377 435816
rect 118982 432112 121698 435792
rect 149102 434728 149422 436194
rect 515362 435544 515730 435568
rect 454905 435514 455225 435538
rect 454905 435242 454929 435514
rect 455201 435242 455225 435514
rect 454905 435218 455225 435242
rect 515362 435212 515386 435544
rect 515706 435538 515730 435544
rect 518241 435538 520957 438218
rect 515706 435218 520957 435538
rect 515706 435212 515730 435218
rect 515362 435188 515730 435212
rect 149102 434408 149964 434728
rect 515362 432544 515730 432568
rect 454905 432514 455225 432538
rect 454905 432242 454929 432514
rect 455201 432242 455225 432514
rect 454905 432218 455225 432242
rect 515362 432212 515386 432544
rect 515706 432538 515730 432544
rect 518241 432538 520957 435218
rect 515706 432218 520957 432538
rect 515706 432212 515730 432218
rect 515362 432188 515730 432212
rect 118982 431792 120252 432112
rect 120572 431792 121698 432112
rect 129057 432088 129377 432112
rect 129057 431816 129081 432088
rect 129353 431816 129377 432088
rect 129057 431792 129377 431816
rect 118982 428112 121698 431792
rect 515362 429544 515730 429568
rect 454905 429514 455225 429538
rect 454905 429242 454929 429514
rect 455201 429242 455225 429514
rect 454905 429218 455225 429242
rect 515362 429212 515386 429544
rect 515706 429538 515730 429544
rect 518241 429538 520957 432218
rect 515706 429218 520957 429538
rect 515706 429212 515730 429218
rect 515362 429188 515730 429212
rect 118982 427792 120252 428112
rect 120572 427792 121698 428112
rect 129057 428088 129377 428112
rect 129057 427816 129081 428088
rect 129353 427816 129377 428088
rect 129057 427792 129377 427816
rect 118982 424112 121698 427792
rect 515362 426544 515730 426568
rect 454905 426514 455225 426538
rect 454905 426242 454929 426514
rect 455201 426242 455225 426514
rect 454905 426218 455225 426242
rect 515362 426212 515386 426544
rect 515706 426538 515730 426544
rect 518241 426538 520957 429218
rect 515706 426218 520957 426538
rect 515706 426212 515730 426218
rect 515362 426188 515730 426212
rect 118982 423792 120252 424112
rect 120572 423792 121698 424112
rect 129057 424088 129377 424112
rect 129057 423816 129081 424088
rect 129353 423816 129377 424088
rect 129057 423792 129377 423816
rect 118982 420112 121698 423792
rect 515362 423544 515730 423568
rect 454905 423514 455225 423538
rect 454905 423242 454929 423514
rect 455201 423242 455225 423514
rect 454905 423218 455225 423242
rect 515362 423212 515386 423544
rect 515706 423538 515730 423544
rect 518241 423538 520957 426218
rect 515706 423218 520957 423538
rect 515706 423212 515730 423218
rect 515362 423188 515730 423212
rect 515362 420544 515730 420568
rect 454905 420514 455225 420538
rect 454905 420242 454929 420514
rect 455201 420242 455225 420514
rect 454905 420218 455225 420242
rect 515362 420212 515386 420544
rect 515706 420538 515730 420544
rect 518241 420538 520957 423218
rect 515706 420218 520957 420538
rect 515706 420212 515730 420218
rect 515362 420188 515730 420212
rect 118982 419792 120252 420112
rect 120572 419792 121698 420112
rect 129057 420088 129377 420112
rect 129057 419816 129081 420088
rect 129353 419816 129377 420088
rect 129057 419792 129377 419816
rect 118982 416112 121698 419792
rect 515362 417544 515730 417568
rect 454905 417514 455225 417538
rect 454905 417242 454929 417514
rect 455201 417242 455225 417514
rect 454905 417218 455225 417242
rect 515362 417212 515386 417544
rect 515706 417538 515730 417544
rect 518241 417538 520957 420218
rect 515706 417218 520957 417538
rect 515706 417212 515730 417218
rect 515362 417188 515730 417212
rect 118982 415792 120252 416112
rect 120572 415792 121698 416112
rect 129057 416088 129377 416112
rect 129057 415816 129081 416088
rect 129353 415816 129377 416088
rect 129057 415792 129377 415816
rect 118982 412112 121698 415792
rect 515362 414544 515730 414568
rect 454905 414514 455225 414538
rect 454905 414242 454929 414514
rect 455201 414242 455225 414514
rect 454905 414218 455225 414242
rect 515362 414212 515386 414544
rect 515706 414538 515730 414544
rect 518241 414538 520957 417218
rect 515706 414218 520957 414538
rect 515706 414212 515730 414218
rect 515362 414188 515730 414212
rect 118982 411792 120252 412112
rect 120572 411792 121698 412112
rect 129057 412088 129377 412112
rect 129057 411816 129081 412088
rect 129353 411816 129377 412088
rect 129057 411792 129377 411816
rect 118982 408112 121698 411792
rect 515362 411544 515730 411568
rect 454905 411514 455225 411538
rect 454905 411242 454929 411514
rect 455201 411242 455225 411514
rect 454905 411218 455225 411242
rect 515362 411212 515386 411544
rect 515706 411538 515730 411544
rect 518241 411538 520957 414218
rect 515706 411218 520957 411538
rect 515706 411212 515730 411218
rect 515362 411188 515730 411212
rect 515362 408544 515730 408568
rect 454905 408514 455225 408538
rect 454905 408242 454929 408514
rect 455201 408242 455225 408514
rect 454905 408218 455225 408242
rect 515362 408212 515386 408544
rect 515706 408538 515730 408544
rect 518241 408538 520957 411218
rect 515706 408218 520957 408538
rect 515706 408212 515730 408218
rect 515362 408188 515730 408212
rect 118982 407792 120252 408112
rect 120572 407792 121698 408112
rect 129057 408088 129377 408112
rect 129057 407816 129081 408088
rect 129353 407816 129377 408088
rect 129057 407792 129377 407816
rect 118982 404112 121698 407792
rect 515362 405544 515730 405568
rect 454905 405514 455225 405538
rect 454905 405242 454929 405514
rect 455201 405242 455225 405514
rect 454905 405218 455225 405242
rect 515362 405212 515386 405544
rect 515706 405538 515730 405544
rect 518241 405538 520957 408218
rect 515706 405218 520957 405538
rect 515706 405212 515730 405218
rect 515362 405188 515730 405212
rect 118982 403792 120252 404112
rect 120572 403792 121698 404112
rect 129057 404088 129377 404112
rect 129057 403816 129081 404088
rect 129353 403816 129377 404088
rect 129057 403792 129377 403816
rect 118982 400112 121698 403792
rect 515362 402544 515730 402568
rect 454905 402514 455225 402538
rect 454905 402242 454929 402514
rect 455201 402242 455225 402514
rect 454905 402218 455225 402242
rect 515362 402212 515386 402544
rect 515706 402538 515730 402544
rect 518241 402538 520957 405218
rect 515706 402218 520957 402538
rect 515706 402212 515730 402218
rect 515362 402188 515730 402212
rect 118982 399792 120252 400112
rect 120572 399792 121698 400112
rect 129057 400088 129377 400112
rect 129057 399816 129081 400088
rect 129353 399816 129377 400088
rect 129057 399792 129377 399816
rect 118982 396112 121698 399792
rect 515362 399544 515730 399568
rect 454905 399514 455225 399538
rect 454905 399242 454929 399514
rect 455201 399242 455225 399514
rect 454905 399218 455225 399242
rect 515362 399212 515386 399544
rect 515706 399538 515730 399544
rect 518241 399538 520957 402218
rect 515706 399218 520957 399538
rect 515706 399212 515730 399218
rect 515362 399188 515730 399212
rect 515362 396544 515730 396568
rect 454905 396514 455225 396538
rect 454905 396242 454929 396514
rect 455201 396242 455225 396514
rect 454905 396218 455225 396242
rect 515362 396212 515386 396544
rect 515706 396538 515730 396544
rect 518241 396538 520957 399218
rect 515706 396218 520957 396538
rect 515706 396212 515730 396218
rect 515362 396188 515730 396212
rect 118982 395792 120252 396112
rect 120572 395792 121698 396112
rect 129057 396088 129377 396112
rect 129057 395816 129081 396088
rect 129353 395816 129377 396088
rect 129057 395792 129377 395816
rect 118982 392112 121698 395792
rect 515362 393544 515730 393568
rect 454905 393514 455225 393538
rect 454905 393242 454929 393514
rect 455201 393242 455225 393514
rect 454905 393218 455225 393242
rect 515362 393212 515386 393544
rect 515706 393538 515730 393544
rect 518241 393538 520957 396218
rect 515706 393218 520957 393538
rect 515706 393212 515730 393218
rect 515362 393188 515730 393212
rect 118982 391792 120252 392112
rect 120572 391792 121698 392112
rect 129057 392088 129377 392112
rect 129057 391816 129081 392088
rect 129353 391816 129377 392088
rect 129057 391792 129377 391816
rect 118982 388112 121698 391792
rect 515362 390544 515730 390568
rect 454905 390514 455225 390538
rect 454905 390242 454929 390514
rect 455201 390242 455225 390514
rect 454905 390218 455225 390242
rect 515362 390212 515386 390544
rect 515706 390538 515730 390544
rect 518241 390538 520957 393218
rect 515706 390218 520957 390538
rect 515706 390212 515730 390218
rect 515362 390188 515730 390212
rect 118982 387792 120252 388112
rect 120572 387792 121698 388112
rect 129057 388088 129377 388112
rect 129057 387816 129081 388088
rect 129353 387816 129377 388088
rect 129057 387792 129377 387816
rect 118982 384112 121698 387792
rect 515362 387544 515730 387568
rect 454905 387514 455225 387538
rect 454905 387242 454929 387514
rect 455201 387242 455225 387514
rect 454905 387218 455225 387242
rect 515362 387212 515386 387544
rect 515706 387538 515730 387544
rect 518241 387538 520957 390218
rect 515706 387218 520957 387538
rect 515706 387212 515730 387218
rect 515362 387188 515730 387212
rect 515362 384544 515730 384568
rect 454905 384514 455225 384538
rect 454905 384242 454929 384514
rect 455201 384242 455225 384514
rect 454905 384218 455225 384242
rect 515362 384212 515386 384544
rect 515706 384538 515730 384544
rect 518241 384538 520957 387218
rect 515706 384218 520957 384538
rect 515706 384212 515730 384218
rect 515362 384188 515730 384212
rect 118982 383792 120252 384112
rect 120572 383792 121698 384112
rect 129057 384088 129377 384112
rect 129057 383816 129081 384088
rect 129353 383816 129377 384088
rect 129057 383792 129377 383816
rect 118982 380112 121698 383792
rect 515362 381544 515730 381568
rect 454905 381514 455225 381538
rect 454905 381242 454929 381514
rect 455201 381242 455225 381514
rect 454905 381218 455225 381242
rect 515362 381212 515386 381544
rect 515706 381538 515730 381544
rect 518241 381538 520957 384218
rect 515706 381218 520957 381538
rect 515706 381212 515730 381218
rect 515362 381188 515730 381212
rect 118982 379792 120252 380112
rect 120572 379792 121698 380112
rect 129057 380088 129377 380112
rect 129057 379816 129081 380088
rect 129353 379816 129377 380088
rect 129057 379792 129377 379816
rect 118982 376112 121698 379792
rect 515362 378544 515730 378568
rect 454905 378514 455225 378538
rect 454905 378242 454929 378514
rect 455201 378242 455225 378514
rect 454905 378218 455225 378242
rect 515362 378212 515386 378544
rect 515706 378538 515730 378544
rect 518241 378538 520957 381218
rect 515706 378218 520957 378538
rect 515706 378212 515730 378218
rect 515362 378188 515730 378212
rect 118982 375792 120252 376112
rect 120572 375792 121698 376112
rect 129057 376088 129377 376112
rect 129057 375816 129081 376088
rect 129353 375816 129377 376088
rect 129057 375792 129377 375816
rect 118982 372112 121698 375792
rect 515362 375544 515730 375568
rect 454905 375514 455225 375538
rect 454905 375242 454929 375514
rect 455201 375242 455225 375514
rect 454905 375218 455225 375242
rect 515362 375212 515386 375544
rect 515706 375538 515730 375544
rect 518241 375538 520957 378218
rect 515706 375218 520957 375538
rect 515706 375212 515730 375218
rect 515362 375188 515730 375212
rect 515362 372544 515730 372568
rect 454905 372514 455225 372538
rect 454905 372242 454929 372514
rect 455201 372242 455225 372514
rect 454905 372218 455225 372242
rect 515362 372212 515386 372544
rect 515706 372538 515730 372544
rect 518241 372538 520957 375218
rect 515706 372218 520957 372538
rect 515706 372212 515730 372218
rect 515362 372188 515730 372212
rect 118982 371792 120252 372112
rect 120572 371792 121698 372112
rect 129057 372088 129377 372112
rect 129057 371816 129081 372088
rect 129353 371816 129377 372088
rect 129057 371792 129377 371816
rect 118982 368112 121698 371792
rect 515362 369544 515730 369568
rect 454905 369514 455225 369538
rect 454905 369242 454929 369514
rect 455201 369242 455225 369514
rect 454905 369218 455225 369242
rect 515362 369212 515386 369544
rect 515706 369538 515730 369544
rect 518241 369538 520957 372218
rect 515706 369218 520957 369538
rect 515706 369212 515730 369218
rect 515362 369188 515730 369212
rect 118982 367792 120252 368112
rect 120572 367792 121698 368112
rect 129057 368088 129377 368112
rect 129057 367816 129081 368088
rect 129353 367816 129377 368088
rect 129057 367792 129377 367816
rect 118982 364112 121698 367792
rect 515362 366544 515730 366568
rect 454905 366514 455225 366538
rect 454905 366242 454929 366514
rect 455201 366242 455225 366514
rect 454905 366218 455225 366242
rect 515362 366212 515386 366544
rect 515706 366538 515730 366544
rect 518241 366538 520957 369218
rect 515706 366218 520957 366538
rect 515706 366212 515730 366218
rect 515362 366188 515730 366212
rect 118982 363792 120252 364112
rect 120572 363792 121698 364112
rect 129057 364088 129377 364112
rect 129057 363816 129081 364088
rect 129353 363816 129377 364088
rect 129057 363792 129377 363816
rect 118982 360112 121698 363792
rect 515362 363544 515730 363568
rect 454905 363514 455225 363538
rect 454905 363242 454929 363514
rect 455201 363242 455225 363514
rect 454905 363218 455225 363242
rect 515362 363212 515386 363544
rect 515706 363538 515730 363544
rect 518241 363538 520957 366218
rect 515706 363218 520957 363538
rect 515706 363212 515730 363218
rect 515362 363188 515730 363212
rect 515362 360544 515730 360568
rect 454905 360514 455225 360538
rect 454905 360242 454929 360514
rect 455201 360242 455225 360514
rect 454905 360218 455225 360242
rect 515362 360212 515386 360544
rect 515706 360538 515730 360544
rect 518241 360538 520957 363218
rect 515706 360218 520957 360538
rect 515706 360212 515730 360218
rect 515362 360188 515730 360212
rect 118982 359792 120252 360112
rect 120572 359792 121698 360112
rect 129057 360088 129377 360112
rect 129057 359816 129081 360088
rect 129353 359816 129377 360088
rect 129057 359792 129377 359816
rect 118982 356112 121698 359792
rect 515362 357544 515730 357568
rect 454905 357514 455225 357538
rect 454905 357242 454929 357514
rect 455201 357242 455225 357514
rect 454905 357218 455225 357242
rect 515362 357212 515386 357544
rect 515706 357538 515730 357544
rect 518241 357538 520957 360218
rect 515706 357218 520957 357538
rect 515706 357212 515730 357218
rect 515362 357188 515730 357212
rect 118982 355792 120252 356112
rect 120572 355792 121698 356112
rect 129057 356088 129377 356112
rect 129057 355816 129081 356088
rect 129353 355816 129377 356088
rect 129057 355792 129377 355816
rect 118982 352112 121698 355792
rect 515362 354544 515730 354568
rect 454905 354514 455225 354538
rect 454905 354242 454929 354514
rect 455201 354242 455225 354514
rect 454905 354218 455225 354242
rect 515362 354212 515386 354544
rect 515706 354538 515730 354544
rect 518241 354538 520957 357218
rect 515706 354218 520957 354538
rect 515706 354212 515730 354218
rect 515362 354188 515730 354212
rect 118982 351792 120252 352112
rect 120572 351792 121698 352112
rect 129057 352088 129377 352112
rect 129057 351816 129081 352088
rect 129353 351816 129377 352088
rect 129057 351792 129377 351816
rect 118982 348112 121698 351792
rect 515362 351544 515730 351568
rect 454905 351514 455225 351538
rect 454905 351242 454929 351514
rect 455201 351242 455225 351514
rect 454905 351218 455225 351242
rect 515362 351212 515386 351544
rect 515706 351538 515730 351544
rect 518241 351538 520957 354218
rect 515706 351218 520957 351538
rect 515706 351212 515730 351218
rect 515362 351188 515730 351212
rect 515362 348544 515730 348568
rect 454905 348514 455225 348538
rect 454905 348242 454929 348514
rect 455201 348242 455225 348514
rect 454905 348218 455225 348242
rect 515362 348212 515386 348544
rect 515706 348538 515730 348544
rect 518241 348538 520957 351218
rect 515706 348218 520957 348538
rect 515706 348212 515730 348218
rect 515362 348188 515730 348212
rect 118982 347792 120252 348112
rect 120572 347792 121698 348112
rect 129057 348088 129377 348112
rect 129057 347816 129081 348088
rect 129353 347816 129377 348088
rect 129057 347792 129377 347816
rect 118982 344112 121698 347792
rect 515362 345544 515730 345568
rect 454905 345514 455225 345538
rect 454905 345242 454929 345514
rect 455201 345242 455225 345514
rect 454905 345218 455225 345242
rect 515362 345212 515386 345544
rect 515706 345538 515730 345544
rect 518241 345538 520957 348218
rect 515706 345218 520957 345538
rect 515706 345212 515730 345218
rect 515362 345188 515730 345212
rect 118982 343792 120252 344112
rect 120572 343792 121698 344112
rect 129057 344088 129377 344112
rect 129057 343816 129081 344088
rect 129353 343816 129377 344088
rect 129057 343792 129377 343816
rect 118982 340112 121698 343792
rect 515362 342544 515730 342568
rect 454905 342514 455225 342538
rect 454905 342242 454929 342514
rect 455201 342242 455225 342514
rect 454905 342218 455225 342242
rect 515362 342212 515386 342544
rect 515706 342538 515730 342544
rect 518241 342538 520957 345218
rect 515706 342218 520957 342538
rect 515706 342212 515730 342218
rect 515362 342188 515730 342212
rect 118982 339792 120252 340112
rect 120572 339792 121698 340112
rect 129057 340088 129377 340112
rect 129057 339816 129081 340088
rect 129353 339816 129377 340088
rect 129057 339792 129377 339816
rect 118982 336112 121698 339792
rect 515362 339544 515730 339568
rect 454905 339514 455225 339538
rect 454905 339242 454929 339514
rect 455201 339242 455225 339514
rect 454905 339218 455225 339242
rect 515362 339212 515386 339544
rect 515706 339538 515730 339544
rect 518241 339538 520957 342218
rect 515706 339218 520957 339538
rect 515706 339212 515730 339218
rect 515362 339188 515730 339212
rect 515362 336544 515730 336568
rect 454905 336514 455225 336538
rect 454905 336242 454929 336514
rect 455201 336242 455225 336514
rect 454905 336218 455225 336242
rect 515362 336212 515386 336544
rect 515706 336538 515730 336544
rect 518241 336538 520957 339218
rect 515706 336218 520957 336538
rect 515706 336212 515730 336218
rect 515362 336188 515730 336212
rect 118982 335792 120252 336112
rect 120572 335792 121698 336112
rect 129057 336088 129377 336112
rect 129057 335816 129081 336088
rect 129353 335816 129377 336088
rect 129057 335792 129377 335816
rect 118982 332112 121698 335792
rect 515362 333544 515730 333568
rect 454905 333514 455225 333538
rect 454905 333242 454929 333514
rect 455201 333242 455225 333514
rect 454905 333218 455225 333242
rect 515362 333212 515386 333544
rect 515706 333538 515730 333544
rect 518241 333538 520957 336218
rect 515706 333218 520957 333538
rect 515706 333212 515730 333218
rect 515362 333188 515730 333212
rect 118982 331792 120252 332112
rect 120572 331792 121698 332112
rect 129057 332088 129377 332112
rect 129057 331816 129081 332088
rect 129353 331816 129377 332088
rect 129057 331792 129377 331816
rect 118982 328112 121698 331792
rect 515362 330544 515730 330568
rect 454905 330514 455225 330538
rect 454905 330242 454929 330514
rect 455201 330242 455225 330514
rect 454905 330218 455225 330242
rect 515362 330212 515386 330544
rect 515706 330538 515730 330544
rect 518241 330538 520957 333218
rect 515706 330218 520957 330538
rect 515706 330212 515730 330218
rect 515362 330188 515730 330212
rect 118982 327792 120252 328112
rect 120572 327792 121698 328112
rect 129057 328088 129377 328112
rect 129057 327816 129081 328088
rect 129353 327816 129377 328088
rect 129057 327792 129377 327816
rect 118982 324112 121698 327792
rect 515362 327544 515730 327568
rect 454905 327514 455225 327538
rect 454905 327242 454929 327514
rect 455201 327242 455225 327514
rect 454905 327218 455225 327242
rect 515362 327212 515386 327544
rect 515706 327538 515730 327544
rect 518241 327538 520957 330218
rect 515706 327218 520957 327538
rect 515706 327212 515730 327218
rect 515362 327188 515730 327212
rect 515362 324544 515730 324568
rect 454905 324514 455225 324538
rect 454905 324242 454929 324514
rect 455201 324242 455225 324514
rect 454905 324218 455225 324242
rect 515362 324212 515386 324544
rect 515706 324538 515730 324544
rect 518241 324538 520957 327218
rect 515706 324218 520957 324538
rect 515706 324212 515730 324218
rect 515362 324188 515730 324212
rect 118982 323792 120252 324112
rect 120572 323792 121698 324112
rect 129057 324088 129377 324112
rect 129057 323816 129081 324088
rect 129353 323816 129377 324088
rect 129057 323792 129377 323816
rect 118982 320112 121698 323792
rect 515362 321544 515730 321568
rect 454905 321514 455225 321538
rect 454905 321242 454929 321514
rect 455201 321242 455225 321514
rect 454905 321218 455225 321242
rect 515362 321212 515386 321544
rect 515706 321538 515730 321544
rect 518241 321538 520957 324218
rect 515706 321218 520957 321538
rect 515706 321212 515730 321218
rect 515362 321188 515730 321212
rect 118982 319792 120252 320112
rect 120572 319792 121698 320112
rect 129057 320088 129377 320112
rect 129057 319816 129081 320088
rect 129353 319816 129377 320088
rect 129057 319792 129377 319816
rect 118982 316112 121698 319792
rect 515362 318544 515730 318568
rect 454905 318514 455225 318538
rect 454905 318242 454929 318514
rect 455201 318242 455225 318514
rect 454905 318218 455225 318242
rect 515362 318212 515386 318544
rect 515706 318538 515730 318544
rect 518241 318538 520957 321218
rect 515706 318218 520957 318538
rect 515706 318212 515730 318218
rect 515362 318188 515730 318212
rect 118982 315792 120252 316112
rect 120572 315792 121698 316112
rect 129057 316088 129377 316112
rect 129057 315816 129081 316088
rect 129353 315816 129377 316088
rect 129057 315792 129377 315816
rect 118982 312112 121698 315792
rect 515362 315544 515730 315568
rect 454905 315514 455225 315538
rect 454905 315242 454929 315514
rect 455201 315242 455225 315514
rect 454905 315218 455225 315242
rect 515362 315212 515386 315544
rect 515706 315538 515730 315544
rect 518241 315538 520957 318218
rect 515706 315218 520957 315538
rect 515706 315212 515730 315218
rect 515362 315188 515730 315212
rect 515362 312544 515730 312568
rect 454905 312514 455225 312538
rect 454905 312242 454929 312514
rect 455201 312242 455225 312514
rect 454905 312218 455225 312242
rect 515362 312212 515386 312544
rect 515706 312538 515730 312544
rect 518241 312538 520957 315218
rect 515706 312218 520957 312538
rect 515706 312212 515730 312218
rect 515362 312188 515730 312212
rect 118982 311792 120252 312112
rect 120572 311792 121698 312112
rect 129057 312088 129377 312112
rect 129057 311816 129081 312088
rect 129353 311816 129377 312088
rect 129057 311792 129377 311816
rect 118982 308112 121698 311792
rect 515362 309544 515730 309568
rect 454905 309514 455225 309538
rect 454905 309242 454929 309514
rect 455201 309242 455225 309514
rect 454905 309218 455225 309242
rect 515362 309212 515386 309544
rect 515706 309538 515730 309544
rect 518241 309538 520957 312218
rect 515706 309218 520957 309538
rect 515706 309212 515730 309218
rect 515362 309188 515730 309212
rect 118982 307792 120252 308112
rect 120572 307792 121698 308112
rect 129057 308088 129377 308112
rect 129057 307816 129081 308088
rect 129353 307816 129377 308088
rect 129057 307792 129377 307816
rect 118982 304112 121698 307792
rect 515362 306544 515730 306568
rect 454905 306514 455225 306538
rect 454905 306242 454929 306514
rect 455201 306242 455225 306514
rect 454905 306218 455225 306242
rect 515362 306212 515386 306544
rect 515706 306538 515730 306544
rect 518241 306538 520957 309218
rect 515706 306218 520957 306538
rect 515706 306212 515730 306218
rect 515362 306188 515730 306212
rect 118982 303792 120252 304112
rect 120572 303792 121698 304112
rect 129057 304088 129377 304112
rect 129057 303816 129081 304088
rect 129353 303816 129377 304088
rect 129057 303792 129377 303816
rect 118982 300112 121698 303792
rect 515362 303544 515730 303568
rect 454905 303514 455225 303538
rect 454905 303242 454929 303514
rect 455201 303242 455225 303514
rect 454905 303218 455225 303242
rect 515362 303212 515386 303544
rect 515706 303538 515730 303544
rect 518241 303538 520957 306218
rect 515706 303218 520957 303538
rect 515706 303212 515730 303218
rect 515362 303188 515730 303212
rect 515362 300544 515730 300568
rect 454905 300514 455225 300538
rect 454905 300242 454929 300514
rect 455201 300242 455225 300514
rect 454905 300218 455225 300242
rect 515362 300212 515386 300544
rect 515706 300538 515730 300544
rect 518241 300538 520957 303218
rect 515706 300218 520957 300538
rect 515706 300212 515730 300218
rect 515362 300188 515730 300212
rect 118982 299792 120252 300112
rect 120572 299792 121698 300112
rect 129057 300088 129377 300112
rect 129057 299816 129081 300088
rect 129353 299816 129377 300088
rect 129057 299792 129377 299816
rect 118982 296112 121698 299792
rect 515362 297544 515730 297568
rect 454905 297514 455225 297538
rect 454905 297242 454929 297514
rect 455201 297242 455225 297514
rect 454905 297218 455225 297242
rect 515362 297212 515386 297544
rect 515706 297538 515730 297544
rect 518241 297538 520957 300218
rect 515706 297218 520957 297538
rect 515706 297212 515730 297218
rect 515362 297188 515730 297212
rect 118982 295792 120252 296112
rect 120572 295792 121698 296112
rect 129057 296088 129377 296112
rect 129057 295816 129081 296088
rect 129353 295816 129377 296088
rect 129057 295792 129377 295816
rect 118982 292112 121698 295792
rect 515362 294544 515730 294568
rect 454905 294514 455225 294538
rect 454905 294242 454929 294514
rect 455201 294242 455225 294514
rect 454905 294218 455225 294242
rect 515362 294212 515386 294544
rect 515706 294538 515730 294544
rect 518241 294538 520957 297218
rect 515706 294218 520957 294538
rect 515706 294212 515730 294218
rect 515362 294188 515730 294212
rect 118982 291792 120252 292112
rect 120572 291792 121698 292112
rect 129057 292088 129377 292112
rect 129057 291816 129081 292088
rect 129353 291816 129377 292088
rect 129057 291792 129377 291816
rect 118982 288112 121698 291792
rect 515362 291544 515730 291568
rect 454905 291514 455225 291538
rect 454905 291242 454929 291514
rect 455201 291242 455225 291514
rect 454905 291218 455225 291242
rect 515362 291212 515386 291544
rect 515706 291538 515730 291544
rect 518241 291538 520957 294218
rect 515706 291218 520957 291538
rect 515706 291212 515730 291218
rect 515362 291188 515730 291212
rect 515362 288544 515730 288568
rect 454905 288514 455225 288538
rect 454905 288242 454929 288514
rect 455201 288242 455225 288514
rect 454905 288218 455225 288242
rect 515362 288212 515386 288544
rect 515706 288538 515730 288544
rect 518241 288538 520957 291218
rect 515706 288218 520957 288538
rect 515706 288212 515730 288218
rect 515362 288188 515730 288212
rect 118982 287792 120252 288112
rect 120572 287792 121698 288112
rect 129057 288088 129377 288112
rect 129057 287816 129081 288088
rect 129353 287816 129377 288088
rect 129057 287792 129377 287816
rect 118982 284112 121698 287792
rect 515362 285544 515730 285568
rect 454905 285514 455225 285538
rect 454905 285242 454929 285514
rect 455201 285242 455225 285514
rect 454905 285218 455225 285242
rect 515362 285212 515386 285544
rect 515706 285538 515730 285544
rect 518241 285538 520957 288218
rect 515706 285218 520957 285538
rect 515706 285212 515730 285218
rect 515362 285188 515730 285212
rect 118982 283792 120252 284112
rect 120572 283792 121698 284112
rect 129057 284088 129377 284112
rect 129057 283816 129081 284088
rect 129353 283816 129377 284088
rect 129057 283792 129377 283816
rect 118982 280112 121698 283792
rect 515362 282544 515730 282568
rect 454905 282514 455225 282538
rect 454905 282242 454929 282514
rect 455201 282242 455225 282514
rect 454905 282218 455225 282242
rect 515362 282212 515386 282544
rect 515706 282538 515730 282544
rect 518241 282538 520957 285218
rect 515706 282218 520957 282538
rect 515706 282212 515730 282218
rect 515362 282188 515730 282212
rect 118982 279792 120252 280112
rect 120572 279792 121698 280112
rect 129057 280088 129377 280112
rect 129057 279816 129081 280088
rect 129353 279816 129377 280088
rect 129057 279792 129377 279816
rect 118982 276112 121698 279792
rect 515362 279544 515730 279568
rect 454905 279514 455225 279538
rect 454905 279242 454929 279514
rect 455201 279242 455225 279514
rect 454905 279218 455225 279242
rect 515362 279212 515386 279544
rect 515706 279538 515730 279544
rect 518241 279538 520957 282218
rect 515706 279218 520957 279538
rect 515706 279212 515730 279218
rect 515362 279188 515730 279212
rect 515362 276544 515730 276568
rect 454905 276514 455225 276538
rect 454905 276242 454929 276514
rect 455201 276242 455225 276514
rect 454905 276218 455225 276242
rect 515362 276212 515386 276544
rect 515706 276538 515730 276544
rect 518241 276538 520957 279218
rect 515706 276218 520957 276538
rect 515706 276212 515730 276218
rect 515362 276188 515730 276212
rect 118982 275792 120252 276112
rect 120572 275792 121698 276112
rect 129057 276088 129377 276112
rect 129057 275816 129081 276088
rect 129353 275816 129377 276088
rect 129057 275792 129377 275816
rect 118982 272112 121698 275792
rect 515362 273544 515730 273568
rect 454905 273514 455225 273538
rect 454905 273242 454929 273514
rect 455201 273242 455225 273514
rect 454905 273218 455225 273242
rect 515362 273212 515386 273544
rect 515706 273538 515730 273544
rect 518241 273538 520957 276218
rect 515706 273218 520957 273538
rect 515706 273212 515730 273218
rect 515362 273188 515730 273212
rect 118982 271792 120252 272112
rect 120572 271792 121698 272112
rect 129057 272088 129377 272112
rect 129057 271816 129081 272088
rect 129353 271816 129377 272088
rect 129057 271792 129377 271816
rect 118982 268112 121698 271792
rect 515362 270544 515730 270568
rect 454905 270514 455225 270538
rect 454905 270242 454929 270514
rect 455201 270242 455225 270514
rect 454905 270218 455225 270242
rect 515362 270212 515386 270544
rect 515706 270538 515730 270544
rect 518241 270538 520957 273218
rect 515706 270218 520957 270538
rect 515706 270212 515730 270218
rect 515362 270188 515730 270212
rect 118982 267792 120252 268112
rect 120572 267792 121698 268112
rect 129057 268088 129377 268112
rect 129057 267816 129081 268088
rect 129353 267816 129377 268088
rect 129057 267792 129377 267816
rect 118982 264112 121698 267792
rect 515362 267544 515730 267568
rect 454905 267514 455225 267538
rect 454905 267242 454929 267514
rect 455201 267242 455225 267514
rect 454905 267218 455225 267242
rect 515362 267212 515386 267544
rect 515706 267538 515730 267544
rect 518241 267538 520957 270218
rect 515706 267218 520957 267538
rect 515706 267212 515730 267218
rect 515362 267188 515730 267212
rect 515362 264544 515730 264568
rect 454905 264514 455225 264538
rect 454905 264242 454929 264514
rect 455201 264242 455225 264514
rect 454905 264218 455225 264242
rect 515362 264212 515386 264544
rect 515706 264538 515730 264544
rect 518241 264538 520957 267218
rect 515706 264218 520957 264538
rect 515706 264212 515730 264218
rect 515362 264188 515730 264212
rect 118982 263792 120252 264112
rect 120572 263792 121698 264112
rect 129057 264088 129377 264112
rect 129057 263816 129081 264088
rect 129353 263816 129377 264088
rect 129057 263792 129377 263816
rect 118982 260112 121698 263792
rect 515362 261544 515730 261568
rect 454905 261514 455225 261538
rect 454905 261242 454929 261514
rect 455201 261242 455225 261514
rect 454905 261218 455225 261242
rect 515362 261212 515386 261544
rect 515706 261538 515730 261544
rect 518241 261538 520957 264218
rect 515706 261218 520957 261538
rect 515706 261212 515730 261218
rect 515362 261188 515730 261212
rect 118982 259792 120252 260112
rect 120572 259792 121698 260112
rect 129057 260088 129377 260112
rect 129057 259816 129081 260088
rect 129353 259816 129377 260088
rect 129057 259792 129377 259816
rect 118982 256112 121698 259792
rect 515362 258544 515730 258568
rect 454905 258514 455225 258538
rect 454905 258242 454929 258514
rect 455201 258242 455225 258514
rect 454905 258218 455225 258242
rect 515362 258212 515386 258544
rect 515706 258538 515730 258544
rect 518241 258538 520957 261218
rect 515706 258218 520957 258538
rect 515706 258212 515730 258218
rect 515362 258188 515730 258212
rect 118982 255792 120252 256112
rect 120572 255792 121698 256112
rect 129057 256088 129377 256112
rect 129057 255816 129081 256088
rect 129353 255816 129377 256088
rect 129057 255792 129377 255816
rect 118982 252112 121698 255792
rect 515362 255544 515730 255568
rect 454905 255514 455225 255538
rect 454905 255242 454929 255514
rect 455201 255242 455225 255514
rect 454905 255218 455225 255242
rect 515362 255212 515386 255544
rect 515706 255538 515730 255544
rect 518241 255538 520957 258218
rect 515706 255218 520957 255538
rect 515706 255212 515730 255218
rect 515362 255188 515730 255212
rect 515362 252544 515730 252568
rect 454905 252514 455225 252538
rect 454905 252242 454929 252514
rect 455201 252242 455225 252514
rect 454905 252218 455225 252242
rect 515362 252212 515386 252544
rect 515706 252538 515730 252544
rect 518241 252538 520957 255218
rect 515706 252218 520957 252538
rect 515706 252212 515730 252218
rect 515362 252188 515730 252212
rect 118982 251792 120252 252112
rect 120572 251792 121698 252112
rect 129057 252088 129377 252112
rect 129057 251816 129081 252088
rect 129353 251816 129377 252088
rect 129057 251792 129377 251816
rect 118982 248112 121698 251792
rect 515362 249544 515730 249568
rect 454905 249514 455225 249538
rect 454905 249242 454929 249514
rect 455201 249242 455225 249514
rect 454905 249218 455225 249242
rect 515362 249212 515386 249544
rect 515706 249538 515730 249544
rect 518241 249538 520957 252218
rect 515706 249218 520957 249538
rect 515706 249212 515730 249218
rect 515362 249188 515730 249212
rect 118982 247792 120252 248112
rect 120572 247792 121698 248112
rect 129057 248088 129377 248112
rect 129057 247816 129081 248088
rect 129353 247816 129377 248088
rect 129057 247792 129377 247816
rect 118982 244112 121698 247792
rect 515362 246544 515730 246568
rect 454905 246514 455225 246538
rect 454905 246242 454929 246514
rect 455201 246242 455225 246514
rect 454905 246218 455225 246242
rect 515362 246212 515386 246544
rect 515706 246538 515730 246544
rect 518241 246538 520957 249218
rect 515706 246218 520957 246538
rect 515706 246212 515730 246218
rect 515362 246188 515730 246212
rect 118982 243792 120252 244112
rect 120572 243792 121698 244112
rect 129057 244088 129377 244112
rect 129057 243816 129081 244088
rect 129353 243816 129377 244088
rect 129057 243792 129377 243816
rect 118982 240112 121698 243792
rect 515362 243544 515730 243568
rect 454905 243514 455225 243538
rect 454905 243242 454929 243514
rect 455201 243242 455225 243514
rect 454905 243218 455225 243242
rect 515362 243212 515386 243544
rect 515706 243538 515730 243544
rect 518241 243538 520957 246218
rect 515706 243218 520957 243538
rect 515706 243212 515730 243218
rect 515362 243188 515730 243212
rect 515362 240544 515730 240568
rect 454905 240514 455225 240538
rect 454905 240242 454929 240514
rect 455201 240242 455225 240514
rect 454905 240218 455225 240242
rect 515362 240212 515386 240544
rect 515706 240538 515730 240544
rect 518241 240538 520957 243218
rect 515706 240218 520957 240538
rect 515706 240212 515730 240218
rect 515362 240188 515730 240212
rect 118982 239792 120252 240112
rect 120572 239792 121698 240112
rect 129057 240088 129377 240112
rect 129057 239816 129081 240088
rect 129353 239816 129377 240088
rect 129057 239792 129377 239816
rect 118982 236112 121698 239792
rect 515362 237544 515730 237568
rect 454905 237514 455225 237538
rect 454905 237242 454929 237514
rect 455201 237242 455225 237514
rect 454905 237218 455225 237242
rect 515362 237212 515386 237544
rect 515706 237538 515730 237544
rect 518241 237538 520957 240218
rect 515706 237218 520957 237538
rect 515706 237212 515730 237218
rect 515362 237188 515730 237212
rect 118982 235792 120252 236112
rect 120572 235792 121698 236112
rect 129057 236088 129377 236112
rect 129057 235816 129081 236088
rect 129353 235816 129377 236088
rect 129057 235792 129377 235816
rect 118982 232112 121698 235792
rect 515362 234544 515730 234568
rect 454905 234514 455225 234538
rect 454905 234242 454929 234514
rect 455201 234242 455225 234514
rect 454905 234218 455225 234242
rect 515362 234212 515386 234544
rect 515706 234538 515730 234544
rect 518241 234538 520957 237218
rect 515706 234218 520957 234538
rect 515706 234212 515730 234218
rect 515362 234188 515730 234212
rect 118982 231792 120252 232112
rect 120572 231792 121698 232112
rect 129057 232088 129377 232112
rect 129057 231816 129081 232088
rect 129353 231816 129377 232088
rect 129057 231792 129377 231816
rect 118982 228112 121698 231792
rect 515362 231544 515730 231568
rect 454905 231514 455225 231538
rect 454905 231242 454929 231514
rect 455201 231242 455225 231514
rect 454905 231218 455225 231242
rect 515362 231212 515386 231544
rect 515706 231538 515730 231544
rect 518241 231538 520957 234218
rect 515706 231218 520957 231538
rect 515706 231212 515730 231218
rect 515362 231188 515730 231212
rect 515362 228544 515730 228568
rect 454905 228514 455225 228538
rect 454905 228242 454929 228514
rect 455201 228242 455225 228514
rect 454905 228218 455225 228242
rect 515362 228212 515386 228544
rect 515706 228538 515730 228544
rect 518241 228538 520957 231218
rect 515706 228218 520957 228538
rect 515706 228212 515730 228218
rect 515362 228188 515730 228212
rect 118982 227792 120252 228112
rect 120572 227792 121698 228112
rect 129057 228088 129377 228112
rect 129057 227816 129081 228088
rect 129353 227816 129377 228088
rect 129057 227792 129377 227816
rect 118982 224112 121698 227792
rect 515362 225544 515730 225568
rect 454905 225514 455225 225538
rect 454905 225242 454929 225514
rect 455201 225242 455225 225514
rect 454905 225218 455225 225242
rect 515362 225212 515386 225544
rect 515706 225538 515730 225544
rect 518241 225538 520957 228218
rect 515706 225218 520957 225538
rect 515706 225212 515730 225218
rect 515362 225188 515730 225212
rect 118982 223792 120252 224112
rect 120572 223792 121698 224112
rect 129057 224088 129377 224112
rect 129057 223816 129081 224088
rect 129353 223816 129377 224088
rect 129057 223792 129377 223816
rect 118982 220112 121698 223792
rect 515362 222544 515730 222568
rect 454905 222514 455225 222538
rect 454905 222242 454929 222514
rect 455201 222242 455225 222514
rect 454905 222218 455225 222242
rect 515362 222212 515386 222544
rect 515706 222538 515730 222544
rect 518241 222538 520957 225218
rect 515706 222218 520957 222538
rect 515706 222212 515730 222218
rect 515362 222188 515730 222212
rect 118982 219792 120252 220112
rect 120572 219792 121698 220112
rect 129057 220088 129377 220112
rect 129057 219816 129081 220088
rect 129353 219816 129377 220088
rect 129057 219792 129377 219816
rect 118982 216112 121698 219792
rect 515362 219544 515730 219568
rect 454905 219514 455225 219538
rect 454905 219242 454929 219514
rect 455201 219242 455225 219514
rect 454905 219218 455225 219242
rect 515362 219212 515386 219544
rect 515706 219538 515730 219544
rect 518241 219538 520957 222218
rect 515706 219218 520957 219538
rect 515706 219212 515730 219218
rect 515362 219188 515730 219212
rect 515362 216544 515730 216568
rect 454905 216514 455225 216538
rect 454905 216242 454929 216514
rect 455201 216242 455225 216514
rect 454905 216218 455225 216242
rect 515362 216212 515386 216544
rect 515706 216538 515730 216544
rect 518241 216538 520957 219218
rect 515706 216218 520957 216538
rect 515706 216212 515730 216218
rect 515362 216188 515730 216212
rect 118982 215792 120252 216112
rect 120572 215792 121698 216112
rect 129057 216088 129377 216112
rect 129057 215816 129081 216088
rect 129353 215816 129377 216088
rect 129057 215792 129377 215816
rect 118982 212112 121698 215792
rect 515362 213544 515730 213568
rect 454905 213514 455225 213538
rect 454905 213242 454929 213514
rect 455201 213242 455225 213514
rect 454905 213218 455225 213242
rect 515362 213212 515386 213544
rect 515706 213538 515730 213544
rect 518241 213538 520957 216218
rect 515706 213218 520957 213538
rect 515706 213212 515730 213218
rect 515362 213188 515730 213212
rect 118982 211792 120252 212112
rect 120572 211792 121698 212112
rect 129057 212088 129377 212112
rect 129057 211816 129081 212088
rect 129353 211816 129377 212088
rect 129057 211792 129377 211816
rect 118982 208112 121698 211792
rect 515362 210544 515730 210568
rect 454905 210514 455225 210538
rect 454905 210242 454929 210514
rect 455201 210242 455225 210514
rect 454905 210218 455225 210242
rect 515362 210212 515386 210544
rect 515706 210538 515730 210544
rect 518241 210538 520957 213218
rect 515706 210218 520957 210538
rect 515706 210212 515730 210218
rect 515362 210188 515730 210212
rect 118982 207792 120252 208112
rect 120572 207792 121698 208112
rect 129057 208088 129377 208112
rect 129057 207816 129081 208088
rect 129353 207816 129377 208088
rect 129057 207792 129377 207816
rect 118982 204112 121698 207792
rect 515362 207544 515730 207568
rect 454905 207514 455225 207538
rect 454905 207242 454929 207514
rect 455201 207242 455225 207514
rect 454905 207218 455225 207242
rect 515362 207212 515386 207544
rect 515706 207538 515730 207544
rect 518241 207538 520957 210218
rect 515706 207218 520957 207538
rect 515706 207212 515730 207218
rect 515362 207188 515730 207212
rect 515362 204544 515730 204568
rect 454905 204514 455225 204538
rect 454905 204242 454929 204514
rect 455201 204242 455225 204514
rect 454905 204218 455225 204242
rect 515362 204212 515386 204544
rect 515706 204538 515730 204544
rect 518241 204538 520957 207218
rect 515706 204218 520957 204538
rect 515706 204212 515730 204218
rect 515362 204188 515730 204212
rect 118982 203792 120252 204112
rect 120572 203792 121698 204112
rect 129057 204088 129377 204112
rect 129057 203816 129081 204088
rect 129353 203816 129377 204088
rect 129057 203792 129377 203816
rect 118982 200112 121698 203792
rect 515362 201544 515730 201568
rect 454905 201514 455225 201538
rect 454905 201242 454929 201514
rect 455201 201242 455225 201514
rect 454905 201218 455225 201242
rect 515362 201212 515386 201544
rect 515706 201538 515730 201544
rect 518241 201538 520957 204218
rect 515706 201218 520957 201538
rect 515706 201212 515730 201218
rect 515362 201188 515730 201212
rect 118982 199792 120252 200112
rect 120572 199792 121698 200112
rect 129057 200088 129377 200112
rect 129057 199816 129081 200088
rect 129353 199816 129377 200088
rect 129057 199792 129377 199816
rect 118982 196112 121698 199792
rect 515362 198544 515730 198568
rect 454905 198514 455225 198538
rect 454905 198242 454929 198514
rect 455201 198242 455225 198514
rect 454905 198218 455225 198242
rect 515362 198212 515386 198544
rect 515706 198538 515730 198544
rect 518241 198538 520957 201218
rect 515706 198218 520957 198538
rect 553276 198242 558076 453196
rect 515706 198212 515730 198218
rect 515362 198188 515730 198212
rect 118982 195792 120252 196112
rect 120572 195792 121698 196112
rect 129057 196088 129377 196112
rect 129057 195816 129081 196088
rect 129353 195816 129377 196088
rect 129057 195792 129377 195816
rect 118982 192112 121698 195792
rect 515362 195544 515730 195568
rect 454905 195514 455225 195538
rect 454905 195242 454929 195514
rect 455201 195242 455225 195514
rect 454905 195218 455225 195242
rect 515362 195212 515386 195544
rect 515706 195538 515730 195544
rect 518241 195538 520957 198218
rect 515706 195218 520957 195538
rect 515706 195212 515730 195218
rect 515362 195188 515730 195212
rect 515362 192544 515730 192568
rect 454905 192514 455225 192538
rect 454905 192242 454929 192514
rect 455201 192242 455225 192514
rect 454905 192218 455225 192242
rect 515362 192212 515386 192544
rect 515706 192538 515730 192544
rect 518241 192538 520957 195218
rect 515706 192218 520957 192538
rect 515706 192212 515730 192218
rect 515362 192188 515730 192212
rect 118982 191792 120252 192112
rect 120572 191792 121698 192112
rect 129057 192088 129377 192112
rect 129057 191816 129081 192088
rect 129353 191816 129377 192088
rect 129057 191792 129377 191816
rect 118982 188112 121698 191792
rect 515362 189544 515730 189568
rect 454905 189514 455225 189538
rect 454905 189242 454929 189514
rect 455201 189242 455225 189514
rect 454905 189218 455225 189242
rect 515362 189212 515386 189544
rect 515706 189538 515730 189544
rect 518241 189538 520957 192218
rect 552812 196966 579468 198242
rect 552812 191768 554140 196966
rect 578296 191768 579468 196966
rect 552812 190928 579468 191768
rect 515706 189218 520957 189538
rect 515706 189212 515730 189218
rect 515362 189188 515730 189212
rect 118982 187792 120252 188112
rect 120572 187792 121698 188112
rect 129057 188088 129377 188112
rect 129057 187816 129081 188088
rect 129353 187816 129377 188088
rect 129057 187792 129377 187816
rect 118982 184112 121698 187792
rect 515362 186544 515730 186568
rect 454905 186514 455225 186538
rect 454905 186242 454929 186514
rect 455201 186242 455225 186514
rect 454905 186218 455225 186242
rect 515362 186212 515386 186544
rect 515706 186538 515730 186544
rect 518241 186538 520957 189218
rect 553276 187154 558076 190928
rect 515706 186218 520957 186538
rect 515706 186212 515730 186218
rect 515362 186188 515730 186212
rect 118982 183792 120252 184112
rect 120572 183792 121698 184112
rect 129057 184088 129377 184112
rect 129057 183816 129081 184088
rect 129353 183816 129377 184088
rect 129057 183792 129377 183816
rect 118982 180112 121698 183792
rect 515362 183544 515730 183568
rect 454905 183514 455225 183538
rect 454905 183242 454929 183514
rect 455201 183242 455225 183514
rect 454905 183218 455225 183242
rect 515362 183212 515386 183544
rect 515706 183538 515730 183544
rect 518241 183538 520957 186218
rect 515706 183218 520957 183538
rect 515706 183212 515730 183218
rect 515362 183188 515730 183212
rect 515362 180544 515730 180568
rect 454905 180514 455225 180538
rect 454905 180242 454929 180514
rect 455201 180242 455225 180514
rect 454905 180218 455225 180242
rect 515362 180212 515386 180544
rect 515706 180538 515730 180544
rect 518241 180538 520957 183218
rect 551320 186340 579660 187154
rect 551320 181150 553050 186340
rect 576862 181150 579660 186340
rect 551320 180540 579660 181150
rect 515706 180218 520957 180538
rect 515706 180212 515730 180218
rect 515362 180188 515730 180212
rect 118982 179792 120252 180112
rect 120572 179792 121698 180112
rect 129057 180088 129377 180112
rect 129057 179816 129081 180088
rect 129353 179816 129377 180088
rect 129057 179792 129377 179816
rect 118982 176112 121698 179792
rect 515362 177544 515730 177568
rect 454905 177514 455225 177538
rect 454905 177242 454929 177514
rect 455201 177242 455225 177514
rect 454905 177218 455225 177242
rect 515362 177212 515386 177544
rect 515706 177538 515730 177544
rect 518241 177538 520957 180218
rect 515706 177218 520957 177538
rect 515706 177212 515730 177218
rect 515362 177188 515730 177212
rect 118982 175792 120252 176112
rect 120572 175792 121698 176112
rect 129057 176088 129377 176112
rect 129057 175816 129081 176088
rect 129353 175816 129377 176088
rect 129057 175792 129377 175816
rect 118982 172112 121698 175792
rect 515362 174544 515730 174568
rect 454905 174514 455225 174538
rect 454905 174242 454929 174514
rect 455201 174242 455225 174514
rect 454905 174218 455225 174242
rect 515362 174212 515386 174544
rect 515706 174538 515730 174544
rect 518241 174538 520957 177218
rect 515706 174218 520957 174538
rect 515706 174212 515730 174218
rect 515362 174188 515730 174212
rect 118982 171792 120252 172112
rect 120572 171792 121698 172112
rect 129057 172088 129377 172112
rect 129057 171816 129081 172088
rect 129353 171816 129377 172088
rect 129057 171792 129377 171816
rect 118982 168112 121698 171792
rect 515362 171544 515730 171568
rect 454905 171514 455225 171538
rect 454905 171242 454929 171514
rect 455201 171242 455225 171514
rect 454905 171218 455225 171242
rect 515362 171212 515386 171544
rect 515706 171538 515730 171544
rect 518241 171538 520957 174218
rect 515706 171218 520957 171538
rect 515706 171212 515730 171218
rect 515362 171188 515730 171212
rect 515362 168544 515730 168568
rect 454905 168514 455225 168538
rect 454905 168242 454929 168514
rect 455201 168242 455225 168514
rect 454905 168218 455225 168242
rect 515362 168212 515386 168544
rect 515706 168538 515730 168544
rect 518241 168538 520957 171218
rect 515706 168218 520957 168538
rect 515706 168212 515730 168218
rect 515362 168188 515730 168212
rect 118982 167792 120252 168112
rect 120572 167792 121698 168112
rect 129057 168088 129377 168112
rect 129057 167816 129081 168088
rect 129353 167816 129377 168088
rect 129057 167792 129377 167816
rect 118982 164112 121698 167792
rect 515362 165544 515730 165568
rect 454905 165514 455225 165538
rect 454905 165242 454929 165514
rect 455201 165242 455225 165514
rect 454905 165218 455225 165242
rect 515362 165212 515386 165544
rect 515706 165538 515730 165544
rect 518241 165538 520957 168218
rect 553276 167476 558076 180540
rect 515706 165218 520957 165538
rect 515706 165212 515730 165218
rect 515362 165188 515730 165212
rect 118982 163792 120252 164112
rect 120572 163792 121698 164112
rect 129057 164088 129377 164112
rect 129057 163816 129081 164088
rect 129353 163816 129377 164088
rect 129057 163792 129377 163816
rect 118982 160112 121698 163792
rect 515362 162544 515730 162568
rect 454905 162514 455225 162538
rect 454905 162242 454929 162514
rect 455201 162242 455225 162514
rect 454905 162218 455225 162242
rect 515362 162212 515386 162544
rect 515706 162538 515730 162544
rect 518241 162538 520957 165218
rect 550944 164186 571790 167476
rect 550944 162676 553300 164186
rect 515706 162218 520957 162538
rect 515706 162212 515730 162218
rect 515362 162188 515730 162212
rect 118982 159792 120252 160112
rect 120572 159792 121698 160112
rect 129057 160088 129377 160112
rect 129057 159816 129081 160088
rect 129353 159816 129377 160088
rect 129057 159792 129377 159816
rect 118982 156112 121698 159792
rect 515362 159544 515730 159568
rect 454905 159514 455225 159538
rect 454905 159242 454929 159514
rect 455201 159242 455225 159514
rect 454905 159218 455225 159242
rect 515362 159212 515386 159544
rect 515706 159538 515730 159544
rect 518241 159538 520957 162218
rect 515706 159218 520957 159538
rect 515706 159212 515730 159218
rect 515362 159188 515730 159212
rect 515362 156544 515730 156568
rect 454905 156514 455225 156538
rect 454905 156242 454929 156514
rect 455201 156242 455225 156514
rect 454905 156218 455225 156242
rect 515362 156212 515386 156544
rect 515706 156538 515730 156544
rect 518241 156538 520957 159218
rect 515706 156218 520957 156538
rect 515706 156212 515730 156218
rect 515362 156188 515730 156212
rect 118982 155792 120252 156112
rect 120572 155792 121698 156112
rect 129057 156088 129377 156112
rect 129057 155816 129081 156088
rect 129353 155816 129377 156088
rect 129057 155792 129377 155816
rect 118982 152112 121698 155792
rect 515362 153544 515730 153568
rect 454905 153514 455225 153538
rect 454905 153242 454929 153514
rect 455201 153242 455225 153514
rect 454905 153218 455225 153242
rect 515362 153212 515386 153544
rect 515706 153538 515730 153544
rect 518241 153538 520957 156218
rect 515706 153218 520957 153538
rect 515706 153212 515730 153218
rect 515362 153188 515730 153212
rect 118982 151792 120252 152112
rect 120572 151792 121698 152112
rect 129057 152088 129377 152112
rect 129057 151816 129081 152088
rect 129353 151816 129377 152088
rect 129057 151792 129377 151816
rect 118982 148112 121698 151792
rect 515362 150544 515730 150568
rect 454905 150514 455225 150538
rect 454905 150242 454929 150514
rect 455201 150242 455225 150514
rect 454905 150218 455225 150242
rect 515362 150212 515386 150544
rect 515706 150538 515730 150544
rect 518241 150538 520957 153218
rect 515706 150218 520957 150538
rect 515706 150212 515730 150218
rect 515362 150188 515730 150212
rect 118982 147792 120252 148112
rect 120572 147792 121698 148112
rect 129057 148088 129377 148112
rect 129057 147816 129081 148088
rect 129353 147816 129377 148088
rect 129057 147792 129377 147816
rect 118982 144112 121698 147792
rect 118982 143792 120252 144112
rect 120572 143792 121698 144112
rect 129057 144088 129377 144112
rect 129057 143816 129081 144088
rect 129353 143816 129377 144088
rect 129057 143792 129377 143816
rect 118982 140112 121698 143792
rect 518241 141320 520957 150218
rect 494530 141266 520957 141320
rect 494530 141242 507515 141266
rect 118982 139792 120252 140112
rect 120572 139792 121698 140112
rect 129057 140088 129377 140112
rect 129057 139816 129081 140088
rect 129353 139816 129377 140088
rect 129057 139792 129377 139816
rect 494530 139876 495525 141242
rect 496891 139876 507515 141242
rect 494530 139852 507515 139876
rect 510119 139852 520957 141266
rect 494530 139799 520957 139852
rect 118982 109188 121698 139792
rect 453395 134620 453715 134644
rect 453395 134348 453419 134620
rect 453691 134348 453715 134620
rect 453395 134324 453715 134348
rect 150296 115072 150616 115096
rect 150296 114800 150320 115072
rect 150592 114800 150616 115072
rect 150296 114776 150616 114800
rect 153296 115072 153616 115096
rect 153296 114800 153320 115072
rect 153592 114800 153616 115072
rect 153296 114776 153616 114800
rect 156296 115072 156616 115096
rect 156296 114800 156320 115072
rect 156592 114800 156616 115072
rect 156296 114776 156616 114800
rect 159296 115072 159616 115096
rect 159296 114800 159320 115072
rect 159592 114800 159616 115072
rect 159296 114776 159616 114800
rect 162296 115072 162616 115096
rect 162296 114800 162320 115072
rect 162592 114800 162616 115072
rect 162296 114776 162616 114800
rect 165296 115072 165616 115096
rect 165296 114800 165320 115072
rect 165592 114800 165616 115072
rect 165296 114776 165616 114800
rect 168296 115072 168616 115096
rect 168296 114800 168320 115072
rect 168592 114800 168616 115072
rect 168296 114776 168616 114800
rect 171296 115072 171616 115096
rect 171296 114800 171320 115072
rect 171592 114800 171616 115072
rect 171296 114776 171616 114800
rect 174296 115072 174616 115096
rect 174296 114800 174320 115072
rect 174592 114800 174616 115072
rect 174296 114776 174616 114800
rect 177296 115072 177616 115096
rect 177296 114800 177320 115072
rect 177592 114800 177616 115072
rect 177296 114776 177616 114800
rect 180296 115072 180616 115096
rect 180296 114800 180320 115072
rect 180592 114800 180616 115072
rect 180296 114776 180616 114800
rect 183296 115072 183616 115096
rect 183296 114800 183320 115072
rect 183592 114800 183616 115072
rect 183296 114776 183616 114800
rect 186296 115072 186616 115096
rect 186296 114800 186320 115072
rect 186592 114800 186616 115072
rect 186296 114776 186616 114800
rect 189296 115072 189616 115096
rect 189296 114800 189320 115072
rect 189592 114800 189616 115072
rect 189296 114776 189616 114800
rect 192296 115072 192616 115096
rect 192296 114800 192320 115072
rect 192592 114800 192616 115072
rect 192296 114776 192616 114800
rect 195296 115072 195616 115096
rect 195296 114800 195320 115072
rect 195592 114800 195616 115072
rect 195296 114776 195616 114800
rect 198296 115072 198616 115096
rect 198296 114800 198320 115072
rect 198592 114800 198616 115072
rect 198296 114776 198616 114800
rect 201296 115072 201616 115096
rect 201296 114800 201320 115072
rect 201592 114800 201616 115072
rect 201296 114776 201616 114800
rect 204296 115072 204616 115096
rect 204296 114800 204320 115072
rect 204592 114800 204616 115072
rect 204296 114776 204616 114800
rect 207296 115072 207616 115096
rect 207296 114800 207320 115072
rect 207592 114800 207616 115072
rect 207296 114776 207616 114800
rect 210296 115072 210616 115096
rect 210296 114800 210320 115072
rect 210592 114800 210616 115072
rect 210296 114776 210616 114800
rect 213296 115072 213616 115096
rect 213296 114800 213320 115072
rect 213592 114800 213616 115072
rect 213296 114776 213616 114800
rect 216296 115072 216616 115096
rect 216296 114800 216320 115072
rect 216592 114800 216616 115072
rect 216296 114776 216616 114800
rect 219296 115072 219616 115096
rect 219296 114800 219320 115072
rect 219592 114800 219616 115072
rect 219296 114776 219616 114800
rect 222296 115072 222616 115096
rect 222296 114800 222320 115072
rect 222592 114800 222616 115072
rect 222296 114776 222616 114800
rect 225296 115072 225616 115096
rect 225296 114800 225320 115072
rect 225592 114800 225616 115072
rect 225296 114776 225616 114800
rect 228296 115072 228616 115096
rect 228296 114800 228320 115072
rect 228592 114800 228616 115072
rect 228296 114776 228616 114800
rect 231296 115072 231616 115096
rect 231296 114800 231320 115072
rect 231592 114800 231616 115072
rect 231296 114776 231616 114800
rect 234296 115072 234616 115096
rect 234296 114800 234320 115072
rect 234592 114800 234616 115072
rect 234296 114776 234616 114800
rect 237296 115072 237616 115096
rect 237296 114800 237320 115072
rect 237592 114800 237616 115072
rect 237296 114776 237616 114800
rect 240296 115072 240616 115096
rect 240296 114800 240320 115072
rect 240592 114800 240616 115072
rect 240296 114776 240616 114800
rect 243296 115072 243616 115096
rect 243296 114800 243320 115072
rect 243592 114800 243616 115072
rect 243296 114776 243616 114800
rect 246296 115072 246616 115096
rect 246296 114800 246320 115072
rect 246592 114800 246616 115072
rect 246296 114776 246616 114800
rect 249296 115072 249616 115096
rect 249296 114800 249320 115072
rect 249592 114800 249616 115072
rect 249296 114776 249616 114800
rect 252296 115072 252616 115096
rect 252296 114800 252320 115072
rect 252592 114800 252616 115072
rect 252296 114776 252616 114800
rect 255296 115072 255616 115096
rect 255296 114800 255320 115072
rect 255592 114800 255616 115072
rect 255296 114776 255616 114800
rect 258296 115072 258616 115096
rect 258296 114800 258320 115072
rect 258592 114800 258616 115072
rect 258296 114776 258616 114800
rect 261296 115072 261616 115096
rect 261296 114800 261320 115072
rect 261592 114800 261616 115072
rect 261296 114776 261616 114800
rect 264296 115072 264616 115096
rect 264296 114800 264320 115072
rect 264592 114800 264616 115072
rect 264296 114776 264616 114800
rect 267296 115072 267616 115096
rect 267296 114800 267320 115072
rect 267592 114800 267616 115072
rect 267296 114776 267616 114800
rect 270296 115072 270616 115096
rect 270296 114800 270320 115072
rect 270592 114800 270616 115072
rect 270296 114776 270616 114800
rect 273296 115072 273616 115096
rect 273296 114800 273320 115072
rect 273592 114800 273616 115072
rect 273296 114776 273616 114800
rect 276296 115072 276616 115096
rect 276296 114800 276320 115072
rect 276592 114800 276616 115072
rect 276296 114776 276616 114800
rect 279296 115072 279616 115096
rect 279296 114800 279320 115072
rect 279592 114800 279616 115072
rect 279296 114776 279616 114800
rect 282296 115072 282616 115096
rect 282296 114800 282320 115072
rect 282592 114800 282616 115072
rect 282296 114776 282616 114800
rect 285296 115072 285616 115096
rect 285296 114800 285320 115072
rect 285592 114800 285616 115072
rect 285296 114776 285616 114800
rect 288296 115072 288616 115096
rect 288296 114800 288320 115072
rect 288592 114800 288616 115072
rect 288296 114776 288616 114800
rect 291296 115072 291616 115096
rect 291296 114800 291320 115072
rect 291592 114800 291616 115072
rect 291296 114776 291616 114800
rect 294296 115072 294616 115096
rect 294296 114800 294320 115072
rect 294592 114800 294616 115072
rect 294296 114776 294616 114800
rect 297296 115072 297616 115096
rect 297296 114800 297320 115072
rect 297592 114800 297616 115072
rect 297296 114776 297616 114800
rect 300296 115072 300616 115096
rect 300296 114800 300320 115072
rect 300592 114800 300616 115072
rect 300296 114776 300616 114800
rect 303296 115072 303616 115096
rect 303296 114800 303320 115072
rect 303592 114800 303616 115072
rect 303296 114776 303616 114800
rect 306296 115072 306616 115096
rect 306296 114800 306320 115072
rect 306592 114800 306616 115072
rect 306296 114776 306616 114800
rect 309296 115072 309616 115096
rect 309296 114800 309320 115072
rect 309592 114800 309616 115072
rect 309296 114776 309616 114800
rect 312296 115072 312616 115096
rect 312296 114800 312320 115072
rect 312592 114800 312616 115072
rect 312296 114776 312616 114800
rect 315296 115072 315616 115096
rect 315296 114800 315320 115072
rect 315592 114800 315616 115072
rect 315296 114776 315616 114800
rect 318296 115072 318616 115096
rect 318296 114800 318320 115072
rect 318592 114800 318616 115072
rect 318296 114776 318616 114800
rect 321296 115072 321616 115096
rect 321296 114800 321320 115072
rect 321592 114800 321616 115072
rect 321296 114776 321616 114800
rect 324296 115072 324616 115096
rect 324296 114800 324320 115072
rect 324592 114800 324616 115072
rect 324296 114776 324616 114800
rect 327296 115072 327616 115096
rect 327296 114800 327320 115072
rect 327592 114800 327616 115072
rect 327296 114776 327616 114800
rect 330296 115072 330616 115096
rect 330296 114800 330320 115072
rect 330592 114800 330616 115072
rect 330296 114776 330616 114800
rect 333296 115072 333616 115096
rect 333296 114800 333320 115072
rect 333592 114800 333616 115072
rect 333296 114776 333616 114800
rect 336296 115072 336616 115096
rect 336296 114800 336320 115072
rect 336592 114800 336616 115072
rect 336296 114776 336616 114800
rect 339296 115072 339616 115096
rect 339296 114800 339320 115072
rect 339592 114800 339616 115072
rect 339296 114776 339616 114800
rect 342296 115072 342616 115096
rect 342296 114800 342320 115072
rect 342592 114800 342616 115072
rect 342296 114776 342616 114800
rect 345296 115072 345616 115096
rect 345296 114800 345320 115072
rect 345592 114800 345616 115072
rect 345296 114776 345616 114800
rect 348296 115072 348616 115096
rect 348296 114800 348320 115072
rect 348592 114800 348616 115072
rect 348296 114776 348616 114800
rect 351296 115072 351616 115096
rect 351296 114800 351320 115072
rect 351592 114800 351616 115072
rect 351296 114776 351616 114800
rect 354296 115072 354616 115096
rect 354296 114800 354320 115072
rect 354592 114800 354616 115072
rect 354296 114776 354616 114800
rect 357296 115072 357616 115096
rect 357296 114800 357320 115072
rect 357592 114800 357616 115072
rect 357296 114776 357616 114800
rect 360296 115072 360616 115096
rect 360296 114800 360320 115072
rect 360592 114800 360616 115072
rect 360296 114776 360616 114800
rect 363296 115072 363616 115096
rect 363296 114800 363320 115072
rect 363592 114800 363616 115072
rect 363296 114776 363616 114800
rect 366296 115072 366616 115096
rect 366296 114800 366320 115072
rect 366592 114800 366616 115072
rect 366296 114776 366616 114800
rect 369296 115072 369616 115096
rect 369296 114800 369320 115072
rect 369592 114800 369616 115072
rect 369296 114776 369616 114800
rect 372296 115072 372616 115096
rect 372296 114800 372320 115072
rect 372592 114800 372616 115072
rect 372296 114776 372616 114800
rect 375296 115072 375616 115096
rect 375296 114800 375320 115072
rect 375592 114800 375616 115072
rect 375296 114776 375616 114800
rect 378296 115072 378616 115096
rect 378296 114800 378320 115072
rect 378592 114800 378616 115072
rect 378296 114776 378616 114800
rect 381296 115072 381616 115096
rect 381296 114800 381320 115072
rect 381592 114800 381616 115072
rect 381296 114776 381616 114800
rect 384296 115072 384616 115096
rect 384296 114800 384320 115072
rect 384592 114800 384616 115072
rect 384296 114776 384616 114800
rect 387296 115072 387616 115096
rect 387296 114800 387320 115072
rect 387592 114800 387616 115072
rect 387296 114776 387616 114800
rect 390296 115072 390616 115096
rect 390296 114800 390320 115072
rect 390592 114800 390616 115072
rect 390296 114776 390616 114800
rect 393296 115072 393616 115096
rect 393296 114800 393320 115072
rect 393592 114800 393616 115072
rect 393296 114776 393616 114800
rect 396296 115072 396616 115096
rect 396296 114800 396320 115072
rect 396592 114800 396616 115072
rect 396296 114776 396616 114800
rect 399296 115072 399616 115096
rect 399296 114800 399320 115072
rect 399592 114800 399616 115072
rect 399296 114776 399616 114800
rect 402296 115072 402616 115096
rect 402296 114800 402320 115072
rect 402592 114800 402616 115072
rect 402296 114776 402616 114800
rect 405296 115072 405616 115096
rect 405296 114800 405320 115072
rect 405592 114800 405616 115072
rect 405296 114776 405616 114800
rect 408296 115072 408616 115096
rect 408296 114800 408320 115072
rect 408592 114800 408616 115072
rect 408296 114776 408616 114800
rect 411296 115072 411616 115096
rect 411296 114800 411320 115072
rect 411592 114800 411616 115072
rect 411296 114776 411616 114800
rect 414296 115072 414616 115096
rect 414296 114800 414320 115072
rect 414592 114800 414616 115072
rect 414296 114776 414616 114800
rect 420296 115072 420616 115096
rect 420296 114800 420320 115072
rect 420592 114800 420616 115072
rect 420296 114776 420616 114800
rect 423296 115072 423616 115096
rect 423296 114800 423320 115072
rect 423592 114800 423616 115072
rect 423296 114776 423616 114800
rect 426296 115072 426616 115096
rect 426296 114800 426320 115072
rect 426592 114800 426616 115072
rect 426296 114776 426616 114800
rect 429296 115072 429616 115096
rect 429296 114800 429320 115072
rect 429592 114800 429616 115072
rect 429296 114776 429616 114800
rect 432296 115072 432616 115096
rect 432296 114800 432320 115072
rect 432592 114800 432616 115072
rect 432296 114776 432616 114800
rect 435296 115072 435616 115096
rect 435296 114800 435320 115072
rect 435592 114800 435616 115072
rect 435296 114776 435616 114800
rect 438296 115072 438616 115096
rect 438296 114800 438320 115072
rect 438592 114800 438616 115072
rect 438296 114776 438616 114800
rect 441296 115072 441616 115096
rect 441296 114800 441320 115072
rect 441592 114800 441616 115072
rect 441296 114776 441616 114800
rect 444296 115072 444616 115096
rect 444296 114800 444320 115072
rect 444592 114800 444616 115072
rect 444296 114776 444616 114800
rect 518241 109188 520957 139799
rect 553276 159434 553300 162676
rect 558052 162676 571790 164186
rect 558052 159434 558076 162676
rect 553276 127150 558076 159434
rect 553276 126465 557323 127150
rect 558008 126465 558076 127150
rect 118982 106472 525544 109188
rect 96516 95142 101386 95166
rect 96516 90342 96540 95142
rect 101340 92376 101386 95142
rect 553276 95118 558076 126465
rect 101340 90342 101364 92376
rect 553276 90366 553300 95118
rect 558052 90366 558076 95118
rect 553276 90342 558076 90366
rect 96516 90318 101364 90342
rect 424324 88506 428724 88906
rect 432124 88506 432724 88906
rect 488924 88506 489924 88906
rect 423524 87906 429724 88506
rect 431924 87906 433124 88506
rect 434524 87906 448124 88506
rect 422724 87506 430324 87906
rect 431524 87506 433124 87906
rect 434324 87506 448124 87906
rect 450124 87906 454924 88506
rect 450124 87506 455124 87906
rect 422324 86906 433124 87506
rect 434524 86906 448324 87506
rect 450124 86906 455324 87506
rect 461924 86906 467808 88506
rect 469706 87906 477924 88506
rect 469706 87506 478924 87906
rect 488924 87506 490124 88506
rect 469706 86906 479924 87506
rect 421724 86306 433124 86906
rect 435724 86306 448324 86906
rect 451324 86306 455524 86906
rect 463124 86306 467324 86906
rect 469724 86306 480324 86906
rect 488724 86306 490324 87506
rect 421524 85906 425324 86306
rect 428324 85906 433124 86306
rect 436124 85906 448324 86306
rect 451724 85906 455924 86306
rect 421124 85306 424924 85906
rect 428924 85306 433124 85906
rect 420724 84906 424124 85306
rect 429524 84906 433124 85306
rect 436324 84906 439524 85906
rect 445524 85306 448324 85906
rect 451924 85306 455924 85906
rect 463724 85906 466724 86306
rect 470524 85906 480524 86306
rect 463724 85306 466324 85906
rect 446524 84906 448324 85306
rect 452324 84906 456124 85306
rect 420524 84306 423924 84906
rect 429924 84306 433124 84906
rect 420324 83706 423524 84306
rect 430124 83706 433124 84306
rect 420124 83306 423124 83706
rect 430324 83306 433124 83706
rect 419924 82706 422924 83306
rect 430724 82706 433124 83306
rect 419524 82306 422724 82706
rect 430924 82306 433124 82706
rect 419324 81706 422524 82306
rect 419124 81106 422524 81706
rect 431124 81106 433124 82306
rect 419124 80706 422324 81106
rect 431324 80706 433124 81106
rect 418924 80106 421924 80706
rect 418724 79706 421924 80106
rect 431524 79706 433124 80706
rect 418724 79106 421724 79706
rect 418324 78106 421524 79106
rect 431924 78506 433124 79706
rect 418124 77506 421524 78106
rect 418124 76506 421324 77506
rect 432124 76906 433324 78506
rect 417924 75906 421324 76506
rect 432324 76506 433324 76906
rect 432324 75906 433124 76506
rect 417924 74906 421124 75906
rect 399524 72426 399924 74706
rect 399404 72106 399924 72426
rect 417724 72906 421124 74906
rect 399124 70506 399724 72106
rect 417724 71306 420724 72906
rect 398924 69226 399524 70506
rect 402324 69906 403524 70506
rect 401924 69820 403524 69906
rect 401924 69506 403724 69820
rect 398804 68906 399524 69226
rect 401524 68906 402324 69506
rect 184686 64156 190686 66356
rect 223686 65756 224286 66356
rect 184686 60556 185686 64156
rect 184686 59556 185486 60556
rect 187486 51756 188086 64156
rect 190086 59556 190686 64156
rect 194286 62156 196086 62556
rect 200646 62156 201086 62196
rect 202286 62156 203886 62556
rect 208686 62156 209686 62556
rect 211086 62156 212286 62556
rect 216686 62156 218686 62556
rect 223486 62156 224286 65756
rect 238086 65156 240686 67356
rect 246486 65756 249086 66356
rect 249486 65756 250086 66356
rect 315198 65900 317598 66300
rect 318798 65900 321198 66300
rect 359598 65900 361398 66300
rect 245886 65156 250286 65756
rect 231886 62156 233486 62556
rect 193886 61556 196686 62156
rect 199086 61876 201086 62156
rect 193486 61156 197286 61556
rect 199086 61156 200966 61876
rect 201486 61556 204486 62156
rect 206686 61556 207966 62156
rect 208286 61556 210286 62156
rect 210686 61556 212886 62156
rect 216286 61556 219086 62156
rect 201286 61156 204886 61556
rect 193086 60556 197486 61156
rect 199086 60556 205086 61156
rect 206286 60556 213086 61556
rect 215686 61156 219486 61556
rect 215486 60556 219886 61156
rect 222286 60556 227486 62156
rect 230886 61556 233886 62156
rect 230286 61156 234486 61556
rect 230286 60556 234686 61156
rect 192886 59956 194686 60556
rect 195886 59956 197686 60556
rect 199486 59956 202486 60556
rect 203686 59956 205486 60556
rect 206686 59956 209086 60556
rect 209486 59956 211486 60556
rect 212086 59956 213286 60556
rect 215286 59956 216886 60556
rect 218286 59956 220086 60556
rect 222486 59956 227286 60556
rect 230286 59956 231886 60556
rect 233286 59956 234686 60556
rect 192686 59556 194086 59956
rect 196286 59556 197886 59956
rect 192686 58956 193886 59556
rect 196686 58956 197886 59556
rect 200086 59556 202086 59956
rect 204286 59556 205686 59956
rect 200086 58956 201886 59556
rect 204486 58956 205686 59556
rect 207086 59556 208486 59956
rect 209686 59556 211086 59956
rect 192486 58556 193686 58956
rect 192486 57956 193486 58556
rect 197086 57956 198286 58956
rect 192286 57356 193486 57956
rect 192286 54756 193086 57356
rect 197286 56956 198286 57956
rect 200086 58556 201486 58956
rect 204686 58556 205886 58956
rect 200086 57956 201286 58556
rect 197286 56356 198486 56956
rect 197486 55356 198486 56356
rect 192286 54356 193486 54756
rect 192486 53756 193486 54356
rect 197286 53756 198286 55356
rect 192486 52756 193686 53756
rect 197086 53156 198286 53756
rect 200086 54756 201086 57956
rect 204886 56956 205886 58556
rect 205086 56356 205886 56956
rect 207086 58556 208286 59556
rect 209686 58556 210886 59556
rect 205086 55756 206086 56356
rect 200086 54356 201286 54756
rect 204886 54356 205886 55756
rect 200086 53156 201486 54356
rect 204686 53756 205886 54356
rect 204486 53156 205686 53756
rect 196686 52756 197886 53156
rect 192686 52156 194086 52756
rect 196486 52156 197886 52756
rect 200086 52756 202086 53156
rect 204286 52756 205686 53156
rect 200086 52156 202286 52756
rect 203686 52156 205486 52756
rect 192886 51756 194286 52156
rect 196086 51756 197686 52156
rect 200086 51756 205086 52156
rect 207086 51756 208086 58556
rect 209686 51756 210686 58556
rect 212286 51756 213286 59956
rect 215086 59556 216486 59956
rect 218886 59556 220286 59956
rect 214686 58956 216286 59556
rect 219086 58956 220286 59556
rect 214686 58556 215886 58956
rect 219286 58556 220486 58956
rect 214686 57956 215686 58556
rect 214486 57356 215686 57956
rect 219486 57356 220486 58556
rect 214486 55356 220686 57356
rect 214486 54356 215686 55356
rect 214686 53756 215686 54356
rect 214686 53156 215886 53756
rect 215086 52756 216286 53156
rect 220086 52756 220486 53156
rect 223486 52756 224286 59956
rect 230286 59556 230886 59956
rect 233686 59556 234886 59956
rect 232086 57356 233486 57956
rect 233886 57356 234886 59556
rect 230886 56956 234886 57356
rect 230286 56356 234886 56956
rect 230086 55756 234886 56356
rect 229886 55356 231886 55756
rect 233486 55356 234886 55756
rect 229886 54756 231286 55356
rect 229686 54356 230886 54756
rect 229686 52756 230686 54356
rect 233886 53156 234886 55356
rect 233486 52756 234886 53156
rect 215086 52156 216486 52756
rect 219486 52156 220686 52756
rect 223486 52156 224686 52756
rect 227486 52156 228286 52756
rect 229686 52156 230886 52756
rect 233286 52156 234886 52756
rect 215286 51756 216886 52156
rect 219086 51756 220686 52156
rect 223686 51756 224886 52156
rect 227086 51756 228286 52156
rect 185686 50156 189886 51756
rect 192886 51156 197486 51756
rect 193086 50556 197286 51156
rect 200086 50836 200966 51756
rect 201286 51156 204886 51756
rect 193686 50156 197086 50556
rect 194086 49556 196486 50156
rect 200086 46556 201086 50836
rect 201486 50556 204686 51156
rect 202086 50156 203886 50556
rect 206286 50156 208686 51756
rect 209686 50156 211486 51756
rect 212286 50156 214086 51756
rect 215486 51156 220486 51756
rect 223686 51156 228286 51756
rect 229886 51756 231086 52156
rect 232686 51756 234886 52156
rect 239686 51756 240686 65156
rect 245686 64756 250286 65156
rect 245486 64156 247486 64756
rect 248086 64156 250286 64756
rect 315198 64700 317798 65900
rect 318798 64700 321398 65900
rect 359598 65300 361598 65900
rect 315398 64300 317598 64700
rect 318798 64300 321198 64700
rect 359598 64300 361998 65300
rect 363598 64700 366398 66300
rect 363798 64300 366398 64700
rect 369798 64300 370998 67900
rect 398924 66906 399244 68906
rect 401124 68306 402124 68906
rect 400924 67906 401524 68306
rect 400724 67626 401324 67906
rect 403324 67626 403724 69506
rect 417524 68106 420724 71306
rect 400604 67306 401324 67626
rect 403204 67306 403724 67626
rect 400124 66906 400924 67306
rect 398924 66306 400724 66906
rect 399124 65706 400124 66306
rect 403124 65706 403524 67306
rect 402724 65306 403524 65706
rect 417724 66106 420724 68106
rect 436724 72306 439524 84906
rect 446724 84306 448324 84906
rect 446924 82706 448324 84306
rect 447124 81706 448324 82706
rect 447524 80106 448324 81706
rect 452524 84306 456324 84906
rect 463924 84306 466124 85306
rect 470724 84306 473924 85906
rect 476524 85306 481124 85906
rect 477524 84906 481524 85306
rect 488524 84906 490724 86306
rect 477924 84306 481524 84906
rect 452524 83706 456524 84306
rect 464324 83706 466124 84306
rect 452524 83306 456724 83706
rect 452524 82306 457124 83306
rect 452524 81706 457324 82306
rect 452524 81106 457524 81706
rect 452524 80706 457724 81106
rect 452524 80106 457924 80706
rect 452524 79386 453804 80106
rect 454124 79706 457924 80106
rect 445924 75906 446924 77506
rect 445724 74306 446924 75906
rect 452524 74906 453924 79386
rect 454324 79106 458324 79706
rect 454724 78506 458524 79106
rect 454924 78106 458724 78506
rect 454924 77506 458924 78106
rect 455124 76906 458924 77506
rect 455324 76506 459124 76906
rect 455524 75906 459524 76506
rect 455924 75506 459724 75906
rect 445524 73306 446924 74306
rect 445324 72906 446924 73306
rect 445124 72306 446924 72906
rect 436724 69706 446924 72306
rect 402724 64306 403324 65306
rect 406124 64706 406924 65306
rect 405724 64306 407324 64706
rect 417724 64506 421124 66106
rect 245486 63756 246686 64156
rect 248686 63756 250286 64156
rect 245286 63156 246486 63756
rect 245286 60556 246286 63156
rect 249086 62556 250286 63756
rect 249286 61156 250286 62556
rect 254086 62156 256086 62556
rect 253686 61556 256486 62156
rect 253086 61156 257086 61556
rect 252886 60556 257286 61156
rect 245286 59956 246486 60556
rect 252686 59956 254286 60556
rect 255886 59956 257486 60556
rect 245486 59556 246886 59956
rect 252486 59556 253886 59956
rect 256286 59556 257686 59956
rect 245486 58956 247886 59556
rect 252286 58956 253686 59556
rect 256486 58956 257686 59556
rect 315798 59500 316598 64300
rect 319598 59500 320598 64300
rect 360398 63100 362198 64300
rect 324798 62100 326398 62700
rect 334598 62100 335198 62700
rect 341998 62100 342798 62700
rect 360398 62100 362398 63100
rect 323798 61700 326798 62100
rect 330798 61700 332598 62100
rect 333798 61700 335998 62100
rect 338198 61700 339998 62100
rect 341198 61700 343398 62100
rect 323198 61100 327398 61700
rect 323198 60500 327598 61100
rect 330398 60500 332598 61700
rect 333598 61100 336198 61700
rect 333198 60500 336398 61100
rect 337998 60500 339998 61700
rect 340998 61100 343598 61700
rect 340598 60500 343998 61100
rect 323198 60100 324798 60500
rect 326198 60100 327598 60500
rect 330798 60100 332598 60500
rect 332918 60100 334678 60500
rect 334998 60100 336398 60500
rect 338198 60100 339998 60500
rect 340398 60100 342198 60500
rect 342518 60100 343998 60500
rect 345198 60500 347598 62100
rect 349198 60500 351598 62100
rect 345198 60100 347198 60500
rect 349398 60100 351598 60500
rect 360398 61700 362598 62100
rect 360398 60180 361278 61700
rect 361598 60500 362798 61700
rect 323198 59500 323798 60100
rect 326598 59500 327798 60100
rect 245686 58556 249086 58956
rect 252286 58556 253486 58956
rect 256686 58556 257886 58956
rect 246286 57956 249486 58556
rect 252286 57956 253086 58556
rect 246886 57356 250086 57956
rect 251886 57356 253086 57956
rect 257086 57356 257886 58556
rect 315798 57500 320598 59500
rect 324998 57500 326398 57900
rect 326798 57500 327798 59500
rect 247886 56956 250286 57356
rect 248886 56356 250286 56956
rect 249286 55756 250486 56356
rect 245086 54356 245686 55356
rect 245086 53156 245886 54356
rect 249486 53156 250486 55756
rect 251886 55356 258286 57356
rect 251886 54356 253086 55356
rect 252286 53756 253086 54356
rect 252286 53156 253486 53756
rect 245086 52756 246286 53156
rect 249286 52756 250486 53156
rect 252486 52756 253686 53156
rect 257486 52756 257886 53156
rect 245086 52156 246486 52756
rect 249086 52156 250286 52756
rect 252486 52156 253886 52756
rect 257086 52156 258286 52756
rect 245086 51756 246686 52156
rect 248686 51756 250286 52156
rect 252686 51756 254286 52156
rect 256486 51756 258286 52156
rect 229886 51156 235886 51756
rect 237486 51156 242886 51756
rect 245086 51156 247686 51756
rect 248006 51156 250086 51756
rect 252886 51156 257886 51756
rect 315798 51700 316598 57500
rect 319598 51700 320598 57500
rect 323798 56900 327798 57500
rect 323198 56500 327798 56900
rect 322998 55900 327798 56500
rect 322798 55300 324798 55900
rect 326398 55300 327798 55900
rect 322798 54900 324198 55300
rect 322598 54300 323798 54900
rect 322598 52700 323598 54300
rect 326798 53300 327798 55300
rect 326398 52700 327798 53300
rect 322598 52300 323798 52700
rect 326198 52300 327798 52700
rect 322798 51700 323998 52300
rect 325598 51700 327798 52300
rect 331998 59500 334398 60100
rect 335598 59500 336198 60100
rect 339398 59500 341798 60100
rect 342998 59500 343598 60100
rect 345598 59500 346798 60100
rect 331998 59100 333798 59500
rect 339398 59100 341198 59500
rect 345798 59100 346798 59500
rect 349998 59500 351198 60100
rect 349998 59100 350798 59500
rect 331998 58500 333598 59100
rect 339398 58500 340998 59100
rect 345798 58500 346998 59100
rect 331998 57900 333398 58500
rect 339398 57900 340798 58500
rect 345998 57900 346998 58500
rect 349598 58500 350798 59100
rect 349598 57900 350598 58500
rect 331998 57500 333198 57900
rect 339398 57500 340598 57900
rect 345998 57500 347198 57900
rect 331998 51700 332598 57500
rect 339398 51700 339998 57500
rect 346398 56900 347198 57500
rect 349398 57500 350598 57900
rect 349398 56900 350398 57500
rect 346398 56500 347598 56900
rect 346598 55900 347598 56500
rect 349198 56500 350398 56900
rect 349198 55900 350198 56500
rect 346598 55300 347798 55900
rect 346798 54900 347798 55300
rect 348998 55300 350198 55900
rect 348998 54900 349998 55300
rect 346798 54300 347998 54900
rect 346998 53900 347998 54300
rect 348798 54300 349998 54900
rect 348798 53900 349598 54300
rect 346998 53300 348198 53900
rect 347198 52700 348198 53300
rect 348518 53300 349598 53900
rect 348518 52700 349398 53300
rect 347198 52300 349398 52700
rect 215686 50556 220286 51156
rect 223886 50556 228286 51156
rect 230086 50556 235886 51156
rect 237286 50556 243086 51156
rect 215886 50156 220086 50556
rect 223886 50156 227686 50556
rect 230286 50156 233566 50556
rect 233886 50156 235886 50556
rect 237486 50156 243086 50556
rect 245086 50556 249886 51156
rect 253086 50556 257686 51156
rect 314798 51100 317598 51700
rect 318798 51100 321398 51700
rect 322798 51100 328798 51700
rect 245086 50156 245566 50556
rect 245886 50156 249486 50556
rect 253486 50156 257486 50556
rect 216486 49556 219286 50156
rect 224286 49556 227086 50156
rect 230686 49556 233086 50156
rect 246486 49556 249086 50156
rect 253886 49556 256686 50156
rect 314798 50100 317798 51100
rect 318798 50100 321598 51100
rect 322998 50700 328798 51100
rect 323198 50100 326598 50700
rect 326918 50100 328798 50700
rect 330198 50100 335198 51700
rect 337598 50100 342798 51700
rect 347598 51100 349198 52300
rect 360398 51700 361398 60180
rect 361998 60100 363198 60500
rect 362198 59500 363198 60100
rect 362198 59100 363398 59500
rect 362398 57900 363598 59100
rect 362598 57500 363798 57900
rect 362798 56900 363798 57500
rect 362798 56500 363998 56900
rect 363198 55300 364398 56500
rect 363398 54900 364478 55300
rect 363598 54300 364478 54900
rect 364798 54300 365798 64300
rect 402524 63706 403324 64306
rect 405524 63706 407524 64306
rect 368398 60100 370998 62100
rect 402524 61106 403124 63706
rect 404924 63106 406324 63706
rect 406724 63106 407524 63706
rect 404724 62706 405924 63106
rect 404524 62106 405524 62706
rect 406924 62106 407524 63106
rect 417924 63506 421124 64506
rect 417924 62906 421324 63506
rect 403924 61706 405124 62106
rect 403724 61106 404924 61706
rect 406724 61106 407524 62106
rect 418124 61906 421324 62906
rect 418124 61306 421524 61906
rect 402524 60506 404524 61106
rect 402724 60106 403924 60506
rect 406724 60106 407324 61106
rect 418324 60906 421524 61306
rect 418324 60306 421724 60906
rect 363598 53900 365798 54300
rect 363798 52700 365798 53900
rect 363998 51700 365798 52700
rect 369998 51700 370998 60100
rect 403124 59506 403524 60106
rect 406324 58906 407124 60106
rect 418724 59706 421724 60306
rect 409524 58906 410924 59506
rect 418724 59306 421924 59706
rect 406124 57506 407124 58906
rect 409324 58506 411124 58906
rect 418924 58706 422324 59306
rect 408724 57906 411124 58506
rect 419124 58306 422324 58706
rect 432524 58306 433324 58706
rect 408524 57506 411524 57906
rect 419124 57706 422524 58306
rect 432324 57706 433524 58306
rect 406124 55906 406924 57506
rect 408324 56906 409724 57506
rect 407924 56306 409524 56906
rect 410524 56306 411524 57506
rect 419324 57106 422724 57706
rect 432124 57106 433524 57706
rect 419524 56706 422924 57106
rect 431924 56706 433324 57106
rect 407524 55906 409124 56306
rect 410324 55906 411524 56306
rect 419924 56106 423124 56706
rect 431324 56106 433124 56706
rect 406124 55306 408724 55906
rect 406124 54906 408324 55306
rect 410324 54906 411124 55906
rect 419924 55706 423524 56106
rect 431124 55706 432724 56106
rect 420124 55106 423924 55706
rect 430724 55106 432524 55706
rect 406124 54306 408124 54906
rect 406724 53706 407524 54306
rect 409924 53706 411124 54906
rect 420324 54506 424124 55106
rect 430124 54506 432324 55106
rect 436724 54506 439524 69706
rect 444124 69106 446924 69706
rect 445124 68706 446924 69106
rect 445324 68106 446924 68706
rect 445524 67106 446924 68106
rect 445724 65506 446924 67106
rect 445924 64506 446924 65506
rect 445924 63906 446724 64506
rect 448924 60906 449524 61306
rect 448724 60306 449524 60906
rect 448324 59306 449524 60306
rect 448124 58706 449524 59306
rect 448124 58306 449324 58706
rect 452724 58306 453924 74906
rect 456124 74306 459924 75506
rect 456324 73906 460124 74306
rect 456524 73306 460324 73906
rect 456724 72906 460724 73306
rect 457124 72306 460724 72906
rect 457124 71706 460924 72306
rect 457324 71306 461124 71706
rect 457524 70706 461324 71306
rect 457724 70306 461524 70706
rect 457924 69106 461924 70306
rect 458324 68706 462124 69106
rect 458524 68106 462324 68706
rect 458724 67706 462524 68106
rect 458924 66506 462724 67706
rect 459124 66106 463124 66506
rect 459524 65506 463324 66106
rect 459724 64906 463324 65506
rect 459924 64506 463524 64906
rect 464324 64506 465924 83706
rect 470924 71706 473924 84306
rect 478124 83706 481724 84306
rect 488324 83706 490924 84906
rect 478324 83306 481924 83706
rect 478724 82706 482324 83306
rect 487924 82706 491124 83706
rect 478924 82306 482324 82706
rect 479124 80706 482524 82306
rect 487724 81106 491324 82706
rect 479324 75506 482724 80706
rect 487524 80106 491524 81106
rect 487324 79106 488604 80106
rect 488924 79106 491924 80106
rect 487324 78506 488524 79106
rect 487124 78106 488524 78506
rect 489124 78106 492124 79106
rect 487124 77506 488324 78106
rect 486724 76506 488324 77506
rect 489524 77506 492124 78106
rect 489524 76506 492324 77506
rect 486524 75506 487924 76506
rect 489724 75506 492524 76506
rect 479324 74906 482524 75506
rect 479124 73906 482524 74906
rect 486324 74906 487924 75506
rect 486324 73906 487724 74906
rect 489924 74306 492724 75506
rect 489924 73906 493124 74306
rect 478924 72906 482324 73906
rect 486124 72906 487524 73906
rect 490124 72906 493124 73906
rect 478724 72306 481924 72906
rect 485924 72306 487524 72906
rect 478324 71706 481724 72306
rect 470924 70306 473524 71706
rect 478124 71306 481524 71706
rect 485924 71306 487324 72306
rect 490324 71706 493324 72906
rect 477724 70706 481324 71306
rect 476924 70306 481124 70706
rect 485524 70306 487124 71306
rect 490724 70706 493524 71706
rect 490724 70306 493724 70706
rect 470924 69706 474524 70306
rect 475124 69706 480524 70306
rect 485324 69706 487124 70306
rect 490924 69706 493724 70306
rect 470924 69106 480124 69706
rect 485324 69106 486724 69706
rect 490924 69106 493924 69706
rect 470924 68706 479924 69106
rect 485124 68706 486724 69106
rect 470924 68106 479124 68706
rect 470924 67706 478124 68106
rect 485124 67706 486524 68706
rect 491124 68106 493924 69106
rect 470924 67106 473924 67706
rect 470924 66106 473524 67106
rect 484924 66506 486324 67706
rect 491324 67106 494324 68106
rect 491324 66506 494524 67106
rect 484724 66106 486324 66506
rect 491524 66106 494524 66506
rect 459924 63906 463724 64506
rect 460124 63506 463724 63906
rect 460324 62906 463924 63506
rect 464324 62906 465724 64506
rect 460724 62306 465724 62906
rect 460924 61906 465724 62306
rect 461124 60906 465724 61906
rect 461324 60306 465724 60906
rect 461524 59706 465724 60306
rect 461924 58706 465724 59706
rect 462124 58306 465724 58706
rect 447924 57706 449324 58306
rect 447724 57106 449324 57706
rect 447724 56706 449124 57106
rect 447524 56106 449124 56706
rect 447124 55706 449124 56106
rect 446724 55106 449124 55706
rect 452524 55106 454124 58306
rect 462324 57706 465724 58306
rect 462524 57106 465724 57706
rect 462724 56706 465724 57106
rect 463124 55706 465724 56706
rect 470924 55706 473924 66106
rect 484724 65506 494724 66106
rect 484324 64906 494724 65506
rect 484324 63906 494924 64906
rect 484124 63506 494924 63906
rect 484124 62906 485524 63506
rect 483924 61906 485524 62906
rect 492124 62306 495124 63506
rect 483724 60306 485324 61906
rect 492324 61306 495524 62306
rect 492524 60906 495524 61306
rect 483524 59306 485124 60306
rect 492524 59706 495724 60906
rect 483124 58706 485124 59306
rect 492724 58706 495924 59706
rect 483124 58306 484924 58706
rect 482924 57706 484924 58306
rect 493124 57706 496124 58706
rect 482924 57106 484724 57706
rect 482724 56706 484724 57106
rect 482724 56106 484324 56706
rect 493324 56106 496324 57706
rect 463324 55106 465724 55706
rect 446324 54506 448924 55106
rect 413524 53706 414524 54306
rect 420724 54106 424724 54506
rect 429724 54106 432124 54506
rect 436324 54106 439724 54506
rect 445324 54106 448924 54506
rect 452324 54106 454324 55106
rect 463524 54506 465724 55106
rect 463724 54106 465724 54506
rect 470724 54506 473924 55706
rect 482524 55106 484324 56106
rect 470724 54106 474124 54506
rect 482324 54106 484324 55106
rect 409924 53306 410924 53706
rect 413124 53306 414724 53706
rect 421124 53506 425524 54106
rect 428724 53506 431524 54106
rect 436124 53506 448924 54106
rect 451924 53506 454724 54106
rect 409724 52306 410924 53306
rect 412724 52706 415124 53306
rect 421324 52906 431324 53506
rect 435924 52906 448724 53506
rect 451524 52906 455124 53506
rect 463924 52906 465724 54106
rect 470524 53506 474124 54106
rect 481924 53506 484324 54106
rect 493524 55106 496724 56106
rect 493524 54506 496924 55106
rect 493524 53506 497124 54506
rect 470324 52906 474524 53506
rect 481524 52906 484724 53506
rect 493324 52906 497524 53506
rect 412324 52306 415124 52706
rect 421724 52506 430924 52906
rect 434524 52506 448724 52906
rect 450324 52506 456324 52906
rect 464324 52506 465724 52906
rect 347798 50700 349198 51100
rect 323598 49700 325998 50100
rect 347798 49700 348998 50700
rect 359798 50100 362598 51700
rect 364398 51100 365798 51700
rect 364598 50100 365798 51100
rect 367998 50100 373398 51700
rect 409724 51106 410724 52306
rect 412124 51706 415324 52306
rect 422324 51906 430324 52506
rect 434324 51906 448724 52506
rect 411724 51106 413524 51706
rect 409524 51026 410724 51106
rect 409524 50106 410604 51026
rect 411524 50706 413324 51106
rect 414124 50706 415324 51706
rect 422724 51506 429924 51906
rect 434524 51506 448724 51906
rect 450124 51506 456324 52506
rect 464524 51906 465724 52506
rect 464724 51506 465724 51906
rect 468724 52506 475924 52906
rect 480724 52506 485924 52906
rect 491924 52506 498324 52906
rect 468724 51506 476324 52506
rect 480524 51506 486124 52506
rect 491924 51506 498524 52506
rect 423524 50906 429124 51506
rect 410924 50106 412924 50706
rect 413924 50106 415324 50706
rect 424724 50306 428324 50906
rect 464924 50306 465724 51506
rect 409524 49706 412724 50106
rect 347598 48500 348798 49700
rect 409724 49106 412324 49706
rect 413924 49106 415124 50106
rect 409724 48506 411924 49106
rect 413524 48506 415124 49106
rect 347198 47500 348398 48500
rect 409924 48106 411524 48506
rect 413524 47506 414724 48506
rect 347198 47100 348198 47500
rect 199086 44956 202486 46556
rect 346998 46500 348198 47100
rect 413324 46506 414724 47506
rect 501724 48106 502124 48506
rect 501724 47506 502724 48106
rect 501724 46906 503324 47506
rect 501924 46506 503924 46906
rect 345198 45900 348998 46500
rect 345198 45500 349198 45900
rect 345198 44900 348998 45500
rect 413324 44906 414524 46506
rect 501924 45906 504324 46506
rect 502124 45506 505124 45906
rect 502124 44906 505524 45506
rect 413324 44306 505924 44906
rect 413324 43906 506524 44306
rect 413124 43306 506324 43906
rect 412724 42906 505724 43306
rect 412324 42306 414124 42906
rect 502124 42306 505124 42906
rect 412124 41706 413924 42306
rect 501924 41706 504524 42306
rect 411924 41306 413524 41706
rect 501924 41306 503924 41706
rect 411524 40706 413124 41306
rect 501724 40706 503324 41306
rect 411124 40306 412924 40706
rect 501724 40306 502924 40706
rect 235886 39756 236886 40156
rect 182686 38156 185286 38556
rect 185686 38156 186486 38556
rect 182286 37556 186486 38156
rect 196686 37556 199486 39756
rect 235086 39156 237486 39756
rect 234886 38556 237886 39156
rect 234686 38156 238086 38556
rect 247686 38156 249486 39756
rect 255286 39156 257086 39756
rect 255086 38156 257086 39156
rect 234486 37556 235886 38156
rect 236686 37556 238286 38156
rect 247886 37556 249486 38156
rect 255286 37556 257086 38156
rect 296198 38100 300198 38700
rect 181886 37156 186486 37556
rect 181686 36556 183486 37156
rect 184286 36556 186486 37156
rect 181686 35956 183086 36556
rect 185086 35956 186486 36556
rect 181486 34956 182686 35956
rect 185286 35556 186486 35956
rect 181486 33356 182286 34956
rect 185486 33956 186486 35556
rect 190486 34556 192286 34956
rect 189886 33956 192886 34556
rect 185686 33356 186486 33956
rect 189286 33356 193086 33956
rect 181486 32956 182686 33356
rect 189086 32956 193686 33356
rect 181486 32356 182886 32956
rect 188886 32356 190686 32956
rect 191886 32356 193886 32956
rect 181686 31756 183086 32356
rect 188886 31756 190286 32356
rect 192486 31756 193886 32356
rect 181886 31356 184086 31756
rect 181886 30756 185286 31356
rect 188686 30756 189886 31756
rect 192886 30756 194086 31756
rect 182286 30356 185886 30756
rect 188286 30356 189486 30756
rect 193086 30356 194286 30756
rect 183086 29756 186286 30356
rect 188286 29756 189286 30356
rect 193486 29756 194286 30356
rect 184286 29156 186486 29756
rect 185086 28756 186486 29156
rect 185486 28156 186686 28756
rect 181086 27156 181886 27756
rect 181086 25556 182086 27156
rect 185686 25556 186686 28156
rect 188286 27756 194286 29756
rect 188286 26556 189286 27756
rect 188286 26156 189486 26556
rect 181086 25156 182286 25556
rect 185486 25156 186686 25556
rect 188686 25156 189886 26156
rect 193686 25156 194086 25556
rect 181086 24556 182686 25156
rect 185286 24556 186686 25156
rect 188886 24556 190286 25156
rect 193486 24556 194286 25156
rect 181086 23956 183086 24556
rect 185086 23956 186486 24556
rect 188886 23956 190486 24556
rect 192686 23956 194286 24556
rect 198486 23956 199486 37556
rect 234286 37156 235686 37556
rect 237086 37156 238486 37556
rect 234286 36556 235486 37156
rect 237286 36556 238486 37156
rect 234286 35956 235086 36556
rect 233886 34956 235086 35956
rect 237486 35956 238486 36556
rect 237486 35556 238686 35956
rect 205486 34556 207086 34956
rect 213286 34556 215086 34956
rect 220486 34556 221886 34956
rect 204686 33956 207886 34556
rect 210886 33956 212286 34556
rect 212886 33956 215486 34556
rect 219486 33956 222686 34556
rect 204486 33356 208286 33956
rect 210686 33356 212286 33956
rect 212686 33356 215686 33956
rect 219086 33356 223086 33956
rect 203886 32956 208486 33356
rect 210686 32956 215886 33356
rect 218886 32956 223086 33356
rect 233886 32956 234886 34956
rect 237886 34556 238686 35556
rect 237886 33956 239086 34556
rect 240486 33956 243286 34556
rect 203886 32356 205686 32956
rect 207086 32356 208686 32956
rect 210886 32356 213486 32956
rect 214686 32356 216286 32956
rect 218886 32356 220486 32956
rect 221886 32356 223486 32956
rect 203686 31756 205086 32356
rect 207286 31756 209086 32356
rect 203486 31356 204886 31756
rect 207886 31356 209086 31756
rect 211686 31756 213286 32356
rect 215086 31756 216286 32356
rect 219086 31756 219486 32356
rect 222486 31756 223486 32356
rect 203486 30756 204686 31356
rect 203286 29756 204486 30756
rect 208086 30356 209286 31356
rect 208286 29756 209286 30356
rect 203286 27756 209286 29756
rect 211686 30756 212886 31756
rect 215286 31356 216286 31756
rect 215286 30756 216486 31356
rect 211686 30356 212686 30756
rect 203286 27156 204286 27756
rect 203286 26156 204486 27156
rect 203486 25556 204686 26156
rect 203486 25156 204886 25556
rect 208686 25156 209286 25556
rect 203686 24556 205086 25156
rect 208286 24556 209286 25156
rect 203886 23956 205686 24556
rect 207886 23956 209286 24556
rect 211686 23956 212286 30356
rect 215486 23956 216486 30756
rect 220686 29756 221886 30356
rect 222686 29756 223686 31756
rect 219486 29156 223686 29756
rect 219086 28756 223686 29156
rect 218886 28156 223686 28756
rect 218686 27756 220486 28156
rect 222286 27756 223686 28156
rect 218686 27156 220086 27756
rect 218286 26556 219486 27156
rect 218286 24556 219286 26556
rect 222686 26156 223686 27756
rect 233886 28156 234686 32956
rect 233886 26556 234886 28156
rect 238086 27756 239086 33956
rect 240286 32956 243286 33956
rect 244486 32956 247486 34556
rect 248686 33356 249486 37556
rect 250686 34556 252486 34956
rect 250286 33956 253086 34556
rect 249886 33356 253486 33956
rect 256286 33356 257086 37556
rect 295998 37700 300998 38100
rect 295998 37100 301398 37700
rect 296198 36500 301598 37100
rect 328598 36500 329798 40300
rect 366198 39700 367198 40300
rect 381398 39700 382398 40300
rect 388798 39700 389798 40300
rect 410924 39706 412724 40306
rect 501724 39706 502124 40306
rect 365198 39100 367998 39700
rect 372198 39100 376398 39700
rect 380598 39100 382998 39700
rect 387998 39100 390398 39700
rect 410524 39106 412324 39706
rect 361398 38700 361838 38740
rect 364998 38700 368398 39100
rect 350598 38100 353198 38700
rect 350198 37700 353678 38100
rect 353998 37700 354798 38700
rect 357998 38100 360798 38700
rect 361398 38420 362198 38700
rect 361518 38100 362198 38420
rect 364798 38100 368598 38700
rect 372198 38100 376598 39100
rect 380398 38700 383198 39100
rect 387798 38700 390998 39100
rect 410324 38706 411924 39106
rect 380198 38100 383598 38700
rect 387598 38100 391198 38700
rect 409924 38106 411724 38706
rect 357598 37700 361198 38100
rect 361518 37700 362398 38100
rect 364598 37700 366198 38100
rect 367198 37700 368798 38100
rect 349998 37100 354798 37700
rect 357398 37100 362398 37700
rect 349598 36500 351598 37100
rect 352398 36500 354798 37100
rect 357198 36500 358998 37100
rect 359798 36500 362398 37100
rect 364398 37100 365798 37700
rect 367598 37100 368798 37700
rect 372198 37700 376398 38100
rect 379998 37700 381398 38100
rect 381998 37700 383798 38100
rect 387598 37700 388998 38100
rect 389798 37700 391398 38100
rect 409724 37706 411524 38106
rect 364398 36500 365598 37100
rect 367998 36500 369198 37100
rect 258486 34556 259886 34956
rect 257686 33956 260686 34556
rect 257486 33356 260886 33956
rect 248686 32956 253686 33356
rect 256286 32956 261286 33356
rect 240486 32356 243086 32956
rect 244686 32356 247086 32956
rect 248686 32356 251086 32956
rect 252286 32356 253886 32956
rect 256286 32356 258686 32956
rect 259686 32356 261286 32956
rect 241086 31756 242286 32356
rect 245486 31756 246486 32356
rect 241486 31356 242286 31756
rect 245286 31356 246486 31756
rect 248686 31756 250686 32356
rect 252686 31756 254086 32356
rect 248686 31356 250286 31756
rect 252886 31356 254086 31756
rect 256286 31756 258286 32356
rect 260086 31756 261486 32356
rect 241486 30756 242686 31356
rect 245286 30756 246286 31356
rect 241686 30356 242686 30756
rect 241686 29756 242886 30356
rect 241886 29156 242886 29756
rect 245086 29756 246286 30756
rect 248686 30356 250086 31356
rect 253086 30756 254286 31356
rect 253486 30356 254286 30756
rect 256286 30756 257686 31756
rect 260286 31356 261886 31756
rect 260686 30756 261886 31356
rect 256286 30356 257486 30756
rect 260886 30356 261886 30756
rect 297198 30900 297798 36500
rect 300198 36100 301598 36500
rect 349398 36100 350798 36500
rect 352998 36100 354798 36500
rect 300398 35500 301998 36100
rect 300998 35100 301998 35500
rect 349198 35500 350598 36100
rect 353198 35500 354798 36100
rect 356798 36100 358598 36500
rect 360398 36100 362398 36500
rect 356798 35500 357998 36100
rect 360998 35500 362398 36100
rect 349198 35100 350398 35500
rect 353598 35100 354798 35500
rect 356598 35100 357798 35500
rect 300998 34500 302198 35100
rect 305998 34500 307598 35100
rect 313598 34500 315198 35100
rect 321398 34500 322998 35100
rect 336398 34500 337998 35100
rect 301198 33500 302198 34500
rect 305198 33900 308398 34500
rect 312998 33900 315798 34500
rect 316118 33900 316798 34500
rect 304798 33500 308598 33900
rect 312398 33500 316798 33900
rect 300998 32900 302198 33500
rect 304598 32900 309198 33500
rect 312198 32900 316798 33500
rect 318198 33500 320198 34500
rect 320598 33900 323598 34500
rect 320518 33500 323998 33900
rect 318198 32900 324198 33500
rect 327198 32900 329798 34500
rect 300998 32500 301998 32900
rect 300798 31900 301998 32500
rect 304398 32500 306198 32900
rect 307398 32500 309398 32900
rect 304398 31900 305798 32500
rect 307998 31900 309398 32500
rect 311998 32500 313598 32900
rect 315198 32500 316798 32900
rect 318398 32500 321598 32900
rect 322798 32500 324398 32900
rect 327398 32500 329798 32900
rect 333798 33900 335198 34500
rect 335798 33900 338398 34500
rect 348998 33900 350198 35100
rect 353798 33900 354798 35100
rect 333798 32900 338798 33900
rect 348798 33500 349998 33900
rect 353998 33500 354798 33900
rect 356398 33900 357598 35100
rect 361198 34500 362398 35500
rect 363998 36100 365198 36500
rect 363998 35100 364998 36100
rect 364398 34500 364798 35100
rect 333798 32500 336398 32900
rect 337598 32500 339198 32900
rect 311998 31900 313198 32500
rect 315598 31900 316798 32500
rect 300198 31300 301998 31900
rect 298998 30900 301598 31300
rect 303998 30900 305198 31900
rect 308398 30900 309598 31900
rect 311998 30900 312998 31900
rect 315798 30900 316798 31900
rect 245086 29156 245886 29756
rect 241886 28756 243086 29156
rect 242086 27756 243086 28756
rect 244686 28756 245886 29156
rect 248686 29156 249886 30356
rect 253486 29156 254686 30356
rect 244686 28156 245686 28756
rect 244486 27756 245686 28156
rect 248686 27756 249486 29156
rect 233886 26156 235086 26556
rect 237886 26156 238686 27756
rect 242086 27156 243286 27756
rect 244486 27156 245486 27756
rect 242286 26556 243286 27156
rect 244286 26556 245486 27156
rect 242286 26156 243486 26556
rect 222486 25556 223686 26156
rect 222286 25156 223686 25556
rect 221886 24556 223686 25156
rect 234286 25556 235086 26156
rect 237486 25556 238686 26156
rect 242686 25556 243486 26156
rect 244286 25556 245286 26556
rect 234286 25156 235486 25556
rect 237486 25156 238486 25556
rect 242686 25156 243886 25556
rect 234286 24556 235686 25156
rect 237286 24556 238486 25156
rect 242886 24556 243886 25156
rect 244206 25156 245286 25556
rect 248686 26156 249886 27756
rect 253686 27156 254686 29156
rect 253486 26556 254686 27156
rect 256286 26556 257286 30356
rect 260886 29756 262086 30356
rect 261086 26556 262086 29756
rect 253486 26156 254286 26556
rect 248686 25556 250086 26156
rect 248686 25156 250286 25556
rect 253086 25156 254286 26156
rect 256286 25556 257486 26556
rect 260886 26156 262086 26556
rect 297198 30300 301398 30900
rect 303798 30300 304998 30900
rect 308598 30300 309798 30900
rect 311998 30300 313198 30900
rect 315998 30300 316798 30900
rect 319198 31900 321198 32500
rect 323198 31900 324798 32500
rect 319198 31300 320798 31900
rect 323598 31300 324798 31900
rect 319198 30900 320598 31300
rect 323798 30900 324998 31300
rect 319198 30300 320398 30900
rect 297198 29900 300998 30300
rect 303798 29900 304798 30300
rect 308798 29900 309798 30300
rect 297198 29300 300798 29900
rect 256286 25156 257686 25556
rect 260686 25156 261886 26156
rect 244206 24556 245086 25156
rect 218286 23956 219486 24556
rect 221486 23956 223686 24556
rect 234486 23956 235886 24556
rect 237086 23956 238286 24556
rect 242886 23956 245086 24556
rect 248686 24556 250486 25156
rect 252686 24556 254086 25156
rect 256286 24556 257886 25156
rect 260286 24556 261486 25156
rect 248686 23956 250686 24556
rect 252486 23956 253886 24556
rect 256286 23956 258286 24556
rect 259886 23956 261486 24556
rect 297198 24100 297798 29300
rect 299198 28700 300998 29300
rect 299798 28300 301198 28700
rect 299998 27700 301398 28300
rect 303798 27700 309798 29900
rect 312198 29900 313998 30300
rect 312198 29300 315598 29900
rect 312398 28700 315998 29300
rect 312998 28300 316598 28700
rect 314198 27700 316798 28300
rect 300198 27100 301598 27700
rect 300398 26700 301598 27100
rect 303798 26700 304798 27700
rect 315398 27100 316998 27700
rect 315798 26700 316998 27100
rect 300798 26100 301998 26700
rect 303798 26100 304998 26700
rect 311798 26100 312398 26700
rect 300998 25100 302198 26100
rect 303998 25100 305198 26100
rect 309198 25100 309598 25700
rect 311798 25100 312798 26100
rect 315998 25100 316998 26700
rect 301198 24100 302398 25100
rect 304398 24500 305798 25100
rect 308798 24500 309798 25100
rect 304398 24100 305998 24500
rect 308198 24100 309798 24500
rect 181086 22956 186286 23956
rect 189086 23556 194286 23956
rect 196286 23556 201486 23956
rect 203886 23556 209286 23956
rect 189286 22956 194086 23556
rect 196086 22956 201886 23556
rect 204486 22956 209086 23556
rect 181086 22556 181766 22956
rect 182086 22556 185686 22956
rect 189886 22556 193686 22956
rect 196286 22556 201886 22956
rect 204686 22556 208486 22956
rect 210686 22556 213286 23956
rect 214686 23556 216886 23956
rect 218686 23556 220286 23956
rect 220606 23556 224686 23956
rect 234486 23556 238286 23956
rect 214686 22556 217086 23556
rect 218686 22956 224686 23556
rect 234686 22956 238086 23556
rect 243086 22956 244686 23956
rect 247686 23556 253886 23956
rect 255286 23556 261286 23956
rect 218886 22556 222286 22956
rect 222686 22556 224686 22956
rect 234886 22556 237886 22956
rect 243086 22556 244486 22956
rect 247686 22556 249486 23556
rect 249886 22956 253686 23556
rect 250086 22556 253086 22956
rect 255086 22556 257086 23556
rect 257406 22956 261086 23556
rect 296198 23500 298998 24100
rect 301398 23500 303198 24100
rect 304598 23500 309798 24100
rect 311798 24500 312998 25100
rect 315798 24500 316998 25100
rect 311798 24100 313198 24500
rect 315598 24100 316998 24500
rect 319198 27100 320198 30300
rect 323998 29300 324998 30900
rect 324198 28700 324998 29300
rect 324198 28300 325198 28700
rect 319198 26700 320398 27100
rect 323998 26700 324998 28300
rect 319198 25700 320598 26700
rect 323798 26100 324998 26700
rect 323598 25700 324798 26100
rect 319198 25100 321198 25700
rect 323198 25100 324798 25700
rect 319198 24500 321398 25100
rect 322798 24500 324398 25100
rect 319198 24100 324198 24500
rect 328998 24100 329798 32500
rect 334598 31900 336198 32500
rect 337998 31900 339198 32500
rect 334598 31300 335998 31900
rect 338198 31300 339398 31900
rect 334598 30900 335798 31300
rect 334598 24100 335598 30900
rect 338398 24100 339398 31300
rect 341598 29300 347198 31300
rect 348798 27700 349598 33500
rect 354198 32900 354518 33500
rect 356398 32900 357398 33900
rect 361398 33500 362398 34500
rect 368198 33500 369198 36500
rect 361598 32900 362198 33500
rect 367998 32900 369198 33500
rect 372198 33500 373198 37700
rect 379598 37100 381198 37700
rect 382598 37100 383798 37700
rect 387398 37100 388598 37700
rect 390198 37100 391398 37700
rect 409324 37106 410924 37706
rect 379598 36500 380798 37100
rect 382798 36500 383998 37100
rect 387398 36500 388398 37100
rect 390398 36500 391598 37100
rect 409124 36506 410724 37106
rect 379398 35500 380598 36500
rect 382998 36100 383998 36500
rect 387198 36100 388398 36500
rect 390798 36100 391598 36500
rect 408724 36106 410524 36506
rect 379398 34500 380398 35500
rect 382998 35100 384198 36100
rect 379198 33900 380398 34500
rect 373598 33500 375398 33900
rect 372198 32900 375798 33500
rect 356198 27700 357198 32900
rect 367598 32500 368798 32900
rect 367398 31900 368798 32500
rect 372198 32500 375998 32900
rect 372198 31900 376398 32500
rect 367198 31300 368598 31900
rect 372198 31300 373598 31900
rect 375198 31300 376598 31900
rect 366998 30900 368398 31300
rect 372198 30900 373198 31300
rect 375398 30900 376798 31300
rect 366798 30300 368198 30900
rect 375598 30300 376798 30900
rect 366398 29900 367998 30300
rect 375798 29900 376798 30300
rect 366198 29300 367598 29900
rect 375998 29300 376798 29900
rect 365998 28700 367398 29300
rect 365798 28300 367198 28700
rect 365598 27700 366998 28300
rect 348798 27100 349998 27700
rect 348998 26700 349998 27100
rect 356398 26700 357398 27700
rect 365198 27100 366798 27700
rect 364998 26700 366398 27100
rect 375998 26700 376998 29300
rect 379198 27700 380198 33900
rect 383198 33500 384198 35100
rect 383598 29300 384198 33500
rect 387198 32500 387998 36100
rect 390798 35500 391998 36100
rect 408524 35506 410324 36106
rect 390998 33900 391998 35500
rect 408124 34906 409724 35506
rect 407924 34506 409524 34906
rect 407524 33906 409324 34506
rect 390998 33500 392198 33900
rect 407124 33506 409124 33906
rect 390798 32500 392198 33500
rect 406924 32906 408524 33506
rect 387198 31900 388398 32500
rect 390398 31900 392198 32500
rect 406724 32306 408324 32906
rect 406324 31906 408124 32306
rect 387398 31300 388598 31900
rect 390198 31300 392198 31900
rect 405924 31306 407524 31906
rect 387398 30900 388798 31300
rect 389998 30900 392198 31300
rect 405724 30906 407324 31306
rect 387598 30300 392198 30900
rect 405524 30306 407124 30906
rect 387598 29900 390998 30300
rect 387998 29300 390798 29900
rect 391318 29580 392198 30300
rect 405124 29706 406924 30306
rect 348998 26100 350198 26700
rect 354198 26100 354998 26700
rect 356398 26100 357598 26700
rect 361998 26100 362398 26700
rect 364798 26100 366198 26700
rect 348998 25700 350398 26100
rect 353998 25700 354998 26100
rect 349198 25100 350398 25700
rect 353798 25100 354998 25700
rect 356598 25700 357798 26100
rect 361398 25700 362398 26100
rect 364598 25700 365998 26100
rect 375798 25700 376798 26700
rect 379398 26100 380398 27700
rect 383198 26700 384198 29300
rect 388398 28700 390198 29300
rect 391198 28700 392198 29580
rect 404924 29306 406724 29706
rect 404524 28706 406124 29306
rect 390998 28300 392198 28700
rect 404324 28306 405924 28706
rect 390998 27100 391998 28300
rect 403924 27706 405724 28306
rect 403724 27106 405124 27706
rect 390798 26700 391998 27100
rect 403324 26706 404924 27106
rect 379398 25700 380598 26100
rect 382998 25700 384198 26700
rect 390398 26100 391598 26700
rect 403124 26106 404724 26706
rect 390198 25700 391598 26100
rect 402724 25706 404524 26106
rect 356598 25100 357998 25700
rect 361198 25100 362398 25700
rect 364398 25100 365798 25700
rect 371598 25100 372398 25700
rect 375598 25100 376798 25700
rect 379598 25100 380598 25700
rect 349398 24500 350798 25100
rect 353598 24500 354998 25100
rect 356798 24500 358398 25100
rect 360998 24500 362398 25100
rect 363998 24500 365598 25100
rect 368398 24500 369198 25100
rect 371598 24500 372998 25100
rect 375398 24500 376598 25100
rect 379598 24500 380798 25100
rect 382798 24500 383998 25700
rect 389998 25100 391398 25700
rect 402324 25106 403924 25706
rect 389798 24500 391198 25100
rect 402124 24506 403724 25106
rect 349598 24100 351198 24500
rect 352998 24100 354798 24500
rect 357198 24100 358798 24500
rect 360798 24100 362198 24500
rect 363798 24100 365198 24500
rect 368398 24100 369398 24500
rect 371598 24100 373198 24500
rect 374798 24100 376598 24500
rect 379998 24100 381198 24500
rect 382598 24100 383798 24500
rect 389198 24100 391198 24500
rect 401924 24106 403524 24506
rect 311798 23500 314398 24100
rect 314718 23500 316798 24100
rect 295998 23100 299198 23500
rect 257486 22556 260886 22956
rect 182686 21956 185286 22556
rect 190286 21956 192886 22556
rect 205086 21956 208086 22556
rect 219286 21956 221686 22556
rect 235486 21956 237286 22556
rect 250486 21956 252686 22556
rect 257886 21956 260286 22556
rect 296198 22500 299198 23100
rect 301598 22500 303398 23500
rect 304798 23100 309598 23500
rect 311798 23100 316598 23500
rect 319198 23180 320078 24100
rect 320398 23500 323998 24100
rect 305198 22500 309198 23100
rect 311798 22500 316398 23100
rect 305798 21900 308398 22500
rect 313198 21900 315798 22500
rect 319198 18900 320198 23180
rect 320598 23100 323798 23500
rect 321198 22500 322998 23100
rect 326598 22500 332198 24100
rect 333598 22500 336198 24100
rect 337598 22500 339998 24100
rect 349998 23500 351998 24100
rect 352398 23500 354398 24100
rect 357398 23500 359598 24100
rect 359918 23500 361998 24100
rect 350198 23100 354198 23500
rect 357598 23100 361598 23500
rect 350398 22500 353798 23100
rect 357798 22500 361398 23100
rect 363798 22500 369398 24100
rect 371798 23500 376398 24100
rect 379998 23500 383598 24100
rect 371998 23100 375998 23500
rect 380198 23100 383598 23500
rect 387198 23500 390798 24100
rect 401524 23506 403124 24106
rect 387198 23100 390398 23500
rect 372398 22500 375798 23100
rect 380398 22500 382998 23100
rect 387198 22500 389998 23100
rect 401124 22906 402724 23506
rect 400924 22506 402524 22906
rect 350798 21900 353198 22500
rect 358398 21900 360998 22500
rect 372998 21900 375398 22500
rect 380798 21900 382798 22500
rect 387398 21900 389598 22500
rect 400724 21906 402324 22506
rect 400124 21506 401924 21906
rect 399924 20906 401524 21506
rect 399724 20306 401324 20906
rect 399524 19906 401124 20306
rect 398924 19306 400724 19906
rect 398724 18906 400324 19306
rect 318198 17300 321598 18900
rect 398524 18306 400124 18906
rect 397924 17706 399724 18306
rect 397724 17306 399524 17706
rect 394924 16306 395324 17306
rect 397524 16706 399124 17306
rect 397324 16306 398924 16706
rect 394724 15106 395324 16306
rect 396724 15706 398524 16306
rect 396524 15106 398324 15706
rect 394324 14106 395524 15106
rect 396324 14706 397924 15106
rect 396124 14106 397724 14706
rect 394124 13706 397324 14106
rect 393924 13106 397124 13706
rect 393924 12506 396724 13106
rect 393724 12106 396324 12506
rect 393724 11506 396524 12106
rect 393524 10906 396724 11506
rect 393524 10506 397324 10906
rect 393124 9906 397524 10506
rect 393124 9506 397324 9906
rect 392924 8906 396524 9506
rect 392724 8306 395524 8906
rect 392724 7906 394724 8306
rect 392524 7306 393924 7906
rect 392524 6906 392924 7306
use array_SR  array_SR_0
timestamp 1758232856
transform 1 0 149469 0 1 114190
box -21072 586 308046 327366
use bias  bias_1
timestamp 1758232856
transform 1 0 289348 0 1 473566
box 790 -2236 7180 -220
use opamp_wrapper  opamp_wrapper_0
timestamp 1758232856
transform 1 0 464481 0 1 129134
box -2280 -2669 27441 13665
use opamp_wrapper  opamp_wrapper_1
timestamp 1758232856
transform 1 0 309932 0 1 580259
box -2280 -2669 27441 13665
use pixel_array  pixel_array_0
timestamp 1758232856
transform 1 0 294314 0 1 588742
box -3720 -8600 11230 5820
use sky130_fd_pr__res_generic_m3_3NNQKJ  sky130_fd_pr__res_generic_m3_3NNQKJ_0
timestamp 1758069660
transform 0 1 582837 -1 0 364836
box -50 -107 50 107
use sky130_fd_pr__res_generic_m3_3NNQKJ  sky130_fd_pr__res_generic_m3_3NNQKJ_1
timestamp 1758069660
transform 0 1 767 -1 0 462426
box -50 -107 50 107
<< labels >>
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
